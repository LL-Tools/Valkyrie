

module b17_C_AntiSAT_k_128_2 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936;

  XNOR2_X1 U11084 ( .A(n14259), .B(n12243), .ZN(n14216) );
  AND2_X1 U11085 ( .A1(n15286), .A2(n9757), .ZN(n16294) );
  CLKBUF_X1 U11086 ( .A(n11500), .Z(n12155) );
  INV_X2 U11087 ( .A(n17770), .ZN(n17758) );
  NAND2_X1 U11088 ( .A1(n11717), .A2(n20108), .ZN(n11748) );
  XNOR2_X1 U11089 ( .A(n11671), .B(n11670), .ZN(n11697) );
  NAND2_X1 U11090 ( .A1(n10460), .A2(n10500), .ZN(n10695) );
  NOR2_X1 U11091 ( .A1(n11704), .A2(n20644), .ZN(n12288) );
  AND2_X1 U11092 ( .A1(n10512), .A2(n12734), .ZN(n12719) );
  INV_X1 U11093 ( .A(n15393), .ZN(n15517) );
  AND2_X1 U11094 ( .A1(n12734), .A2(n10513), .ZN(n10580) );
  CLKBUF_X1 U11096 ( .A(n15339), .Z(n17187) );
  CLKBUF_X2 U11097 ( .A(n11870), .Z(n12221) );
  CLKBUF_X2 U11098 ( .A(n11911), .Z(n12223) );
  CLKBUF_X2 U11099 ( .A(n11473), .Z(n12069) );
  BUF_X1 U11100 ( .A(n10390), .Z(n13931) );
  CLKBUF_X2 U11101 ( .A(n10637), .Z(n9665) );
  INV_X2 U11102 ( .A(n13763), .ZN(n10374) );
  OR2_X1 U11103 ( .A1(n11432), .A2(n11431), .ZN(n13278) );
  BUF_X1 U11104 ( .A(n11474), .Z(n12199) );
  NAND4_X2 U11105 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(
        n11548) );
  AND2_X1 U11106 ( .A1(n13261), .A2(n14751), .ZN(n11595) );
  AND2_X1 U11107 ( .A1(n13258), .A2(n14751), .ZN(n11579) );
  AND2_X1 U11108 ( .A1(n13258), .A2(n11420), .ZN(n11911) );
  AND2_X1 U11109 ( .A1(n11418), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13258) );
  INV_X2 U11110 ( .A(n12882), .ZN(n9668) );
  AND2_X2 U11111 ( .A1(n10519), .A2(n13614), .ZN(n9644) );
  NAND3_X1 U11112 ( .A1(n9847), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12861) );
  NAND2_X1 U11113 ( .A1(n20143), .A2(n11548), .ZN(n12295) );
  INV_X1 U11114 ( .A(n10175), .ZN(n10181) );
  AND2_X2 U11115 ( .A1(n10519), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10524) );
  NOR2_X1 U11116 ( .A1(n17847), .A2(n15530), .ZN(n15531) );
  OR2_X1 U11117 ( .A1(n18649), .A2(n14180), .ZN(n17140) );
  AND3_X1 U11118 ( .A1(n10646), .A2(n10684), .A3(n10034), .ZN(n10791) );
  INV_X1 U11119 ( .A(n13559), .ZN(n12724) );
  AND2_X1 U11120 ( .A1(n10524), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10763) );
  INV_X1 U11121 ( .A(n12714), .ZN(n12697) );
  INV_X1 U11122 ( .A(n9665), .ZN(n13227) );
  XNOR2_X1 U11123 ( .A(n10986), .B(n10985), .ZN(n10984) );
  INV_X1 U11124 ( .A(n15393), .ZN(n9642) );
  CLKBUF_X3 U11125 ( .A(n15485), .Z(n9647) );
  INV_X1 U11126 ( .A(n14256), .ZN(n12421) );
  AND4_X1 U11127 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n11518) );
  NAND2_X1 U11128 ( .A1(n20124), .A2(n13402), .ZN(n20739) );
  INV_X1 U11129 ( .A(n13402), .ZN(n20107) );
  NAND2_X2 U11130 ( .A1(n10294), .A2(n13763), .ZN(n12987) );
  NAND2_X1 U11131 ( .A1(n11201), .A2(n11200), .ZN(n12546) );
  OR2_X1 U11132 ( .A1(n15059), .A2(n14841), .ZN(n14843) );
  NAND2_X1 U11133 ( .A1(n15258), .A2(n13753), .ZN(n13777) );
  NAND2_X1 U11134 ( .A1(n10374), .A2(n9667), .ZN(n11106) );
  XNOR2_X1 U11135 ( .A(n9885), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16352) );
  NAND2_X1 U11136 ( .A1(n20913), .A2(n18815), .ZN(n16905) );
  OR2_X1 U11137 ( .A1(n14951), .A2(n14939), .ZN(n14941) );
  NOR2_X1 U11138 ( .A1(n15257), .A2(n15256), .ZN(n15258) );
  INV_X1 U11139 ( .A(n19989), .ZN(n19995) );
  AOI211_X1 U11140 ( .C1(n15871), .C2(n14613), .A(n14612), .B(n14611), .ZN(
        n14614) );
  AOI21_X1 U11141 ( .B1(n16202), .B2(n9895), .A(n9893), .ZN(n15626) );
  INV_X1 U11142 ( .A(n13827), .ZN(n10500) );
  BUF_X1 U11143 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n18649) );
  INV_X2 U11144 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18798) );
  AND2_X2 U11145 ( .A1(n13255), .A2(n13273), .ZN(n13397) );
  NAND3_X2 U11146 ( .A1(n11554), .A2(n11549), .A3(n20124), .ZN(n13255) );
  BUF_X4 U11147 ( .A(n14106), .Z(n17188) );
  NAND2_X2 U11148 ( .A1(n14455), .A2(n9762), .ZN(n12063) );
  AND2_X4 U11149 ( .A1(n14329), .A2(n11993), .ZN(n14455) );
  NAND2_X2 U11150 ( .A1(n9944), .A2(n10742), .ZN(n10959) );
  NOR2_X4 U11151 ( .A1(n15009), .A2(n9971), .ZN(n14966) );
  XNOR2_X2 U11152 ( .A(n12315), .B(n12316), .ZN(n13377) );
  NOR2_X2 U11153 ( .A1(n16251), .A2(n9858), .ZN(n16228) );
  AND2_X2 U11155 ( .A1(n10519), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9640) );
  AND2_X4 U11156 ( .A1(n13258), .A2(n14752), .ZN(n11500) );
  NOR2_X2 U11157 ( .A1(n16209), .A2(n16277), .ZN(n16203) );
  BUF_X2 U11158 ( .A(n14999), .Z(n9641) );
  XNOR2_X2 U11159 ( .A(n12610), .B(n12607), .ZN(n13373) );
  AOI21_X2 U11160 ( .B1(n10181), .B2(n10178), .A(n9712), .ZN(n10177) );
  BUF_X4 U11161 ( .A(n10443), .Z(n10993) );
  OAI211_X2 U11162 ( .C1(n11061), .C2(n10638), .A(n10445), .B(n10444), .ZN(
        n10985) );
  AOI211_X2 U11163 ( .C1(n20068), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14631), .B(n14630), .ZN(n14632) );
  XNOR2_X1 U11164 ( .A(n10459), .B(n10458), .ZN(n13827) );
  XNOR2_X2 U11165 ( .A(n10783), .B(n15313), .ZN(n15111) );
  NAND2_X2 U11166 ( .A1(n10782), .A2(n19025), .ZN(n10783) );
  AND2_X1 U11167 ( .A1(n10519), .A2(n13614), .ZN(n9643) );
  INV_X1 U11168 ( .A(n9643), .ZN(n9645) );
  AND2_X1 U11169 ( .A1(n10519), .A2(n13614), .ZN(n10518) );
  NOR2_X2 U11170 ( .A1(n9789), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13617) );
  OAI21_X1 U11171 ( .B1(n16360), .B2(n9816), .A(n9815), .ZN(n9814) );
  OR2_X1 U11172 ( .A1(n17551), .A2(n17758), .ZN(n17545) );
  XNOR2_X1 U11173 ( .A(n12520), .B(n12519), .ZN(n14711) );
  NAND2_X1 U11174 ( .A1(n16294), .A2(n15253), .ZN(n15254) );
  AND2_X1 U11175 ( .A1(n11698), .A2(n11697), .ZN(n11717) );
  XNOR2_X1 U11176 ( .A(n11681), .B(n12314), .ZN(n20185) );
  BUF_X1 U11177 ( .A(n13827), .Z(n13613) );
  NOR2_X1 U11178 ( .A1(n17239), .A2(n17370), .ZN(n17312) );
  INV_X4 U11179 ( .A(n16861), .ZN(n16909) );
  OAI21_X2 U11180 ( .B1(n15697), .B2(n17428), .A(n15696), .ZN(n17384) );
  INV_X2 U11181 ( .A(n17997), .ZN(n18657) );
  CLKBUF_X2 U11182 ( .A(n17455), .Z(n9649) );
  AND2_X1 U11183 ( .A1(n10654), .A2(n10655), .ZN(n10653) );
  AND2_X2 U11184 ( .A1(n12940), .A2(n10150), .ZN(n10973) );
  NAND2_X1 U11185 ( .A1(n10405), .A2(n10389), .ZN(n10407) );
  INV_X1 U11186 ( .A(n10386), .ZN(n11186) );
  NAND2_X1 U11187 ( .A1(n11106), .A2(n12987), .ZN(n13049) );
  AOI21_X1 U11188 ( .B1(n10134), .B2(n9695), .A(n17848), .ZN(n17847) );
  BUF_X1 U11189 ( .A(n10370), .Z(n13936) );
  CLKBUF_X1 U11190 ( .A(n10373), .Z(n12586) );
  NOR2_X1 U11191 ( .A1(n18195), .A2(n18841), .ZN(n15603) );
  NAND2_X1 U11192 ( .A1(n10369), .A2(n10368), .ZN(n13941) );
  NAND2_X1 U11193 ( .A1(n12951), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12952) );
  INV_X1 U11194 ( .A(n10373), .ZN(n9646) );
  NAND2_X1 U11195 ( .A1(n10307), .A2(n10306), .ZN(n10637) );
  BUF_X2 U11196 ( .A(n11941), .Z(n11927) );
  BUF_X2 U11197 ( .A(n11479), .Z(n9659) );
  BUF_X2 U11198 ( .A(n12215), .Z(n12068) );
  BUF_X2 U11199 ( .A(n11579), .Z(n12222) );
  CLKBUF_X2 U11200 ( .A(n11611), .Z(n12214) );
  INV_X4 U11201 ( .A(n17140), .ZN(n17181) );
  CLKBUF_X3 U11202 ( .A(n15484), .Z(n9654) );
  CLKBUF_X2 U11203 ( .A(n12887), .Z(n12915) );
  CLKBUF_X1 U11204 ( .A(n12814), .Z(n9671) );
  CLKBUF_X2 U11205 ( .A(n15355), .Z(n17097) );
  CLKBUF_X2 U11206 ( .A(n15482), .Z(n17110) );
  CLKBUF_X3 U11207 ( .A(n12739), .Z(n9661) );
  NAND3_X2 U11208 ( .A1(n9847), .A2(n9846), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12882) );
  AND3_X2 U11209 ( .A1(n9789), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12739) );
  INV_X2 U11210 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11419) );
  INV_X2 U11211 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9789) );
  OAI211_X1 U11212 ( .C1(n10217), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n12541) );
  OR2_X1 U11213 ( .A1(n12584), .A2(n16317), .ZN(n10252) );
  XNOR2_X1 U11214 ( .A(n14234), .B(n14233), .ZN(n14240) );
  NAND2_X1 U11215 ( .A1(n10217), .A2(n10212), .ZN(n10214) );
  AOI22_X1 U11216 ( .A1(n15931), .A2(n20090), .B1(n20089), .B2(n15930), .ZN(
        n15937) );
  OR2_X1 U11217 ( .A1(n10904), .A2(n11091), .ZN(n10905) );
  NAND2_X1 U11218 ( .A1(n12574), .A2(n10213), .ZN(n10217) );
  OR2_X1 U11219 ( .A1(n14968), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15121) );
  NAND2_X1 U11220 ( .A1(n9874), .A2(n10027), .ZN(n12574) );
  OR2_X1 U11221 ( .A1(n11072), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10233) );
  OR2_X1 U11222 ( .A1(n15067), .A2(n9760), .ZN(n9914) );
  OAI21_X1 U11223 ( .B1(n16290), .B2(n16330), .A(n9863), .ZN(n9862) );
  AND2_X1 U11224 ( .A1(n11072), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12558) );
  NOR2_X1 U11225 ( .A1(n9704), .A2(n9922), .ZN(n9921) );
  XNOR2_X1 U11226 ( .A(n10903), .B(n11091), .ZN(n14968) );
  NAND2_X1 U11227 ( .A1(n11090), .A2(n9718), .ZN(n10903) );
  OR2_X1 U11228 ( .A1(n11090), .A2(n10026), .ZN(n9874) );
  NAND2_X1 U11229 ( .A1(n15269), .A2(n9860), .ZN(n16241) );
  INV_X1 U11230 ( .A(n14500), .ZN(n14580) );
  NAND2_X1 U11231 ( .A1(n10069), .A2(n10070), .ZN(n14500) );
  AND2_X1 U11232 ( .A1(n9941), .A2(n9943), .ZN(n15088) );
  AND2_X1 U11233 ( .A1(n9798), .A2(n9726), .ZN(n14589) );
  NAND2_X1 U11234 ( .A1(n14974), .A2(n14976), .ZN(n11090) );
  CLKBUF_X1 U11235 ( .A(n15009), .Z(n15187) );
  NOR2_X1 U11236 ( .A1(n9726), .A2(n14586), .ZN(n14574) );
  OAI21_X1 U11237 ( .B1(n9799), .B2(n9784), .A(n15874), .ZN(n9798) );
  OAI21_X1 U11238 ( .B1(n15001), .B2(n19236), .A(n9851), .ZN(n9850) );
  INV_X1 U11239 ( .A(n10070), .ZN(n14259) );
  XNOR2_X1 U11240 ( .A(n12852), .B(n12849), .ZN(n14803) );
  CLKBUF_X1 U11241 ( .A(n15035), .Z(n15036) );
  OR2_X1 U11242 ( .A1(n14413), .A2(n14294), .ZN(n15817) );
  AND2_X1 U11243 ( .A1(n10815), .A2(n16232), .ZN(n10873) );
  INV_X1 U11244 ( .A(n15837), .ZN(n15732) );
  NAND2_X1 U11245 ( .A1(n9926), .A2(n9927), .ZN(n10815) );
  NAND2_X1 U11247 ( .A1(n9817), .A2(n9814), .ZN(n16398) );
  NAND2_X1 U11248 ( .A1(n10075), .A2(n10071), .ZN(n16172) );
  OR2_X1 U11249 ( .A1(n12761), .A2(n12782), .ZN(n10245) );
  NAND2_X1 U11250 ( .A1(n10182), .A2(n10184), .ZN(n15886) );
  AND2_X1 U11251 ( .A1(n10185), .A2(n15890), .ZN(n10184) );
  NAND2_X1 U11252 ( .A1(n9900), .A2(n9721), .ZN(n10175) );
  NAND2_X1 U11253 ( .A1(n12976), .A2(n12977), .ZN(n14245) );
  NOR2_X1 U11254 ( .A1(n10964), .A2(n10801), .ZN(n10963) );
  NOR2_X1 U11255 ( .A1(n16114), .A2(n16113), .ZN(n16112) );
  NAND2_X1 U11256 ( .A1(n10012), .A2(n10011), .ZN(n13794) );
  OR2_X1 U11257 ( .A1(n10959), .A2(n10958), .ZN(n10964) );
  XNOR2_X1 U11258 ( .A(n12977), .B(n12548), .ZN(n16102) );
  AND2_X1 U11259 ( .A1(n15891), .A2(n15898), .ZN(n10183) );
  NAND2_X1 U11260 ( .A1(n9901), .A2(n16056), .ZN(n12388) );
  AND2_X1 U11261 ( .A1(n10172), .A2(n10171), .ZN(n16120) );
  XNOR2_X1 U11262 ( .A(n12356), .B(n12355), .ZN(n15898) );
  INV_X1 U11263 ( .A(n10945), .ZN(n9944) );
  OR2_X1 U11264 ( .A1(n15849), .A2(n15846), .ZN(n9906) );
  NOR2_X2 U11265 ( .A1(n9693), .A2(n14865), .ZN(n14867) );
  AND2_X1 U11266 ( .A1(n9969), .A2(n10941), .ZN(n9968) );
  NAND2_X1 U11267 ( .A1(n9796), .A2(n12354), .ZN(n12356) );
  NAND2_X1 U11268 ( .A1(n10230), .A2(n10231), .ZN(n10694) );
  INV_X1 U11269 ( .A(n9855), .ZN(n10742) );
  NOR2_X1 U11270 ( .A1(n9833), .A2(n9830), .ZN(n15949) );
  NAND2_X1 U11271 ( .A1(n9853), .A2(n10735), .ZN(n9855) );
  AND2_X1 U11272 ( .A1(n10004), .A2(n16232), .ZN(n9883) );
  NAND2_X1 U11273 ( .A1(n12350), .A2(n12378), .ZN(n9796) );
  NAND2_X1 U11274 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  AND2_X1 U11275 ( .A1(n10781), .A2(n10780), .ZN(n10957) );
  AND2_X1 U11276 ( .A1(n11766), .A2(n11794), .ZN(n12350) );
  OAI21_X1 U11277 ( .B1(n10532), .B2(n9722), .A(n10531), .ZN(n10612) );
  NOR2_X1 U11278 ( .A1(n16153), .A2(n16154), .ZN(n16152) );
  NAND2_X1 U11279 ( .A1(n13306), .A2(n9790), .ZN(n13453) );
  XNOR2_X1 U11280 ( .A(n12382), .B(n11797), .ZN(n12372) );
  AND3_X1 U11281 ( .A1(n10483), .A2(n10482), .A3(n10481), .ZN(n10484) );
  AND2_X1 U11282 ( .A1(n10717), .A2(n10716), .ZN(n9854) );
  INV_X1 U11283 ( .A(n14702), .ZN(n20079) );
  OR2_X1 U11284 ( .A1(n10538), .A2(n10537), .ZN(n10267) );
  OAI22_X1 U11285 ( .A1(n10699), .A2(n10539), .B1(n13930), .B2(n10695), .ZN(
        n10540) );
  OR2_X1 U11286 ( .A1(n19361), .A2(n12858), .ZN(n10716) );
  OR2_X1 U11287 ( .A1(n14706), .A2(n20097), .ZN(n14702) );
  XNOR2_X1 U11288 ( .A(n12329), .B(n20082), .ZN(n13499) );
  XNOR2_X1 U11289 ( .A(n13294), .B(n13293), .ZN(n19872) );
  AND2_X1 U11290 ( .A1(n12606), .A2(n12605), .ZN(n13374) );
  OR2_X1 U11291 ( .A1(n19361), .A2(n12808), .ZN(n10485) );
  OR2_X1 U11292 ( .A1(n10707), .A2(n10549), .ZN(n10551) );
  OR2_X1 U11293 ( .A1(n10137), .A2(n17603), .ZN(n10136) );
  NAND2_X1 U11294 ( .A1(n9714), .A2(n10500), .ZN(n10699) );
  AND2_X1 U11295 ( .A1(n14423), .A2(n9984), .ZN(n14284) );
  AND2_X1 U11296 ( .A1(n13414), .A2(n13409), .ZN(n14706) );
  AND2_X1 U11297 ( .A1(n13414), .A2(n13400), .ZN(n20097) );
  AND2_X1 U11298 ( .A1(n15551), .A2(n17919), .ZN(n10137) );
  OAI21_X1 U11299 ( .B1(n13292), .B2(n13291), .A(n13293), .ZN(n12606) );
  OR2_X2 U11300 ( .A1(n10477), .A2(n10476), .ZN(n10541) );
  NAND2_X1 U11301 ( .A1(n12318), .A2(n12317), .ZN(n12329) );
  NOR2_X1 U11302 ( .A1(n17658), .A2(n15548), .ZN(n17654) );
  AND2_X1 U11303 ( .A1(n9703), .A2(n10454), .ZN(n10460) );
  INV_X2 U11304 ( .A(n14567), .ZN(n9648) );
  NAND2_X1 U11305 ( .A1(n9703), .A2(n10475), .ZN(n19301) );
  AND2_X1 U11306 ( .A1(n13311), .A2(n13310), .ZN(n13469) );
  NOR2_X1 U11307 ( .A1(n10464), .A2(n10461), .ZN(n9925) );
  NOR2_X1 U11308 ( .A1(n17779), .A2(n18090), .ZN(n17778) );
  NAND2_X1 U11309 ( .A1(n11626), .A2(n11639), .ZN(n11681) );
  AND2_X1 U11310 ( .A1(n10825), .A2(n10826), .ZN(n18917) );
  NAND2_X1 U11311 ( .A1(n10500), .A2(n19068), .ZN(n10476) );
  AOI21_X1 U11312 ( .B1(n13827), .B2(n10099), .A(n12604), .ZN(n13293) );
  NAND2_X1 U11313 ( .A1(n11716), .A2(n11715), .ZN(n20108) );
  NAND2_X1 U11314 ( .A1(n10102), .A2(n10468), .ZN(n19068) );
  NAND2_X1 U11315 ( .A1(n15545), .A2(n18090), .ZN(n17759) );
  AND2_X1 U11316 ( .A1(n10470), .A2(n10469), .ZN(n10493) );
  NAND2_X1 U11317 ( .A1(n17706), .A2(n17975), .ZN(n17659) );
  NAND2_X1 U11318 ( .A1(n9845), .A2(n12293), .ZN(n13386) );
  AND2_X1 U11319 ( .A1(n10468), .A2(n9737), .ZN(n10101) );
  NAND2_X1 U11320 ( .A1(n10098), .A2(n12591), .ZN(n12594) );
  XNOR2_X1 U11321 ( .A(n13530), .B(n20247), .ZN(n20711) );
  INV_X1 U11322 ( .A(n9826), .ZN(n15545) );
  NAND2_X1 U11323 ( .A1(n10459), .A2(n10438), .ZN(n9792) );
  CLKBUF_X1 U11324 ( .A(n10451), .Z(n10468) );
  NAND2_X1 U11325 ( .A1(n11243), .A2(n11242), .ZN(n15317) );
  OR2_X1 U11326 ( .A1(n17791), .A2(n15543), .ZN(n9826) );
  NAND2_X1 U11327 ( .A1(n10188), .A2(n10193), .ZN(n10189) );
  NAND2_X2 U11328 ( .A1(n12926), .A2(n16343), .ZN(n19078) );
  CLKBUF_X1 U11329 ( .A(n10450), .Z(n10453) );
  NAND2_X1 U11330 ( .A1(n10449), .A2(n10448), .ZN(n10469) );
  CLKBUF_X1 U11331 ( .A(n11688), .Z(n11689) );
  NAND2_X1 U11332 ( .A1(n19029), .A2(n18931), .ZN(n18916) );
  OR2_X1 U11333 ( .A1(n11650), .A2(n11651), .ZN(n11648) );
  AND2_X1 U11334 ( .A1(n9896), .A2(n11632), .ZN(n11635) );
  NOR2_X1 U11335 ( .A1(n11232), .A2(n10116), .ZN(n10119) );
  INV_X1 U11336 ( .A(n18623), .ZN(n18660) );
  XNOR2_X1 U11337 ( .A(n9896), .B(n11578), .ZN(n11688) );
  NAND2_X1 U11338 ( .A1(n10434), .A2(n10433), .ZN(n10457) );
  NOR2_X1 U11339 ( .A1(n15588), .A2(n17808), .ZN(n15590) );
  AND2_X1 U11340 ( .A1(n13973), .A2(n13972), .ZN(n14027) );
  NAND2_X1 U11341 ( .A1(n9795), .A2(n11565), .ZN(n9896) );
  INV_X2 U11342 ( .A(n17233), .ZN(n17219) );
  XNOR2_X1 U11343 ( .A(n11086), .B(n11085), .ZN(n12932) );
  INV_X2 U11344 ( .A(n11082), .ZN(n11079) );
  NAND2_X2 U11345 ( .A1(n18841), .A2(n17430), .ZN(n17478) );
  NAND2_X1 U11346 ( .A1(n10791), .A2(n10790), .ZN(n10799) );
  NAND2_X1 U11347 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  AND2_X1 U11348 ( .A1(n10653), .A2(n10032), .ZN(n10034) );
  NAND2_X1 U11349 ( .A1(n9805), .A2(n9701), .ZN(n9804) );
  INV_X1 U11350 ( .A(n11051), .ZN(n11061) );
  NAND2_X1 U11351 ( .A1(n15540), .A2(n17354), .ZN(n17770) );
  NOR3_X1 U11352 ( .A1(n15695), .A2(n18224), .A3(n14206), .ZN(n16516) );
  AND2_X2 U11353 ( .A1(n11169), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11051) );
  NAND2_X1 U11354 ( .A1(n10413), .A2(n11186), .ZN(n11028) );
  NOR2_X1 U11355 ( .A1(n14177), .A2(n15559), .ZN(n16515) );
  NOR2_X1 U11356 ( .A1(n10785), .A2(n10033), .ZN(n10032) );
  AND2_X1 U11357 ( .A1(n10645), .A2(n10650), .ZN(n10655) );
  MUX2_X1 U11358 ( .A(n10329), .B(n11137), .S(n13936), .Z(n10357) );
  XNOR2_X1 U11359 ( .A(n15531), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9805) );
  OR2_X1 U11360 ( .A1(n17363), .A2(n15516), .ZN(n15537) );
  NAND2_X1 U11361 ( .A1(n11202), .A2(n9665), .ZN(n11381) );
  AND2_X1 U11362 ( .A1(n13049), .A2(n10356), .ZN(n9892) );
  NOR2_X1 U11363 ( .A1(n12296), .A2(n11556), .ZN(n11572) );
  NAND2_X1 U11364 ( .A1(n11499), .A2(n11498), .ZN(n13244) );
  INV_X1 U11365 ( .A(n20739), .ZN(n13319) );
  AND3_X1 U11366 ( .A1(n11163), .A2(n10105), .A3(n10294), .ZN(n10106) );
  AND2_X1 U11367 ( .A1(n10395), .A2(n13763), .ZN(n10105) );
  NOR2_X1 U11368 ( .A1(n12987), .A2(n12960), .ZN(n10413) );
  INV_X1 U11369 ( .A(n13941), .ZN(n11163) );
  XOR2_X1 U11370 ( .A(n17380), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17859) );
  AND2_X2 U11371 ( .A1(n13402), .A2(n13422), .ZN(n13362) );
  AND3_X1 U11372 ( .A1(n10608), .A2(n10254), .A3(n10607), .ZN(n11228) );
  NAND2_X1 U11373 ( .A1(n20135), .A2(n11548), .ZN(n13088) );
  INV_X1 U11374 ( .A(n12295), .ZN(n11545) );
  OR2_X1 U11375 ( .A1(n11543), .A2(n20135), .ZN(n13087) );
  INV_X1 U11376 ( .A(n11672), .ZN(n13584) );
  NOR2_X4 U11377 ( .A1(n13402), .A2(n13422), .ZN(n14364) );
  AND2_X1 U11378 ( .A1(n13346), .A2(n13580), .ZN(n11672) );
  NAND2_X1 U11379 ( .A1(n10210), .A2(n10208), .ZN(n10373) );
  CLKBUF_X1 U11380 ( .A(n17611), .Z(n18570) );
  OR2_X2 U11381 ( .A1(n11452), .A2(n11451), .ZN(n11556) );
  OR2_X2 U11382 ( .A1(n11497), .A2(n11496), .ZN(n13580) );
  CLKBUF_X2 U11383 ( .A(n11542), .Z(n13346) );
  AND4_X1 U11384 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11521) );
  AND4_X1 U11385 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11540) );
  NOR2_X2 U11386 ( .A1(n20104), .A2(n20103), .ZN(n20105) );
  AND4_X1 U11387 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11539) );
  AND4_X1 U11388 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11538) );
  AND4_X1 U11389 ( .A1(n11513), .A2(n11512), .A3(n11511), .A4(n11510), .ZN(
        n11519) );
  AND4_X1 U11390 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11520) );
  AND4_X1 U11391 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11541) );
  AND4_X1 U11392 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n11472) );
  AND4_X1 U11393 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11471) );
  AND4_X1 U11394 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11469) );
  BUF_X2 U11395 ( .A(n9662), .Z(n17115) );
  NAND2_X2 U11396 ( .A1(n18832), .A2(n18718), .ZN(n18775) );
  INV_X2 U11397 ( .A(n18724), .ZN(n9650) );
  AND2_X2 U11398 ( .A1(n9671), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12700) );
  NAND2_X2 U11399 ( .A1(n19835), .A2(n19784), .ZN(n19838) );
  NAND2_X2 U11400 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19835), .ZN(n19834) );
  INV_X1 U11401 ( .A(n10300), .ZN(n9669) );
  CLKBUF_X2 U11402 ( .A(n15344), .Z(n16937) );
  INV_X1 U11403 ( .A(n9699), .ZN(n17053) );
  BUF_X2 U11404 ( .A(n15424), .Z(n9662) );
  BUF_X2 U11405 ( .A(n15339), .Z(n17092) );
  INV_X1 U11407 ( .A(n9671), .ZN(n9651) );
  AND2_X2 U11408 ( .A1(n18859), .A2(n12960), .ZN(n19044) );
  INV_X2 U11409 ( .A(n16507), .ZN(U215) );
  INV_X2 U11410 ( .A(n9657), .ZN(n9658) );
  BUF_X4 U11411 ( .A(n14111), .Z(n9653) );
  NOR2_X1 U11412 ( .A1(n17799), .A2(n17806), .ZN(n16745) );
  CLKBUF_X3 U11413 ( .A(n11474), .Z(n12216) );
  OR2_X1 U11414 ( .A1(n16905), .A2(n14085), .ZN(n15393) );
  INV_X1 U11415 ( .A(n18696), .ZN(n16908) );
  INV_X2 U11416 ( .A(n16511), .ZN(n16513) );
  NOR2_X1 U11417 ( .A1(n12961), .A2(n19228), .ZN(n12962) );
  AND2_X2 U11418 ( .A1(n11425), .A2(n11426), .ZN(n11479) );
  AND2_X2 U11419 ( .A1(n11420), .A2(n11426), .ZN(n11491) );
  NOR2_X1 U11420 ( .A1(n18801), .A2(n18700), .ZN(n18838) );
  INV_X2 U11421 ( .A(n12882), .ZN(n12887) );
  NAND2_X2 U11422 ( .A1(n10512), .A2(n13614), .ZN(n10300) );
  BUF_X2 U11423 ( .A(n12739), .Z(n9660) );
  INV_X2 U11424 ( .A(n12861), .ZN(n12814) );
  AND2_X2 U11425 ( .A1(n13257), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13261) );
  NAND2_X1 U11426 ( .A1(n18798), .A2(n18808), .ZN(n14089) );
  NAND2_X1 U11427 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20913), .ZN(
        n14088) );
  NAND2_X1 U11428 ( .A1(n18815), .A2(n18649), .ZN(n14086) );
  NAND2_X1 U11429 ( .A1(n18798), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14087) );
  AND2_X2 U11430 ( .A1(n14751), .A2(n13526), .ZN(n11474) );
  INV_X1 U11431 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19228) );
  AND2_X1 U11432 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13526) );
  AND2_X2 U11433 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10519) );
  INV_X2 U11434 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13614) );
  NAND2_X2 U11435 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18661) );
  AND2_X1 U11436 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18638) );
  INV_X2 U11437 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11673) );
  AND2_X1 U11438 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16859) );
  NAND2_X1 U11439 ( .A1(n9925), .A2(n13728), .ZN(n19656) );
  INV_X1 U11440 ( .A(n11446), .ZN(n9657) );
  NAND2_X1 U11441 ( .A1(n10460), .A2(n13613), .ZN(n19361) );
  INV_X2 U11442 ( .A(n12947), .ZN(n19047) );
  NAND2_X2 U11443 ( .A1(n12612), .A2(n12611), .ZN(n13306) );
  INV_X1 U11444 ( .A(n9891), .ZN(n10950) );
  XNOR2_X1 U11445 ( .A(n10945), .B(n9855), .ZN(n9891) );
  AND2_X1 U11446 ( .A1(n13261), .A2(n14752), .ZN(n9655) );
  NOR2_X1 U11447 ( .A1(n14088), .A2(n14087), .ZN(n9656) );
  NOR2_X1 U11448 ( .A1(n14088), .A2(n14087), .ZN(n15344) );
  NOR2_X2 U11449 ( .A1(n9829), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11420) );
  NOR2_X2 U11450 ( .A1(n10611), .A2(n11206), .ZN(n9856) );
  AND2_X2 U11451 ( .A1(n14966), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11072) );
  AND2_X1 U11452 ( .A1(n11425), .A2(n13526), .ZN(n11941) );
  AND2_X1 U11453 ( .A1(n14752), .A2(n11426), .ZN(n11446) );
  NAND2_X1 U11454 ( .A1(n9902), .A2(n10179), .ZN(n14650) );
  AND2_X2 U11455 ( .A1(n14593), .A2(n15950), .ZN(n9723) );
  OR2_X2 U11456 ( .A1(n10487), .A2(n10500), .ZN(n10708) );
  BUF_X2 U11457 ( .A(n11550), .Z(n13410) );
  NAND2_X1 U11458 ( .A1(n10400), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9875) );
  AND2_X1 U11459 ( .A1(n13261), .A2(n11420), .ZN(n12215) );
  NAND2_X2 U11460 ( .A1(n11552), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11630) );
  AND2_X4 U11461 ( .A1(n11169), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9674) );
  NAND2_X2 U11462 ( .A1(n13786), .A2(n13785), .ZN(n13784) );
  AND2_X2 U11463 ( .A1(n14615), .A2(n15834), .ZN(n14593) );
  AND2_X1 U11464 ( .A1(n14752), .A2(n13526), .ZN(n11473) );
  NOR2_X1 U11465 ( .A1(n14088), .A2(n14084), .ZN(n15424) );
  NAND2_X2 U11466 ( .A1(n9877), .A2(n10784), .ZN(n15104) );
  NOR2_X2 U11467 ( .A1(n13779), .A2(n13832), .ZN(n13830) );
  NAND2_X1 U11468 ( .A1(n11629), .A2(n11628), .ZN(n11631) );
  NAND2_X4 U11469 ( .A1(n20157), .A2(n11655), .ZN(n13545) );
  NAND2_X2 U11470 ( .A1(n11634), .A2(n11633), .ZN(n20157) );
  INV_X1 U11471 ( .A(n10300), .ZN(n9663) );
  INV_X1 U11472 ( .A(n12740), .ZN(n9664) );
  NOR2_X2 U11473 ( .A1(n10391), .A2(n10392), .ZN(n11135) );
  AOI21_X2 U11474 ( .B1(n10442), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10423), .ZN(n10429) );
  NAND2_X2 U11475 ( .A1(n10416), .A2(n10379), .ZN(n10442) );
  AND2_X1 U11476 ( .A1(n10177), .A2(n9905), .ZN(n9902) );
  NAND2_X1 U11477 ( .A1(n14824), .A2(n14823), .ZN(n14822) );
  NAND2_X2 U11478 ( .A1(n13530), .A2(n11656), .ZN(n13515) );
  NAND2_X2 U11479 ( .A1(n11649), .A2(n11648), .ZN(n13530) );
  NAND2_X2 U11480 ( .A1(n11545), .A2(n10265), .ZN(n11557) );
  XNOR2_X2 U11481 ( .A(n12336), .B(n13592), .ZN(n13590) );
  AOI21_X2 U11482 ( .B1(n14070), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14069), .ZN(n14629) );
  BUF_X4 U11484 ( .A(n10637), .Z(n9666) );
  NOR2_X2 U11485 ( .A1(n14034), .A2(n10054), .ZN(n14329) );
  NAND2_X2 U11486 ( .A1(n11906), .A2(n11905), .ZN(n14034) );
  INV_X1 U11487 ( .A(n10294), .ZN(n9667) );
  NAND2_X4 U11488 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  INV_X4 U11489 ( .A(n10378), .ZN(n11215) );
  INV_X2 U11490 ( .A(n10490), .ZN(n13728) );
  INV_X1 U11491 ( .A(n9665), .ZN(n9670) );
  NOR2_X2 U11492 ( .A1(n14285), .A2(n14286), .ZN(n14269) );
  NAND2_X1 U11493 ( .A1(n10490), .A2(n10499), .ZN(n10711) );
  NAND2_X1 U11494 ( .A1(n10494), .A2(n10490), .ZN(n19330) );
  AND2_X2 U11495 ( .A1(n14421), .A2(n10060), .ZN(n14294) );
  NOR2_X4 U11496 ( .A1(n12063), .A2(n14430), .ZN(n14421) );
  BUF_X1 U11497 ( .A(n12319), .Z(n9672) );
  AND2_X1 U11498 ( .A1(n11169), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U11499 ( .A1(n9955), .A2(n9951), .ZN(n10386) );
  AND2_X1 U11500 ( .A1(n10385), .A2(n11139), .ZN(n9951) );
  OAI21_X1 U11501 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18808), .A(
        n14183), .ZN(n14184) );
  OR2_X1 U11502 ( .A1(n14187), .A2(n14188), .ZN(n14183) );
  NAND2_X1 U11503 ( .A1(n12387), .A2(n12388), .ZN(n9900) );
  OR2_X1 U11504 ( .A1(n12281), .A2(n11604), .ZN(n11609) );
  NAND2_X1 U11505 ( .A1(n11556), .A2(n13402), .ZN(n11704) );
  AND2_X1 U11506 ( .A1(n11704), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12272) );
  MUX2_X1 U11507 ( .A(n12586), .B(n10390), .S(n10393), .Z(n10394) );
  NAND2_X1 U11508 ( .A1(n11137), .A2(n19245), .ZN(n10403) );
  INV_X1 U11509 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9909) );
  AND2_X1 U11510 ( .A1(n10924), .A2(n10632), .ZN(n10640) );
  AND2_X1 U11511 ( .A1(n12253), .A2(n12252), .ZN(n12413) );
  OR2_X1 U11512 ( .A1(n12284), .A2(n12251), .ZN(n12253) );
  NAND2_X1 U11513 ( .A1(n15779), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U11514 ( .A1(n14294), .A2(n14296), .ZN(n14285) );
  AND2_X1 U11515 ( .A1(n14449), .A2(n14316), .ZN(n10066) );
  NOR2_X1 U11516 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  INV_X1 U11517 ( .A(n14465), .ZN(n10057) );
  NOR2_X1 U11518 ( .A1(n10051), .A2(n9772), .ZN(n10050) );
  NAND2_X1 U11519 ( .A1(n11750), .A2(n11749), .ZN(n11765) );
  NOR2_X1 U11520 ( .A1(n13346), .A2(n11673), .ZN(n11830) );
  OR2_X1 U11521 ( .A1(n13580), .A2(n11673), .ZN(n12146) );
  NOR2_X1 U11522 ( .A1(n12393), .A2(n12396), .ZN(n10205) );
  INV_X1 U11523 ( .A(n15847), .ZN(n10207) );
  INV_X1 U11524 ( .A(n13844), .ZN(n9977) );
  AND2_X1 U11525 ( .A1(n14256), .A2(n13362), .ZN(n12505) );
  NOR2_X1 U11526 ( .A1(n11092), .A2(n9781), .ZN(n10028) );
  INV_X1 U11527 ( .A(n9718), .ZN(n10029) );
  AOI21_X1 U11528 ( .B1(n9929), .B2(n9932), .A(n9928), .ZN(n9927) );
  INV_X1 U11529 ( .A(n16233), .ZN(n9928) );
  AND2_X1 U11530 ( .A1(n10088), .A2(n11011), .ZN(n10087) );
  INV_X1 U11531 ( .A(n13510), .ZN(n11011) );
  OAI211_X1 U11532 ( .C1(n9954), .C2(n10387), .A(n9952), .B(n10386), .ZN(
        n11194) );
  NAND2_X1 U11533 ( .A1(n9953), .A2(n9956), .ZN(n9952) );
  AND2_X1 U11534 ( .A1(n13931), .A2(n19888), .ZN(n11200) );
  AND2_X1 U11535 ( .A1(n9646), .A2(n12590), .ZN(n13307) );
  AND2_X1 U11536 ( .A1(n11215), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12590) );
  NOR2_X1 U11537 ( .A1(n14084), .A2(n18661), .ZN(n14111) );
  INV_X1 U11538 ( .A(n13362), .ZN(n13349) );
  AND2_X1 U11539 ( .A1(n11673), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12241) );
  INV_X1 U11540 ( .A(n12146), .ZN(n12242) );
  AND2_X1 U11541 ( .A1(n13395), .A2(n13578), .ZN(n13414) );
  NAND2_X1 U11542 ( .A1(n10041), .A2(n10042), .ZN(n10804) );
  INV_X1 U11543 ( .A(n10799), .ZN(n10041) );
  NOR2_X1 U11544 ( .A1(n12928), .A2(n10077), .ZN(n10076) );
  INV_X1 U11545 ( .A(n12563), .ZN(n10077) );
  NAND2_X1 U11546 ( .A1(n13752), .A2(n9785), .ZN(n13779) );
  AND2_X1 U11547 ( .A1(n13751), .A2(n13780), .ZN(n9785) );
  OR2_X1 U11548 ( .A1(n15104), .A2(n10792), .ZN(n10228) );
  NOR2_X1 U11549 ( .A1(n16905), .A2(n14087), .ZN(n15355) );
  INV_X1 U11550 ( .A(n9699), .ZN(n17098) );
  AND2_X1 U11551 ( .A1(n13421), .A2(n13058), .ZN(n20733) );
  OAI21_X1 U11552 ( .B1(n14711), .B2(n16079), .A(n14712), .ZN(n9828) );
  NAND2_X1 U11553 ( .A1(n10933), .A2(n16343), .ZN(n13051) );
  NAND2_X1 U11554 ( .A1(n9865), .A2(n16209), .ZN(n16290) );
  OR2_X1 U11555 ( .A1(n16208), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9865) );
  AND2_X1 U11556 ( .A1(n12276), .A2(n12277), .ZN(n9842) );
  INV_X1 U11557 ( .A(n12280), .ZN(n9841) );
  OR2_X1 U11558 ( .A1(n11739), .A2(n11738), .ZN(n12351) );
  INV_X1 U11559 ( .A(n12380), .ZN(n11636) );
  AND2_X1 U11560 ( .A1(n12288), .A2(n12378), .ZN(n12283) );
  NAND2_X1 U11561 ( .A1(n11564), .A2(n11630), .ZN(n11643) );
  OAI21_X1 U11562 ( .B1(n11563), .B2(n13247), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11564) );
  AND2_X1 U11563 ( .A1(n13249), .A2(n12418), .ZN(n13081) );
  NOR2_X1 U11564 ( .A1(n10393), .A2(n13941), .ZN(n10385) );
  AND2_X1 U11565 ( .A1(n16126), .A2(n10045), .ZN(n10044) );
  INV_X1 U11566 ( .A(n10906), .ZN(n10045) );
  NOR2_X1 U11567 ( .A1(n14988), .A2(n10152), .ZN(n10151) );
  NAND2_X1 U11568 ( .A1(n10020), .A2(n10022), .ZN(n10017) );
  AND4_X1 U11569 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10630) );
  NAND2_X1 U11570 ( .A1(n9724), .A2(n10357), .ZN(n10416) );
  INV_X1 U11571 ( .A(n11159), .ZN(n10405) );
  AOI22_X1 U11572 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U11573 ( .A1(n10634), .A2(n10633), .ZN(n10641) );
  INV_X1 U11574 ( .A(n10640), .ZN(n10634) );
  OR2_X1 U11575 ( .A1(n11108), .A2(n10909), .ZN(n10924) );
  NOR2_X1 U11576 ( .A1(n13278), .A2(n11556), .ZN(n9800) );
  NAND2_X1 U11577 ( .A1(n9997), .A2(n14445), .ZN(n9996) );
  NOR2_X1 U11578 ( .A1(n10063), .A2(n14306), .ZN(n10062) );
  INV_X1 U11579 ( .A(n14422), .ZN(n10063) );
  NAND2_X1 U11580 ( .A1(n11838), .A2(n10052), .ZN(n10051) );
  INV_X1 U11581 ( .A(n13838), .ZN(n10052) );
  NAND2_X1 U11582 ( .A1(n14645), .A2(n12397), .ZN(n10203) );
  OR2_X1 U11583 ( .A1(n11601), .A2(n11600), .ZN(n12377) );
  INV_X1 U11584 ( .A(n11793), .ZN(n9908) );
  INV_X1 U11585 ( .A(n12357), .ZN(n10186) );
  NAND2_X1 U11586 ( .A1(n12421), .A2(n13362), .ZN(n12510) );
  NAND2_X1 U11587 ( .A1(n13386), .A2(n13385), .ZN(n13387) );
  NAND2_X1 U11588 ( .A1(n11686), .A2(n10195), .ZN(n10194) );
  NAND2_X1 U11589 ( .A1(n10193), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10192) );
  NOR2_X1 U11590 ( .A1(n10196), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10191) );
  INV_X1 U11591 ( .A(n11686), .ZN(n10196) );
  NAND2_X1 U11592 ( .A1(n9898), .A2(n9802), .ZN(n11639) );
  AND2_X1 U11593 ( .A1(n9897), .A2(n11610), .ZN(n9802) );
  INV_X1 U11594 ( .A(n11624), .ZN(n9897) );
  AND2_X1 U11595 ( .A1(n11701), .A2(n20119), .ZN(n11651) );
  NAND2_X1 U11596 ( .A1(n20711), .A2(n20644), .ZN(n11716) );
  AOI21_X1 U11597 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19869), .A(
        n10666), .ZN(n10916) );
  NOR2_X1 U11598 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  INV_X1 U11599 ( .A(n10663), .ZN(n10665) );
  AND2_X1 U11600 ( .A1(n9743), .A2(n11033), .ZN(n10035) );
  NAND2_X1 U11601 ( .A1(n10877), .A2(n11100), .ZN(n10874) );
  NAND2_X1 U11602 ( .A1(n10834), .A2(n11100), .ZN(n10819) );
  OR2_X1 U11603 ( .A1(n10833), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10834) );
  AND2_X1 U11604 ( .A1(n10810), .A2(n10038), .ZN(n10037) );
  INV_X1 U11605 ( .A(n10849), .ZN(n10038) );
  NAND2_X1 U11606 ( .A1(n10791), .A2(n9866), .ZN(n10806) );
  AND2_X1 U11607 ( .A1(n10790), .A2(n10039), .ZN(n9866) );
  AND2_X1 U11608 ( .A1(n10042), .A2(n10040), .ZN(n10039) );
  NAND2_X1 U11609 ( .A1(n11156), .A2(n10413), .ZN(n10000) );
  NAND2_X1 U11610 ( .A1(n14815), .A2(n12806), .ZN(n12829) );
  INV_X1 U11611 ( .A(n12802), .ZN(n12805) );
  INV_X1 U11612 ( .A(n14935), .ZN(n10108) );
  INV_X1 U11613 ( .A(n14849), .ZN(n12658) );
  NAND2_X1 U11614 ( .A1(n13830), .A2(n16186), .ZN(n14849) );
  OAI21_X1 U11615 ( .B1(n10490), .B2(n12592), .A(n12589), .ZN(n12610) );
  NOR2_X1 U11616 ( .A1(n10158), .A2(n10157), .ZN(n10156) );
  INV_X1 U11617 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10157) );
  NAND2_X1 U11618 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U11619 ( .A1(n14995), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10220) );
  OR2_X1 U11620 ( .A1(n15636), .A2(n10801), .ZN(n10879) );
  INV_X1 U11621 ( .A(n15035), .ZN(n9848) );
  AND2_X1 U11622 ( .A1(n16210), .A2(n15019), .ZN(n9942) );
  AND2_X1 U11623 ( .A1(n10127), .A2(n15278), .ZN(n10126) );
  NOR2_X1 U11624 ( .A1(n11007), .A2(n10089), .ZN(n10088) );
  INV_X1 U11625 ( .A(n13485), .ZN(n10089) );
  OR2_X1 U11626 ( .A1(n11006), .A2(n13463), .ZN(n11007) );
  NAND2_X1 U11627 ( .A1(n9876), .A2(n19037), .ZN(n10740) );
  NAND2_X1 U11628 ( .A1(n10950), .A2(n10801), .ZN(n9876) );
  NAND2_X1 U11629 ( .A1(n10016), .A2(n10019), .ZN(n10013) );
  NAND2_X1 U11630 ( .A1(n9703), .A2(n10463), .ZN(n19413) );
  NAND2_X1 U11631 ( .A1(n10211), .A2(n10273), .ZN(n10210) );
  NAND2_X1 U11632 ( .A1(n10209), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10208) );
  NAND2_X1 U11633 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14085) );
  INV_X1 U11634 ( .A(n15493), .ZN(n9820) );
  AND2_X1 U11635 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9819) );
  INV_X1 U11636 ( .A(n15494), .ZN(n9822) );
  INV_X1 U11637 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n20889) );
  OR2_X1 U11638 ( .A1(n14089), .A2(n14088), .ZN(n15479) );
  XNOR2_X1 U11639 ( .A(n17380), .B(n15576), .ZN(n15529) );
  NOR2_X1 U11640 ( .A1(n17342), .A2(n18213), .ZN(n15606) );
  NOR2_X1 U11641 ( .A1(n17360), .A2(n15537), .ZN(n15540) );
  NOR2_X1 U11642 ( .A1(n17801), .A2(n15539), .ZN(n15542) );
  XOR2_X1 U11643 ( .A(n15537), .B(n17360), .Z(n15538) );
  NAND2_X1 U11644 ( .A1(n17821), .A2(n9808), .ZN(n9807) );
  NAND2_X1 U11645 ( .A1(n9809), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9808) );
  INV_X1 U11646 ( .A(n17822), .ZN(n9809) );
  NAND2_X1 U11647 ( .A1(n17822), .A2(n15535), .ZN(n9806) );
  INV_X1 U11648 ( .A(n17802), .ZN(n10147) );
  AOI21_X1 U11649 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18191), .A(
        n14191), .ZN(n14205) );
  NOR2_X1 U11650 ( .A1(n18635), .A2(n14206), .ZN(n15604) );
  NOR2_X1 U11651 ( .A1(n14095), .A2(n14094), .ZN(n15415) );
  NOR2_X1 U11652 ( .A1(n14147), .A2(n14146), .ZN(n14168) );
  INV_X1 U11653 ( .A(n16515), .ZN(n16524) );
  NAND2_X1 U11654 ( .A1(n12421), .A2(n12513), .ZN(n13082) );
  NOR2_X1 U11655 ( .A1(n11548), .A2(n11556), .ZN(n13348) );
  AND2_X1 U11656 ( .A1(n13276), .A2(n13275), .ZN(n13577) );
  NOR2_X1 U11657 ( .A1(n14260), .A2(n10068), .ZN(n10067) );
  INV_X1 U11658 ( .A(n14271), .ZN(n10068) );
  NOR2_X1 U11659 ( .A1(n14593), .A2(n10253), .ZN(n14597) );
  OR2_X1 U11660 ( .A1(n12152), .A2(n12151), .ZN(n14412) );
  AND2_X1 U11661 ( .A1(n12027), .A2(n12026), .ZN(n14449) );
  AND2_X1 U11662 ( .A1(n12008), .A2(n12007), .ZN(n14316) );
  NAND2_X1 U11663 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  INV_X1 U11664 ( .A(n14330), .ZN(n10055) );
  NOR2_X1 U11665 ( .A1(n11956), .A2(n14669), .ZN(n11957) );
  NAND2_X1 U11666 ( .A1(n11957), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U11667 ( .A1(n10053), .A2(n10056), .ZN(n14467) );
  INV_X1 U11668 ( .A(n14034), .ZN(n10053) );
  AOI21_X1 U11669 ( .B1(n12350), .B2(n11830), .A(n11772), .ZN(n13704) );
  AND2_X1 U11670 ( .A1(n13360), .A2(n11695), .ZN(n10048) );
  NAND2_X1 U11671 ( .A1(n13361), .A2(n13360), .ZN(n13359) );
  AND2_X1 U11672 ( .A1(n14707), .A2(n16048), .ZN(n14710) );
  NOR2_X1 U11673 ( .A1(n9985), .A2(n9990), .ZN(n9984) );
  INV_X1 U11674 ( .A(n14282), .ZN(n9990) );
  INV_X1 U11675 ( .A(n9986), .ZN(n9985) );
  INV_X1 U11676 ( .A(n13989), .ZN(n9901) );
  AND3_X1 U11677 ( .A1(n12450), .A2(n12461), .A3(n12449), .ZN(n13844) );
  INV_X1 U11678 ( .A(n12442), .ZN(n9975) );
  NAND2_X1 U11679 ( .A1(n9981), .A2(n9978), .ZN(n13843) );
  NOR2_X1 U11680 ( .A1(n9982), .A2(n13788), .ZN(n9978) );
  AND2_X1 U11681 ( .A1(n13252), .A2(n13390), .ZN(n13401) );
  OAI21_X1 U11682 ( .B1(n11681), .B2(n12314), .A(n11639), .ZN(n11696) );
  INV_X1 U11683 ( .A(n13386), .ZN(n13391) );
  INV_X1 U11684 ( .A(n20708), .ZN(n20445) );
  NOR2_X1 U11685 ( .A1(n20254), .A2(n20253), .ZN(n20541) );
  OAI221_X2 U11686 ( .B1(n16088), .B2(n15671), .C1(n16092), .C2(n15671), .A(
        n20644), .ZN(n20254) );
  NOR2_X1 U11687 ( .A1(n14771), .A2(n16122), .ZN(n10170) );
  NOR2_X1 U11688 ( .A1(n19047), .A2(n16152), .ZN(n16141) );
  INV_X1 U11689 ( .A(n15034), .ZN(n10161) );
  AND2_X1 U11690 ( .A1(n11363), .A2(n11362), .ZN(n13961) );
  AND2_X1 U11691 ( .A1(n11265), .A2(n11264), .ZN(n13874) );
  OR2_X1 U11692 ( .A1(n13636), .A2(n12970), .ZN(n13040) );
  NAND2_X1 U11693 ( .A1(n14867), .A2(n10121), .ZN(n12977) );
  NOR2_X1 U11694 ( .A1(n9773), .A2(n10122), .ZN(n10121) );
  INV_X1 U11695 ( .A(n11409), .ZN(n10122) );
  OAI21_X1 U11696 ( .B1(n14790), .B2(n10096), .A(n9691), .ZN(n10094) );
  NAND2_X1 U11697 ( .A1(n14796), .A2(n12874), .ZN(n10090) );
  XNOR2_X1 U11698 ( .A(n14835), .B(n12782), .ZN(n14824) );
  NOR2_X1 U11699 ( .A1(n16307), .A2(n10128), .ZN(n10127) );
  INV_X1 U11700 ( .A(n15287), .ZN(n10128) );
  NAND2_X1 U11701 ( .A1(n10120), .A2(n9768), .ZN(n13801) );
  INV_X1 U11702 ( .A(n11232), .ZN(n10115) );
  OR2_X1 U11703 ( .A1(n10164), .A2(n16198), .ZN(n10163) );
  NOR2_X1 U11704 ( .A1(n11073), .A2(n10239), .ZN(n10238) );
  NOR2_X1 U11705 ( .A1(n10025), .A2(n14230), .ZN(n10213) );
  NOR2_X2 U11706 ( .A1(n14985), .A2(n14984), .ZN(n14974) );
  NAND2_X1 U11707 ( .A1(n10006), .A2(n10880), .ZN(n10005) );
  INV_X1 U11708 ( .A(n10007), .ZN(n10006) );
  NOR2_X1 U11709 ( .A1(n10261), .A2(n10008), .ZN(n10007) );
  INV_X1 U11710 ( .A(n15011), .ZN(n10008) );
  NOR2_X1 U11711 ( .A1(n16212), .A2(n9940), .ZN(n9939) );
  INV_X1 U11712 ( .A(n15085), .ZN(n9940) );
  AND2_X1 U11713 ( .A1(n9942), .A2(n15086), .ZN(n9938) );
  INV_X1 U11714 ( .A(n15264), .ZN(n15241) );
  NAND2_X1 U11715 ( .A1(n16221), .A2(n16312), .ZN(n9963) );
  OR2_X1 U11716 ( .A1(n19094), .A2(n16324), .ZN(n9962) );
  AND2_X1 U11717 ( .A1(n11327), .A2(n11326), .ZN(n16296) );
  NAND2_X1 U11718 ( .A1(n15286), .A2(n10126), .ZN(n16295) );
  AOI21_X1 U11719 ( .B1(n10227), .B2(n10223), .A(n9681), .ZN(n10222) );
  NOR2_X1 U11720 ( .A1(n10224), .A2(n16248), .ZN(n10223) );
  INV_X1 U11721 ( .A(n16246), .ZN(n10229) );
  AND2_X1 U11722 ( .A1(n10227), .A2(n10226), .ZN(n10225) );
  INV_X1 U11723 ( .A(n16248), .ZN(n10226) );
  AND2_X1 U11724 ( .A1(n10796), .A2(n15095), .ZN(n10227) );
  OR2_X1 U11725 ( .A1(n10803), .A2(n15292), .ZN(n16246) );
  NAND2_X1 U11726 ( .A1(n15112), .A2(n15111), .ZN(n9877) );
  NAND2_X1 U11727 ( .A1(n9891), .A2(n10739), .ZN(n13856) );
  INV_X1 U11728 ( .A(n10694), .ZN(n10946) );
  NAND2_X1 U11729 ( .A1(n13732), .A2(n13888), .ZN(n10014) );
  NAND2_X1 U11730 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  INV_X1 U11731 ( .A(n10452), .ZN(n10103) );
  INV_X1 U11732 ( .A(n10453), .ZN(n10104) );
  AND2_X1 U11733 ( .A1(n11198), .A2(n11170), .ZN(n15240) );
  NAND2_X1 U11734 ( .A1(n13230), .A2(n12597), .ZN(n13292) );
  NAND2_X1 U11735 ( .A1(n10347), .A2(n10273), .ZN(n10355) );
  NOR2_X1 U11736 ( .A1(n19698), .A2(n19411), .ZN(n19415) );
  NAND2_X1 U11737 ( .A1(n19113), .A2(n19142), .ZN(n19450) );
  NAND2_X1 U11738 ( .A1(n19872), .A2(n19854), .ZN(n19502) );
  NAND2_X1 U11739 ( .A1(n19872), .A2(n19883), .ZN(n19859) );
  OR2_X1 U11740 ( .A1(n19872), .A2(n19883), .ZN(n19624) );
  NAND2_X1 U11741 ( .A1(n10299), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10307) );
  OR2_X1 U11742 ( .A1(n19872), .A2(n19854), .ZN(n19698) );
  AOI22_X2 U11743 ( .A1(n12960), .A2(n15328), .B1(n13758), .B2(n16338), .ZN(
        n19447) );
  NOR2_X1 U11744 ( .A1(n14137), .A2(n14136), .ZN(n17239) );
  NAND2_X1 U11745 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15475) );
  XNOR2_X1 U11746 ( .A(n15529), .B(n18154), .ZN(n17848) );
  NOR2_X2 U11747 ( .A1(n14167), .A2(n14166), .ZN(n18841) );
  AND2_X1 U11748 ( .A1(n16357), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9816) );
  NAND2_X1 U11749 ( .A1(n17593), .A2(n17920), .ZN(n15550) );
  AND2_X1 U11750 ( .A1(n17570), .A2(n10137), .ZN(n17551) );
  NAND2_X1 U11751 ( .A1(n17570), .A2(n17603), .ZN(n17604) );
  XNOR2_X1 U11752 ( .A(n15542), .B(n15541), .ZN(n17792) );
  NAND2_X1 U11753 ( .A1(n17812), .A2(n10148), .ZN(n10144) );
  NAND2_X1 U11754 ( .A1(n10145), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10146) );
  OAI21_X1 U11755 ( .B1(n17821), .B2(n17822), .A(n15535), .ZN(n15536) );
  NAND2_X1 U11756 ( .A1(n17821), .A2(n17822), .ZN(n17820) );
  INV_X1 U11757 ( .A(n18688), .ZN(n18836) );
  NAND2_X1 U11758 ( .A1(n18852), .A2(n15604), .ZN(n18665) );
  AOI211_X1 U11759 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n14124), .B(n14123), .ZN(n14125) );
  INV_X1 U11760 ( .A(n18841), .ZN(n18203) );
  INV_X1 U11761 ( .A(n14168), .ZN(n18224) );
  NAND2_X1 U11762 ( .A1(n20733), .A2(n12416), .ZN(n15779) );
  AND2_X1 U11763 ( .A1(n15902), .A2(n20067), .ZN(n15871) );
  XNOR2_X1 U11764 ( .A(n9794), .B(n14758), .ZN(n12404) );
  NAND2_X1 U11765 ( .A1(n10174), .A2(n10173), .ZN(n9794) );
  NAND2_X1 U11766 ( .A1(n14574), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10173) );
  NAND2_X1 U11767 ( .A1(n14589), .A2(n12403), .ZN(n10174) );
  AND2_X1 U11768 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15925), .ZN(
        n15918) );
  OAI21_X1 U11769 ( .B1(n14704), .B2(n16048), .A(n20078), .ZN(n9833) );
  INV_X1 U11770 ( .A(n14743), .ZN(n9832) );
  AND2_X1 U11771 ( .A1(n13414), .A2(n13413), .ZN(n20089) );
  OR2_X1 U11772 ( .A1(n12564), .A2(n11083), .ZN(n10075) );
  NOR2_X1 U11773 ( .A1(n10076), .A2(n11083), .ZN(n10072) );
  NAND2_X1 U11774 ( .A1(n10111), .A2(n10110), .ZN(n10109) );
  INV_X1 U11775 ( .A(n19077), .ZN(n10110) );
  INV_X1 U11776 ( .A(n10112), .ZN(n10111) );
  OR2_X1 U11777 ( .A1(n13453), .A2(n10112), .ZN(n19076) );
  AND2_X1 U11778 ( .A1(n9915), .A2(n19222), .ZN(n9910) );
  NAND2_X1 U11779 ( .A1(n16203), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16202) );
  NAND2_X1 U11780 ( .A1(n13051), .A2(n10969), .ZN(n19229) );
  AND2_X1 U11781 ( .A1(n19229), .A2(n19877), .ZN(n19239) );
  OR2_X1 U11782 ( .A1(n13051), .A2(n11215), .ZN(n19234) );
  NAND2_X1 U11783 ( .A1(n9881), .A2(n9879), .ZN(n11151) );
  NOR2_X1 U11784 ( .A1(n9731), .A2(n11183), .ZN(n9882) );
  NAND2_X1 U11785 ( .A1(n9852), .A2(n14990), .ZN(n15164) );
  OR2_X1 U11786 ( .A1(n9641), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9852) );
  NOR2_X1 U11787 ( .A1(n9913), .A2(n9924), .ZN(n9912) );
  INV_X1 U11788 ( .A(n9918), .ZN(n9913) );
  OAI21_X1 U11789 ( .B1(n9924), .B2(n9918), .A(n9916), .ZN(n9915) );
  NAND2_X1 U11790 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  NAND2_X1 U11791 ( .A1(n9920), .A2(n15030), .ZN(n9917) );
  AOI21_X1 U11792 ( .B1(n16291), .B2(n16334), .A(n9864), .ZN(n9863) );
  NOR2_X1 U11793 ( .A1(n16289), .A2(n16329), .ZN(n9864) );
  NAND2_X1 U11794 ( .A1(n11198), .A2(n11197), .ZN(n16324) );
  INV_X1 U11795 ( .A(n16312), .ZN(n16329) );
  AND2_X1 U11796 ( .A1(n11198), .A2(n19901), .ZN(n16334) );
  INV_X1 U11797 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19896) );
  INV_X1 U11798 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19888) );
  INV_X1 U11799 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19869) );
  AND2_X1 U11800 ( .A1(n13641), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15328) );
  NOR2_X1 U11801 ( .A1(n19450), .A2(n19859), .ZN(n19364) );
  INV_X1 U11802 ( .A(n16887), .ZN(n16910) );
  INV_X1 U11803 ( .A(n16923), .ZN(n16907) );
  NOR2_X2 U11804 ( .A1(n17232), .A2(n17342), .ZN(n17233) );
  NOR2_X1 U11805 ( .A1(n18234), .A2(n17277), .ZN(n17272) );
  INV_X1 U11806 ( .A(n16409), .ZN(n17354) );
  NOR2_X1 U11807 ( .A1(n15470), .A2(n15469), .ZN(n17371) );
  INV_X2 U11808 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18808) );
  NAND2_X1 U11809 ( .A1(n9840), .A2(n9839), .ZN(n9838) );
  NAND2_X1 U11810 ( .A1(n12278), .A2(n12260), .ZN(n9839) );
  INV_X1 U11811 ( .A(n12320), .ZN(n11606) );
  OR2_X1 U11812 ( .A1(n10708), .A2(n10548), .ZN(n10552) );
  AND2_X1 U11813 ( .A1(n20504), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12267) );
  CLKBUF_X1 U11814 ( .A(n11491), .Z(n12224) );
  NAND2_X1 U11815 ( .A1(n11741), .A2(n11740), .ZN(n11749) );
  AND2_X1 U11816 ( .A1(n11749), .A2(n11763), .ZN(n9907) );
  INV_X1 U11817 ( .A(n12288), .ZN(n12281) );
  INV_X1 U11818 ( .A(n11603), .ZN(n10195) );
  OR2_X1 U11819 ( .A1(n11621), .A2(n11620), .ZN(n12321) );
  OR2_X1 U11820 ( .A1(n11714), .A2(n11713), .ZN(n12340) );
  NAND2_X1 U11821 ( .A1(n10641), .A2(n10635), .ZN(n10663) );
  NOR2_X1 U11822 ( .A1(n10779), .A2(n9873), .ZN(n9872) );
  NAND2_X1 U11823 ( .A1(n10776), .A2(n10778), .ZN(n9873) );
  OR2_X1 U11824 ( .A1(n13931), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U11825 ( .A1(n19361), .A2(n12763), .ZN(n10556) );
  AOI22_X1 U11826 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10313) );
  NAND2_X1 U11827 ( .A1(n13728), .A2(n10493), .ZN(n10471) );
  AND2_X1 U11828 ( .A1(n17366), .A2(n15585), .ZN(n15571) );
  AND2_X1 U11829 ( .A1(n14203), .A2(n14201), .ZN(n14182) );
  AND2_X1 U11830 ( .A1(n16515), .A2(n15603), .ZN(n14181) );
  NOR2_X1 U11831 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20913), .ZN(
        n14201) );
  NOR2_X1 U11832 ( .A1(n14318), .A2(n9998), .ZN(n9997) );
  INV_X1 U11833 ( .A(n14071), .ZN(n9998) );
  INV_X1 U11834 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12057) );
  AND2_X1 U11835 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  INV_X1 U11836 ( .A(n14443), .ZN(n10065) );
  INV_X1 U11837 ( .A(n12237), .ZN(n12206) );
  OR2_X1 U11838 ( .A1(n14035), .A2(n10059), .ZN(n10058) );
  INV_X1 U11839 ( .A(n14475), .ZN(n10059) );
  INV_X1 U11840 ( .A(n12241), .ZN(n11935) );
  NAND2_X1 U11841 ( .A1(n14593), .A2(n9797), .ZN(n9799) );
  NOR2_X1 U11842 ( .A1(n9782), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9797) );
  NOR2_X1 U11843 ( .A1(n14297), .A2(n9987), .ZN(n9986) );
  INV_X1 U11844 ( .A(n9988), .ZN(n9987) );
  NOR2_X1 U11845 ( .A1(n9989), .A2(n14414), .ZN(n9988) );
  INV_X1 U11846 ( .A(n14308), .ZN(n9989) );
  NOR2_X1 U11847 ( .A1(n9992), .A2(n14468), .ZN(n9991) );
  INV_X1 U11848 ( .A(n9993), .ZN(n9992) );
  NOR2_X1 U11849 ( .A1(n14476), .A2(n9994), .ZN(n9993) );
  INV_X1 U11850 ( .A(n14038), .ZN(n9994) );
  INV_X1 U11851 ( .A(n12388), .ZN(n10178) );
  INV_X1 U11852 ( .A(n12393), .ZN(n12400) );
  INV_X1 U11853 ( .A(n12505), .ZN(n12518) );
  NAND2_X1 U11854 ( .A1(n12426), .A2(n12425), .ZN(n12428) );
  AND2_X1 U11855 ( .A1(n13085), .A2(n13084), .ZN(n13252) );
  NAND2_X1 U11856 ( .A1(n11643), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9795) );
  NAND2_X1 U11857 ( .A1(n20135), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12380) );
  NAND2_X1 U11858 ( .A1(n9898), .A2(n11610), .ZN(n11625) );
  INV_X1 U11859 ( .A(n13091), .ZN(n11499) );
  NAND2_X1 U11860 ( .A1(n12291), .A2(n12292), .ZN(n9845) );
  INV_X1 U11861 ( .A(n20254), .ZN(n20115) );
  INV_X1 U11862 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20412) );
  OR2_X1 U11863 ( .A1(n10530), .A2(n10529), .ZN(n10636) );
  AND2_X1 U11864 ( .A1(n10044), .A2(n11094), .ZN(n10043) );
  INV_X1 U11865 ( .A(n10844), .ZN(n10036) );
  NAND2_X1 U11866 ( .A1(n18982), .A2(n10810), .ZN(n10850) );
  NOR2_X1 U11867 ( .A1(n10806), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10809) );
  NOR2_X1 U11868 ( .A1(n10788), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10042) );
  INV_X1 U11869 ( .A(n10737), .ZN(n10033) );
  NOR2_X1 U11870 ( .A1(n10686), .A2(n10685), .ZN(n10738) );
  NAND2_X1 U11871 ( .A1(n10646), .A2(n10653), .ZN(n10685) );
  NAND2_X1 U11872 ( .A1(n11156), .A2(n9709), .ZN(n9999) );
  NOR2_X1 U11873 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U11874 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12607) );
  INV_X1 U11875 ( .A(n12975), .ZN(n10123) );
  NAND2_X1 U11876 ( .A1(n11402), .A2(n10131), .ZN(n10130) );
  AND2_X1 U11877 ( .A1(n14880), .A2(n14879), .ZN(n11402) );
  INV_X1 U11878 ( .A(n13307), .ZN(n12846) );
  NOR2_X1 U11879 ( .A1(n10132), .A2(n14909), .ZN(n10131) );
  INV_X1 U11880 ( .A(n14901), .ZN(n10132) );
  AND2_X1 U11881 ( .A1(n9689), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10150) );
  NAND2_X1 U11882 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  INV_X1 U11883 ( .A(n13778), .ZN(n10080) );
  NOR2_X1 U11884 ( .A1(n10082), .A2(n15078), .ZN(n10081) );
  NAND2_X1 U11885 ( .A1(n10165), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10164) );
  INV_X1 U11886 ( .A(n10166), .ZN(n10165) );
  NAND2_X1 U11887 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10166) );
  NAND2_X1 U11888 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10239) );
  AND2_X1 U11889 ( .A1(n9783), .A2(n9973), .ZN(n9972) );
  INV_X1 U11890 ( .A(n9974), .ZN(n9973) );
  NOR2_X1 U11891 ( .A1(n15146), .A2(n15154), .ZN(n10240) );
  OR3_X1 U11892 ( .A1(n10898), .A2(n10801), .A3(n15146), .ZN(n14973) );
  INV_X1 U11893 ( .A(n14830), .ZN(n10084) );
  AND2_X1 U11894 ( .A1(n9702), .A2(n15002), .ZN(n10004) );
  INV_X1 U11895 ( .A(n15002), .ZN(n10003) );
  NAND2_X1 U11896 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9974) );
  AND2_X1 U11897 ( .A1(n15202), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10241) );
  INV_X1 U11898 ( .A(n13834), .ZN(n10082) );
  INV_X1 U11899 ( .A(n12546), .ZN(n12547) );
  INV_X1 U11900 ( .A(n10792), .ZN(n10224) );
  AOI21_X1 U11901 ( .B1(n10961), .B2(n9949), .A(n9948), .ZN(n9946) );
  INV_X1 U11902 ( .A(n15103), .ZN(n9949) );
  INV_X1 U11903 ( .A(n16266), .ZN(n9948) );
  INV_X1 U11904 ( .A(n10961), .ZN(n9950) );
  NAND2_X1 U11905 ( .A1(n13738), .A2(n10117), .ZN(n10116) );
  INV_X1 U11906 ( .A(n13802), .ZN(n10117) );
  NAND2_X1 U11907 ( .A1(n10954), .A2(n13857), .ZN(n10952) );
  NAND2_X1 U11908 ( .A1(n10441), .A2(n10440), .ZN(n10986) );
  INV_X1 U11909 ( .A(n10612), .ZN(n10231) );
  OR2_X1 U11910 ( .A1(n13185), .A2(n10940), .ZN(n10942) );
  NOR2_X1 U11911 ( .A1(n11215), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11202) );
  INV_X1 U11912 ( .A(n10351), .ZN(n10352) );
  NAND2_X1 U11913 ( .A1(n10342), .A2(n10341), .ZN(n10393) );
  NAND2_X1 U11914 ( .A1(n10334), .A2(n10273), .ZN(n10342) );
  OAI21_X1 U11915 ( .B1(n10340), .B2(n10339), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U11916 ( .A1(n10490), .A2(n10502), .ZN(n19442) );
  NOR2_X1 U11917 ( .A1(n10501), .A2(n10500), .ZN(n10502) );
  INV_X1 U11918 ( .A(n10493), .ZN(n10501) );
  NAND2_X1 U11919 ( .A1(n13728), .A2(n14013), .ZN(n10477) );
  AOI22_X1 U11920 ( .A1(n12739), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U11921 ( .A1(n19876), .A2(n19702), .ZN(n13762) );
  AND2_X1 U11922 ( .A1(n10642), .A2(n10641), .ZN(n11107) );
  AND2_X1 U11923 ( .A1(n10922), .A2(n10921), .ZN(n11120) );
  INV_X1 U11924 ( .A(n14085), .ZN(n10133) );
  NOR2_X1 U11925 ( .A1(n14089), .A2(n18661), .ZN(n15485) );
  NAND2_X1 U11926 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18808), .ZN(
        n14084) );
  NOR2_X1 U11927 ( .A1(n17787), .A2(n16746), .ZN(n17697) );
  OR2_X1 U11928 ( .A1(n17516), .A2(n17770), .ZN(n10135) );
  OR2_X1 U11929 ( .A1(n14181), .A2(n16516), .ZN(n15605) );
  AND2_X1 U11930 ( .A1(n15574), .A2(n15573), .ZN(n15585) );
  INV_X1 U11931 ( .A(n15609), .ZN(n18656) );
  NAND2_X1 U11932 ( .A1(n18638), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14180) );
  INV_X1 U11933 ( .A(n16516), .ZN(n17429) );
  INV_X1 U11934 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14385) );
  AND2_X1 U11935 ( .A1(n12490), .A2(n12489), .ZN(n14445) );
  NOR2_X1 U11936 ( .A1(n14460), .A2(n9995), .ZN(n14446) );
  INV_X1 U11937 ( .A(n9997), .ZN(n9995) );
  AND2_X1 U11938 ( .A1(n12453), .A2(n12452), .ZN(n13972) );
  NAND2_X1 U11939 ( .A1(n12172), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12212) );
  NOR2_X1 U11940 ( .A1(n12149), .A2(n14620), .ZN(n12150) );
  NAND2_X1 U11941 ( .A1(n12150), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12170) );
  AND2_X1 U11942 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  INV_X1 U11943 ( .A(n14412), .ZN(n10061) );
  NAND2_X1 U11944 ( .A1(n14421), .A2(n14422), .ZN(n14303) );
  NOR2_X1 U11945 ( .A1(n12109), .A2(n15729), .ZN(n12110) );
  NOR2_X1 U11946 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  NAND2_X1 U11947 ( .A1(n12059), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12109) );
  NOR2_X1 U11948 ( .A1(n12024), .A2(n14637), .ZN(n12025) );
  NAND2_X1 U11949 ( .A1(n12025), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12058) );
  NOR2_X1 U11950 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  NAND2_X1 U11951 ( .A1(n11990), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12024) );
  AND2_X1 U11952 ( .A1(n11959), .A2(n11958), .ZN(n14465) );
  NAND2_X1 U11953 ( .A1(n11934), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11956) );
  NOR2_X1 U11954 ( .A1(n20886), .A2(n11897), .ZN(n11934) );
  INV_X1 U11955 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20886) );
  NOR2_X1 U11956 ( .A1(n11904), .A2(n14490), .ZN(n11905) );
  INV_X1 U11957 ( .A(n11882), .ZN(n11897) );
  NAND2_X1 U11958 ( .A1(n11857), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11896) );
  CLKBUF_X1 U11959 ( .A(n14024), .Z(n14042) );
  AOI21_X1 U11960 ( .B1(n11837), .B2(n11674), .A(n11836), .ZN(n13971) );
  INV_X1 U11961 ( .A(n11798), .ZN(n11799) );
  NAND2_X1 U11962 ( .A1(n11799), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U11963 ( .A1(n11786), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11798) );
  INV_X1 U11964 ( .A(n13704), .ZN(n11773) );
  NAND2_X1 U11965 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11720) );
  NOR2_X1 U11966 ( .A1(n11720), .A2(n14385), .ZN(n11745) );
  NAND2_X1 U11967 ( .A1(n13502), .A2(n11695), .ZN(n13566) );
  NAND2_X1 U11968 ( .A1(n9844), .A2(n9843), .ZN(n14709) );
  NAND2_X1 U11969 ( .A1(n14708), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9844) );
  NAND2_X1 U11970 ( .A1(n14423), .A2(n9988), .ZN(n14417) );
  NAND2_X1 U11971 ( .A1(n14423), .A2(n14308), .ZN(n14415) );
  OR2_X1 U11972 ( .A1(n9697), .A2(n14432), .ZN(n14434) );
  NAND2_X1 U11973 ( .A1(n9801), .A2(n10202), .ZN(n12398) );
  NAND2_X1 U11974 ( .A1(n14650), .A2(n10204), .ZN(n9801) );
  AOI21_X1 U11975 ( .B1(n10204), .B2(n10206), .A(n10203), .ZN(n10202) );
  NAND2_X1 U11976 ( .A1(n10201), .A2(n14645), .ZN(n10200) );
  OR2_X1 U11977 ( .A1(n10204), .A2(n10199), .ZN(n10198) );
  INV_X1 U11978 ( .A(n14645), .ZN(n10199) );
  NOR2_X1 U11979 ( .A1(n14460), .A2(n14318), .ZN(n14320) );
  OR2_X1 U11980 ( .A1(n14458), .A2(n14457), .ZN(n14460) );
  AND2_X1 U11981 ( .A1(n14345), .A2(n9991), .ZN(n14469) );
  NAND2_X1 U11982 ( .A1(n14345), .A2(n9993), .ZN(n14479) );
  NAND2_X1 U11983 ( .A1(n14345), .A2(n14038), .ZN(n14477) );
  AND2_X1 U11984 ( .A1(n15858), .A2(n12395), .ZN(n15846) );
  NOR2_X1 U11985 ( .A1(n14488), .A2(n14346), .ZN(n14345) );
  OR2_X1 U11986 ( .A1(n14486), .A2(n14485), .ZN(n14488) );
  NAND2_X1 U11987 ( .A1(n14027), .A2(n14026), .ZN(n14047) );
  OR2_X1 U11988 ( .A1(n14047), .A2(n14048), .ZN(n14486) );
  NAND2_X1 U11989 ( .A1(n10176), .A2(n10181), .ZN(n14689) );
  NAND2_X1 U11990 ( .A1(n13991), .A2(n12388), .ZN(n10176) );
  AND2_X1 U11991 ( .A1(n9981), .A2(n9979), .ZN(n13973) );
  NOR2_X1 U11992 ( .A1(n9976), .A2(n12442), .ZN(n9979) );
  NAND2_X1 U11993 ( .A1(n15891), .A2(n10186), .ZN(n10185) );
  NAND2_X1 U11994 ( .A1(n12310), .A2(n12309), .ZN(n20064) );
  INV_X1 U11995 ( .A(n13082), .ZN(n13345) );
  INV_X1 U11996 ( .A(n11557), .ZN(n14755) );
  AND2_X1 U11997 ( .A1(n20710), .A2(n20106), .ZN(n20214) );
  AND2_X1 U11998 ( .A1(n20185), .A2(n20109), .ZN(n20444) );
  AND2_X1 U11999 ( .A1(n9672), .A2(n20108), .ZN(n20584) );
  AOI21_X1 U12000 ( .B1(n20504), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20254), 
        .ZN(n20588) );
  NAND2_X1 U12001 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20115), .ZN(n20148) );
  AND2_X1 U12002 ( .A1(n20643), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12294) );
  OR2_X1 U12003 ( .A1(n16140), .A2(n19047), .ZN(n10172) );
  NOR2_X1 U12004 ( .A1(n10889), .A2(n10046), .ZN(n16127) );
  NAND2_X1 U12005 ( .A1(n10893), .A2(n10047), .ZN(n10046) );
  NOR2_X1 U12006 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(P2_EBX_REG_26__SCAN_IN), 
        .ZN(n10047) );
  OR2_X1 U12007 ( .A1(n16127), .A2(n10831), .ZN(n10902) );
  AND2_X1 U12008 ( .A1(n10149), .A2(n19029), .ZN(n16153) );
  OR2_X1 U12009 ( .A1(n14786), .A2(n14997), .ZN(n10149) );
  NAND2_X1 U12010 ( .A1(n9869), .A2(n9868), .ZN(n10889) );
  INV_X1 U12011 ( .A(n10882), .ZN(n9868) );
  INV_X1 U12012 ( .A(n10883), .ZN(n9869) );
  NAND2_X1 U12013 ( .A1(n10819), .A2(n9690), .ZN(n10877) );
  NAND2_X1 U12014 ( .A1(n10874), .A2(n10875), .ZN(n10883) );
  INV_X1 U12015 ( .A(n10819), .ZN(n10838) );
  NAND2_X1 U12016 ( .A1(n18982), .A2(n10037), .ZN(n10852) );
  AND2_X1 U12017 ( .A1(n18982), .A2(n9739), .ZN(n10845) );
  NOR2_X1 U12018 ( .A1(n9665), .A2(n10998), .ZN(n10788) );
  NOR2_X1 U12019 ( .A1(n10799), .A2(n10788), .ZN(n10798) );
  INV_X1 U12020 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13824) );
  NOR2_X1 U12021 ( .A1(n10074), .A2(n10078), .ZN(n10073) );
  INV_X1 U12022 ( .A(n10076), .ZN(n10074) );
  NAND2_X1 U12023 ( .A1(n10113), .A2(n10114), .ZN(n10112) );
  XNOR2_X1 U12024 ( .A(n12829), .B(n9788), .ZN(n9787) );
  XNOR2_X1 U12025 ( .A(n12802), .B(n12804), .ZN(n14817) );
  NAND2_X1 U12026 ( .A1(n14817), .A2(n14816), .ZN(n14815) );
  NOR2_X1 U12027 ( .A1(n14908), .A2(n10129), .ZN(n14899) );
  INV_X1 U12028 ( .A(n10131), .ZN(n10129) );
  INV_X1 U12029 ( .A(n14920), .ZN(n10107) );
  AND2_X1 U12030 ( .A1(n12658), .A2(n9765), .ZN(n14938) );
  NAND2_X1 U12031 ( .A1(n12658), .A2(n12657), .ZN(n14936) );
  CLKBUF_X1 U12032 ( .A(n14849), .Z(n16185) );
  NAND2_X1 U12033 ( .A1(n15286), .A2(n15287), .ZN(n16306) );
  AND2_X1 U12034 ( .A1(n19151), .A2(n19150), .ZN(n19184) );
  OR2_X1 U12035 ( .A1(n13636), .A2(n12979), .ZN(n13052) );
  INV_X1 U12036 ( .A(n13132), .ZN(n14220) );
  NOR2_X1 U12037 ( .A1(n14806), .A2(n11063), .ZN(n12564) );
  NOR3_X2 U12038 ( .A1(n13777), .A2(n10079), .A3(n14847), .ZN(n15057) );
  NAND2_X1 U12039 ( .A1(n10156), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10155) );
  INV_X1 U12040 ( .A(n12955), .ZN(n10154) );
  NAND2_X1 U12041 ( .A1(n12959), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12961) );
  NAND2_X1 U12042 ( .A1(n11073), .A2(n10239), .ZN(n10236) );
  NOR2_X1 U12043 ( .A1(n9733), .A2(n11103), .ZN(n10212) );
  AOI21_X1 U12044 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(n10024) );
  AND2_X1 U12045 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11182), .ZN(
        n12562) );
  NOR2_X1 U12046 ( .A1(n10905), .A2(n9731), .ZN(n9880) );
  NAND2_X1 U12047 ( .A1(n14810), .A2(n14804), .ZN(n14806) );
  NAND2_X1 U12048 ( .A1(n9972), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9971) );
  NAND2_X1 U12049 ( .A1(n10221), .A2(n15154), .ZN(n10219) );
  NAND2_X1 U12050 ( .A1(n14994), .A2(n10220), .ZN(n10218) );
  NOR3_X1 U12051 ( .A1(n14831), .A2(n10085), .A3(n14830), .ZN(n14827) );
  NOR2_X1 U12052 ( .A1(n14908), .A2(n14909), .ZN(n14910) );
  NOR2_X1 U12053 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  AOI21_X1 U12054 ( .B1(n9919), .B2(n15027), .A(n15040), .ZN(n9918) );
  INV_X1 U12055 ( .A(n15025), .ZN(n9919) );
  INV_X1 U12056 ( .A(n15027), .ZN(n9920) );
  NAND2_X1 U12057 ( .A1(n16271), .A2(n9676), .ZN(n14949) );
  INV_X1 U12058 ( .A(n13950), .ZN(n10124) );
  AOI21_X1 U12059 ( .B1(n15251), .B2(n9937), .A(n9935), .ZN(n15075) );
  AND2_X1 U12060 ( .A1(n9938), .A2(n15621), .ZN(n9937) );
  OAI21_X1 U12061 ( .B1(n9686), .B2(n9936), .A(n9741), .ZN(n9935) );
  INV_X1 U12062 ( .A(n15621), .ZN(n9936) );
  AND2_X1 U12063 ( .A1(n15021), .A2(n15022), .ZN(n15076) );
  NAND2_X1 U12064 ( .A1(n16271), .A2(n16272), .ZN(n16273) );
  NAND2_X1 U12065 ( .A1(n15082), .A2(n15239), .ZN(n16209) );
  NOR2_X1 U12066 ( .A1(n13777), .A2(n13778), .ZN(n13833) );
  NAND2_X1 U12067 ( .A1(n15251), .A2(n9942), .ZN(n9941) );
  AND2_X1 U12068 ( .A1(n15251), .A2(n15019), .ZN(n16214) );
  AOI21_X1 U12069 ( .B1(n9931), .B2(n9930), .A(n9750), .ZN(n9929) );
  INV_X1 U12070 ( .A(n10225), .ZN(n9930) );
  INV_X1 U12071 ( .A(n13658), .ZN(n10086) );
  INV_X1 U12072 ( .A(n16296), .ZN(n10125) );
  OR2_X1 U12073 ( .A1(n15274), .A2(n16252), .ZN(n9858) );
  NAND2_X1 U12074 ( .A1(n13484), .A2(n10087), .ZN(n13659) );
  NAND2_X1 U12075 ( .A1(n9857), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9861) );
  INV_X1 U12076 ( .A(n16251), .ZN(n9857) );
  NAND2_X1 U12077 ( .A1(n13484), .A2(n13485), .ZN(n13483) );
  NAND2_X1 U12078 ( .A1(n13854), .A2(n13853), .ZN(n9878) );
  XNOR2_X1 U12079 ( .A(n10740), .B(n10739), .ZN(n13854) );
  AOI21_X1 U12080 ( .B1(n10015), .B2(n10021), .A(n9752), .ZN(n10011) );
  OR2_X1 U12081 ( .A1(n11210), .A2(n11215), .ZN(n13170) );
  NAND2_X1 U12082 ( .A1(n10097), .A2(n10100), .ZN(n13231) );
  NAND2_X1 U12083 ( .A1(n9737), .A2(n12592), .ZN(n10100) );
  NAND2_X1 U12084 ( .A1(n10101), .A2(n10102), .ZN(n10097) );
  XNOR2_X1 U12085 ( .A(n12594), .B(n12595), .ZN(n13232) );
  NOR2_X1 U12086 ( .A1(n13183), .A2(n11232), .ZN(n13739) );
  NAND2_X1 U12087 ( .A1(n12587), .A2(n19888), .ZN(n12602) );
  NAND2_X1 U12088 ( .A1(n9640), .A2(n10273), .ZN(n13559) );
  NAND2_X1 U12089 ( .A1(n11127), .A2(n11125), .ZN(n13641) );
  NAND2_X1 U12090 ( .A1(n10367), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10368) );
  NOR2_X1 U12091 ( .A1(n13827), .A2(n10498), .ZN(n10499) );
  INV_X1 U12092 ( .A(n10476), .ZN(n10475) );
  INV_X1 U12093 ( .A(n19330), .ZN(n19333) );
  NOR2_X1 U12094 ( .A1(n10500), .A2(n10498), .ZN(n10492) );
  NOR2_X2 U12095 ( .A1(n14220), .A2(n13762), .ZN(n19261) );
  NOR2_X2 U12096 ( .A1(n14221), .A2(n13762), .ZN(n19262) );
  AND2_X1 U12097 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19702), .ZN(n19258) );
  AND2_X1 U12098 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19692), .ZN(
        n12598) );
  INV_X1 U12099 ( .A(n19447), .ZN(n19702) );
  NAND2_X1 U12100 ( .A1(n15606), .A2(n14176), .ZN(n14206) );
  NAND2_X1 U12101 ( .A1(n15601), .A2(n18656), .ZN(n18623) );
  INV_X1 U12102 ( .A(n15605), .ZN(n18624) );
  OR2_X1 U12103 ( .A1(n18661), .A2(n14085), .ZN(n9694) );
  OR2_X1 U12104 ( .A1(n9887), .A2(n9886), .ZN(n9885) );
  INV_X1 U12105 ( .A(n15492), .ZN(n9823) );
  NOR2_X1 U12106 ( .A1(n15491), .A2(n9822), .ZN(n9821) );
  NOR2_X1 U12107 ( .A1(n9820), .A2(n9819), .ZN(n9818) );
  INV_X1 U12108 ( .A(n18195), .ZN(n15695) );
  INV_X1 U12109 ( .A(n14194), .ZN(n18645) );
  NOR2_X1 U12110 ( .A1(n17427), .A2(n17389), .ZN(n17406) );
  NAND2_X1 U12111 ( .A1(n16379), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16353) );
  NOR2_X1 U12112 ( .A1(n17628), .A2(n17629), .ZN(n17610) );
  NOR2_X1 U12113 ( .A1(n17662), .A2(n17663), .ZN(n17648) );
  NAND2_X1 U12114 ( .A1(n17688), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17662) );
  AND2_X1 U12115 ( .A1(n17697), .A2(n17702), .ZN(n17688) );
  AOI21_X1 U12116 ( .B1(n17615), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18570), .ZN(n17700) );
  INV_X1 U12117 ( .A(n16859), .ZN(n17830) );
  INV_X1 U12118 ( .A(n17868), .ZN(n17829) );
  NAND2_X1 U12119 ( .A1(n9824), .A2(n17504), .ZN(n15556) );
  NAND2_X1 U12120 ( .A1(n10135), .A2(n9825), .ZN(n9824) );
  NAND2_X1 U12121 ( .A1(n17514), .A2(n17500), .ZN(n9825) );
  NOR2_X1 U12122 ( .A1(n15515), .A2(n15514), .ZN(n16409) );
  INV_X1 U12123 ( .A(n10135), .ZN(n16408) );
  NOR2_X1 U12124 ( .A1(n17912), .A2(n17919), .ZN(n17544) );
  NAND2_X1 U12125 ( .A1(n17591), .A2(n17920), .ZN(n17912) );
  NAND2_X1 U12126 ( .A1(n17920), .A2(n18014), .ZN(n17910) );
  OR2_X1 U12127 ( .A1(n18087), .A2(n18203), .ZN(n18629) );
  INV_X1 U12128 ( .A(n17659), .ZN(n17593) );
  NAND2_X1 U12129 ( .A1(n17659), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15547) );
  AND2_X1 U12130 ( .A1(n17999), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17975) );
  NAND2_X1 U12131 ( .A1(n17734), .A2(n17975), .ZN(n18009) );
  INV_X1 U12132 ( .A(n18051), .ZN(n17734) );
  INV_X1 U12133 ( .A(n18639), .ZN(n18648) );
  NOR2_X1 U12134 ( .A1(n17792), .A2(n18104), .ZN(n17791) );
  NAND2_X1 U12135 ( .A1(n10147), .A2(n10143), .ZN(n10142) );
  INV_X1 U12136 ( .A(n10146), .ZN(n10143) );
  INV_X1 U12137 ( .A(n18629), .ZN(n18054) );
  NOR2_X1 U12138 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18194), .ZN(n18543) );
  NOR2_X1 U12139 ( .A1(n14105), .A2(n14104), .ZN(n18213) );
  INV_X1 U12140 ( .A(n18543), .ZN(n18265) );
  OAI22_X1 U12141 ( .A1(n16349), .A2(n18629), .B1(n18625), .B2(n16407), .ZN(
        n18631) );
  CLKBUF_X1 U12142 ( .A(n13132), .Z(n14221) );
  INV_X1 U12143 ( .A(n15771), .ZN(n15803) );
  AND2_X1 U12144 ( .A1(n15779), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19977) );
  AND2_X1 U12145 ( .A1(n15779), .A2(n13841), .ZN(n19989) );
  AND2_X1 U12146 ( .A1(n12533), .A2(n12521), .ZN(n19994) );
  INV_X1 U12147 ( .A(n14494), .ZN(n20003) );
  INV_X1 U12148 ( .A(n20008), .ZN(n14483) );
  AND2_X2 U12149 ( .A1(n13352), .A2(n13578), .ZN(n20008) );
  NAND2_X1 U12150 ( .A1(n14270), .A2(n14260), .ZN(n10069) );
  AND2_X1 U12151 ( .A1(n9648), .A2(n13583), .ZN(n14503) );
  INV_X1 U12152 ( .A(n14503), .ZN(n14559) );
  INV_X1 U12153 ( .A(n14508), .ZN(n14561) );
  NAND2_X1 U12154 ( .A1(n13579), .A2(n13578), .ZN(n14567) );
  NAND2_X1 U12155 ( .A1(n13577), .A2(n13576), .ZN(n13579) );
  INV_X1 U12156 ( .A(n14568), .ZN(n14571) );
  INV_X2 U12157 ( .A(n20010), .ZN(n20030) );
  XNOR2_X1 U12158 ( .A(n14600), .B(n14599), .ZN(n15907) );
  NAND2_X1 U12159 ( .A1(n10249), .A2(n14598), .ZN(n14600) );
  AND2_X1 U12160 ( .A1(n14455), .A2(n14316), .ZN(n14450) );
  INV_X1 U12161 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14637) );
  INV_X1 U12162 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19964) );
  NAND2_X1 U12163 ( .A1(n19920), .A2(n12301), .ZN(n15902) );
  NAND2_X1 U12164 ( .A1(n11680), .A2(n11695), .ZN(n13500) );
  INV_X1 U12165 ( .A(n15902), .ZN(n20068) );
  OAI21_X1 U12166 ( .B1(n15907), .B2(n16073), .A(n15906), .ZN(n15908) );
  NAND2_X1 U12167 ( .A1(n15919), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15906) );
  OR2_X1 U12168 ( .A1(n14284), .A2(n14283), .ZN(n15911) );
  AND2_X1 U12169 ( .A1(n16049), .A2(n15960), .ZN(n9830) );
  NAND2_X1 U12170 ( .A1(n10180), .A2(n12388), .ZN(n13999) );
  OR2_X1 U12171 ( .A1(n13991), .A2(n12387), .ZN(n10180) );
  NAND2_X1 U12172 ( .A1(n9981), .A2(n9980), .ZN(n13789) );
  INV_X1 U12173 ( .A(n9982), .ZN(n9980) );
  NAND2_X1 U12174 ( .A1(n10187), .A2(n12357), .ZN(n15893) );
  OR2_X1 U12175 ( .A1(n12305), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16057) );
  INV_X1 U12176 ( .A(n20097), .ZN(n14699) );
  INV_X1 U12177 ( .A(n14706), .ZN(n20092) );
  NAND2_X1 U12178 ( .A1(n13414), .A2(n13401), .ZN(n20093) );
  INV_X1 U12179 ( .A(n20718), .ZN(n20590) );
  INV_X1 U12180 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20101) );
  NOR2_X1 U12181 ( .A1(n20479), .A2(n13391), .ZN(n15671) );
  NOR2_X1 U12182 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16083) );
  OAI21_X1 U12183 ( .B1(n20272), .B2(n20255), .A(n20541), .ZN(n20274) );
  AND2_X1 U12184 ( .A1(n20337), .A2(n20534), .ZN(n20349) );
  NOR2_X1 U12185 ( .A1(n20504), .A2(n20335), .ZN(n20356) );
  OAI211_X1 U12186 ( .C1(n20381), .C2(n20479), .A(n20416), .B(n20365), .ZN(
        n20383) );
  INV_X1 U12187 ( .A(n20443), .ZN(n20435) );
  OAI22_X1 U12188 ( .A1(n20422), .A2(n20421), .B1(n20420), .B2(n20533), .ZN(
        n20439) );
  OAI21_X1 U12189 ( .B1(n20422), .B2(n20419), .A(n20418), .ZN(n20440) );
  INV_X1 U12190 ( .A(n20467), .ZN(n20470) );
  NOR2_X1 U12191 ( .A1(n20504), .A2(n20581), .ZN(n20634) );
  AND2_X1 U12192 ( .A1(n20584), .A2(n20534), .ZN(n20637) );
  INV_X1 U12193 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20643) );
  NAND2_X1 U12194 ( .A1(n19047), .A2(n10168), .ZN(n10167) );
  INV_X1 U12195 ( .A(n14771), .ZN(n10168) );
  NOR2_X1 U12196 ( .A1(n16163), .A2(n19047), .ZN(n14786) );
  INV_X1 U12197 ( .A(n10149), .ZN(n14785) );
  NAND2_X1 U12198 ( .A1(n19047), .A2(n10161), .ZN(n10159) );
  NOR2_X1 U12199 ( .A1(n18890), .A2(n18891), .ZN(n18889) );
  NOR2_X1 U12200 ( .A1(n18906), .A2(n19047), .ZN(n18890) );
  INV_X1 U12201 ( .A(n19024), .ZN(n19062) );
  AND2_X1 U12202 ( .A1(n13040), .A2(n12991), .ZN(n19045) );
  INV_X1 U12203 ( .A(n18958), .ZN(n19067) );
  CLKBUF_X1 U12204 ( .A(n13779), .Z(n13831) );
  AND2_X1 U12205 ( .A1(n9736), .A2(n12616), .ZN(n9790) );
  INV_X1 U12206 ( .A(n16181), .ZN(n19079) );
  XNOR2_X1 U12207 ( .A(n13373), .B(n13374), .ZN(n19113) );
  NAND2_X1 U12208 ( .A1(n13154), .A2(n12925), .ZN(n12926) );
  NOR2_X1 U12209 ( .A1(n12566), .A2(n12565), .ZN(n12974) );
  OAI211_X1 U12210 ( .C1(n14791), .C2(n10095), .A(n10093), .B(n10092), .ZN(
        n14227) );
  NAND2_X1 U12211 ( .A1(n9691), .A2(n12923), .ZN(n10095) );
  NAND2_X1 U12212 ( .A1(n10094), .A2(n9774), .ZN(n10093) );
  AND2_X1 U12213 ( .A1(n19111), .A2(n13228), .ZN(n16190) );
  AND2_X1 U12214 ( .A1(n15286), .A2(n10127), .ZN(n15277) );
  NAND2_X1 U12215 ( .A1(n19111), .A2(n13238), .ZN(n14962) );
  INV_X1 U12216 ( .A(n19890), .ZN(n19142) );
  INV_X1 U12217 ( .A(n19111), .ZN(n19137) );
  INV_X1 U12218 ( .A(n14962), .ZN(n19138) );
  NOR2_X1 U12219 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13758), .ZN(n19215) );
  INV_X2 U12220 ( .A(n19147), .ZN(n13147) );
  NOR2_X1 U12221 ( .A1(n19234), .A2(n10235), .ZN(n10234) );
  INV_X1 U12222 ( .A(n10236), .ZN(n10235) );
  INV_X1 U12223 ( .A(n16202), .ZN(n15237) );
  INV_X1 U12224 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16198) );
  NAND2_X1 U12225 ( .A1(n15102), .A2(n15103), .ZN(n9947) );
  INV_X1 U12226 ( .A(n19234), .ZN(n19224) );
  INV_X1 U12227 ( .A(n19239), .ZN(n16206) );
  INV_X1 U12228 ( .A(n19229), .ZN(n19230) );
  XOR2_X1 U12229 ( .A(n12928), .B(n12927), .Z(n14250) );
  NAND2_X1 U12230 ( .A1(n10001), .A2(n10005), .ZN(n15003) );
  NAND2_X1 U12231 ( .A1(n10873), .A2(n9702), .ZN(n10001) );
  NAND2_X1 U12232 ( .A1(n10009), .A2(n10007), .ZN(n15010) );
  NAND2_X1 U12233 ( .A1(n10873), .A2(n10262), .ZN(n10009) );
  NAND2_X1 U12234 ( .A1(n16330), .A2(n15238), .ZN(n9895) );
  INV_X1 U12235 ( .A(n9894), .ZN(n9893) );
  AOI21_X1 U12236 ( .B1(n16277), .B2(n15240), .A(n16276), .ZN(n9894) );
  NAND2_X1 U12237 ( .A1(n9934), .A2(n9686), .ZN(n15620) );
  NAND2_X1 U12238 ( .A1(n15251), .A2(n9938), .ZN(n9934) );
  AND2_X1 U12239 ( .A1(n15267), .A2(n9960), .ZN(n9959) );
  AOI21_X1 U12240 ( .B1(n15262), .B2(n15261), .A(n9961), .ZN(n9960) );
  NAND2_X1 U12241 ( .A1(n15104), .A2(n10225), .ZN(n9933) );
  NAND2_X1 U12242 ( .A1(n10228), .A2(n10227), .ZN(n16247) );
  INV_X1 U12243 ( .A(n15082), .ZN(n15098) );
  AND2_X1 U12244 ( .A1(n10949), .A2(n10948), .ZN(n9967) );
  OAI21_X1 U12245 ( .B1(n13732), .B2(n11098), .A(n10018), .ZN(n13725) );
  NAND2_X1 U12246 ( .A1(n10014), .A2(n10020), .ZN(n13724) );
  AND2_X1 U12247 ( .A1(n11198), .A2(n11192), .ZN(n16312) );
  INV_X1 U12248 ( .A(n16324), .ZN(n16301) );
  INV_X1 U12249 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19886) );
  AND2_X1 U12250 ( .A1(n19864), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19876) );
  NAND2_X1 U12251 ( .A1(n13230), .A2(n13233), .ZN(n19883) );
  OR2_X1 U12252 ( .A1(n13232), .A2(n13231), .ZN(n13233) );
  INV_X1 U12253 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12599) );
  XNOR2_X1 U12254 ( .A(n13292), .B(n13291), .ZN(n13294) );
  INV_X1 U12255 ( .A(n19883), .ZN(n19854) );
  INV_X1 U12256 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13168) );
  INV_X1 U12257 ( .A(n19351), .ZN(n19353) );
  OAI21_X1 U12258 ( .B1(n19383), .B2(n19888), .A(n19368), .ZN(n19385) );
  INV_X1 U12259 ( .A(n19420), .ZN(n19438) );
  INV_X1 U12260 ( .A(n19523), .ZN(n19547) );
  INV_X1 U12261 ( .A(n19737), .ZN(n19606) );
  INV_X1 U12262 ( .A(n19743), .ZN(n19639) );
  NOR2_X1 U12263 ( .A1(n19648), .A2(n19624), .ZN(n19644) );
  INV_X1 U12264 ( .A(n19753), .ZN(n19678) );
  OAI21_X1 U12265 ( .B1(n19660), .B2(n19659), .A(n19658), .ZN(n19685) );
  INV_X1 U12266 ( .A(n19681), .ZN(n19683) );
  INV_X1 U12267 ( .A(n19242), .ZN(n19695) );
  INV_X1 U12268 ( .A(n19597), .ZN(n19710) );
  INV_X1 U12269 ( .A(n19274), .ZN(n19708) );
  INV_X1 U12270 ( .A(n19669), .ZN(n19716) );
  INV_X1 U12271 ( .A(n19280), .ZN(n19720) );
  INV_X1 U12272 ( .A(n19605), .ZN(n19728) );
  AND2_X1 U12273 ( .A1(n19245), .A2(n19258), .ZN(n19726) );
  OAI22_X1 U12274 ( .A1(n19254), .A2(n19253), .B1(n19252), .B2(n19251), .ZN(
        n19734) );
  AND2_X1 U12275 ( .A1(n9665), .A2(n19258), .ZN(n19732) );
  AND2_X1 U12276 ( .A1(n12598), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19745) );
  NOR2_X2 U12277 ( .A1(n19625), .A2(n19698), .ZN(n19749) );
  INV_X1 U12278 ( .A(n19289), .ZN(n19744) );
  INV_X1 U12279 ( .A(n13163), .ZN(n16343) );
  AND3_X1 U12280 ( .A1(n13654), .A2(n13653), .A3(n13652), .ZN(n16342) );
  NAND2_X1 U12281 ( .A1(n18631), .A2(n18836), .ZN(n16525) );
  NAND2_X1 U12282 ( .A1(n16666), .A2(n16909), .ZN(n16659) );
  NAND2_X1 U12283 ( .A1(n16674), .A2(n16909), .ZN(n16667) );
  NAND2_X1 U12284 ( .A1(n16667), .A2(n17598), .ZN(n16666) );
  NOR2_X1 U12285 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16740), .ZN(n16720) );
  NOR2_X2 U12286 ( .A1(n18791), .A2(n16907), .ZN(n16887) );
  NOR2_X2 U12287 ( .A1(n16544), .A2(n16547), .ZN(n16900) );
  OAI211_X1 U12288 ( .C1(n18788), .C2(n18684), .A(n16541), .B(n18853), .ZN(
        n16923) );
  INV_X1 U12289 ( .A(n17356), .ZN(n17352) );
  INV_X1 U12290 ( .A(n17261), .ZN(n17258) );
  NOR2_X1 U12291 ( .A1(n17281), .A2(n17307), .ZN(n17297) );
  NOR2_X2 U12292 ( .A1(n14117), .A2(n14116), .ZN(n17342) );
  NOR2_X1 U12293 ( .A1(n15450), .A2(n15449), .ZN(n17360) );
  NOR2_X1 U12294 ( .A1(n17462), .A2(n17352), .ZN(n17374) );
  INV_X1 U12295 ( .A(n15480), .ZN(n15481) );
  NOR2_X1 U12296 ( .A1(n18645), .A2(n15699), .ZN(n17381) );
  INV_X1 U12297 ( .A(n17384), .ZN(n15699) );
  NOR2_X1 U12298 ( .A1(n15699), .A2(n15698), .ZN(n17382) );
  INV_X1 U12299 ( .A(n17381), .ZN(n17376) );
  NOR2_X1 U12300 ( .A1(n18838), .A2(n17406), .ZN(n17416) );
  CLKBUF_X1 U12301 ( .A(n17416), .Z(n17423) );
  NOR2_X1 U12303 ( .A1(n17540), .A2(n17541), .ZN(n17530) );
  INV_X1 U12304 ( .A(n17780), .ZN(n17733) );
  NAND2_X1 U12305 ( .A1(n17633), .A2(n17920), .ZN(n17562) );
  NOR2_X1 U12306 ( .A1(n17585), .A2(n17586), .ZN(n17568) );
  AND2_X1 U12307 ( .A1(n17766), .A2(n17975), .ZN(n17633) );
  INV_X1 U12308 ( .A(n17633), .ZN(n17670) );
  INV_X1 U12309 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17721) );
  INV_X1 U12310 ( .A(n17672), .ZN(n17730) );
  NOR2_X1 U12311 ( .A1(n17871), .A2(n17354), .ZN(n17780) );
  INV_X1 U12312 ( .A(n16745), .ZN(n17787) );
  INV_X1 U12313 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17806) );
  NAND2_X1 U12314 ( .A1(n16859), .A2(n9720), .ZN(n17799) );
  INV_X1 U12315 ( .A(n17611), .ZN(n18266) );
  NOR2_X1 U12316 ( .A1(n17831), .A2(n17829), .ZN(n17865) );
  NAND2_X1 U12317 ( .A1(n17672), .A2(n17617), .ZN(n17860) );
  INV_X1 U12318 ( .A(n17871), .ZN(n17861) );
  OR2_X1 U12319 ( .A1(n16525), .A2(n18841), .ZN(n17871) );
  INV_X1 U12320 ( .A(n17842), .ZN(n17872) );
  OAI21_X1 U12321 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18835), .A(n16525), 
        .ZN(n17868) );
  NAND2_X1 U12322 ( .A1(n16361), .A2(n16362), .ZN(n9817) );
  INV_X1 U12323 ( .A(n16362), .ZN(n9815) );
  NAND2_X1 U12324 ( .A1(n17570), .A2(n15551), .ZN(n17552) );
  NAND2_X1 U12325 ( .A1(n17604), .A2(n15552), .ZN(n17571) );
  NAND2_X1 U12326 ( .A1(n18061), .A2(n18657), .ZN(n18087) );
  NOR2_X1 U12327 ( .A1(n17706), .A2(n17739), .ZN(n18094) );
  NAND2_X1 U12328 ( .A1(n15536), .A2(n17820), .ZN(n17813) );
  AND3_X1 U12329 ( .A1(n15536), .A2(n17820), .A3(n10145), .ZN(n17811) );
  INV_X1 U12330 ( .A(n9803), .ZN(n18140) );
  OAI221_X2 U12331 ( .B1(n15570), .B2(n16348), .C1(n15570), .C2(n15569), .A(
        n18836), .ZN(n18167) );
  INV_X1 U12332 ( .A(n18167), .ZN(n18175) );
  INV_X1 U12333 ( .A(n18172), .ZN(n18178) );
  INV_X1 U12334 ( .A(n18638), .ZN(n18640) );
  NOR2_X1 U12335 ( .A1(n18788), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18692) );
  AND2_X1 U12336 ( .A1(n13011), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20102)
         );
  NOR3_X1 U12338 ( .A1(n14715), .A2(n14714), .A3(n9828), .ZN(n9827) );
  INV_X1 U12339 ( .A(n12404), .ZN(n9793) );
  AOI21_X1 U12340 ( .B1(n9833), .B2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n9780), .ZN(n15964) );
  AND2_X1 U12341 ( .A1(n9832), .A2(n9831), .ZN(n14745) );
  NAND2_X1 U12342 ( .A1(n9833), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9831) );
  OAI21_X1 U12343 ( .B1(n15164), .B2(n19234), .A(n9849), .ZN(P2_U2990) );
  INV_X1 U12344 ( .A(n9850), .ZN(n9849) );
  AOI21_X1 U12345 ( .B1(n16173), .B2(n19239), .A(n15000), .ZN(n9851) );
  INV_X1 U12346 ( .A(n15037), .ZN(n9922) );
  NAND2_X1 U12347 ( .A1(n12541), .A2(n16334), .ZN(n12557) );
  AND2_X1 U12348 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  INV_X1 U12349 ( .A(n9862), .ZN(n16292) );
  NAND2_X1 U12350 ( .A1(n9964), .A2(n9957), .ZN(P2_U3033) );
  INV_X1 U12351 ( .A(n9958), .ZN(n9957) );
  NAND2_X1 U12352 ( .A1(n16223), .A2(n16313), .ZN(n9964) );
  OAI21_X1 U12353 ( .B1(n15268), .B2(n16317), .A(n9959), .ZN(n9958) );
  OR2_X1 U12354 ( .A1(n16577), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9884) );
  OAI21_X1 U12355 ( .B1(n16376), .B2(n17783), .A(n9888), .ZN(P3_U2800) );
  NOR2_X1 U12356 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  NOR3_X1 U12357 ( .A1(n17523), .A2(n16371), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9890) );
  OAI21_X1 U12358 ( .B1(n16374), .B2(n16393), .A(n16375), .ZN(n9889) );
  NAND2_X1 U12359 ( .A1(n9813), .A2(n9811), .ZN(P3_U2831) );
  AOI21_X1 U12360 ( .B1(n16399), .B2(n18178), .A(n9812), .ZN(n9811) );
  NAND2_X1 U12361 ( .A1(n16398), .A2(n18076), .ZN(n9813) );
  OAI21_X1 U12362 ( .B1(n16401), .B2(n17974), .A(n16400), .ZN(n9812) );
  NAND2_X1 U12363 ( .A1(n12658), .A2(n9687), .ZN(n14839) );
  OR2_X1 U12364 ( .A1(n14774), .A2(n10801), .ZN(n11092) );
  INV_X1 U12365 ( .A(n10684), .ZN(n10686) );
  AND2_X1 U12366 ( .A1(n9680), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9675) );
  NAND2_X1 U12367 ( .A1(n12943), .A2(n9680), .ZN(n12941) );
  AND2_X1 U12368 ( .A1(n9688), .A2(n15244), .ZN(n9676) );
  INV_X2 U12369 ( .A(n12733), .ZN(n10511) );
  AND2_X2 U12370 ( .A1(n11215), .A2(n19888), .ZN(n11211) );
  NAND2_X1 U12371 ( .A1(n15082), .A2(n10241), .ZN(n15055) );
  NAND2_X1 U12372 ( .A1(n9641), .A2(n10240), .ZN(n14977) );
  NAND2_X1 U12373 ( .A1(n10154), .A2(n10156), .ZN(n12954) );
  OR2_X1 U12374 ( .A1(n12952), .A2(n10164), .ZN(n9677) );
  OR2_X1 U12375 ( .A1(n15009), .A2(n15179), .ZN(n9678) );
  OR2_X1 U12376 ( .A1(n13784), .A2(n13838), .ZN(n9679) );
  AND2_X1 U12377 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U12378 ( .A1(n9878), .A2(n10741), .ZN(n15112) );
  OR2_X1 U12379 ( .A1(n9766), .A2(n10229), .ZN(n9681) );
  AOI21_X1 U12380 ( .B1(n11092), .B2(n12561), .A(n9749), .ZN(n10030) );
  INV_X1 U12381 ( .A(n10030), .ZN(n10026) );
  AND2_X1 U12382 ( .A1(n10119), .A2(n13862), .ZN(n9682) );
  INV_X1 U12383 ( .A(n10031), .ZN(n11137) );
  OAI21_X1 U12384 ( .B1(n15104), .B2(n9932), .A(n9929), .ZN(n16231) );
  AND2_X1 U12385 ( .A1(n10192), .A2(n10194), .ZN(n9683) );
  NAND2_X1 U12386 ( .A1(n11163), .A2(n10395), .ZN(n11158) );
  INV_X1 U12387 ( .A(n11158), .ZN(n11161) );
  AND2_X1 U12388 ( .A1(n9675), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9684) );
  OAI21_X1 U12389 ( .B1(n10005), .B2(n10003), .A(n9751), .ZN(n10002) );
  INV_X1 U12390 ( .A(n13183), .ZN(n10120) );
  INV_X1 U12391 ( .A(n12393), .ZN(n15874) );
  AND2_X1 U12392 ( .A1(n12943), .A2(n9675), .ZN(n9685) );
  OR2_X1 U12393 ( .A1(n9939), .A2(n15020), .ZN(n9686) );
  NAND2_X1 U12394 ( .A1(n12940), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12936) );
  AND2_X1 U12395 ( .A1(n9765), .A2(n14840), .ZN(n9687) );
  AND2_X1 U12396 ( .A1(n10124), .A2(n16272), .ZN(n9688) );
  AND2_X1 U12397 ( .A1(n10151), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9689) );
  INV_X1 U12398 ( .A(n10021), .ZN(n10020) );
  OAI21_X1 U12399 ( .B1(n10022), .B2(n10801), .A(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10021) );
  AND2_X1 U12400 ( .A1(n10035), .A2(n10821), .ZN(n9690) );
  INV_X1 U12401 ( .A(n10019), .ZN(n10018) );
  NAND2_X1 U12402 ( .A1(n13888), .A2(n10662), .ZN(n10019) );
  INV_X1 U12403 ( .A(n13675), .ZN(n9981) );
  NAND2_X1 U12404 ( .A1(n12904), .A2(n12903), .ZN(n9691) );
  NOR2_X1 U12405 ( .A1(n14084), .A2(n14086), .ZN(n15339) );
  AND2_X1 U12406 ( .A1(n10241), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9692) );
  BUF_X1 U12407 ( .A(n12814), .Z(n12910) );
  INV_X1 U12408 ( .A(n13507), .ZN(n10113) );
  OR3_X1 U12409 ( .A1(n14908), .A2(n10130), .A3(n14873), .ZN(n9693) );
  NAND2_X1 U12410 ( .A1(n10179), .A2(n10177), .ZN(n14661) );
  OR2_X1 U12411 ( .A1(n17380), .A2(n18802), .ZN(n9695) );
  OR3_X1 U12412 ( .A1(n14831), .A2(n10083), .A3(n14819), .ZN(n9696) );
  NAND2_X1 U12413 ( .A1(n9641), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14990) );
  OR3_X1 U12414 ( .A1(n14460), .A2(n9996), .A3(n14439), .ZN(n9697) );
  AND2_X1 U12415 ( .A1(n15082), .A2(n9692), .ZN(n15046) );
  NAND2_X1 U12416 ( .A1(n14455), .A2(n10066), .ZN(n14442) );
  NOR2_X1 U12417 ( .A1(n12957), .A2(n15115), .ZN(n12958) );
  NOR2_X1 U12418 ( .A1(n12955), .A2(n16270), .ZN(n12956) );
  AND2_X1 U12419 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12959) );
  NOR2_X1 U12420 ( .A1(n14089), .A2(n16905), .ZN(n15484) );
  INV_X1 U12421 ( .A(n17812), .ZN(n10145) );
  AND2_X1 U12422 ( .A1(n9970), .A2(n9972), .ZN(n9698) );
  NAND2_X1 U12423 ( .A1(n10453), .A2(n10469), .ZN(n14013) );
  OR2_X1 U12424 ( .A1(n14084), .A2(n16905), .ZN(n9699) );
  NOR2_X1 U12425 ( .A1(n14034), .A2(n14035), .ZN(n14036) );
  NAND2_X1 U12426 ( .A1(n14455), .A2(n10064), .ZN(n9700) );
  NAND2_X1 U12427 ( .A1(n10218), .A2(n10219), .ZN(n14985) );
  XOR2_X1 U12428 ( .A(n15532), .B(n17371), .Z(n9701) );
  AND2_X1 U12429 ( .A1(n10262), .A2(n10880), .ZN(n9702) );
  NAND2_X1 U12430 ( .A1(n9947), .A2(n10961), .ZN(n16265) );
  AND2_X1 U12431 ( .A1(n10490), .A2(n14013), .ZN(n9703) );
  AND3_X1 U12432 ( .A1(n15187), .A2(n19224), .A3(n15186), .ZN(n9704) );
  AND2_X1 U12433 ( .A1(n13258), .A2(n11425), .ZN(n11501) );
  AND2_X1 U12434 ( .A1(n15067), .A2(n15025), .ZN(n9705) );
  NOR2_X1 U12435 ( .A1(n12955), .A2(n10158), .ZN(n12953) );
  OR2_X1 U12436 ( .A1(n14908), .A2(n10130), .ZN(n9706) );
  NOR3_X1 U12437 ( .A1(n17562), .A2(n17919), .A3(n17898), .ZN(n9707) );
  AND2_X1 U12438 ( .A1(n10819), .A2(n10035), .ZN(n9708) );
  NAND2_X1 U12439 ( .A1(n10373), .A2(n9666), .ZN(n10391) );
  AND2_X1 U12440 ( .A1(n10413), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9709) );
  NOR2_X1 U12441 ( .A1(n15009), .A2(n9974), .ZN(n14999) );
  AND2_X1 U12442 ( .A1(n11163), .A2(n10391), .ZN(n9710) );
  NOR2_X1 U12443 ( .A1(n10207), .A2(n10205), .ZN(n10204) );
  OR2_X1 U12444 ( .A1(n13857), .A2(n10957), .ZN(n9711) );
  NOR2_X1 U12445 ( .A1(n14034), .A2(n10058), .ZN(n14464) );
  NOR2_X1 U12446 ( .A1(n11686), .A2(n10195), .ZN(n10193) );
  AND2_X1 U12447 ( .A1(n15858), .A2(n20884), .ZN(n9712) );
  AND2_X1 U12448 ( .A1(n11089), .A2(n10232), .ZN(n9713) );
  NOR2_X1 U12449 ( .A1(n10477), .A2(n19068), .ZN(n9714) );
  AND3_X1 U12450 ( .A1(n10237), .A2(n10236), .A3(n10233), .ZN(n9715) );
  OR2_X1 U12451 ( .A1(n10699), .A2(n12816), .ZN(n9716) );
  AND2_X1 U12452 ( .A1(n11161), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12453 ( .A1(n14421), .A2(n10062), .ZN(n14304) );
  AND2_X1 U12454 ( .A1(n14973), .A2(n10901), .ZN(n9718) );
  OR2_X1 U12455 ( .A1(n19556), .A2(n10550), .ZN(n9719) );
  AND2_X1 U12456 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U12457 ( .A1(n15874), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9721) );
  OR2_X1 U12458 ( .A1(n10509), .A2(n10508), .ZN(n9722) );
  INV_X1 U12459 ( .A(n15009), .ZN(n9970) );
  INV_X1 U12460 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9846) );
  OAI211_X1 U12461 ( .C1(n9875), .C2(n9789), .A(n9999), .B(n10427), .ZN(n10428) );
  AOI21_X1 U12462 ( .B1(n10815), .B2(n9883), .A(n10002), .ZN(n14994) );
  NAND2_X1 U12463 ( .A1(n15082), .A2(n15202), .ZN(n15068) );
  INV_X1 U12464 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9847) );
  INV_X1 U12465 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10268) );
  AND2_X1 U12466 ( .A1(n9892), .A2(n9717), .ZN(n9724) );
  NAND2_X1 U12467 ( .A1(n9933), .A2(n10222), .ZN(n15270) );
  OR2_X1 U12468 ( .A1(n10774), .A2(n10773), .ZN(n9725) );
  NOR2_X1 U12469 ( .A1(n10029), .A2(n10028), .ZN(n10027) );
  NAND2_X1 U12470 ( .A1(n14606), .A2(n14729), .ZN(n9726) );
  AND2_X1 U12471 ( .A1(n12393), .A2(n14654), .ZN(n10206) );
  INV_X1 U12472 ( .A(n10206), .ZN(n10201) );
  INV_X1 U12473 ( .A(n11126), .ZN(n19245) );
  INV_X1 U12474 ( .A(n10393), .ZN(n11126) );
  AND2_X1 U12475 ( .A1(n10087), .A2(n10086), .ZN(n9727) );
  AND2_X1 U12476 ( .A1(n10144), .A2(n9806), .ZN(n9728) );
  AOI21_X1 U12477 ( .B1(n14890), .B2(n14891), .A(n12783), .ZN(n12802) );
  AND2_X1 U12478 ( .A1(n10719), .A2(n9854), .ZN(n9729) );
  AND2_X1 U12479 ( .A1(n9683), .A2(n12378), .ZN(n9730) );
  INV_X1 U12480 ( .A(n13788), .ZN(n9983) );
  NOR2_X1 U12481 ( .A1(n12952), .A2(n10163), .ZN(n12945) );
  INV_X1 U12482 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n12960) );
  AND2_X1 U12483 ( .A1(n11159), .A2(n10106), .ZN(n11169) );
  XNOR2_X1 U12484 ( .A(n11092), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9731) );
  AND2_X1 U12485 ( .A1(n14423), .A2(n9986), .ZN(n9732) );
  NOR2_X1 U12486 ( .A1(n12955), .A2(n10155), .ZN(n12951) );
  NOR2_X1 U12487 ( .A1(n12952), .A2(n12965), .ZN(n12948) );
  INV_X1 U12488 ( .A(n12573), .ZN(n10025) );
  NAND2_X1 U12489 ( .A1(n14231), .A2(n14228), .ZN(n9733) );
  NOR2_X1 U12490 ( .A1(n20185), .A2(n20184), .ZN(n9734) );
  INV_X1 U12491 ( .A(n9932), .ZN(n9931) );
  NAND2_X1 U12492 ( .A1(n10222), .A2(n9745), .ZN(n9932) );
  INV_X1 U12493 ( .A(n10801), .ZN(n11098) );
  AND2_X1 U12494 ( .A1(n11554), .A2(n11549), .ZN(n9735) );
  AND2_X1 U12495 ( .A1(n12945), .A2(n10971), .ZN(n12943) );
  AND2_X1 U12496 ( .A1(n12614), .A2(n12615), .ZN(n9736) );
  AND2_X1 U12497 ( .A1(n13671), .A2(n11773), .ZN(n13706) );
  INV_X1 U12498 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19058) );
  INV_X1 U12499 ( .A(n13278), .ZN(n13249) );
  INV_X1 U12500 ( .A(n10790), .ZN(n9867) );
  AND2_X1 U12501 ( .A1(n10243), .A2(n10242), .ZN(n15114) );
  AND2_X1 U12502 ( .A1(n12593), .A2(n19298), .ZN(n9737) );
  AND2_X1 U12503 ( .A1(n16271), .A2(n9688), .ZN(n9738) );
  AND2_X1 U12504 ( .A1(n10037), .A2(n10036), .ZN(n9739) );
  OR3_X1 U12505 ( .A1(n13777), .A2(n13778), .A3(n10082), .ZN(n9740) );
  OR2_X1 U12506 ( .A1(n13960), .A2(n10864), .ZN(n9741) );
  NAND2_X1 U12507 ( .A1(n17653), .A2(n17770), .ZN(n17570) );
  AND2_X1 U12508 ( .A1(n12943), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12942) );
  NOR2_X1 U12509 ( .A1(n12952), .A2(n10166), .ZN(n12949) );
  OR2_X1 U12510 ( .A1(n9665), .A2(n10820), .ZN(n9742) );
  AND2_X1 U12511 ( .A1(n10818), .A2(n9742), .ZN(n9743) );
  NAND2_X1 U12512 ( .A1(n10694), .A2(n9969), .ZN(n13732) );
  OR2_X1 U12513 ( .A1(n14831), .A2(n10083), .ZN(n9744) );
  OR2_X1 U12514 ( .A1(n15271), .A2(n15274), .ZN(n9745) );
  OR2_X1 U12515 ( .A1(n14460), .A2(n9996), .ZN(n9746) );
  OR2_X1 U12516 ( .A1(n10799), .A2(n13227), .ZN(n11100) );
  NAND2_X1 U12517 ( .A1(n13231), .A2(n13232), .ZN(n13230) );
  AND2_X1 U12518 ( .A1(n9907), .A2(n9908), .ZN(n9747) );
  OR2_X1 U12519 ( .A1(n17770), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9748) );
  AND2_X1 U12520 ( .A1(n11091), .A2(n11183), .ZN(n9749) );
  INV_X1 U12521 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15031) );
  INV_X1 U12522 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16245) );
  AND2_X1 U12523 ( .A1(n15271), .A2(n15274), .ZN(n9750) );
  AND2_X1 U12524 ( .A1(n12658), .A2(n9770), .ZN(n14834) );
  INV_X1 U12525 ( .A(n15030), .ZN(n9924) );
  OR2_X1 U12526 ( .A1(n16167), .A2(n10886), .ZN(n9751) );
  AND2_X1 U12527 ( .A1(n10018), .A2(n11098), .ZN(n9752) );
  OR2_X1 U12528 ( .A1(n13777), .A2(n10079), .ZN(n9753) );
  NOR2_X1 U12529 ( .A1(n13784), .A2(n10051), .ZN(n13970) );
  AND2_X1 U12530 ( .A1(n20093), .A2(n20079), .ZN(n16048) );
  INV_X1 U12531 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16270) );
  INV_X1 U12532 ( .A(n10016), .ZN(n10015) );
  NAND2_X1 U12533 ( .A1(n13726), .A2(n10017), .ZN(n10016) );
  INV_X1 U12534 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12965) );
  NAND2_X1 U12535 ( .A1(n14822), .A2(n10245), .ZN(n14890) );
  OR2_X1 U12536 ( .A1(n12288), .A2(n12286), .ZN(n9754) );
  AND2_X1 U12537 ( .A1(n9991), .A2(n14331), .ZN(n9755) );
  AND2_X1 U12538 ( .A1(n10653), .A2(n10737), .ZN(n9756) );
  AND2_X1 U12539 ( .A1(n10126), .A2(n10125), .ZN(n9757) );
  AND2_X1 U12540 ( .A1(n10161), .A2(n15045), .ZN(n9758) );
  AND2_X1 U12541 ( .A1(n9739), .A2(n10842), .ZN(n9759) );
  OR2_X1 U12542 ( .A1(n9920), .A2(n15030), .ZN(n9760) );
  AND2_X1 U12543 ( .A1(n9676), .A2(n11388), .ZN(n9761) );
  AND2_X1 U12544 ( .A1(n12062), .A2(n10064), .ZN(n9762) );
  INV_X1 U12545 ( .A(n10261), .ZN(n10010) );
  INV_X1 U12546 ( .A(n10524), .ZN(n13603) );
  NAND2_X1 U12547 ( .A1(n9975), .A2(n13775), .ZN(n9982) );
  AND2_X1 U12548 ( .A1(n10934), .A2(n11215), .ZN(n19222) );
  OR2_X1 U12549 ( .A1(n16353), .A2(n17864), .ZN(n9887) );
  NAND2_X1 U12550 ( .A1(n10357), .A2(n9892), .ZN(n11193) );
  NAND2_X1 U12551 ( .A1(n13306), .A2(n12614), .ZN(n13459) );
  NAND2_X1 U12552 ( .A1(n13306), .A2(n9736), .ZN(n13451) );
  OR2_X1 U12553 ( .A1(n13453), .A2(n13507), .ZN(n13508) );
  NOR2_X1 U12554 ( .A1(n13675), .A2(n12442), .ZN(n9763) );
  AND2_X1 U12555 ( .A1(n13469), .A2(n13468), .ZN(n13368) );
  NAND2_X1 U12556 ( .A1(n12940), .A2(n9689), .ZN(n12933) );
  INV_X1 U12557 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9829) );
  OR2_X1 U12558 ( .A1(n13569), .A2(n12435), .ZN(n13675) );
  NAND2_X1 U12559 ( .A1(n10694), .A2(n9968), .ZN(n13731) );
  INV_X1 U12560 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20644) );
  NAND2_X1 U12561 ( .A1(n13484), .A2(n10088), .ZN(n9764) );
  AND2_X1 U12562 ( .A1(n12657), .A2(n10108), .ZN(n9765) );
  NOR3_X1 U12563 ( .A1(n18992), .A2(n10801), .A3(n16252), .ZN(n9766) );
  OR2_X1 U12564 ( .A1(n13316), .A2(n15658), .ZN(n19920) );
  INV_X1 U12565 ( .A(n19920), .ZN(n20070) );
  BUF_X1 U12566 ( .A(n12947), .Z(n19029) );
  AND2_X1 U12567 ( .A1(n13752), .A2(n13751), .ZN(n13749) );
  INV_X1 U12568 ( .A(n16122), .ZN(n10171) );
  OR2_X1 U12569 ( .A1(n10682), .A2(n10681), .ZN(n11203) );
  AND2_X1 U12570 ( .A1(n10141), .A2(n10146), .ZN(n9767) );
  AND2_X1 U12571 ( .A1(n10115), .A2(n13738), .ZN(n9768) );
  INV_X1 U12572 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10148) );
  INV_X1 U12573 ( .A(n12592), .ZN(n10099) );
  AND2_X1 U12574 ( .A1(n12940), .A2(n10151), .ZN(n9769) );
  INV_X1 U12575 ( .A(n10118), .ZN(n13861) );
  AND2_X1 U12576 ( .A1(n9687), .A2(n10107), .ZN(n9770) );
  INV_X1 U12577 ( .A(n14825), .ZN(n10085) );
  INV_X1 U12578 ( .A(n16212), .ZN(n9943) );
  NOR2_X1 U12579 ( .A1(n11084), .A2(n12579), .ZN(n12577) );
  AND2_X1 U12580 ( .A1(n10378), .A2(n12828), .ZN(n9771) );
  OAI21_X1 U12581 ( .B1(n12872), .B2(n12871), .A(n12870), .ZN(n14797) );
  AND2_X1 U12582 ( .A1(n11855), .A2(n11854), .ZN(n9772) );
  OR2_X1 U12583 ( .A1(n12565), .A2(n10123), .ZN(n9773) );
  OR2_X1 U12584 ( .A1(n9691), .A2(n10096), .ZN(n9774) );
  AND2_X1 U12585 ( .A1(n14790), .A2(n10096), .ZN(n9775) );
  NAND2_X1 U12586 ( .A1(n15552), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9776) );
  AND2_X1 U12587 ( .A1(n14802), .A2(n12874), .ZN(n9777) );
  AND2_X1 U12588 ( .A1(n10134), .A2(n9695), .ZN(n9778) );
  AND2_X1 U12589 ( .A1(n9692), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9779) );
  INV_X1 U12590 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10152) );
  INV_X1 U12591 ( .A(n13656), .ZN(n10114) );
  AND2_X1 U12592 ( .A1(n20074), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n9780) );
  INV_X1 U12593 ( .A(n12923), .ZN(n10096) );
  AND2_X1 U12594 ( .A1(n11183), .A2(n12561), .ZN(n9781) );
  OR2_X1 U12595 ( .A1(n14594), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9782) );
  AND2_X1 U12596 ( .A1(n10240), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9783) );
  INV_X1 U12597 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10139) );
  INV_X1 U12598 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10140) );
  INV_X1 U12599 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9886) );
  INV_X1 U12600 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10040) );
  OR2_X1 U12601 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9784) );
  NOR3_X4 U12602 ( .A1(n18650), .A2(n18378), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18464) );
  AND2_X2 U12603 ( .A1(n9787), .A2(n9771), .ZN(n14812) );
  NOR2_X1 U12604 ( .A1(n14812), .A2(n9786), .ZN(n14872) );
  NOR2_X1 U12605 ( .A1(n9787), .A2(n9771), .ZN(n9786) );
  INV_X1 U12606 ( .A(n10259), .ZN(n9788) );
  AND2_X4 U12607 ( .A1(n13617), .A2(n13614), .ZN(n10510) );
  OAI21_X1 U12608 ( .B1(n14858), .B2(n14947), .A(n9791), .ZN(P2_U2890) );
  AND2_X1 U12609 ( .A1(n14857), .A2(n14856), .ZN(n9791) );
  XNOR2_X2 U12610 ( .A(n9965), .B(n10984), .ZN(n10490) );
  NAND2_X2 U12611 ( .A1(n9792), .A2(n10439), .ZN(n9965) );
  NAND2_X2 U12612 ( .A1(n10451), .A2(n10431), .ZN(n10459) );
  AND2_X2 U12613 ( .A1(n14834), .A2(n12712), .ZN(n14835) );
  NOR2_X4 U12614 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11426) );
  AND2_X4 U12615 ( .A1(n11426), .A2(n14751), .ZN(n11490) );
  AND2_X4 U12616 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14751) );
  OAI21_X1 U12617 ( .B1(n9793), .B2(n16073), .A(n9827), .ZN(P1_U3000) );
  INV_X1 U12618 ( .A(n9799), .ZN(n14607) );
  NAND3_X1 U12619 ( .A1(n20139), .A2(n9800), .A3(n12418), .ZN(n13091) );
  NAND2_X2 U12620 ( .A1(n11441), .A2(n10266), .ZN(n12418) );
  OR2_X2 U12621 ( .A1(n13991), .A2(n10175), .ZN(n10179) );
  INV_X2 U12622 ( .A(n11748), .ZN(n11750) );
  INV_X1 U12623 ( .A(n9804), .ZN(n17837) );
  OAI21_X1 U12624 ( .B1(n9805), .B2(n9701), .A(n9804), .ZN(n9803) );
  NAND3_X1 U12625 ( .A1(n9807), .A2(n10147), .A3(n9728), .ZN(n9810) );
  NAND2_X1 U12626 ( .A1(n9810), .A2(n10142), .ZN(n17801) );
  NAND3_X1 U12627 ( .A1(n9823), .A2(n9821), .A3(n9818), .ZN(n15576) );
  NOR2_X2 U12628 ( .A1(n17529), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17528) );
  OAI211_X2 U12629 ( .C1(n17546), .C2(n17898), .A(n9748), .B(n17545), .ZN(
        n17529) );
  NOR2_X2 U12630 ( .A1(n15555), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17514) );
  AND2_X2 U12631 ( .A1(n9826), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17706) );
  INV_X2 U12632 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18815) );
  INV_X4 U12633 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20913) );
  NAND2_X1 U12634 ( .A1(n9834), .A2(n12289), .ZN(n12290) );
  NAND2_X1 U12635 ( .A1(n9835), .A2(n9754), .ZN(n9834) );
  NAND2_X1 U12636 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  NAND2_X1 U12637 ( .A1(n12283), .A2(n12410), .ZN(n9836) );
  NAND2_X1 U12638 ( .A1(n9838), .A2(n12282), .ZN(n9837) );
  OAI21_X1 U12639 ( .B1(n12275), .B2(n9842), .A(n9841), .ZN(n9840) );
  INV_X1 U12640 ( .A(n14707), .ZN(n15935) );
  INV_X1 U12641 ( .A(n14709), .ZN(n15919) );
  INV_X1 U12642 ( .A(n14710), .ZN(n9843) );
  NAND2_X2 U12643 ( .A1(n9848), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15009) );
  NAND2_X1 U12644 ( .A1(n15082), .A2(n9779), .ZN(n15035) );
  NAND2_X1 U12645 ( .A1(n9729), .A2(n10718), .ZN(n9853) );
  INV_X1 U12646 ( .A(n10611), .ZN(n10230) );
  NAND2_X2 U12647 ( .A1(n10231), .A2(n9856), .ZN(n10945) );
  AND2_X1 U12648 ( .A1(n9861), .A2(n9859), .ZN(n16314) );
  NAND2_X1 U12649 ( .A1(n16251), .A2(n16252), .ZN(n9859) );
  NAND2_X1 U12650 ( .A1(n9861), .A2(n15274), .ZN(n9860) );
  NOR2_X1 U12651 ( .A1(n9725), .A2(n9870), .ZN(n11241) );
  NAND3_X1 U12652 ( .A1(n10777), .A2(n9872), .A3(n9871), .ZN(n9870) );
  NAND2_X1 U12653 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n9871) );
  NAND2_X1 U12654 ( .A1(n10000), .A2(n9875), .ZN(n10432) );
  NAND2_X1 U12655 ( .A1(n10408), .A2(n9875), .ZN(n10409) );
  AOI21_X1 U12656 ( .B1(n14968), .B2(n9882), .A(n9880), .ZN(n9879) );
  NAND3_X1 U12657 ( .A1(n10905), .A2(n15120), .A3(n9731), .ZN(n9881) );
  NAND2_X1 U12658 ( .A1(n14968), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15120) );
  INV_X1 U12659 ( .A(n10873), .ZN(n15017) );
  NAND3_X1 U12660 ( .A1(n16576), .A2(n16575), .A3(n9884), .ZN(P3_U2641) );
  NOR2_X2 U12661 ( .A1(n18648), .A2(n18148), .ZN(n18061) );
  NAND2_X1 U12662 ( .A1(n15082), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16251) );
  NAND3_X1 U12663 ( .A1(n9711), .A2(n10951), .A3(n10952), .ZN(n10243) );
  NAND3_X1 U12664 ( .A1(n13856), .A2(n10948), .A3(n10949), .ZN(n10954) );
  NOR2_X1 U12665 ( .A1(n11193), .A2(n11158), .ZN(n11185) );
  AND2_X2 U12666 ( .A1(n10401), .A2(n10380), .ZN(n11159) );
  NAND2_X1 U12667 ( .A1(n9899), .A2(n11686), .ZN(n9898) );
  NAND2_X1 U12668 ( .A1(n10197), .A2(n11603), .ZN(n9899) );
  INV_X1 U12669 ( .A(n10179), .ZN(n9903) );
  OAI21_X1 U12670 ( .B1(n9904), .B2(n9903), .A(n10204), .ZN(n14644) );
  NAND3_X1 U12671 ( .A1(n10177), .A2(n9905), .A3(n10201), .ZN(n9904) );
  NOR2_X2 U12672 ( .A1(n14662), .A2(n9906), .ZN(n9905) );
  NAND2_X1 U12673 ( .A1(n11750), .A2(n9907), .ZN(n11794) );
  NAND2_X2 U12674 ( .A1(n11750), .A2(n9747), .ZN(n12382) );
  NAND2_X2 U12675 ( .A1(n12382), .A2(n12381), .ZN(n12393) );
  AND3_X4 U12676 ( .A1(n10268), .A2(n9846), .A3(n9909), .ZN(n12911) );
  NAND3_X1 U12677 ( .A1(n9914), .A2(n9911), .A3(n9910), .ZN(n9923) );
  NAND2_X1 U12678 ( .A1(n15067), .A2(n9912), .ZN(n9911) );
  NAND3_X1 U12679 ( .A1(n9914), .A2(n9911), .A3(n9915), .ZN(n15200) );
  NAND2_X1 U12680 ( .A1(n9923), .A2(n9921), .ZN(P2_U2993) );
  OAI22_X1 U12681 ( .A1(n19301), .A2(n12863), .B1(n10702), .B2(n19656), .ZN(
        n10703) );
  NAND2_X1 U12682 ( .A1(n15104), .A2(n9929), .ZN(n9926) );
  INV_X1 U12683 ( .A(n10951), .ZN(n10953) );
  NAND2_X1 U12684 ( .A1(n10952), .A2(n10951), .ZN(n10955) );
  XNOR2_X2 U12685 ( .A(n10959), .B(n10957), .ZN(n10951) );
  NAND2_X2 U12686 ( .A1(n9945), .A2(n10966), .ZN(n15082) );
  OAI21_X1 U12687 ( .B1(n9950), .B2(n15102), .A(n9946), .ZN(n9945) );
  NOR2_X1 U12688 ( .A1(n9956), .A2(n10391), .ZN(n10918) );
  INV_X1 U12689 ( .A(n11194), .ZN(n10388) );
  INV_X1 U12690 ( .A(n10387), .ZN(n9953) );
  INV_X1 U12691 ( .A(n10391), .ZN(n9954) );
  NOR2_X1 U12692 ( .A1(n9666), .A2(n10373), .ZN(n9955) );
  NAND2_X1 U12693 ( .A1(n10385), .A2(n11139), .ZN(n9956) );
  NAND3_X1 U12694 ( .A1(n9963), .A2(n16224), .A3(n9962), .ZN(n9961) );
  AOI21_X1 U12695 ( .B1(n9965), .B2(n10988), .A(n10987), .ZN(n13311) );
  OAI21_X1 U12696 ( .B1(n14253), .B2(n19234), .A(n9966), .ZN(P2_U2984) );
  AND2_X1 U12697 ( .A1(n14239), .A2(n14238), .ZN(n9966) );
  XNOR2_X1 U12698 ( .A(n9967), .B(n13858), .ZN(n13899) );
  NAND2_X1 U12699 ( .A1(n10611), .A2(n10612), .ZN(n9969) );
  NOR2_X4 U12700 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14752) );
  NAND3_X1 U12701 ( .A1(n9977), .A2(n13775), .A3(n9983), .ZN(n9976) );
  NAND2_X1 U12702 ( .A1(n14345), .A2(n9755), .ZN(n14458) );
  NOR2_X2 U12703 ( .A1(n9646), .A2(n9666), .ZN(n10401) );
  AND2_X1 U12704 ( .A1(n10009), .A2(n10010), .ZN(n15012) );
  NAND2_X1 U12705 ( .A1(n13732), .A2(n10013), .ZN(n10012) );
  INV_X1 U12706 ( .A(n13888), .ZN(n10022) );
  NAND2_X1 U12707 ( .A1(n11090), .A2(n10027), .ZN(n10023) );
  NAND2_X1 U12708 ( .A1(n10023), .A2(n10024), .ZN(n14229) );
  NAND2_X1 U12709 ( .A1(n9646), .A2(n10637), .ZN(n10031) );
  NAND3_X1 U12710 ( .A1(n10646), .A2(n10684), .A3(n9756), .ZN(n10786) );
  NAND2_X1 U12711 ( .A1(n10819), .A2(n9743), .ZN(n10829) );
  NAND2_X1 U12712 ( .A1(n10819), .A2(n10818), .ZN(n10839) );
  NAND2_X1 U12713 ( .A1(n18982), .A2(n9759), .ZN(n10833) );
  NAND2_X1 U12714 ( .A1(n10902), .A2(n10044), .ZN(n11093) );
  NAND2_X1 U12715 ( .A1(n10902), .A2(n10043), .ZN(n11099) );
  NAND2_X1 U12716 ( .A1(n10902), .A2(n16126), .ZN(n16125) );
  OR3_X1 U12717 ( .A1(n10889), .A2(P2_EBX_REG_24__SCAN_IN), .A3(
        P2_EBX_REG_25__SCAN_IN), .ZN(n10895) );
  NOR2_X1 U12718 ( .A1(n10889), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10894) );
  NAND3_X1 U12719 ( .A1(n11680), .A2(n10048), .A3(n13361), .ZN(n13502) );
  INV_X1 U12720 ( .A(n13784), .ZN(n10049) );
  NAND2_X1 U12721 ( .A1(n10049), .A2(n10050), .ZN(n14024) );
  INV_X1 U12722 ( .A(n14024), .ZN(n11906) );
  NAND2_X1 U12723 ( .A1(n14269), .A2(n14271), .ZN(n14270) );
  NAND2_X1 U12724 ( .A1(n14269), .A2(n10067), .ZN(n10070) );
  NAND3_X1 U12725 ( .A1(n12556), .A2(n12555), .A3(n12557), .ZN(P2_U3015) );
  AOI21_X1 U12726 ( .B1(n12564), .B2(n10073), .A(n10072), .ZN(n10071) );
  NOR2_X1 U12727 ( .A1(n16172), .A2(n16329), .ZN(n12553) );
  NAND2_X1 U12728 ( .A1(n12564), .A2(n12563), .ZN(n12927) );
  INV_X1 U12729 ( .A(n11083), .ZN(n10078) );
  NAND3_X1 U12730 ( .A1(n14825), .A2(n10084), .A3(n14779), .ZN(n10083) );
  NAND2_X1 U12731 ( .A1(n13484), .A2(n9727), .ZN(n15257) );
  NAND2_X1 U12732 ( .A1(n14803), .A2(n9777), .ZN(n10091) );
  NAND2_X1 U12733 ( .A1(n14791), .A2(n9775), .ZN(n10092) );
  NAND2_X2 U12734 ( .A1(n10091), .A2(n10090), .ZN(n14791) );
  NAND3_X1 U12735 ( .A1(n10453), .A2(n10469), .A3(n10099), .ZN(n10098) );
  NOR2_X2 U12736 ( .A1(n13453), .A2(n10109), .ZN(n13752) );
  NAND2_X1 U12737 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  NAND2_X1 U12738 ( .A1(n9682), .A2(n10120), .ZN(n11243) );
  NAND2_X1 U12739 ( .A1(n14867), .A2(n11409), .ZN(n12566) );
  NAND2_X1 U12740 ( .A1(n16271), .A2(n9761), .ZN(n14951) );
  INV_X2 U12741 ( .A(n17156), .ZN(n15518) );
  NAND3_X1 U12742 ( .A1(n18815), .A2(n18649), .A3(n10133), .ZN(n17156) );
  AOI22_X1 U12743 ( .A1(n15486), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15487) );
  OR2_X1 U12744 ( .A1(n17859), .A2(n17866), .ZN(n10134) );
  INV_X1 U12745 ( .A(n10134), .ZN(n17858) );
  NAND2_X1 U12746 ( .A1(n15555), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17516) );
  NOR2_X1 U12747 ( .A1(n17528), .A2(n15554), .ZN(n15555) );
  AOI21_X2 U12748 ( .B1(n17570), .B2(n10136), .A(n9776), .ZN(n17546) );
  NOR2_X2 U12749 ( .A1(n17759), .A2(n10138), .ZN(n17710) );
  NAND3_X1 U12750 ( .A1(n17744), .A2(n10140), .A3(n10139), .ZN(n10138) );
  NAND3_X1 U12751 ( .A1(n15536), .A2(n17820), .A3(n10144), .ZN(n10141) );
  NAND2_X1 U12752 ( .A1(n12943), .A2(n9684), .ZN(n12939) );
  INV_X1 U12753 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10153) );
  AOI21_X1 U12754 ( .B1(n18906), .B2(n15045), .A(n19047), .ZN(n10162) );
  NAND2_X1 U12755 ( .A1(n10160), .A2(n10159), .ZN(n13024) );
  NAND2_X1 U12756 ( .A1(n18906), .A2(n9758), .ZN(n10160) );
  AOI21_X1 U12757 ( .B1(n16140), .B2(n10171), .A(n19047), .ZN(n14770) );
  NAND2_X1 U12758 ( .A1(n10169), .A2(n10167), .ZN(n14769) );
  NAND2_X1 U12759 ( .A1(n16140), .A2(n10170), .ZN(n10169) );
  INV_X1 U12760 ( .A(n10172), .ZN(n16121) );
  NAND2_X1 U12761 ( .A1(n15835), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14615) );
  NAND2_X1 U12762 ( .A1(n15897), .A2(n15898), .ZN(n10187) );
  NAND2_X1 U12763 ( .A1(n15897), .A2(n10183), .ZN(n10182) );
  NAND3_X1 U12764 ( .A1(n10189), .A2(n9730), .A3(n10190), .ZN(n12310) );
  NAND2_X1 U12765 ( .A1(n11688), .A2(n10191), .ZN(n10190) );
  INV_X1 U12766 ( .A(n11688), .ZN(n10188) );
  NAND3_X1 U12767 ( .A1(n10190), .A2(n9683), .A3(n10189), .ZN(n20184) );
  NAND2_X1 U12768 ( .A1(n11688), .A2(n20644), .ZN(n10197) );
  OAI21_X1 U12769 ( .B1(n14650), .B2(n10200), .A(n10198), .ZN(n14065) );
  NAND4_X1 U12770 ( .A1(n10314), .A2(n10313), .A3(n10315), .A4(n10312), .ZN(
        n10209) );
  NAND4_X1 U12771 ( .A1(n10311), .A2(n10308), .A3(n10309), .A4(n10310), .ZN(
        n10211) );
  NAND2_X1 U12772 ( .A1(n11103), .A2(n9733), .ZN(n10215) );
  INV_X1 U12773 ( .A(n11103), .ZN(n10216) );
  INV_X1 U12774 ( .A(n14995), .ZN(n10221) );
  AND2_X1 U12775 ( .A1(n10228), .A2(n10796), .ZN(n15096) );
  OR2_X2 U12776 ( .A1(n10471), .A2(n13613), .ZN(n19556) );
  NAND3_X1 U12777 ( .A1(n10233), .A2(n10234), .A3(n10237), .ZN(n10232) );
  NAND2_X1 U12778 ( .A1(n11072), .A2(n10238), .ZN(n10237) );
  NAND3_X1 U12779 ( .A1(n10243), .A2(n10242), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10956) );
  NAND3_X1 U12780 ( .A1(n10953), .A2(n9711), .A3(n10954), .ZN(n10242) );
  XNOR2_X1 U12781 ( .A(n11696), .B(n11697), .ZN(n12319) );
  NOR2_X2 U12782 ( .A1(n13245), .A2(n13584), .ZN(n13411) );
  NOR2_X2 U12783 ( .A1(n13244), .A2(n20107), .ZN(n11550) );
  INV_X1 U12784 ( .A(n14834), .ZN(n14919) );
  AND2_X1 U12785 ( .A1(n11069), .A2(n11068), .ZN(n11070) );
  OR2_X1 U12786 ( .A1(n11152), .A2(n16330), .ZN(n11415) );
  OR2_X1 U12787 ( .A1(n11152), .A2(n19234), .ZN(n11069) );
  INV_X1 U12788 ( .A(n20184), .ZN(n20109) );
  OR2_X1 U12789 ( .A1(n12594), .A2(n13235), .ZN(n19890) );
  OR2_X1 U12790 ( .A1(n12594), .A2(n12596), .ZN(n12597) );
  AND2_X1 U12791 ( .A1(n12829), .A2(n10259), .ZN(n10244) );
  NOR2_X1 U12792 ( .A1(n18700), .A2(n17829), .ZN(n17615) );
  INV_X1 U12793 ( .A(n11674), .ZN(n12240) );
  AND2_X1 U12794 ( .A1(n20008), .A2(n13580), .ZN(n20004) );
  NAND2_X1 U12795 ( .A1(n20008), .A2(n20147), .ZN(n14494) );
  INV_X1 U12796 ( .A(n16073), .ZN(n20090) );
  NOR2_X1 U12797 ( .A1(n20185), .A2(n20109), .ZN(n10246) );
  INV_X1 U12798 ( .A(n19759), .ZN(n12968) );
  NAND2_X2 U12799 ( .A1(n9648), .A2(n13582), .ZN(n14572) );
  AND4_X1 U12800 ( .A1(n15820), .A2(n15917), .A3(n15950), .A4(n14595), .ZN(
        n10247) );
  AND4_X1 U12801 ( .A1(n15474), .A2(n15473), .A3(n15472), .A4(n15471), .ZN(
        n10248) );
  OR2_X1 U12802 ( .A1(n14597), .A2(n10247), .ZN(n10249) );
  AND3_X1 U12803 ( .A1(n15477), .A2(n15476), .A3(n15475), .ZN(n10250) );
  AND4_X1 U12804 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10251) );
  AND2_X1 U12805 ( .A1(n15858), .A2(n15818), .ZN(n10253) );
  AND4_X1 U12806 ( .A1(n10602), .A2(n10601), .A3(n10600), .A4(n10599), .ZN(
        n10254) );
  AND2_X1 U12807 ( .A1(n17758), .A2(n17879), .ZN(n10255) );
  INV_X1 U12808 ( .A(n18849), .ZN(n18832) );
  OR2_X1 U12809 ( .A1(n10699), .A2(n10760), .ZN(n10256) );
  INV_X1 U12810 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13976) );
  AND2_X1 U12811 ( .A1(n20718), .A2(n12244), .ZN(n15894) );
  INV_X1 U12812 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15535) );
  AND4_X1 U12813 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10257) );
  OR2_X1 U12814 ( .A1(n13147), .A2(n13053), .ZN(n13108) );
  NAND2_X1 U12815 ( .A1(n9660), .A2(n10273), .ZN(n10258) );
  INV_X1 U12816 ( .A(n16352), .ZN(n16861) );
  AND2_X1 U12817 ( .A1(n12827), .A2(n12847), .ZN(n10259) );
  INV_X1 U12818 ( .A(n12987), .ZN(n10683) );
  INV_X1 U12819 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10662) );
  OR2_X1 U12820 ( .A1(n12584), .A2(n19236), .ZN(n10260) );
  NAND4_X1 U12821 ( .A1(n15029), .A2(n10872), .A3(n15025), .A4(n15026), .ZN(
        n10261) );
  AND4_X1 U12822 ( .A1(n15028), .A2(n15027), .A3(n15621), .A4(n10853), .ZN(
        n10262) );
  OR3_X1 U12823 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17592), .ZN(n10263) );
  INV_X1 U12824 ( .A(n11211), .ZN(n11293) );
  INV_X1 U12825 ( .A(n13460), .ZN(n12615) );
  INV_X1 U12826 ( .A(n13452), .ZN(n12616) );
  AND2_X1 U12827 ( .A1(n11198), .A2(n19903), .ZN(n16313) );
  INV_X1 U12828 ( .A(n11595), .ZN(n11580) );
  AND2_X1 U12829 ( .A1(n11556), .A2(n13580), .ZN(n10265) );
  AND4_X1 U12830 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n10266) );
  INV_X1 U12831 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11027) );
  AND2_X1 U12832 ( .A1(n12272), .A2(n12258), .ZN(n12278) );
  OR2_X1 U12833 ( .A1(n12272), .A2(n12271), .ZN(n12285) );
  AND2_X1 U12834 ( .A1(n19245), .A2(n10390), .ZN(n10356) );
  INV_X1 U12835 ( .A(n12285), .ZN(n12287) );
  NAND2_X1 U12836 ( .A1(n19886), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10632) );
  AOI22_X1 U12837 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10312) );
  OR3_X1 U12838 ( .A1(n12284), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20101), .ZN(n12286) );
  INV_X1 U12839 ( .A(n14436), .ZN(n12062) );
  OR2_X1 U12840 ( .A1(n11783), .A2(n11782), .ZN(n12368) );
  OR2_X1 U12841 ( .A1(n11760), .A2(n11759), .ZN(n12359) );
  OR2_X1 U12842 ( .A1(n11590), .A2(n11589), .ZN(n12320) );
  OR2_X1 U12843 ( .A1(n11667), .A2(n11666), .ZN(n11668) );
  OAI211_X1 U12844 ( .C1(n10386), .C2(n11123), .A(n10377), .B(n10376), .ZN(
        n10426) );
  AND4_X1 U12845 ( .A1(n10256), .A2(n10750), .A3(n10749), .A4(n10748), .ZN(
        n10759) );
  OR2_X1 U12846 ( .A1(n10457), .A2(n10455), .ZN(n10439) );
  AOI22_X1 U12847 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10358) );
  INV_X1 U12848 ( .A(n11543), .ZN(n11498) );
  OR2_X1 U12849 ( .A1(n12281), .A2(n11728), .ZN(n11741) );
  INV_X1 U12850 ( .A(n11668), .ZN(n12323) );
  INV_X1 U12851 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13257) );
  OR2_X1 U12852 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20101), .ZN(
        n12252) );
  XNOR2_X1 U12853 ( .A(n10273), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U12854 ( .A1(n10426), .A2(n10378), .ZN(n10379) );
  NAND2_X1 U12855 ( .A1(n10442), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10412) );
  INV_X1 U12856 ( .A(n12803), .ZN(n12804) );
  NOR2_X1 U12857 ( .A1(n10390), .A2(n10393), .ZN(n10380) );
  INV_X1 U12858 ( .A(n10464), .ZN(n10463) );
  NAND2_X1 U12859 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19896), .ZN(
        n10909) );
  INV_X1 U12861 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11988) );
  INV_X1 U12862 ( .A(n13971), .ZN(n11838) );
  INV_X1 U12863 ( .A(n12510), .ZN(n12471) );
  AND2_X1 U12864 ( .A1(n13422), .A2(n11548), .ZN(n12378) );
  INV_X1 U12865 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11418) );
  AND4_X1 U12866 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11470) );
  NAND2_X1 U12867 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12595) );
  NAND2_X1 U12868 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  AND2_X1 U12869 ( .A1(n12778), .A2(n14892), .ZN(n12799) );
  AND2_X1 U12870 ( .A1(n12754), .A2(n12759), .ZN(n12778) );
  AND2_X1 U12871 ( .A1(n11395), .A2(n11394), .ZN(n14909) );
  AND2_X1 U12872 ( .A1(n11144), .A2(n11143), .ZN(n11173) );
  AOI21_X1 U12873 ( .B1(n18651), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14182), .ZN(n14188) );
  NAND2_X1 U12874 ( .A1(n15550), .A2(n10263), .ZN(n15551) );
  AND2_X1 U12875 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15538), .ZN(
        n15539) );
  INV_X1 U12876 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20869) );
  AND4_X1 U12877 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n11441) );
  INV_X1 U12878 ( .A(n11820), .ZN(n11821) );
  INV_X1 U12879 ( .A(n12415), .ZN(n12416) );
  OR2_X1 U12880 ( .A1(n13575), .A2(n13574), .ZN(n13576) );
  AND2_X1 U12881 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12171), .ZN(
        n12172) );
  NAND2_X1 U12882 ( .A1(n14755), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12237) );
  NOR2_X1 U12883 ( .A1(n20780), .A2(n11896), .ZN(n11882) );
  AND2_X1 U12884 ( .A1(n12480), .A2(n12479), .ZN(n14331) );
  NAND2_X1 U12885 ( .A1(n12283), .A2(n12413), .ZN(n12293) );
  NAND2_X1 U12886 ( .A1(n11609), .A2(n11608), .ZN(n11686) );
  INV_X1 U12887 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20474) );
  INV_X1 U12888 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15115) );
  INV_X1 U12889 ( .A(n10446), .ZN(n10449) );
  AND2_X1 U12890 ( .A1(n12798), .A2(n12797), .ZN(n12800) );
  INV_X1 U12891 ( .A(n10973), .ZN(n12934) );
  INV_X1 U12892 ( .A(n12953), .ZN(n12963) );
  AND2_X1 U12893 ( .A1(n12549), .A2(n12562), .ZN(n14242) );
  NOR2_X1 U12894 ( .A1(n16319), .A2(n16320), .ZN(n15273) );
  AND2_X1 U12895 ( .A1(n11173), .A2(n11172), .ZN(n13553) );
  MUX2_X1 U12896 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11122), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11127) );
  NOR2_X1 U12897 ( .A1(n17508), .A2(n17509), .ZN(n16379) );
  OR2_X1 U12898 ( .A1(n15553), .A2(n10255), .ZN(n15554) );
  NAND2_X1 U12899 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  INV_X1 U12900 ( .A(n18665), .ZN(n18148) );
  AOI21_X1 U12901 ( .B1(n16516), .B2(n18203), .A(n18660), .ZN(n15697) );
  NAND2_X1 U12902 ( .A1(n16083), .A2(n20644), .ZN(n12305) );
  INV_X1 U12903 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20780) );
  NAND2_X1 U12904 ( .A1(n11821), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11839) );
  NAND2_X1 U12905 ( .A1(n11703), .A2(n11702), .ZN(n20247) );
  INV_X1 U12906 ( .A(n19997), .ZN(n19984) );
  AND3_X1 U12907 ( .A1(n11819), .A2(n11818), .A3(n11817), .ZN(n13838) );
  OAI21_X1 U12908 ( .B1(n20710), .B2(n11939), .A(n11727), .ZN(n13567) );
  NAND2_X1 U12909 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  INV_X1 U12910 ( .A(n14453), .ZN(n11993) );
  INV_X1 U12911 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14669) );
  INV_X1 U12912 ( .A(n11830), .ZN(n11939) );
  NOR2_X1 U12913 ( .A1(n11839), .A2(n13976), .ZN(n11856) );
  NAND2_X1 U12914 ( .A1(n11745), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11767) );
  AND3_X1 U12915 ( .A1(n13403), .A2(n13081), .A3(n12299), .ZN(n13277) );
  AND2_X1 U12916 ( .A1(n12502), .A2(n12501), .ZN(n14424) );
  AND2_X1 U12917 ( .A1(n12478), .A2(n12477), .ZN(n14468) );
  AND3_X1 U12918 ( .A1(n12462), .A2(n12461), .A3(n12460), .ZN(n14485) );
  OAI21_X1 U12919 ( .B1(n12314), .B2(n20124), .A(n12313), .ZN(n12316) );
  AND2_X1 U12920 ( .A1(n20159), .A2(n20158), .ZN(n20161) );
  INV_X1 U12921 ( .A(n20187), .ZN(n20416) );
  OR2_X1 U12922 ( .A1(n20710), .A2(n9672), .ZN(n20708) );
  INV_X1 U12923 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20504) );
  INV_X1 U12924 ( .A(n12294), .ZN(n15667) );
  AOI221_X1 U12925 ( .B1(n10916), .B2(n13168), .C1(n10916), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n10915), .ZN(n11124) );
  OAI22_X1 U12926 ( .A1(n12932), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12960), 
        .B2(n11073), .ZN(n12947) );
  NOR2_X1 U12927 ( .A1(n19047), .A2(n13024), .ZN(n15633) );
  AND2_X1 U12928 ( .A1(n11385), .A2(n11384), .ZN(n13950) );
  NAND2_X1 U12929 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13291) );
  NOR2_X1 U12930 ( .A1(n12852), .A2(n12851), .ZN(n14796) );
  AND2_X1 U12931 ( .A1(n11209), .A2(n11208), .ZN(n13802) );
  NAND2_X1 U12932 ( .A1(n13763), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11123) );
  INV_X1 U12933 ( .A(n10944), .ZN(n13797) );
  AND2_X1 U12934 ( .A1(n11150), .A2(n16343), .ZN(n11198) );
  OR2_X1 U12935 ( .A1(n19450), .A2(n19624), .ZN(n19389) );
  AND2_X1 U12936 ( .A1(n19442), .A2(n19441), .ZN(n19446) );
  OR2_X1 U12937 ( .A1(n19648), .A2(n19859), .ZN(n13909) );
  INV_X1 U12938 ( .A(n19864), .ZN(n19652) );
  INV_X1 U12939 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19693) );
  INV_X1 U12940 ( .A(n16522), .ZN(n18622) );
  OAI21_X1 U12941 ( .B1(n14192), .B2(n15566), .A(n14205), .ZN(n16522) );
  NOR2_X1 U12942 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16646), .ZN(n16633) );
  NOR2_X1 U12943 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16787), .ZN(n16770) );
  INV_X1 U12944 ( .A(n16900), .ZN(n16913) );
  AOI21_X1 U12945 ( .B1(n15417), .B2(n15416), .A(n18688), .ZN(n15694) );
  INV_X1 U12946 ( .A(n17370), .ZN(n17296) );
  NAND2_X1 U12947 ( .A1(n17544), .A2(n15611), .ZN(n17883) );
  NAND2_X1 U12948 ( .A1(n17648), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17628) );
  INV_X1 U12949 ( .A(n18009), .ZN(n17591) );
  INV_X1 U12950 ( .A(n18053), .ZN(n17732) );
  INV_X1 U12951 ( .A(n17860), .ZN(n17852) );
  NOR2_X1 U12952 ( .A1(n17883), .A2(n16371), .ZN(n16372) );
  NAND2_X1 U12953 ( .A1(n14179), .A2(n18624), .ZN(n15609) );
  NOR2_X1 U12954 ( .A1(n17758), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17643) );
  INV_X1 U12955 ( .A(n17932), .ZN(n18014) );
  NAND2_X1 U12956 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17769), .ZN(
        n18051) );
  NOR2_X1 U12957 ( .A1(n18105), .A2(n17798), .ZN(n17797) );
  INV_X1 U12958 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18651) );
  NOR2_X2 U12959 ( .A1(n14157), .A2(n14156), .ZN(n15559) );
  NOR2_X1 U12960 ( .A1(n18816), .A2(n18697), .ZN(n18194) );
  AND2_X2 U12961 ( .A1(n12418), .A2(n13422), .ZN(n14256) );
  OAI21_X1 U12962 ( .B1(n14711), .B2(n19985), .A(n12537), .ZN(n12538) );
  AND2_X1 U12963 ( .A1(n12533), .A2(n12531), .ZN(n15771) );
  AND2_X1 U12964 ( .A1(n15779), .A2(n12417), .ZN(n19958) );
  INV_X1 U12965 ( .A(n19963), .ZN(n19955) );
  AND2_X1 U12966 ( .A1(n12533), .A2(n12532), .ZN(n19997) );
  INV_X1 U12967 ( .A(n19913), .ZN(n13578) );
  NOR2_X2 U12968 ( .A1(n14217), .A2(n20102), .ZN(n14562) );
  INV_X1 U12969 ( .A(n13449), .ZN(n20048) );
  INV_X1 U12970 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U12971 ( .A1(n12110), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12149) );
  AND2_X1 U12972 ( .A1(n11856), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11857) );
  NOR2_X1 U12973 ( .A1(n11767), .A2(n19964), .ZN(n11786) );
  OR2_X1 U12974 ( .A1(n13391), .A2(n19913), .ZN(n13316) );
  NOR2_X1 U12975 ( .A1(n14713), .A2(n15970), .ZN(n15961) );
  OAI21_X1 U12976 ( .B1(n14058), .B2(n15938), .A(n20093), .ZN(n16036) );
  INV_X1 U12977 ( .A(n16048), .ZN(n16049) );
  AND2_X1 U12978 ( .A1(n13591), .A2(n16036), .ZN(n16070) );
  INV_X1 U12979 ( .A(n20093), .ZN(n20075) );
  INV_X1 U12980 ( .A(n20641), .ZN(n20150) );
  OAI21_X1 U12981 ( .B1(n20192), .B2(n20190), .A(n20189), .ZN(n20211) );
  INV_X1 U12982 ( .A(n20195), .ZN(n20208) );
  AND2_X1 U12983 ( .A1(n20214), .A2(n20444), .ZN(n20273) );
  AND2_X1 U12984 ( .A1(n20337), .A2(n9734), .ZN(n20325) );
  AND2_X1 U12985 ( .A1(n9672), .A2(n20250), .ZN(n20337) );
  INV_X1 U12986 ( .A(n20352), .ZN(n20382) );
  AND2_X1 U12987 ( .A1(n20185), .A2(n20184), .ZN(n20534) );
  OAI22_X1 U12988 ( .A1(n20483), .A2(n20482), .B1(n20532), .B2(n20481), .ZN(
        n20499) );
  AND2_X1 U12989 ( .A1(n20584), .A2(n10246), .ZN(n20527) );
  OAI211_X1 U12990 ( .C1(n20572), .C2(n20542), .A(n20541), .B(n20540), .ZN(
        n20574) );
  INV_X1 U12991 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20660) );
  INV_X1 U12992 ( .A(n20683), .ZN(n20933) );
  INV_X1 U12993 ( .A(n12564), .ZN(n11065) );
  INV_X1 U12994 ( .A(n19045), .ZN(n19059) );
  NAND2_X1 U12995 ( .A1(n16099), .A2(n12983), .ZN(n19055) );
  INV_X1 U12996 ( .A(n19057), .ZN(n19038) );
  INV_X1 U12997 ( .A(n14947), .ZN(n19139) );
  OAI21_X1 U12998 ( .B1(n13022), .B2(n13021), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13132) );
  INV_X1 U12999 ( .A(n12949), .ZN(n12950) );
  AND2_X1 U13000 ( .A1(n19229), .A2(n19231), .ZN(n19220) );
  CLKBUF_X1 U13001 ( .A(n13854), .Z(n13855) );
  NAND2_X1 U13002 ( .A1(n11174), .A2(n15238), .ZN(n15264) );
  NOR2_X2 U13003 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19864) );
  OAI21_X1 U13004 ( .B1(n13926), .B2(n13925), .A(n13924), .ZN(n19263) );
  NOR2_X1 U13005 ( .A1(n19502), .A2(n19450), .ZN(n19319) );
  NAND2_X1 U13006 ( .A1(n19113), .A2(n19890), .ZN(n19411) );
  INV_X1 U13007 ( .A(n19389), .ZN(n19437) );
  INV_X1 U13008 ( .A(n19500), .ZN(n19492) );
  INV_X1 U13009 ( .A(n19531), .ZN(n19520) );
  OAI21_X1 U13010 ( .B1(n13914), .B2(n13913), .A(n13912), .ZN(n19548) );
  INV_X1 U13011 ( .A(n13909), .ZN(n19579) );
  NOR2_X1 U13012 ( .A1(n19625), .A2(n19859), .ZN(n19614) );
  INV_X1 U13013 ( .A(n19725), .ZN(n19670) );
  OR2_X1 U13014 ( .A1(n19113), .A2(n19890), .ZN(n19625) );
  INV_X1 U13015 ( .A(n19277), .ZN(n19714) );
  AND2_X1 U13016 ( .A1(n12586), .A2(n19258), .ZN(n19738) );
  OR2_X1 U13017 ( .A1(n19113), .A2(n19142), .ZN(n19648) );
  INV_X1 U13018 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19765) );
  NAND2_X1 U13019 ( .A1(n18836), .A2(n18622), .ZN(n17427) );
  NOR2_X1 U13020 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16662), .ZN(n16654) );
  NOR2_X1 U13021 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16692), .ZN(n16673) );
  NOR2_X1 U13022 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16715), .ZN(n16699) );
  NOR2_X1 U13023 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16756), .ZN(n16749) );
  NOR2_X1 U13024 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16792), .ZN(n16791) );
  NOR2_X1 U13025 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16832), .ZN(n16812) );
  NOR2_X1 U13026 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16855), .ZN(n16838) );
  NAND3_X1 U13027 ( .A1(n15694), .A2(n18203), .A3(n18195), .ZN(n17232) );
  NAND2_X1 U13028 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17258), .ZN(n17257) );
  NOR3_X1 U13029 ( .A1(n17314), .A2(n17281), .A3(n17238), .ZN(n17278) );
  NAND2_X1 U13030 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17318), .ZN(n17314) );
  NOR2_X1 U13031 ( .A1(n17479), .A2(n17348), .ZN(n17347) );
  NOR2_X1 U13032 ( .A1(n17429), .A2(n17427), .ZN(n17430) );
  AND2_X1 U13033 ( .A1(n16399), .A2(n17842), .ZN(n16364) );
  NOR2_X1 U13034 ( .A1(n17919), .A2(n17910), .ZN(n17538) );
  NAND2_X1 U13035 ( .A1(n17732), .A2(n17975), .ZN(n17932) );
  INV_X1 U13036 ( .A(n17783), .ZN(n17752) );
  NOR2_X1 U13037 ( .A1(n18265), .A2(n18540), .ZN(n17611) );
  OAI21_X1 U13038 ( .B1(n18634), .B2(n15609), .A(n18633), .ZN(n17997) );
  INV_X1 U13039 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17718) );
  INV_X1 U13040 ( .A(n18098), .ZN(n18076) );
  NAND2_X1 U13041 ( .A1(n18094), .A2(n17770), .ZN(n17769) );
  INV_X1 U13042 ( .A(n18130), .ZN(n18169) );
  INV_X1 U13043 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18650) );
  NOR2_X1 U13044 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18791), .ZN(
        n18816) );
  INV_X1 U13045 ( .A(n18264), .ZN(n18327) );
  INV_X1 U13046 ( .A(n18491), .ZN(n18560) );
  NOR2_X1 U13047 ( .A1(n14208), .A2(n14207), .ZN(n18678) );
  INV_X1 U13048 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18788) );
  INV_X1 U13049 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n20897) );
  NOR2_X1 U13050 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13023), .ZN(n16496)
         );
  INV_X1 U13051 ( .A(U212), .ZN(n16469) );
  OR2_X1 U13052 ( .A1(n13316), .A2(n12407), .ZN(n13421) );
  INV_X1 U13053 ( .A(n12538), .ZN(n12539) );
  INV_X1 U13054 ( .A(n19977), .ZN(n19996) );
  INV_X1 U13055 ( .A(n19994), .ZN(n19985) );
  INV_X1 U13056 ( .A(n19958), .ZN(n19944) );
  AND2_X1 U13057 ( .A1(n19944), .A2(n14365), .ZN(n20002) );
  NAND2_X1 U13058 ( .A1(n20033), .A2(n20735), .ZN(n20010) );
  OAI211_X2 U13059 ( .C1(n13319), .C2(n13400), .A(n13318), .B(n13317), .ZN(
        n20033) );
  NOR2_X1 U13060 ( .A1(n13421), .A2(n13420), .ZN(n13448) );
  INV_X1 U13061 ( .A(n15871), .ZN(n15899) );
  INV_X1 U13062 ( .A(n15894), .ZN(n20104) );
  INV_X1 U13063 ( .A(n20089), .ZN(n16079) );
  NAND2_X1 U13064 ( .A1(n13414), .A2(n13399), .ZN(n16073) );
  INV_X1 U13065 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20722) );
  INV_X1 U13066 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16086) );
  NAND2_X1 U13067 ( .A1(n20214), .A2(n10246), .ZN(n20183) );
  NAND2_X1 U13068 ( .A1(n20214), .A2(n20534), .ZN(n20246) );
  NAND2_X1 U13069 ( .A1(n20337), .A2(n10246), .ZN(n20296) );
  INV_X1 U13070 ( .A(n20325), .ZN(n20324) );
  INV_X1 U13071 ( .A(n20349), .ZN(n20360) );
  NAND2_X1 U13072 ( .A1(n20445), .A2(n10246), .ZN(n20411) );
  NAND2_X1 U13073 ( .A1(n20445), .A2(n9734), .ZN(n20443) );
  NAND2_X1 U13074 ( .A1(n20445), .A2(n20534), .ZN(n20467) );
  NAND2_X1 U13075 ( .A1(n20445), .A2(n20444), .ZN(n20503) );
  NAND2_X1 U13076 ( .A1(n20584), .A2(n9734), .ZN(n20577) );
  NAND2_X1 U13077 ( .A1(n20584), .A2(n20444), .ZN(n20641) );
  INV_X1 U13078 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20479) );
  INV_X1 U13079 ( .A(n20707), .ZN(n20647) );
  INV_X1 U13080 ( .A(n13040), .ZN(n18862) );
  AND2_X1 U13081 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  NAND2_X1 U13082 ( .A1(n18862), .A2(n12971), .ZN(n18958) );
  NAND2_X1 U13083 ( .A1(n18862), .A2(n12988), .ZN(n19024) );
  INV_X1 U13084 ( .A(n18972), .ZN(n19065) );
  AND2_X1 U13085 ( .A1(n12930), .A2(n12929), .ZN(n12931) );
  NAND2_X1 U13086 ( .A1(n14844), .A2(n13931), .ZN(n16181) );
  NAND2_X1 U13087 ( .A1(n19111), .A2(n11137), .ZN(n14947) );
  AND2_X1 U13088 ( .A1(n13225), .A2(n16343), .ZN(n19111) );
  NOR2_X1 U13089 ( .A1(n19139), .A2(n19138), .ZN(n19123) );
  INV_X1 U13090 ( .A(n19096), .ZN(n19145) );
  NAND2_X1 U13091 ( .A1(n19184), .A2(n19152), .ZN(n19182) );
  INV_X1 U13092 ( .A(n19184), .ZN(n19217) );
  OR2_X1 U13093 ( .A1(n13052), .A2(n11215), .ZN(n19147) );
  INV_X1 U13094 ( .A(n19220), .ZN(n16256) );
  INV_X1 U13095 ( .A(n19222), .ZN(n19236) );
  INV_X1 U13096 ( .A(n16334), .ZN(n16317) );
  INV_X1 U13097 ( .A(n16313), .ZN(n16330) );
  INV_X1 U13098 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15693) );
  AOI21_X1 U13099 ( .B1(n13921), .B2(n13925), .A(n13920), .ZN(n19266) );
  INV_X1 U13100 ( .A(n19319), .ZN(n19327) );
  OR2_X1 U13101 ( .A1(n19411), .A2(n19859), .ZN(n19351) );
  INV_X1 U13102 ( .A(n19364), .ZN(n19388) );
  AOI21_X1 U13103 ( .B1(n13761), .B2(n19362), .A(n13760), .ZN(n19410) );
  INV_X1 U13104 ( .A(n19415), .ZN(n19469) );
  OR2_X1 U13105 ( .A1(n19450), .A2(n19698), .ZN(n19500) );
  OR2_X1 U13106 ( .A1(n19625), .A2(n19502), .ZN(n19523) );
  OR2_X1 U13107 ( .A1(n19648), .A2(n19502), .ZN(n19531) );
  AOI21_X1 U13108 ( .B1(n13907), .B2(n13913), .A(n13906), .ZN(n19552) );
  INV_X1 U13109 ( .A(n19614), .ZN(n19583) );
  INV_X1 U13110 ( .A(n19734), .ZN(n19609) );
  INV_X1 U13111 ( .A(n19644), .ZN(n19638) );
  OR2_X1 U13112 ( .A1(n19625), .A2(n19624), .ZN(n19681) );
  OR2_X1 U13113 ( .A1(n19648), .A2(n19698), .ZN(n19753) );
  INV_X1 U13114 ( .A(n19845), .ZN(n19763) );
  INV_X1 U13115 ( .A(n16886), .ZN(n16920) );
  INV_X1 U13116 ( .A(n16897), .ZN(n16919) );
  AND2_X1 U13117 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17108), .ZN(n17123) );
  NOR2_X1 U13118 ( .A1(n17450), .A2(n17271), .ZN(n17270) );
  NOR2_X1 U13119 ( .A1(n18234), .A2(n15699), .ZN(n17356) );
  NOR2_X1 U13120 ( .A1(n15460), .A2(n15459), .ZN(n17363) );
  INV_X1 U13121 ( .A(n17374), .ZN(n17388) );
  INV_X1 U13122 ( .A(n17406), .ZN(n17426) );
  AOI21_X1 U13123 ( .B1(n16398), .B2(n17752), .A(n16364), .ZN(n16365) );
  NAND2_X1 U13124 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17865), .ZN(n17672) );
  INV_X1 U13125 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17716) );
  NAND2_X1 U13126 ( .A1(n17354), .A2(n17861), .ZN(n17783) );
  INV_X1 U13127 ( .A(n18093), .ZN(n17974) );
  NAND3_X1 U13128 ( .A1(n17354), .A2(n18627), .A3(n18175), .ZN(n18098) );
  INV_X1 U13129 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18192) );
  INV_X1 U13130 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18191) );
  NAND2_X1 U13131 ( .A1(n18692), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18688) );
  INV_X1 U13132 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18791) );
  INV_X1 U13133 ( .A(n18787), .ZN(n18701) );
  INV_X1 U13134 ( .A(n18777), .ZN(n18849) );
  INV_X1 U13135 ( .A(n16473), .ZN(n16472) );
  INV_X1 U13136 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13940) );
  NOR2_X2 U13137 ( .A1(n10268), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10512) );
  AOI22_X1 U13138 ( .A1(n12814), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13139 ( .A1(n9668), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13140 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13141 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10269) );
  NAND4_X1 U13142 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10274) );
  INV_X2 U13143 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U13144 ( .A1(n10274), .A2(n10273), .ZN(n10281) );
  AOI22_X1 U13145 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13146 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13147 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13148 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10275) );
  NAND4_X1 U13149 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10279) );
  NAND2_X1 U13150 ( .A1(n10279), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10280) );
  AOI22_X1 U13151 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10285) );
  INV_X1 U13152 ( .A(n10300), .ZN(n10316) );
  AOI22_X1 U13153 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13154 ( .A1(n9668), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13155 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10282) );
  NAND4_X1 U13156 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  NAND2_X1 U13157 ( .A1(n10286), .A2(n10273), .ZN(n10293) );
  AOI22_X1 U13158 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13159 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13160 ( .A1(n12814), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13161 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10287) );
  NAND4_X1 U13162 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10291) );
  NAND2_X1 U13163 ( .A1(n10291), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10292) );
  INV_X2 U13164 ( .A(n10294), .ZN(n10378) );
  AOI22_X1 U13165 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13166 ( .A1(n9668), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13167 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13168 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10295) );
  NAND4_X1 U13169 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10299) );
  AOI22_X1 U13170 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13171 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10303) );
  INV_X1 U13172 ( .A(n10300), .ZN(n12740) );
  AOI22_X1 U13173 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10302) );
  NAND4_X1 U13174 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NAND2_X1 U13175 ( .A1(n10305), .A2(n10273), .ZN(n10306) );
  NAND2_X1 U13176 ( .A1(n9670), .A2(n9667), .ZN(n11199) );
  AOI22_X1 U13177 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13178 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13179 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13180 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13181 ( .A1(n9668), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13182 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U13183 ( .A1(n11199), .A2(n12586), .ZN(n10329) );
  AOI22_X1 U13184 ( .A1(n12814), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13185 ( .A1(n9668), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13186 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13187 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10317) );
  NAND4_X1 U13188 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10321) );
  NAND2_X1 U13189 ( .A1(n10321), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10328) );
  AOI22_X1 U13190 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13191 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13192 ( .A1(n9669), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13193 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13194 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  NAND2_X1 U13195 ( .A1(n10326), .A2(n10273), .ZN(n10327) );
  NAND2_X1 U13196 ( .A1(n10328), .A2(n10327), .ZN(n10370) );
  AOI22_X1 U13197 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13198 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9668), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13199 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10331) );
  NAND4_X1 U13200 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10334) );
  AOI22_X1 U13201 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13202 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U13203 ( .A1(n10336), .A2(n10335), .ZN(n10340) );
  AOI22_X1 U13204 ( .A1(n9668), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13205 ( .A1(n9669), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U13206 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  AOI22_X1 U13207 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13208 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13209 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13210 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10343) );
  NAND4_X1 U13211 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10347) );
  AOI22_X1 U13212 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13213 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13214 ( .A1(n12739), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10348) );
  NAND3_X1 U13215 ( .A1(n10350), .A2(n10349), .A3(n10348), .ZN(n10353) );
  AOI22_X1 U13216 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10351) );
  NAND2_X2 U13218 ( .A1(n10355), .A2(n10354), .ZN(n10390) );
  AOI22_X1 U13219 ( .A1(n9669), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13220 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13221 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10359) );
  NAND4_X1 U13222 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  NAND2_X1 U13223 ( .A1(n10362), .A2(n10273), .ZN(n10369) );
  AOI22_X1 U13224 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12814), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13225 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13226 ( .A1(n9669), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13227 ( .A1(n10510), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13228 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10367) );
  INV_X1 U13229 ( .A(n10370), .ZN(n10395) );
  AND2_X2 U13230 ( .A1(n10390), .A2(n10370), .ZN(n11139) );
  INV_X1 U13231 ( .A(n11106), .ZN(n10372) );
  AND2_X1 U13232 ( .A1(n10390), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U13233 ( .A1(n11161), .A2(n10372), .A3(n10401), .A4(n10371), .ZN(
        n10377) );
  AND4_X1 U13234 ( .A1(n11126), .A2(n10395), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n13941), .ZN(n10375) );
  NAND4_X1 U13235 ( .A1(n10375), .A2(n9954), .A3(n10374), .A4(n13931), .ZN(
        n10376) );
  NAND2_X1 U13236 ( .A1(n9674), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10384) );
  INV_X2 U13237 ( .A(n11028), .ZN(n10443) );
  NAND2_X1 U13238 ( .A1(n12960), .A2(n11027), .ZN(n10424) );
  NAND2_X1 U13239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10381) );
  NAND2_X1 U13240 ( .A1(n10424), .A2(n10381), .ZN(n10382) );
  AOI21_X1 U13241 ( .B1(n10443), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10382), .ZN(
        n10383) );
  NAND2_X1 U13242 ( .A1(n10384), .A2(n10383), .ZN(n10410) );
  NAND2_X1 U13243 ( .A1(n11163), .A2(n10294), .ZN(n10387) );
  NAND2_X1 U13244 ( .A1(n10388), .A2(n13763), .ZN(n10399) );
  NOR2_X1 U13245 ( .A1(n11137), .A2(n10294), .ZN(n10389) );
  NAND2_X1 U13246 ( .A1(n10407), .A2(n10374), .ZN(n10398) );
  NAND4_X1 U13247 ( .A1(n11126), .A2(n10395), .A3(n10390), .A4(n13941), .ZN(
        n10392) );
  NOR2_X1 U13248 ( .A1(n11135), .A2(n13763), .ZN(n10397) );
  OAI211_X1 U13249 ( .C1(n11137), .C2(n10395), .A(n10394), .B(n9710), .ZN(
        n10396) );
  NAND2_X1 U13250 ( .A1(n10397), .A2(n10396), .ZN(n11157) );
  NAND3_X1 U13251 ( .A1(n10399), .A2(n10398), .A3(n11157), .ZN(n10400) );
  INV_X1 U13252 ( .A(n10401), .ZN(n10402) );
  NAND3_X1 U13253 ( .A1(n10031), .A2(n10402), .A3(n11126), .ZN(n10404) );
  NAND2_X1 U13254 ( .A1(n10404), .A2(n10403), .ZN(n11134) );
  NOR2_X1 U13255 ( .A1(n10405), .A2(n13936), .ZN(n10406) );
  AOI21_X2 U13256 ( .B1(n11134), .B2(n11139), .A(n10406), .ZN(n11156) );
  NAND3_X1 U13257 ( .A1(n11156), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10407), 
        .ZN(n10408) );
  NOR2_X1 U13258 ( .A1(n10410), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U13259 ( .A1(n10412), .A2(n10411), .ZN(n10446) );
  AND2_X1 U13260 ( .A1(n10413), .A2(n11161), .ZN(n10414) );
  OAI22_X1 U13261 ( .A1(n10432), .A2(n10414), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11051), .ZN(n10418) );
  INV_X1 U13262 ( .A(n10424), .ZN(n13039) );
  NAND2_X1 U13263 ( .A1(n13039), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10415) );
  AND2_X1 U13264 ( .A1(n10416), .A2(n10415), .ZN(n10417) );
  NAND2_X1 U13265 ( .A1(n10418), .A2(n10417), .ZN(n10447) );
  NAND2_X1 U13266 ( .A1(n10446), .A2(n10447), .ZN(n10450) );
  NAND2_X1 U13267 ( .A1(n9673), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10422) );
  INV_X1 U13268 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10419) );
  OAI22_X1 U13269 ( .A1(n11028), .A2(n10419), .B1(n11027), .B2(n19058), .ZN(
        n10420) );
  INV_X1 U13270 ( .A(n10420), .ZN(n10421) );
  NOR2_X1 U13271 ( .A1(n10424), .A2(n19886), .ZN(n10425) );
  NOR2_X1 U13272 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  XNOR2_X1 U13273 ( .A(n10429), .B(n10428), .ZN(n10452) );
  NAND2_X1 U13274 ( .A1(n10450), .A2(n10452), .ZN(n10451) );
  INV_X1 U13275 ( .A(n10428), .ZN(n10430) );
  NAND2_X1 U13276 ( .A1(n10430), .A2(n10429), .ZN(n10431) );
  NAND2_X1 U13277 ( .A1(n10432), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10434) );
  AOI21_X1 U13278 ( .B1(n12960), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U13279 ( .A1(n10442), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10437) );
  AOI22_X1 U13280 ( .A1(n10443), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10436) );
  NAND2_X1 U13281 ( .A1(n11051), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10435) );
  NAND3_X1 U13282 ( .A1(n10437), .A2(n10436), .A3(n10435), .ZN(n10455) );
  NAND2_X1 U13283 ( .A1(n10457), .A2(n10455), .ZN(n10438) );
  NAND2_X1 U13284 ( .A1(n10432), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10441) );
  NAND2_X1 U13285 ( .A1(n13039), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10440) );
  INV_X1 U13286 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10638) );
  NAND2_X1 U13287 ( .A1(n10442), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10445) );
  AOI22_X1 U13288 ( .A1(n10993), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10444) );
  INV_X1 U13289 ( .A(n10447), .ZN(n10448) );
  INV_X1 U13290 ( .A(n19068), .ZN(n10454) );
  INV_X1 U13291 ( .A(n10455), .ZN(n10456) );
  XNOR2_X1 U13292 ( .A(n10457), .B(n10456), .ZN(n10458) );
  INV_X1 U13293 ( .A(n14013), .ZN(n10461) );
  NAND2_X1 U13294 ( .A1(n9714), .A2(n13613), .ZN(n10696) );
  INV_X1 U13295 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10522) );
  OAI22_X1 U13296 ( .A1(n13940), .A2(n10695), .B1(n10696), .B2(n10522), .ZN(
        n10462) );
  INV_X1 U13297 ( .A(n10462), .ZN(n10486) );
  INV_X1 U13298 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12808) );
  INV_X1 U13299 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U13300 ( .A1(n13827), .A2(n19068), .ZN(n10464) );
  INV_X1 U13301 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10465) );
  OAI22_X1 U13302 ( .A1(n10466), .A2(n19413), .B1(n19656), .B2(n10465), .ZN(
        n10467) );
  INV_X1 U13303 ( .A(n10467), .ZN(n10483) );
  INV_X1 U13304 ( .A(n10468), .ZN(n10470) );
  OR2_X2 U13305 ( .A1(n10471), .A2(n10500), .ZN(n19691) );
  INV_X1 U13306 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10473) );
  INV_X1 U13307 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10472) );
  OAI22_X1 U13308 ( .A1(n19691), .A2(n10473), .B1(n19556), .B2(n10472), .ZN(
        n10474) );
  INV_X1 U13309 ( .A(n10474), .ZN(n10482) );
  INV_X1 U13310 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10479) );
  INV_X1 U13311 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10478) );
  OAI22_X1 U13312 ( .A1(n10479), .A2(n19301), .B1(n10541), .B2(n10478), .ZN(
        n10480) );
  INV_X1 U13313 ( .A(n10480), .ZN(n10481) );
  INV_X1 U13314 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U13315 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n9716), .ZN(
        n10532) );
  INV_X1 U13316 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10489) );
  NOR2_X1 U13317 ( .A1(n14013), .A2(n10452), .ZN(n10491) );
  NAND2_X1 U13318 ( .A1(n13728), .A2(n10491), .ZN(n10487) );
  OR2_X2 U13319 ( .A1(n10487), .A2(n13613), .ZN(n10707) );
  INV_X1 U13320 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10488) );
  OAI22_X1 U13321 ( .A1(n10489), .A2(n10707), .B1(n10708), .B2(n10488), .ZN(
        n10509) );
  INV_X1 U13322 ( .A(n10491), .ZN(n10498) );
  NAND2_X1 U13323 ( .A1(n10490), .A2(n10492), .ZN(n13766) );
  INV_X1 U13324 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10496) );
  INV_X1 U13325 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10495) );
  AND2_X1 U13326 ( .A1(n10500), .A2(n10493), .ZN(n10494) );
  OAI22_X1 U13327 ( .A1(n13766), .A2(n10496), .B1(n10495), .B2(n19330), .ZN(
        n10497) );
  INV_X1 U13328 ( .A(n10497), .ZN(n10507) );
  INV_X1 U13329 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10504) );
  INV_X1 U13330 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10503) );
  OAI22_X1 U13331 ( .A1(n10711), .A2(n10504), .B1(n10503), .B2(n19442), .ZN(
        n10505) );
  INV_X1 U13332 ( .A(n10505), .ZN(n10506) );
  NAND2_X1 U13333 ( .A1(n10507), .A2(n10506), .ZN(n10508) );
  NAND2_X1 U13334 ( .A1(n12910), .A2(n10273), .ZN(n12714) );
  INV_X1 U13335 ( .A(n10510), .ZN(n12733) );
  AND2_X2 U13336 ( .A1(n10511), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12705) );
  AOI22_X1 U13337 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12697), .B1(
        n12705), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10517) );
  AND2_X2 U13338 ( .A1(n12915), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10676) );
  AND2_X1 U13339 ( .A1(n12911), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10582) );
  AOI22_X1 U13340 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10516) );
  NOR2_X1 U13341 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13342 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12719), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10515) );
  AND2_X2 U13343 ( .A1(n12915), .A2(n10273), .ZN(n12690) );
  NAND2_X1 U13344 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10514) );
  NAND4_X1 U13345 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10530) );
  AOI22_X1 U13346 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12683), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10528) );
  AND2_X2 U13347 ( .A1(n10518), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10768) );
  INV_X1 U13348 ( .A(n10768), .ZN(n10619) );
  AND2_X1 U13349 ( .A1(n12734), .A2(n10519), .ZN(n10581) );
  NAND2_X1 U13350 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10521) );
  AND2_X1 U13351 ( .A1(n13617), .A2(n12734), .ZN(n10613) );
  NAND2_X1 U13352 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10520) );
  OAI211_X1 U13353 ( .C1(n10619), .C2(n10522), .A(n10521), .B(n10520), .ZN(
        n10523) );
  INV_X1 U13354 ( .A(n10523), .ZN(n10527) );
  AND2_X1 U13355 ( .A1(n9661), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10667) );
  AOI22_X1 U13356 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10526) );
  AND2_X2 U13357 ( .A1(n9663), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10762) );
  AOI22_X1 U13358 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10525) );
  NAND4_X1 U13359 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n10525), .ZN(
        n10529) );
  INV_X1 U13360 ( .A(n10636), .ZN(n11235) );
  NAND2_X1 U13361 ( .A1(n11235), .A2(n10378), .ZN(n10531) );
  INV_X1 U13362 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10534) );
  INV_X1 U13363 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10533) );
  OAI22_X1 U13364 ( .A1(n10534), .A2(n19301), .B1(n19656), .B2(n10533), .ZN(
        n10538) );
  INV_X1 U13365 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10536) );
  INV_X1 U13366 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10535) );
  OAI22_X1 U13367 ( .A1(n10536), .A2(n19413), .B1(n19691), .B2(n10535), .ZN(
        n10537) );
  INV_X1 U13368 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10539) );
  INV_X1 U13369 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13930) );
  NOR2_X1 U13370 ( .A1(n10267), .A2(n10540), .ZN(n10560) );
  INV_X1 U13371 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12630) );
  AOI21_X1 U13372 ( .B1(n19333), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n10378), .ZN(n10544) );
  INV_X1 U13373 ( .A(n13766), .ZN(n10542) );
  NAND2_X1 U13374 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10543) );
  OAI211_X1 U13375 ( .C1(n10541), .C2(n12630), .A(n10544), .B(n10543), .ZN(
        n10555) );
  INV_X1 U13376 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10571) );
  NOR2_X1 U13377 ( .A1(n19442), .A2(n10571), .ZN(n10547) );
  INV_X1 U13378 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10545) );
  NOR2_X1 U13379 ( .A1(n10711), .A2(n10545), .ZN(n10546) );
  NOR2_X1 U13380 ( .A1(n10547), .A2(n10546), .ZN(n10553) );
  INV_X1 U13381 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10548) );
  INV_X1 U13382 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10549) );
  INV_X1 U13383 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10550) );
  NAND4_X1 U13384 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n9719), .ZN(
        n10554) );
  NOR2_X1 U13385 ( .A1(n10555), .A2(n10554), .ZN(n10559) );
  INV_X1 U13386 ( .A(n10696), .ZN(n10557) );
  INV_X1 U13387 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12770) );
  INV_X1 U13388 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12763) );
  AOI21_X1 U13389 ( .B1(n10557), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n10556), .ZN(n10558) );
  NAND3_X1 U13390 ( .A1(n10560), .A2(n10559), .A3(n10558), .ZN(n10610) );
  AOI22_X1 U13391 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13392 ( .A1(n12724), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13393 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13394 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U13395 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10570) );
  AOI22_X1 U13396 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13397 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13398 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13399 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10565) );
  NAND4_X1 U13400 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10569) );
  NOR2_X1 U13401 ( .A1(n10570), .A2(n10569), .ZN(n11210) );
  INV_X1 U13402 ( .A(n13170), .ZN(n10591) );
  OR2_X1 U13403 ( .A1(n12714), .A2(n10571), .ZN(n10575) );
  NAND2_X1 U13404 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10574) );
  NAND2_X1 U13405 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10573) );
  NAND2_X1 U13406 ( .A1(n10763), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10572) );
  AND4_X1 U13407 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(
        n10590) );
  AOI22_X1 U13408 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12719), .B1(
        n10613), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10579) );
  INV_X2 U13409 ( .A(n10258), .ZN(n12683) );
  NAND2_X1 U13410 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10578) );
  NAND2_X1 U13411 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13412 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10576) );
  AND4_X1 U13413 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10589) );
  AOI22_X1 U13414 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13415 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13416 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10585) );
  NAND2_X1 U13417 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10584) );
  NAND2_X1 U13418 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10583) );
  AND4_X1 U13419 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10587) );
  NAND4_X1 U13420 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n11220) );
  NAND2_X1 U13421 ( .A1(n10591), .A2(n11220), .ZN(n10935) );
  AOI22_X1 U13422 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13423 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10594) );
  NAND2_X1 U13424 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10593) );
  NAND2_X1 U13425 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10592) );
  NAND4_X1 U13426 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10598) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10596) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12791) );
  OAI22_X1 U13429 ( .A1(n12714), .A2(n10596), .B1(n13559), .B2(n12791), .ZN(
        n10597) );
  NOR2_X1 U13430 ( .A1(n10598), .A2(n10597), .ZN(n10608) );
  AOI22_X1 U13431 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12719), .B1(
        n10613), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13432 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10601) );
  NAND2_X1 U13433 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U13434 ( .A1(n10763), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U13435 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10606) );
  NAND2_X1 U13436 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10605) );
  NAND2_X1 U13437 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10604) );
  NAND2_X1 U13438 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10603) );
  AND4_X1 U13439 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10607) );
  NAND2_X1 U13440 ( .A1(n10935), .A2(n11228), .ZN(n10609) );
  AOI22_X1 U13441 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10613), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13442 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10616) );
  NAND2_X1 U13443 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10615) );
  NAND2_X1 U13444 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10614) );
  INV_X1 U13445 ( .A(n12700), .ZN(n10621) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10620) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10618) );
  OAI22_X1 U13448 ( .A1(n10621), .A2(n10620), .B1(n10619), .B2(n10618), .ZN(
        n10623) );
  INV_X1 U13449 ( .A(n10667), .ZN(n10761) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12918) );
  INV_X1 U13451 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11369) );
  OAI22_X1 U13452 ( .A1(n10761), .A2(n12918), .B1(n13559), .B2(n11369), .ZN(
        n10622) );
  NOR2_X1 U13453 ( .A1(n10623), .A2(n10622), .ZN(n10629) );
  AOI22_X1 U13454 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13455 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10627) );
  NAND2_X1 U13456 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10626) );
  NAND2_X1 U13457 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13458 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10624) );
  NAND4_X1 U13459 ( .A1(n10630), .A2(n10629), .A3(n10628), .A4(n10251), .ZN(
        n10787) );
  INV_X1 U13460 ( .A(n10787), .ZN(n10801) );
  NAND2_X1 U13461 ( .A1(n9789), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10631) );
  NAND2_X1 U13462 ( .A1(n10632), .A2(n10631), .ZN(n11108) );
  MUX2_X1 U13463 ( .A(n12599), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n13614), .Z(n10639) );
  INV_X1 U13464 ( .A(n10639), .ZN(n10633) );
  NAND2_X1 U13465 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12599), .ZN(
        n10635) );
  XNOR2_X1 U13466 ( .A(n10663), .B(n10664), .ZN(n10921) );
  MUX2_X1 U13467 ( .A(n10636), .B(n10921), .S(n12987), .Z(n10910) );
  MUX2_X1 U13468 ( .A(n10910), .B(n10638), .S(n13227), .Z(n10646) );
  NAND2_X1 U13469 ( .A1(n10640), .A2(n10639), .ZN(n10642) );
  NAND2_X1 U13470 ( .A1(n12987), .A2(n11107), .ZN(n11105) );
  OAI21_X1 U13471 ( .B1(n12987), .B2(n11228), .A(n11105), .ZN(n10911) );
  INV_X1 U13472 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13295) );
  MUX2_X1 U13473 ( .A(n10911), .B(n13295), .S(n13227), .Z(n10654) );
  INV_X1 U13474 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13475 ( .A1(n13227), .A2(n10643), .ZN(n10647) );
  NAND2_X1 U13476 ( .A1(n11220), .A2(n9666), .ZN(n10644) );
  NAND2_X1 U13477 ( .A1(n10647), .A2(n10644), .ZN(n10645) );
  NAND2_X1 U13478 ( .A1(n13227), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10650) );
  OAI21_X1 U13479 ( .B1(n10646), .B2(n10653), .A(n10685), .ZN(n13888) );
  OAI21_X1 U13480 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19896), .A(
        n10909), .ZN(n11109) );
  MUX2_X1 U13481 ( .A(n11210), .B(n11109), .S(n12987), .Z(n10649) );
  INV_X1 U13482 ( .A(n10647), .ZN(n10648) );
  AOI21_X1 U13483 ( .B1(n10649), .B2(n9665), .A(n10648), .ZN(n14017) );
  NAND2_X1 U13484 ( .A1(n14017), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13171) );
  NOR2_X1 U13485 ( .A1(n10650), .A2(n10643), .ZN(n10651) );
  OR2_X1 U13486 ( .A1(n10655), .A2(n10651), .ZN(n19056) );
  NOR2_X1 U13487 ( .A1(n13171), .A2(n19056), .ZN(n10652) );
  NAND2_X1 U13488 ( .A1(n13171), .A2(n19056), .ZN(n13104) );
  OAI21_X1 U13489 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10652), .A(
        n13104), .ZN(n13191) );
  INV_X1 U13490 ( .A(n10653), .ZN(n10659) );
  INV_X1 U13491 ( .A(n10654), .ZN(n10657) );
  INV_X1 U13492 ( .A(n10655), .ZN(n10656) );
  NAND2_X1 U13493 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  NAND2_X1 U13494 ( .A1(n10659), .A2(n10658), .ZN(n10660) );
  INV_X1 U13495 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13197) );
  XNOR2_X1 U13496 ( .A(n10660), .B(n13197), .ZN(n13190) );
  OR2_X1 U13497 ( .A1(n13191), .A2(n13190), .ZN(n13218) );
  INV_X1 U13498 ( .A(n10660), .ZN(n13822) );
  NAND2_X1 U13499 ( .A1(n13822), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10661) );
  AND2_X1 U13500 ( .A1(n13218), .A2(n10661), .ZN(n13726) );
  INV_X1 U13501 ( .A(n13794), .ZN(n10690) );
  NAND3_X1 U13502 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10916), .A3(
        n13168), .ZN(n10922) );
  AOI22_X1 U13503 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10762), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10675) );
  INV_X1 U13504 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U13505 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10669) );
  NAND2_X1 U13506 ( .A1(n12719), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10668) );
  OAI211_X1 U13507 ( .C1(n10258), .C2(n10670), .A(n10669), .B(n10668), .ZN(
        n10671) );
  INV_X1 U13508 ( .A(n10671), .ZN(n10674) );
  AOI22_X1 U13509 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10673) );
  INV_X1 U13510 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19249) );
  AOI22_X1 U13511 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10672) );
  NAND4_X1 U13512 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(
        n10682) );
  AOI22_X1 U13513 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13514 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13515 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13516 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10677) );
  NAND4_X1 U13517 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  MUX2_X1 U13518 ( .A(n10922), .B(n11203), .S(n10683), .Z(n10908) );
  INV_X1 U13519 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13313) );
  MUX2_X1 U13520 ( .A(n10908), .B(n13313), .S(n13227), .Z(n10684) );
  INV_X1 U13521 ( .A(n10738), .ZN(n10688) );
  NAND2_X1 U13522 ( .A1(n10686), .A2(n10685), .ZN(n10687) );
  NAND2_X1 U13523 ( .A1(n10688), .A2(n10687), .ZN(n13815) );
  INV_X1 U13524 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13860) );
  XNOR2_X1 U13525 ( .A(n13815), .B(n13860), .ZN(n13793) );
  INV_X1 U13526 ( .A(n13793), .ZN(n10689) );
  NAND2_X1 U13527 ( .A1(n10690), .A2(n10689), .ZN(n10693) );
  INV_X1 U13528 ( .A(n13815), .ZN(n10691) );
  NAND2_X1 U13529 ( .A1(n10691), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10692) );
  NAND2_X1 U13530 ( .A1(n10693), .A2(n10692), .ZN(n13853) );
  INV_X1 U13531 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19257) );
  INV_X1 U13532 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10697) );
  OAI22_X1 U13533 ( .A1(n19257), .A2(n10695), .B1(n10696), .B2(n10697), .ZN(
        n10698) );
  INV_X1 U13534 ( .A(n10698), .ZN(n10719) );
  INV_X1 U13535 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10724) );
  NOR2_X1 U13536 ( .A1(n10699), .A2(n10724), .ZN(n10706) );
  INV_X1 U13537 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10701) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10700) );
  OAI22_X1 U13539 ( .A1(n10701), .A2(n19413), .B1(n10541), .B2(n10700), .ZN(
        n10705) );
  INV_X1 U13540 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10725) );
  INV_X1 U13541 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12857) );
  OAI22_X1 U13542 ( .A1(n10725), .A2(n19556), .B1(n19691), .B2(n12857), .ZN(
        n10704) );
  INV_X1 U13543 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12863) );
  INV_X1 U13544 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10702) );
  NOR4_X1 U13545 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10718) );
  INV_X1 U13546 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10710) );
  INV_X1 U13547 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10709) );
  OAI22_X1 U13548 ( .A1(n10710), .A2(n10707), .B1(n10708), .B2(n10709), .ZN(
        n10715) );
  INV_X1 U13549 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12859) );
  INV_X1 U13550 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12864) );
  OAI22_X1 U13551 ( .A1(n12859), .A2(n10711), .B1(n19442), .B2(n12864), .ZN(
        n10713) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12862) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12865) );
  OAI22_X1 U13554 ( .A1(n12862), .A2(n13766), .B1(n19330), .B2(n12865), .ZN(
        n10712) );
  OR2_X1 U13555 ( .A1(n10713), .A2(n10712), .ZN(n10714) );
  NOR2_X1 U13556 ( .A1(n10715), .A2(n10714), .ZN(n10717) );
  INV_X1 U13557 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U13558 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U13559 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U13560 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U13561 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10720) );
  NAND4_X1 U13562 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10727) );
  INV_X1 U13563 ( .A(n12705), .ZN(n10775) );
  OAI22_X1 U13564 ( .A1(n10775), .A2(n10725), .B1(n13559), .B2(n10724), .ZN(
        n10726) );
  NOR2_X1 U13565 ( .A1(n10727), .A2(n10726), .ZN(n10734) );
  AOI22_X1 U13566 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U13567 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U13568 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10729) );
  NAND2_X1 U13569 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10728) );
  AOI22_X1 U13570 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13571 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10732) );
  NAND4_X1 U13572 ( .A1(n10734), .A2(n10257), .A3(n10733), .A4(n10732), .ZN(
        n10736) );
  INV_X1 U13573 ( .A(n10736), .ZN(n11238) );
  NAND2_X1 U13574 ( .A1(n11238), .A2(n10378), .ZN(n10735) );
  INV_X1 U13575 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19041) );
  MUX2_X1 U13576 ( .A(n19041), .B(n10736), .S(n9665), .Z(n10737) );
  OAI21_X1 U13577 ( .B1(n10738), .B2(n10737), .A(n10786), .ZN(n19037) );
  INV_X1 U13578 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13579 ( .A1(n10740), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10741) );
  INV_X1 U13580 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10760) );
  INV_X1 U13581 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10743) );
  INV_X1 U13582 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12890) );
  OAI22_X1 U13583 ( .A1(n10743), .A2(n19413), .B1(n19656), .B2(n12890), .ZN(
        n10744) );
  INV_X1 U13584 ( .A(n10744), .ZN(n10750) );
  INV_X1 U13585 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12893) );
  INV_X1 U13586 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10745) );
  OAI22_X1 U13587 ( .A1(n12893), .A2(n10707), .B1(n19691), .B2(n10745), .ZN(
        n10746) );
  INV_X1 U13588 ( .A(n10746), .ZN(n10749) );
  INV_X1 U13589 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12878) );
  INV_X1 U13590 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12896) );
  OAI22_X1 U13591 ( .A1(n12878), .A2(n19301), .B1(n10541), .B2(n12896), .ZN(
        n10747) );
  INV_X1 U13592 ( .A(n10747), .ZN(n10748) );
  INV_X1 U13593 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13474) );
  INV_X1 U13594 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12891) );
  OAI22_X1 U13595 ( .A1(n13474), .A2(n10695), .B1(n10696), .B2(n12891), .ZN(
        n10751) );
  INV_X1 U13596 ( .A(n10751), .ZN(n10758) );
  INV_X1 U13597 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12875) );
  NOR2_X1 U13598 ( .A1(n19361), .A2(n12875), .ZN(n10756) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12877) );
  INV_X1 U13600 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12879) );
  OAI22_X1 U13601 ( .A1(n12877), .A2(n19330), .B1(n19442), .B2(n12879), .ZN(
        n10755) );
  INV_X1 U13602 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12876) );
  INV_X1 U13603 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12880) );
  OAI22_X1 U13604 ( .A1(n12876), .A2(n10711), .B1(n13766), .B2(n12880), .ZN(
        n10754) );
  INV_X1 U13605 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12895) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10752) );
  OAI22_X1 U13607 ( .A1(n12895), .A2(n19556), .B1(n10708), .B2(n10752), .ZN(
        n10753) );
  NOR4_X1 U13608 ( .A1(n10756), .A2(n10755), .A3(n10754), .A4(n10753), .ZN(
        n10757) );
  NAND3_X1 U13609 ( .A1(n10759), .A2(n10758), .A3(n10757), .ZN(n10781) );
  OAI22_X1 U13610 ( .A1(n10761), .A2(n12890), .B1(n13559), .B2(n10760), .ZN(
        n10767) );
  INV_X1 U13611 ( .A(n10762), .ZN(n10765) );
  INV_X1 U13612 ( .A(n10763), .ZN(n10764) );
  OAI22_X1 U13613 ( .A1(n10765), .A2(n12896), .B1(n10764), .B2(n13474), .ZN(
        n10766) );
  OR2_X1 U13614 ( .A1(n10767), .A2(n10766), .ZN(n10774) );
  NAND2_X1 U13615 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10772) );
  NAND2_X1 U13616 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10771) );
  AOI22_X1 U13617 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U13618 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10769) );
  NAND4_X1 U13619 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10773) );
  OAI22_X1 U13620 ( .A1(n10775), .A2(n12895), .B1(n12714), .B2(n12879), .ZN(
        n10779) );
  AOI22_X1 U13621 ( .A1(n12719), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U13622 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10777) );
  NAND2_X1 U13623 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10776) );
  NAND2_X1 U13624 ( .A1(n10378), .A2(n11241), .ZN(n10780) );
  NAND2_X1 U13625 ( .A1(n10951), .A2(n10801), .ZN(n10782) );
  MUX2_X1 U13626 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11241), .S(n9666), .Z(n10785) );
  XNOR2_X1 U13627 ( .A(n10786), .B(n10785), .ZN(n19025) );
  INV_X1 U13628 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15313) );
  NAND2_X1 U13629 ( .A1(n10783), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10784) );
  INV_X1 U13630 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13482) );
  MUX2_X1 U13631 ( .A(n13482), .B(n10787), .S(n9666), .Z(n10790) );
  INV_X1 U13632 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10998) );
  AND2_X1 U13633 ( .A1(n10799), .A2(n10788), .ZN(n10789) );
  OR2_X1 U13634 ( .A1(n10798), .A2(n10789), .ZN(n13881) );
  NOR2_X1 U13635 ( .A1(n13881), .A2(n10801), .ZN(n10793) );
  NAND2_X1 U13636 ( .A1(n10793), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16259) );
  XNOR2_X1 U13637 ( .A(n10791), .B(n9867), .ZN(n19013) );
  NAND2_X1 U13638 ( .A1(n19013), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16260) );
  NAND2_X1 U13639 ( .A1(n16259), .A2(n16260), .ZN(n10792) );
  INV_X1 U13640 ( .A(n10793), .ZN(n10794) );
  INV_X1 U13641 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U13642 ( .A1(n10794), .A2(n10962), .ZN(n16258) );
  INV_X1 U13643 ( .A(n19013), .ZN(n10795) );
  INV_X1 U13644 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16322) );
  NAND2_X1 U13645 ( .A1(n10795), .A2(n16322), .ZN(n16262) );
  AND2_X1 U13646 ( .A1(n16258), .A2(n16262), .ZN(n10796) );
  INV_X1 U13647 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13466) );
  NOR2_X1 U13648 ( .A1(n9666), .A2(n13466), .ZN(n10797) );
  XNOR2_X1 U13649 ( .A(n10798), .B(n10797), .ZN(n19002) );
  NAND2_X1 U13650 ( .A1(n19002), .A2(n11098), .ZN(n10803) );
  INV_X1 U13651 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15292) );
  NAND2_X1 U13652 ( .A1(n10803), .A2(n15292), .ZN(n15095) );
  NAND3_X1 U13653 ( .A1(n10804), .A2(n13227), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n10800) );
  OAI211_X1 U13654 ( .C1(n10804), .C2(P2_EBX_REG_10__SCAN_IN), .A(n11100), .B(
        n10800), .ZN(n18992) );
  OR2_X1 U13655 ( .A1(n18992), .A2(n10801), .ZN(n10802) );
  AND2_X1 U13656 ( .A1(n10802), .A2(n16252), .ZN(n16248) );
  INV_X1 U13657 ( .A(n10809), .ZN(n10805) );
  NAND2_X2 U13658 ( .A1(n11100), .A2(n10805), .ZN(n18982) );
  AND2_X1 U13659 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10806), .ZN(n10807) );
  NAND2_X1 U13660 ( .A1(n13227), .A2(n10807), .ZN(n18980) );
  NAND2_X1 U13661 ( .A1(n18980), .A2(n11098), .ZN(n10808) );
  OR2_X1 U13662 ( .A1(n18982), .A2(n10808), .ZN(n15271) );
  INV_X1 U13663 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15274) );
  NAND2_X1 U13664 ( .A1(n13227), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10810) );
  OR2_X1 U13665 ( .A1(n10809), .A2(n10810), .ZN(n10811) );
  NAND2_X1 U13666 ( .A1(n10811), .A2(n10850), .ZN(n18970) );
  NOR2_X1 U13667 ( .A1(n18970), .A2(n10801), .ZN(n10812) );
  NAND2_X1 U13668 ( .A1(n10812), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16233) );
  INV_X1 U13669 ( .A(n10812), .ZN(n10814) );
  INV_X1 U13670 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U13671 ( .A1(n10814), .A2(n10813), .ZN(n16232) );
  INV_X1 U13672 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10816) );
  NOR2_X1 U13673 ( .A1(n9665), .A2(n10816), .ZN(n10849) );
  INV_X1 U13674 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11020) );
  NOR2_X1 U13675 ( .A1(n9666), .A2(n11020), .ZN(n10844) );
  NAND2_X1 U13676 ( .A1(n13227), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10842) );
  INV_X1 U13677 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10817) );
  NOR2_X1 U13678 ( .A1(n9666), .A2(n10817), .ZN(n10837) );
  INV_X1 U13679 ( .A(n10837), .ZN(n10818) );
  NOR2_X1 U13680 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10820) );
  INV_X1 U13681 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10821) );
  NAND2_X1 U13682 ( .A1(n13227), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10822) );
  NOR2_X1 U13683 ( .A1(n9708), .A2(n10822), .ZN(n10823) );
  NOR2_X1 U13684 ( .A1(n10874), .A2(n10823), .ZN(n13025) );
  NAND2_X1 U13685 ( .A1(n13025), .A2(n11098), .ZN(n10854) );
  INV_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15196) );
  NAND2_X1 U13687 ( .A1(n10854), .A2(n15196), .ZN(n15028) );
  NAND2_X1 U13688 ( .A1(n13227), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10824) );
  MUX2_X1 U13689 ( .A(n13227), .B(n10824), .S(n10839), .Z(n10825) );
  OR2_X1 U13690 ( .A1(n10839), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13691 ( .A1(n18917), .A2(n11098), .ZN(n10866) );
  INV_X1 U13692 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15203) );
  NAND2_X1 U13693 ( .A1(n10866), .A2(n15203), .ZN(n15064) );
  NAND3_X1 U13694 ( .A1(n10826), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n13227), 
        .ZN(n10827) );
  AND2_X1 U13695 ( .A1(n10827), .A2(n10829), .ZN(n18897) );
  NAND2_X1 U13696 ( .A1(n18897), .A2(n11098), .ZN(n10868) );
  INV_X1 U13697 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15220) );
  NAND2_X1 U13698 ( .A1(n10868), .A2(n15220), .ZN(n15050) );
  NAND2_X1 U13699 ( .A1(n15064), .A2(n15050), .ZN(n15038) );
  NAND2_X1 U13700 ( .A1(n13227), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10828) );
  XNOR2_X1 U13701 ( .A(n10829), .B(n10828), .ZN(n18885) );
  NAND2_X1 U13702 ( .A1(n18885), .A2(n11098), .ZN(n10870) );
  INV_X1 U13703 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15204) );
  AND2_X1 U13704 ( .A1(n10870), .A2(n15204), .ZN(n15039) );
  NOR2_X1 U13705 ( .A1(n15038), .A2(n15039), .ZN(n15027) );
  INV_X1 U13706 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10830) );
  NOR2_X1 U13707 ( .A1(n9665), .A2(n10830), .ZN(n10832) );
  INV_X1 U13708 ( .A(n11100), .ZN(n10831) );
  AOI21_X1 U13709 ( .B1(n10833), .B2(n10832), .A(n10831), .ZN(n10835) );
  AND2_X1 U13710 ( .A1(n10835), .A2(n10834), .ZN(n10863) );
  NAND2_X1 U13711 ( .A1(n10863), .A2(n11098), .ZN(n10836) );
  XNOR2_X1 U13712 ( .A(n10836), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15621) );
  NAND2_X1 U13713 ( .A1(n10838), .A2(n10837), .ZN(n10840) );
  NAND2_X1 U13714 ( .A1(n10840), .A2(n10839), .ZN(n18927) );
  INV_X1 U13715 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10841) );
  OAI21_X1 U13716 ( .B1(n18927), .B2(n10801), .A(n10841), .ZN(n15021) );
  INV_X1 U13717 ( .A(n10842), .ZN(n10843) );
  XNOR2_X1 U13718 ( .A(n10845), .B(n10843), .ZN(n18947) );
  AOI21_X1 U13719 ( .B1(n18947), .B2(n11098), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15020) );
  INV_X1 U13720 ( .A(n15020), .ZN(n15086) );
  AND2_X1 U13721 ( .A1(n10852), .A2(n10844), .ZN(n10846) );
  OR2_X1 U13722 ( .A1(n10846), .A2(n10845), .ZN(n13969) );
  NOR2_X1 U13723 ( .A1(n13969), .A2(n10801), .ZN(n10858) );
  INV_X1 U13724 ( .A(n10858), .ZN(n10848) );
  INV_X1 U13725 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13726 ( .A1(n10848), .A2(n10847), .ZN(n16210) );
  NAND2_X1 U13727 ( .A1(n10850), .A2(n10849), .ZN(n10851) );
  NAND2_X1 U13728 ( .A1(n10852), .A2(n10851), .ZN(n10859) );
  OAI21_X1 U13729 ( .B1(n10859), .B2(n10801), .A(n15261), .ZN(n15019) );
  AND4_X1 U13730 ( .A1(n15021), .A2(n15086), .A3(n16210), .A4(n15019), .ZN(
        n10853) );
  INV_X1 U13731 ( .A(n10854), .ZN(n10855) );
  NAND2_X1 U13732 ( .A1(n10855), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15029) );
  INV_X1 U13733 ( .A(n18927), .ZN(n10857) );
  AND2_X1 U13734 ( .A1(n11098), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10856) );
  NAND2_X1 U13735 ( .A1(n10857), .A2(n10856), .ZN(n15022) );
  AND2_X1 U13736 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16212) );
  INV_X1 U13737 ( .A(n10859), .ZN(n18960) );
  AND2_X1 U13738 ( .A1(n11098), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10860) );
  NAND2_X1 U13739 ( .A1(n18960), .A2(n10860), .ZN(n15018) );
  INV_X1 U13740 ( .A(n15018), .ZN(n10861) );
  NOR2_X1 U13741 ( .A1(n16212), .A2(n10861), .ZN(n10865) );
  AND2_X1 U13742 ( .A1(n11098), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10862) );
  NAND2_X1 U13743 ( .A1(n18947), .A2(n10862), .ZN(n15085) );
  INV_X1 U13744 ( .A(n10863), .ZN(n13960) );
  NAND2_X1 U13745 ( .A1(n11098), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10864) );
  AND4_X1 U13746 ( .A1(n15022), .A2(n10865), .A3(n15085), .A4(n9741), .ZN(
        n10872) );
  INV_X1 U13747 ( .A(n10866), .ZN(n10867) );
  NAND2_X1 U13748 ( .A1(n10867), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15065) );
  INV_X1 U13749 ( .A(n10868), .ZN(n10869) );
  NAND2_X1 U13750 ( .A1(n10869), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15051) );
  AND2_X1 U13751 ( .A1(n15065), .A2(n15051), .ZN(n15025) );
  INV_X1 U13752 ( .A(n10870), .ZN(n10871) );
  NAND2_X1 U13753 ( .A1(n10871), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15026) );
  NAND2_X1 U13754 ( .A1(n13227), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10875) );
  INV_X1 U13755 ( .A(n10875), .ZN(n10876) );
  NAND2_X1 U13756 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  NAND2_X1 U13757 ( .A1(n10883), .A2(n10878), .ZN(n15636) );
  XNOR2_X1 U13758 ( .A(n10879), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15011) );
  INV_X1 U13759 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15179) );
  NAND2_X1 U13760 ( .A1(n10879), .A2(n15179), .ZN(n10880) );
  INV_X1 U13761 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10881) );
  NOR2_X1 U13762 ( .A1(n9666), .A2(n10881), .ZN(n10882) );
  NAND2_X1 U13763 ( .A1(n10883), .A2(n10882), .ZN(n10884) );
  NAND2_X1 U13764 ( .A1(n10889), .A2(n10884), .ZN(n16167) );
  OR2_X1 U13765 ( .A1(n16167), .A2(n10801), .ZN(n10885) );
  XNOR2_X1 U13766 ( .A(n10885), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15002) );
  NAND2_X1 U13767 ( .A1(n11098), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10886) );
  INV_X1 U13768 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15154) );
  NAND2_X1 U13769 ( .A1(n13227), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10887) );
  MUX2_X1 U13770 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10887), .S(n10889), .Z(
        n10888) );
  NAND2_X1 U13771 ( .A1(n10888), .A2(n11100), .ZN(n14781) );
  NOR2_X1 U13772 ( .A1(n14781), .A2(n10801), .ZN(n14995) );
  INV_X1 U13773 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10893) );
  NOR2_X1 U13774 ( .A1(n10894), .A2(n10893), .ZN(n10890) );
  NAND2_X1 U13775 ( .A1(n13227), .A2(n10890), .ZN(n10891) );
  NAND2_X1 U13776 ( .A1(n11100), .A2(n10891), .ZN(n10892) );
  AOI21_X1 U13777 ( .B1(n10894), .B2(n10893), .A(n10892), .ZN(n16148) );
  AOI21_X1 U13778 ( .B1(n16148), .B2(n11098), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14984) );
  NAND2_X1 U13779 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10895), .ZN(n10896) );
  NOR2_X1 U13780 ( .A1(n9666), .A2(n10896), .ZN(n10897) );
  NOR2_X1 U13781 ( .A1(n10902), .A2(n10897), .ZN(n16135) );
  NAND2_X1 U13782 ( .A1(n16135), .A2(n11098), .ZN(n10899) );
  XNOR2_X1 U13783 ( .A(n10899), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14976) );
  INV_X1 U13784 ( .A(n16148), .ZN(n10898) );
  INV_X1 U13785 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15146) );
  INV_X1 U13786 ( .A(n10899), .ZN(n10900) );
  NAND2_X1 U13787 ( .A1(n10900), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10901) );
  NAND2_X1 U13788 ( .A1(n13227), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U13789 ( .A1(n16125), .A2(n11098), .ZN(n11091) );
  INV_X1 U13790 ( .A(n10903), .ZN(n10904) );
  INV_X1 U13791 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11060) );
  NOR2_X1 U13792 ( .A1(n9665), .A2(n11060), .ZN(n10906) );
  NAND2_X1 U13793 ( .A1(n16125), .A2(n10906), .ZN(n10907) );
  NAND2_X1 U13794 ( .A1(n11093), .A2(n10907), .ZN(n14774) );
  INV_X1 U13795 ( .A(n10908), .ZN(n10914) );
  NAND2_X1 U13796 ( .A1(n11108), .A2(n10909), .ZN(n10923) );
  INV_X1 U13797 ( .A(n11109), .ZN(n11112) );
  AND2_X1 U13798 ( .A1(n10923), .A2(n11112), .ZN(n10912) );
  OAI21_X1 U13799 ( .B1(n10912), .B2(n10911), .A(n10910), .ZN(n10913) );
  NOR2_X1 U13800 ( .A1(n10914), .A2(n10913), .ZN(n10917) );
  NOR2_X1 U13801 ( .A1(n15693), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10915) );
  OR2_X1 U13802 ( .A1(n10917), .A2(n11124), .ZN(n19904) );
  INV_X1 U13803 ( .A(n19904), .ZN(n10919) );
  AND2_X1 U13804 ( .A1(n10378), .A2(n13763), .ZN(n12972) );
  AND2_X1 U13805 ( .A1(n10918), .A2(n12972), .ZN(n19903) );
  NAND2_X1 U13806 ( .A1(n10919), .A2(n19903), .ZN(n11131) );
  INV_X1 U13807 ( .A(n10918), .ZN(n10920) );
  NOR2_X1 U13808 ( .A1(n10920), .A2(n12987), .ZN(n19901) );
  NAND2_X1 U13809 ( .A1(n11107), .A2(n11120), .ZN(n10927) );
  NAND2_X1 U13810 ( .A1(n10924), .A2(n10923), .ZN(n11110) );
  NOR2_X1 U13811 ( .A1(n11110), .A2(n10927), .ZN(n10925) );
  OR2_X1 U13812 ( .A1(n11124), .A2(n10925), .ZN(n13636) );
  INV_X1 U13813 ( .A(n13636), .ZN(n10926) );
  OAI21_X1 U13814 ( .B1(n11109), .B2(n10927), .A(n10926), .ZN(n10928) );
  INV_X1 U13815 ( .A(n10928), .ZN(n10930) );
  NAND3_X1 U13816 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10929) );
  NAND2_X1 U13817 ( .A1(n13168), .A2(n10929), .ZN(n13165) );
  INV_X1 U13818 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n15692) );
  OAI21_X1 U13819 ( .B1(n10667), .B2(n13165), .A(n15692), .ZN(n19892) );
  MUX2_X1 U13820 ( .A(n10930), .B(n19892), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19900) );
  NAND2_X1 U13821 ( .A1(n19901), .A2(n19900), .ZN(n10931) );
  NAND2_X1 U13822 ( .A1(n11131), .A2(n10931), .ZN(n10933) );
  NAND2_X1 U13823 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11027), .ZN(n19762) );
  INV_X1 U13824 ( .A(n19762), .ZN(n10932) );
  NAND2_X1 U13825 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10932), .ZN(n13163) );
  INV_X1 U13826 ( .A(n13051), .ZN(n10934) );
  NAND2_X1 U13827 ( .A1(n11151), .A2(n19222), .ZN(n11071) );
  XOR2_X1 U13828 ( .A(n11228), .B(n10935), .Z(n13187) );
  NAND2_X1 U13829 ( .A1(n13170), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13169) );
  XOR2_X1 U13830 ( .A(n11210), .B(n11220), .Z(n10936) );
  NOR2_X1 U13831 ( .A1(n13169), .A2(n10936), .ZN(n10938) );
  INV_X1 U13832 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15334) );
  INV_X1 U13833 ( .A(n13169), .ZN(n10937) );
  XOR2_X1 U13834 ( .A(n10937), .B(n10936), .Z(n13100) );
  NOR2_X1 U13835 ( .A1(n15334), .A2(n13100), .ZN(n13099) );
  NOR2_X1 U13836 ( .A1(n10938), .A2(n13099), .ZN(n10939) );
  XOR2_X1 U13837 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10939), .Z(
        n13186) );
  NOR2_X1 U13838 ( .A1(n13187), .A2(n13186), .ZN(n13185) );
  NOR2_X1 U13839 ( .A1(n10939), .A2(n13197), .ZN(n10940) );
  XNOR2_X1 U13840 ( .A(n10942), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13733) );
  INV_X1 U13841 ( .A(n13733), .ZN(n10941) );
  NAND2_X1 U13842 ( .A1(n10942), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10943) );
  NAND2_X1 U13843 ( .A1(n13731), .A2(n10943), .ZN(n10944) );
  NAND2_X1 U13844 ( .A1(n13797), .A2(n13860), .ZN(n10949) );
  NAND2_X1 U13845 ( .A1(n10944), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10947) );
  OAI21_X1 U13846 ( .B1(n10946), .B2(n11203), .A(n10945), .ZN(n13795) );
  NAND2_X1 U13847 ( .A1(n10947), .A2(n13795), .ZN(n10948) );
  NAND2_X1 U13848 ( .A1(n10950), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13857) );
  NAND2_X1 U13849 ( .A1(n10956), .A2(n10955), .ZN(n10960) );
  XNOR2_X1 U13850 ( .A(n10960), .B(n16322), .ZN(n15102) );
  INV_X1 U13851 ( .A(n10957), .ZN(n10958) );
  XNOR2_X1 U13852 ( .A(n10964), .B(n11098), .ZN(n15103) );
  NAND2_X1 U13853 ( .A1(n10960), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10961) );
  XNOR2_X1 U13854 ( .A(n10963), .B(n10962), .ZN(n16266) );
  INV_X1 U13855 ( .A(n10964), .ZN(n10965) );
  NAND3_X1 U13856 ( .A1(n10965), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11098), .ZN(n10966) );
  INV_X1 U13857 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16252) );
  NOR3_X1 U13858 ( .A1(n15292), .A2(n16252), .A3(n15274), .ZN(n15242) );
  INV_X1 U13859 ( .A(n15242), .ZN(n15265) );
  INV_X1 U13860 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15261) );
  NOR3_X1 U13861 ( .A1(n10847), .A2(n10813), .A3(n15261), .ZN(n16283) );
  INV_X1 U13862 ( .A(n16283), .ZN(n15243) );
  NOR2_X1 U13863 ( .A1(n15265), .A2(n15243), .ZN(n15239) );
  AND3_X1 U13864 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10967) );
  AND2_X1 U13865 ( .A1(n15239), .A2(n10967), .ZN(n15202) );
  INV_X1 U13866 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15132) );
  INV_X1 U13867 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11183) );
  INV_X1 U13868 ( .A(n11072), .ZN(n10968) );
  OAI21_X1 U13869 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14966), .A(
        n10968), .ZN(n11152) );
  NAND2_X1 U13870 ( .A1(n11027), .A2(n19888), .ZN(n19861) );
  INV_X1 U13871 ( .A(n19861), .ZN(n19850) );
  OR2_X1 U13872 ( .A1(n19864), .A2(n19850), .ZN(n19887) );
  NAND2_X1 U13873 ( .A1(n19887), .A2(n12960), .ZN(n10969) );
  NAND2_X1 U13874 ( .A1(n12960), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12592) );
  INV_X1 U13875 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19470) );
  NAND2_X1 U13876 ( .A1(n19470), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U13877 ( .A1(n12592), .A2(n10970), .ZN(n19231) );
  INV_X1 U13878 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U13879 ( .A1(n12962), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12957) );
  NAND2_X1 U13880 ( .A1(n12958), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12955) );
  AND2_X1 U13881 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10971) );
  INV_X1 U13882 ( .A(n12939), .ZN(n10972) );
  AND2_X2 U13883 ( .A1(n10972), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12940) );
  INV_X1 U13884 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14988) );
  INV_X1 U13885 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U13886 ( .A1(n10973), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11084) );
  INV_X1 U13887 ( .A(n11084), .ZN(n10974) );
  AOI21_X1 U13888 ( .B1(n10975), .B2(n12934), .A(n10974), .ZN(n14771) );
  NOR2_X1 U13889 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19861), .ZN(n18859) );
  NAND2_X1 U13890 ( .A1(n19044), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11411) );
  OAI21_X1 U13891 ( .B1(n19229), .B2(n10975), .A(n11411), .ZN(n11067) );
  INV_X1 U13892 ( .A(n10442), .ZN(n11082) );
  NAND2_X1 U13893 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10979) );
  NAND2_X1 U13894 ( .A1(n9674), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U13895 ( .A1(n10993), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10976) );
  AND2_X1 U13896 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13897 ( .A1(n10979), .A2(n10978), .ZN(n13834) );
  INV_X1 U13898 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18940) );
  AOI22_X1 U13899 ( .A1(n10993), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10980) );
  OAI21_X1 U13900 ( .B1(n11061), .B2(n18940), .A(n10980), .ZN(n10981) );
  AOI21_X1 U13901 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11079), .A(
        n10981), .ZN(n13778) );
  AOI22_X1 U13902 ( .A1(n10993), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10982) );
  OAI21_X1 U13903 ( .B1(n11061), .B2(n13482), .A(n10982), .ZN(n10983) );
  AOI21_X1 U13904 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n11079), .A(
        n10983), .ZN(n13479) );
  INV_X1 U13905 ( .A(n10984), .ZN(n10988) );
  NOR2_X1 U13906 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  NAND2_X1 U13907 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10990) );
  AOI22_X1 U13908 ( .A1(n10993), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10989) );
  OAI211_X1 U13909 ( .C1(n13313), .C2(n11061), .A(n10990), .B(n10989), .ZN(
        n13310) );
  AOI22_X1 U13910 ( .A1(n10993), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10992) );
  NAND2_X1 U13911 ( .A1(n9674), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10991) );
  OAI211_X1 U13912 ( .C1(n11082), .C2(n10739), .A(n10992), .B(n10991), .ZN(
        n13468) );
  AOI22_X1 U13913 ( .A1(n10993), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10995) );
  NAND2_X1 U13914 ( .A1(n11051), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10994) );
  OAI211_X1 U13915 ( .C1(n11082), .C2(n15313), .A(n10995), .B(n10994), .ZN(
        n13369) );
  NAND2_X1 U13916 ( .A1(n13368), .A2(n13369), .ZN(n13478) );
  NOR2_X2 U13917 ( .A1(n13479), .A2(n13478), .ZN(n13484) );
  NAND2_X1 U13918 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10997) );
  AOI22_X1 U13919 ( .A1(n10993), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10996) );
  OAI211_X1 U13920 ( .C1(n10998), .C2(n11061), .A(n10997), .B(n10996), .ZN(
        n13485) );
  NAND2_X1 U13921 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U13922 ( .A1(n9674), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13923 ( .A1(n10993), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10999) );
  AND2_X1 U13924 ( .A1(n11000), .A2(n10999), .ZN(n11001) );
  NAND2_X1 U13925 ( .A1(n11002), .A2(n11001), .ZN(n13455) );
  INV_X1 U13926 ( .A(n13455), .ZN(n11006) );
  AOI22_X1 U13927 ( .A1(n10993), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11004) );
  NAND2_X1 U13928 ( .A1(n11051), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11003) );
  NAND2_X1 U13929 ( .A1(n11004), .A2(n11003), .ZN(n11005) );
  AOI21_X1 U13930 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11005), .ZN(n13463) );
  AOI22_X1 U13931 ( .A1(n10993), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11009) );
  NAND2_X1 U13932 ( .A1(n9674), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U13933 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  AOI21_X1 U13934 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11010), .ZN(n13510) );
  AOI22_X1 U13935 ( .A1(n10993), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11013) );
  NAND2_X1 U13936 ( .A1(n11051), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U13937 ( .A1(n11013), .A2(n11012), .ZN(n11014) );
  AOI21_X1 U13938 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11014), .ZN(n13658) );
  AOI22_X1 U13939 ( .A1(n10993), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11016) );
  NAND2_X1 U13940 ( .A1(n11051), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U13941 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  AOI21_X1 U13942 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11017), .ZN(n15256) );
  NAND2_X1 U13943 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11019) );
  AOI22_X1 U13944 ( .A1(n10993), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11018) );
  OAI211_X1 U13945 ( .C1(n11020), .C2(n11061), .A(n11019), .B(n11018), .ZN(
        n13753) );
  AOI22_X1 U13946 ( .A1(n10993), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11022) );
  NAND2_X1 U13947 ( .A1(n9674), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U13948 ( .A1(n11022), .A2(n11021), .ZN(n11023) );
  AOI21_X1 U13949 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11023), .ZN(n15078) );
  INV_X1 U13950 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13951 ( .A1(n10993), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11024) );
  OAI21_X1 U13952 ( .B1(n11061), .B2(n11025), .A(n11024), .ZN(n11026) );
  AOI21_X1 U13953 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11026), .ZN(n14847) );
  NAND2_X1 U13954 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11031) );
  INV_X1 U13955 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19813) );
  INV_X1 U13956 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18902) );
  OAI22_X1 U13957 ( .A1(n11028), .A2(n19813), .B1(n11027), .B2(n18902), .ZN(
        n11029) );
  AOI21_X1 U13958 ( .B1(n11051), .B2(P2_EBX_REG_19__SCAN_IN), .A(n11029), .ZN(
        n11030) );
  NAND2_X1 U13959 ( .A1(n11031), .A2(n11030), .ZN(n15056) );
  NAND2_X1 U13960 ( .A1(n15057), .A2(n15056), .ZN(n15059) );
  INV_X1 U13961 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U13962 ( .A1(n10993), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11032) );
  OAI21_X1 U13963 ( .B1(n11061), .B2(n11033), .A(n11032), .ZN(n11034) );
  AOI21_X1 U13964 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11034), .ZN(n14841) );
  AOI22_X1 U13965 ( .A1(n10993), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11036) );
  NAND2_X1 U13966 ( .A1(n9674), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U13967 ( .A1(n11036), .A2(n11035), .ZN(n11037) );
  AOI21_X1 U13968 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11037), .ZN(n13027) );
  OR2_X2 U13969 ( .A1(n14843), .A2(n13027), .ZN(n14831) );
  INV_X1 U13970 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U13971 ( .A1(n10993), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11038) );
  OAI21_X1 U13972 ( .B1(n11061), .B2(n15635), .A(n11038), .ZN(n11039) );
  AOI21_X1 U13973 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11039), .ZN(n14830) );
  NAND2_X1 U13974 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U13975 ( .A1(n11051), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U13976 ( .A1(n10993), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11040) );
  AND2_X1 U13977 ( .A1(n11041), .A2(n11040), .ZN(n11042) );
  NAND2_X1 U13978 ( .A1(n11043), .A2(n11042), .ZN(n14825) );
  NAND2_X1 U13979 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11047) );
  NAND2_X1 U13980 ( .A1(n11051), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13981 ( .A1(n10993), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11044) );
  AND2_X1 U13982 ( .A1(n11045), .A2(n11044), .ZN(n11046) );
  NAND2_X1 U13983 ( .A1(n11047), .A2(n11046), .ZN(n14779) );
  AOI22_X1 U13984 ( .A1(n10443), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11049) );
  NAND2_X1 U13985 ( .A1(n11051), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11048) );
  NAND2_X1 U13986 ( .A1(n11049), .A2(n11048), .ZN(n11050) );
  AOI21_X1 U13987 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11050), .ZN(n14819) );
  AOI22_X1 U13988 ( .A1(n10443), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11053) );
  NAND2_X1 U13989 ( .A1(n9674), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U13990 ( .A1(n11053), .A2(n11052), .ZN(n11054) );
  AOI21_X1 U13991 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11054), .ZN(n14809) );
  NOR2_X2 U13992 ( .A1(n9696), .A2(n14809), .ZN(n14810) );
  NAND2_X1 U13993 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11058) );
  NAND2_X1 U13994 ( .A1(n9674), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U13995 ( .A1(n10443), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11055) );
  AND2_X1 U13996 ( .A1(n11056), .A2(n11055), .ZN(n11057) );
  NAND2_X1 U13997 ( .A1(n11058), .A2(n11057), .ZN(n14804) );
  AOI22_X1 U13998 ( .A1(n10443), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11059) );
  OAI21_X1 U13999 ( .B1(n11061), .B2(n11060), .A(n11059), .ZN(n11062) );
  AOI21_X1 U14000 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11062), .ZN(n11063) );
  NAND2_X1 U14001 ( .A1(n14806), .A2(n11063), .ZN(n11064) );
  NAND2_X1 U14002 ( .A1(n11065), .A2(n11064), .ZN(n14799) );
  AND2_X1 U14003 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19877) );
  NOR2_X1 U14004 ( .A1(n14799), .A2(n16206), .ZN(n11066) );
  AOI211_X1 U14005 ( .C1(n19220), .C2(n14771), .A(n11067), .B(n11066), .ZN(
        n11068) );
  NAND2_X1 U14006 ( .A1(n11071), .A2(n11070), .ZN(P2_U2986) );
  INV_X1 U14007 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11073) );
  INV_X1 U14008 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U14009 ( .A1(n10443), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11075) );
  NAND2_X1 U14010 ( .A1(n9674), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11074) );
  OAI211_X1 U14011 ( .C1(n11082), .C2(n12570), .A(n11075), .B(n11074), .ZN(
        n12563) );
  AOI22_X1 U14012 ( .A1(n10443), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11077) );
  NAND2_X1 U14013 ( .A1(n11051), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U14014 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  AOI21_X1 U14015 ( .B1(n11079), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11078), .ZN(n12928) );
  AOI22_X1 U14016 ( .A1(n10443), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11081) );
  NAND2_X1 U14017 ( .A1(n9674), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11080) );
  OAI211_X1 U14018 ( .C1(n11082), .C2(n11073), .A(n11081), .B(n11080), .ZN(
        n11083) );
  INV_X1 U14019 ( .A(n16172), .ZN(n16103) );
  INV_X1 U14020 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U14021 ( .A1(n12577), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11086) );
  INV_X1 U14022 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U14023 ( .A1(n19044), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U14024 ( .A1(n19230), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11087) );
  OAI211_X1 U14025 ( .C1(n16256), .C2(n12932), .A(n12551), .B(n11087), .ZN(
        n11088) );
  AOI21_X1 U14026 ( .B1(n16103), .B2(n19239), .A(n11088), .ZN(n11089) );
  NAND2_X1 U14027 ( .A1(n13227), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11094) );
  XOR2_X1 U14028 ( .A(n11094), .B(n11093), .Z(n11097) );
  OAI21_X1 U14029 ( .B1(n11097), .B2(n10801), .A(n12570), .ZN(n12573) );
  NAND2_X1 U14030 ( .A1(n13227), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11095) );
  XNOR2_X1 U14031 ( .A(n11099), .B(n11095), .ZN(n12984) );
  AOI21_X1 U14032 ( .B1(n12984), .B2(n11098), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14230) );
  AND2_X1 U14033 ( .A1(n11098), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11096) );
  NAND2_X1 U14034 ( .A1(n12984), .A2(n11096), .ZN(n14231) );
  INV_X1 U14035 ( .A(n11097), .ZN(n16109) );
  NAND3_X1 U14036 ( .A1(n16109), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11098), .ZN(n14228) );
  OAI21_X1 U14037 ( .B1(n11099), .B2(P2_EBX_REG_30__SCAN_IN), .A(n13227), .ZN(
        n11101) );
  NAND2_X1 U14038 ( .A1(n11101), .A2(n11100), .ZN(n16098) );
  NOR2_X1 U14039 ( .A1(n16098), .A2(n10801), .ZN(n11102) );
  XNOR2_X1 U14040 ( .A(n11102), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11103) );
  NAND2_X1 U14041 ( .A1(n12541), .A2(n19222), .ZN(n11104) );
  NAND2_X1 U14042 ( .A1(n9713), .A2(n11104), .ZN(P2_U2983) );
  INV_X1 U14043 ( .A(n11105), .ZN(n11118) );
  AOI21_X1 U14044 ( .B1(n11123), .B2(n11215), .A(n11107), .ZN(n11117) );
  INV_X1 U14045 ( .A(n11107), .ZN(n11115) );
  OAI21_X1 U14046 ( .B1(n11109), .B2(n11108), .A(n10683), .ZN(n11114) );
  INV_X1 U14047 ( .A(n11110), .ZN(n11111) );
  OAI211_X1 U14048 ( .C1(n11215), .C2(n11112), .A(n10374), .B(n11111), .ZN(
        n11113) );
  OAI211_X1 U14049 ( .C1(n11106), .C2(n11115), .A(n11114), .B(n11113), .ZN(
        n11116) );
  OAI211_X1 U14050 ( .C1(n11118), .C2(n11117), .A(n11116), .B(n11120), .ZN(
        n11119) );
  OAI21_X1 U14051 ( .B1(n11120), .B2(n12987), .A(n11119), .ZN(n11121) );
  OR2_X1 U14052 ( .A1(n11124), .A2(n11121), .ZN(n11122) );
  INV_X1 U14053 ( .A(n11123), .ZN(n19152) );
  NAND2_X1 U14054 ( .A1(n11124), .A2(n19152), .ZN(n11125) );
  NAND2_X1 U14055 ( .A1(n13641), .A2(n11215), .ZN(n19149) );
  NOR2_X1 U14056 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19775) );
  AOI211_X1 U14057 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19775), .ZN(n19150) );
  INV_X1 U14058 ( .A(n19150), .ZN(n19770) );
  NAND2_X1 U14059 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19764) );
  INV_X1 U14060 ( .A(n19764), .ZN(n19778) );
  NOR2_X1 U14061 ( .A1(n19770), .A2(n19778), .ZN(n13158) );
  NAND2_X1 U14062 ( .A1(n13941), .A2(n13158), .ZN(n11149) );
  AOI21_X1 U14063 ( .B1(n11127), .B2(n10374), .A(n11126), .ZN(n11128) );
  NAND2_X1 U14064 ( .A1(n19149), .A2(n11128), .ZN(n11148) );
  MUX2_X1 U14065 ( .A(n11186), .B(n13941), .S(n10378), .Z(n11129) );
  NAND2_X1 U14066 ( .A1(n11129), .A2(n19764), .ZN(n11132) );
  NAND3_X1 U14067 ( .A1(n10918), .A2(n11215), .A3(n19900), .ZN(n11130) );
  OAI211_X1 U14068 ( .C1(n13636), .C2(n11132), .A(n11131), .B(n11130), .ZN(
        n11146) );
  NAND2_X1 U14069 ( .A1(n11186), .A2(n13158), .ZN(n11133) );
  OR2_X1 U14070 ( .A1(n13636), .A2(n11133), .ZN(n11145) );
  NAND2_X1 U14071 ( .A1(n11134), .A2(n11163), .ZN(n11136) );
  NAND2_X1 U14072 ( .A1(n11135), .A2(n10374), .ZN(n13157) );
  NAND2_X1 U14073 ( .A1(n11136), .A2(n13157), .ZN(n11144) );
  INV_X1 U14074 ( .A(n13931), .ZN(n13238) );
  NOR2_X1 U14075 ( .A1(n11137), .A2(n13238), .ZN(n11218) );
  NAND2_X1 U14076 ( .A1(n11218), .A2(n10402), .ZN(n11138) );
  NAND2_X1 U14077 ( .A1(n11138), .A2(n12972), .ZN(n11154) );
  NAND2_X1 U14078 ( .A1(n10378), .A2(n19245), .ZN(n11171) );
  NAND2_X1 U14079 ( .A1(n11171), .A2(n10374), .ZN(n11140) );
  NAND2_X1 U14080 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  NAND2_X1 U14081 ( .A1(n11141), .A2(n11163), .ZN(n11142) );
  AND2_X1 U14082 ( .A1(n11154), .A2(n11142), .ZN(n11143) );
  NAND2_X1 U14083 ( .A1(n11145), .A2(n11173), .ZN(n13152) );
  NOR2_X1 U14084 ( .A1(n11146), .A2(n13152), .ZN(n11147) );
  OAI211_X1 U14085 ( .C1(n19149), .C2(n11149), .A(n11148), .B(n11147), .ZN(
        n11150) );
  NAND2_X1 U14086 ( .A1(n11151), .A2(n16334), .ZN(n11417) );
  NAND2_X1 U14087 ( .A1(n11134), .A2(n13931), .ZN(n11153) );
  NAND2_X1 U14088 ( .A1(n11153), .A2(n11215), .ZN(n13616) );
  NAND2_X1 U14089 ( .A1(n13616), .A2(n11154), .ZN(n11155) );
  NAND2_X1 U14090 ( .A1(n11155), .A2(n13936), .ZN(n11168) );
  NAND3_X1 U14091 ( .A1(n11156), .A2(n11161), .A3(n10407), .ZN(n11167) );
  INV_X1 U14092 ( .A(n11157), .ZN(n11165) );
  OR2_X1 U14093 ( .A1(n11106), .A2(n11158), .ZN(n11188) );
  INV_X1 U14094 ( .A(n11188), .ZN(n11160) );
  NAND2_X1 U14095 ( .A1(n11160), .A2(n11159), .ZN(n13223) );
  INV_X1 U14096 ( .A(n13049), .ZN(n13044) );
  OAI21_X1 U14097 ( .B1(n11161), .B2(n19245), .A(n13044), .ZN(n11162) );
  OAI211_X1 U14098 ( .C1(n11163), .C2(n10374), .A(n13223), .B(n11162), .ZN(
        n11164) );
  NOR2_X1 U14099 ( .A1(n11165), .A2(n11164), .ZN(n11166) );
  NAND3_X1 U14100 ( .A1(n11168), .A2(n11167), .A3(n11166), .ZN(n13612) );
  OR2_X1 U14101 ( .A1(n13612), .A2(n11169), .ZN(n11170) );
  INV_X1 U14102 ( .A(n15240), .ZN(n11174) );
  INV_X1 U14103 ( .A(n11171), .ZN(n11172) );
  NAND2_X1 U14104 ( .A1(n11198), .A2(n13553), .ZN(n15238) );
  NOR2_X1 U14105 ( .A1(n15132), .A2(n15146), .ZN(n15131) );
  INV_X1 U14106 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15172) );
  NOR2_X1 U14107 ( .A1(n15172), .A2(n15179), .ZN(n15165) );
  AND2_X1 U14108 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15205) );
  NAND2_X1 U14109 ( .A1(n15205), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11181) );
  INV_X1 U14110 ( .A(n11181), .ZN(n11175) );
  AND2_X1 U14111 ( .A1(n15202), .A2(n11175), .ZN(n15188) );
  AOI21_X1 U14112 ( .B1(n15188), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15241), .ZN(n11179) );
  NAND2_X1 U14113 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16319) );
  NAND3_X1 U14114 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11180) );
  INV_X1 U14115 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13177) );
  NOR2_X1 U14116 ( .A1(n15334), .A2(n13177), .ZN(n11176) );
  NOR2_X1 U14117 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11176), .ZN(
        n13189) );
  INV_X1 U14118 ( .A(n13189), .ZN(n11178) );
  NOR2_X1 U14119 ( .A1(n19044), .A2(n11198), .ZN(n13195) );
  INV_X1 U14120 ( .A(n13195), .ZN(n13209) );
  INV_X1 U14121 ( .A(n11176), .ZN(n13206) );
  NOR2_X1 U14122 ( .A1(n13197), .A2(n13206), .ZN(n13737) );
  INV_X1 U14123 ( .A(n13737), .ZN(n11177) );
  NAND2_X1 U14124 ( .A1(n15240), .A2(n11177), .ZN(n13196) );
  OAI211_X1 U14125 ( .C1(n15238), .C2(n11178), .A(n13209), .B(n13196), .ZN(
        n13799) );
  AOI221_X1 U14126 ( .B1(n15313), .B2(n15264), .C1(n11180), .C2(n15264), .A(
        n13799), .ZN(n16337) );
  INV_X1 U14127 ( .A(n16337), .ZN(n15312) );
  AOI21_X1 U14128 ( .B1(n15264), .B2(n16319), .A(n15312), .ZN(n15293) );
  INV_X1 U14129 ( .A(n15293), .ZN(n15263) );
  NOR2_X1 U14130 ( .A1(n11179), .A2(n15263), .ZN(n15197) );
  OAI21_X1 U14131 ( .B1(n15241), .B2(n15165), .A(n15197), .ZN(n15160) );
  AOI21_X1 U14132 ( .B1(n15154), .B2(n15264), .A(n15160), .ZN(n15147) );
  OAI21_X1 U14133 ( .B1(n15241), .B2(n15131), .A(n15147), .ZN(n15127) );
  INV_X1 U14134 ( .A(n15127), .ZN(n11184) );
  NOR2_X1 U14135 ( .A1(n13189), .A2(n15238), .ZN(n13736) );
  AOI21_X1 U14136 ( .B1(n15240), .B2(n13737), .A(n13736), .ZN(n13798) );
  NOR2_X1 U14137 ( .A1(n11180), .A2(n13798), .ZN(n15314) );
  NAND2_X1 U14138 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15314), .ZN(
        n16320) );
  NAND2_X1 U14139 ( .A1(n15273), .A2(n15202), .ZN(n15232) );
  NOR3_X1 U14140 ( .A1(n15196), .A2(n11181), .A3(n15232), .ZN(n15177) );
  AND3_X1 U14141 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15177), .ZN(n15153) );
  AND2_X1 U14142 ( .A1(n15153), .A2(n15131), .ZN(n11182) );
  NAND2_X1 U14143 ( .A1(n12562), .A2(n11183), .ZN(n15123) );
  NAND2_X1 U14144 ( .A1(n11184), .A2(n15123), .ZN(n12560) );
  INV_X1 U14145 ( .A(n11185), .ZN(n11191) );
  NAND2_X1 U14146 ( .A1(n11186), .A2(n13763), .ZN(n13599) );
  NAND2_X1 U14147 ( .A1(n13599), .A2(n13157), .ZN(n13635) );
  NAND2_X1 U14148 ( .A1(n10401), .A2(n13931), .ZN(n11187) );
  NOR2_X1 U14149 ( .A1(n11188), .A2(n11187), .ZN(n11189) );
  OR2_X1 U14150 ( .A1(n13635), .A2(n11189), .ZN(n13621) );
  NAND2_X1 U14151 ( .A1(n13621), .A2(n10378), .ZN(n11190) );
  NAND2_X1 U14152 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  NOR2_X1 U14153 ( .A1(n14799), .A2(n16329), .ZN(n11413) );
  INV_X1 U14154 ( .A(n11193), .ZN(n11195) );
  NAND2_X1 U14155 ( .A1(n11195), .A2(n11194), .ZN(n13554) );
  NAND2_X1 U14156 ( .A1(n13635), .A2(n11215), .ZN(n11196) );
  NAND2_X1 U14157 ( .A1(n13554), .A2(n11196), .ZN(n11197) );
  INV_X1 U14158 ( .A(n11199), .ZN(n11201) );
  NAND2_X1 U14159 ( .A1(n12547), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11209) );
  INV_X1 U14160 ( .A(n11203), .ZN(n11206) );
  NAND2_X1 U14161 ( .A1(n11400), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U14162 ( .A1(n11211), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11204) );
  OAI211_X1 U14163 ( .C1(n11381), .C2(n11206), .A(n11205), .B(n11204), .ZN(
        n11207) );
  INV_X1 U14164 ( .A(n11207), .ZN(n11208) );
  OR2_X1 U14165 ( .A1(n11210), .A2(n11381), .ZN(n11214) );
  MUX2_X1 U14166 ( .A(n13931), .B(n19896), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11212) );
  NAND2_X1 U14167 ( .A1(n11137), .A2(n11211), .ZN(n11226) );
  AND2_X1 U14168 ( .A1(n11212), .A2(n11226), .ZN(n11213) );
  NAND2_X1 U14169 ( .A1(n11214), .A2(n11213), .ZN(n13174) );
  INV_X1 U14170 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18877) );
  AOI21_X1 U14171 ( .B1(n11215), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U14172 ( .A1(n13238), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11216) );
  OAI211_X1 U14173 ( .C1(n12546), .C2(n18877), .A(n11217), .B(n11216), .ZN(
        n13173) );
  AND2_X2 U14174 ( .A1(n13174), .A2(n13173), .ZN(n13176) );
  INV_X1 U14175 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19214) );
  OAI222_X1 U14176 ( .A1(n11293), .A2(n15334), .B1(n10264), .B2(n19214), .C1(
        n12546), .C2(n10419), .ZN(n11224) );
  XNOR2_X1 U14177 ( .A(n13176), .B(n11224), .ZN(n13203) );
  MUX2_X1 U14178 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n11218), .S(
        n19888), .Z(n11219) );
  INV_X1 U14179 ( .A(n11219), .ZN(n11223) );
  INV_X1 U14180 ( .A(n11220), .ZN(n11221) );
  OR2_X1 U14181 ( .A1(n11221), .A2(n11381), .ZN(n11222) );
  NAND2_X1 U14182 ( .A1(n11223), .A2(n11222), .ZN(n13204) );
  NOR2_X1 U14183 ( .A1(n13203), .A2(n13204), .ZN(n13202) );
  NOR2_X1 U14184 ( .A1(n13176), .A2(n11224), .ZN(n11225) );
  NOR2_X2 U14185 ( .A1(n13202), .A2(n11225), .ZN(n11231) );
  NAND2_X1 U14186 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11227) );
  OAI211_X1 U14187 ( .C1(n11381), .C2(n11228), .A(n11227), .B(n11226), .ZN(
        n11230) );
  XNOR2_X1 U14188 ( .A(n11231), .B(n11230), .ZN(n13182) );
  INV_X1 U14189 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19786) );
  AOI22_X1 U14190 ( .A1(n11400), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11211), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11229) );
  OAI21_X1 U14191 ( .B1(n12546), .B2(n19786), .A(n11229), .ZN(n13181) );
  NOR2_X1 U14192 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  NOR2_X1 U14193 ( .A1(n11231), .A2(n11230), .ZN(n11232) );
  INV_X1 U14194 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13729) );
  AOI22_X1 U14195 ( .A1(n11211), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11233) );
  OAI21_X1 U14196 ( .B1(n12546), .B2(n13729), .A(n11233), .ZN(n11237) );
  NAND2_X1 U14197 ( .A1(n11400), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11234) );
  OAI21_X1 U14198 ( .B1(n11381), .B2(n11235), .A(n11234), .ZN(n11236) );
  OR2_X1 U14199 ( .A1(n11237), .A2(n11236), .ZN(n13738) );
  INV_X1 U14200 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13863) );
  INV_X2 U14201 ( .A(n10264), .ZN(n11400) );
  AOI22_X1 U14202 ( .A1(n11400), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11211), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11240) );
  OR2_X1 U14203 ( .A1(n11381), .A2(n11238), .ZN(n11239) );
  OAI211_X1 U14204 ( .C1(n12546), .C2(n13863), .A(n11240), .B(n11239), .ZN(
        n13862) );
  OR2_X1 U14205 ( .A1(n11381), .A2(n11241), .ZN(n11242) );
  INV_X1 U14206 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U14207 ( .A1(n11400), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11211), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11244) );
  OAI21_X1 U14208 ( .B1(n12546), .B2(n19792), .A(n11244), .ZN(n15316) );
  NAND2_X1 U14209 ( .A1(n15317), .A2(n15316), .ZN(n11246) );
  OR2_X1 U14210 ( .A1(n11381), .A2(n10801), .ZN(n11245) );
  NAND2_X1 U14211 ( .A1(n11246), .A2(n11245), .ZN(n15300) );
  INV_X1 U14212 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19794) );
  OR2_X1 U14213 ( .A1(n12546), .A2(n19794), .ZN(n11248) );
  AOI22_X1 U14214 ( .A1(n11400), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11211), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11247) );
  NAND2_X1 U14215 ( .A1(n11248), .A2(n11247), .ZN(n15299) );
  NAND2_X1 U14216 ( .A1(n15300), .A2(n15299), .ZN(n15301) );
  NAND2_X1 U14217 ( .A1(n12547), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14218 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14219 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14220 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11250) );
  NAND2_X1 U14221 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11249) );
  AND2_X1 U14222 ( .A1(n11250), .A2(n11249), .ZN(n11252) );
  AOI22_X1 U14223 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14224 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11260) );
  AOI22_X1 U14225 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14226 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14227 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U14228 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11255) );
  NAND4_X1 U14229 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n11259) );
  NOR2_X1 U14230 ( .A1(n11260), .A2(n11259), .ZN(n13486) );
  NAND2_X1 U14231 ( .A1(n11400), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U14232 ( .A1(n11211), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11261) );
  OAI211_X1 U14233 ( .C1(n11381), .C2(n13486), .A(n11262), .B(n11261), .ZN(
        n11263) );
  INV_X1 U14234 ( .A(n11263), .ZN(n11264) );
  NOR2_X2 U14235 ( .A1(n15301), .A2(n13874), .ZN(n15286) );
  INV_X1 U14236 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14237 ( .A1(n11400), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11211), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14238 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12705), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14239 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14240 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12719), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11267) );
  NAND2_X1 U14241 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11266) );
  NAND4_X1 U14242 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11277) );
  NAND2_X1 U14243 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11271) );
  AOI22_X1 U14244 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10613), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11270) );
  AND2_X1 U14245 ( .A1(n11271), .A2(n11270), .ZN(n11275) );
  AOI22_X1 U14246 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14247 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14248 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11272) );
  NAND4_X1 U14249 ( .A1(n11275), .A2(n11274), .A3(n11273), .A4(n11272), .ZN(
        n11276) );
  NOR2_X1 U14250 ( .A1(n11277), .A2(n11276), .ZN(n13460) );
  OR2_X1 U14251 ( .A1(n11381), .A2(n13460), .ZN(n11278) );
  OAI211_X1 U14252 ( .C1(n12546), .C2(n11280), .A(n11279), .B(n11278), .ZN(
        n15287) );
  AOI22_X1 U14253 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10762), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14254 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10763), .ZN(n11285) );
  AOI22_X1 U14255 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10613), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U14256 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11281) );
  AND2_X1 U14257 ( .A1(n11282), .A2(n11281), .ZN(n11284) );
  AOI22_X1 U14258 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14259 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11292) );
  AOI22_X1 U14260 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14261 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14262 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U14263 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11287) );
  NAND4_X1 U14264 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n11291) );
  NOR2_X1 U14265 ( .A1(n11292), .A2(n11291), .ZN(n13452) );
  AOI22_X1 U14266 ( .A1(n11400), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11294) );
  OAI21_X1 U14267 ( .B1(n13452), .B2(n11381), .A(n11294), .ZN(n11295) );
  AOI21_X1 U14268 ( .B1(n12547), .B2(P2_REIP_REG_10__SCAN_IN), .A(n11295), 
        .ZN(n16307) );
  INV_X1 U14269 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14270 ( .A1(n11400), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14271 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14272 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12719), .B1(
        n10613), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11297) );
  NAND2_X1 U14273 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11296) );
  AND2_X1 U14274 ( .A1(n11297), .A2(n11296), .ZN(n11300) );
  AOI22_X1 U14275 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14276 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14277 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11307) );
  AOI22_X1 U14278 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14279 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14280 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U14281 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11302) );
  NAND4_X1 U14282 ( .A1(n11305), .A2(n11304), .A3(n11303), .A4(n11302), .ZN(
        n11306) );
  NOR2_X1 U14283 ( .A1(n11307), .A2(n11306), .ZN(n13507) );
  OR2_X1 U14284 ( .A1(n11381), .A2(n13507), .ZN(n11308) );
  OAI211_X1 U14285 ( .C1(n12546), .C2(n11310), .A(n11309), .B(n11308), .ZN(
        n15278) );
  NAND2_X1 U14286 ( .A1(n12547), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14287 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10762), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14288 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n10763), .ZN(n11315) );
  AOI22_X1 U14289 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10613), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11312) );
  NAND2_X1 U14290 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11311) );
  AND2_X1 U14291 ( .A1(n11312), .A2(n11311), .ZN(n11314) );
  AOI22_X1 U14292 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11313) );
  NAND4_X1 U14293 ( .A1(n11316), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n11322) );
  AOI22_X1 U14294 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14295 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14296 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11318) );
  NAND2_X1 U14297 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11317) );
  NAND4_X1 U14298 ( .A1(n11320), .A2(n11319), .A3(n11318), .A4(n11317), .ZN(
        n11321) );
  NOR2_X1 U14299 ( .A1(n11322), .A2(n11321), .ZN(n13656) );
  NAND2_X1 U14300 ( .A1(n11400), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14301 ( .A1(n11211), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11323) );
  OAI211_X1 U14302 ( .C1(n11381), .C2(n13656), .A(n11324), .B(n11323), .ZN(
        n11325) );
  INV_X1 U14303 ( .A(n11325), .ZN(n11326) );
  INV_X1 U14304 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14305 ( .A1(n11400), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14306 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12683), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14307 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U14308 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11328) );
  AND2_X1 U14309 ( .A1(n11329), .A2(n11328), .ZN(n11332) );
  AOI22_X1 U14310 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14311 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11330) );
  NAND4_X1 U14312 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11339) );
  AOI22_X1 U14313 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14314 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14315 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U14316 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11334) );
  NAND4_X1 U14317 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  NOR2_X1 U14318 ( .A1(n11339), .A2(n11338), .ZN(n19077) );
  OR2_X1 U14319 ( .A1(n11381), .A2(n19077), .ZN(n11340) );
  OAI211_X1 U14320 ( .C1(n12546), .C2(n11342), .A(n11341), .B(n11340), .ZN(
        n15253) );
  NAND2_X1 U14321 ( .A1(n12547), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U14322 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11343) );
  OAI21_X1 U14323 ( .B1(n12893), .B2(n13559), .A(n11343), .ZN(n11349) );
  AOI22_X1 U14324 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U14325 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14326 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11345) );
  NAND2_X1 U14327 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11344) );
  NAND4_X1 U14328 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11348) );
  NOR2_X1 U14329 ( .A1(n11349), .A2(n11348), .ZN(n11357) );
  AOI22_X1 U14330 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11353) );
  NAND2_X1 U14331 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14332 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14333 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11350) );
  AND4_X1 U14334 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11356) );
  AOI22_X1 U14335 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14336 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11354) );
  NAND4_X1 U14337 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n13751) );
  INV_X1 U14338 ( .A(n13751), .ZN(n11360) );
  NAND2_X1 U14339 ( .A1(n11400), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U14340 ( .A1(n11211), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11358) );
  OAI211_X1 U14341 ( .C1(n11381), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        n11361) );
  INV_X1 U14342 ( .A(n11361), .ZN(n11362) );
  NOR2_X4 U14343 ( .A1(n15254), .A2(n13961), .ZN(n16271) );
  INV_X1 U14344 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15090) );
  AOI22_X1 U14345 ( .A1(n11400), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14346 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U14347 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11366) );
  NAND2_X1 U14348 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11365) );
  NAND2_X1 U14349 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11364) );
  NAND4_X1 U14350 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11371) );
  NAND2_X1 U14351 ( .A1(n10763), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11368) );
  OAI21_X1 U14352 ( .B1(n12714), .B2(n11369), .A(n11368), .ZN(n11370) );
  NOR2_X1 U14353 ( .A1(n11371), .A2(n11370), .ZN(n11379) );
  AOI22_X1 U14354 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12719), .B1(
        n10613), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11375) );
  NAND2_X1 U14355 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11374) );
  NAND2_X1 U14356 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14357 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11372) );
  AND4_X1 U14358 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11378) );
  AOI22_X1 U14359 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10762), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14360 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14361 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n13780) );
  INV_X1 U14362 ( .A(n13780), .ZN(n11380) );
  OR2_X1 U14363 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  OAI211_X1 U14364 ( .C1(n12546), .C2(n15090), .A(n11383), .B(n11382), .ZN(
        n16272) );
  NAND2_X1 U14365 ( .A1(n12547), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14366 ( .A1(n11400), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11384) );
  INV_X1 U14367 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U14368 ( .A1(n11400), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11386) );
  OAI21_X1 U14369 ( .B1(n12546), .B2(n19810), .A(n11386), .ZN(n15244) );
  INV_X1 U14370 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U14371 ( .A1(n11400), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11387) );
  OAI21_X1 U14372 ( .B1(n12546), .B2(n15070), .A(n11387), .ZN(n11388) );
  INV_X1 U14373 ( .A(n11388), .ZN(n14948) );
  AOI22_X1 U14374 ( .A1(n11400), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11389) );
  OAI21_X1 U14375 ( .B1(n12546), .B2(n19813), .A(n11389), .ZN(n11390) );
  INV_X1 U14376 ( .A(n11390), .ZN(n14939) );
  INV_X1 U14377 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U14378 ( .A1(n11400), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11391) );
  OAI21_X1 U14379 ( .B1(n12546), .B2(n15043), .A(n11391), .ZN(n11392) );
  INV_X1 U14380 ( .A(n11392), .ZN(n14926) );
  NOR2_X2 U14381 ( .A1(n14941), .A2(n14926), .ZN(n14927) );
  INV_X1 U14382 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19816) );
  AOI22_X1 U14383 ( .A1(n11400), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11393) );
  OAI21_X1 U14384 ( .B1(n12546), .B2(n19816), .A(n11393), .ZN(n13029) );
  NAND2_X1 U14385 ( .A1(n14927), .A2(n13029), .ZN(n14908) );
  NAND2_X1 U14386 ( .A1(n12547), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14387 ( .A1(n11400), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11394) );
  INV_X1 U14388 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19820) );
  OR2_X1 U14389 ( .A1(n12546), .A2(n19820), .ZN(n11397) );
  AOI22_X1 U14390 ( .A1(n11400), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11396) );
  NAND2_X1 U14391 ( .A1(n11397), .A2(n11396), .ZN(n14901) );
  NAND2_X1 U14392 ( .A1(n12547), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14393 ( .A1(n11400), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U14394 ( .A1(n11399), .A2(n11398), .ZN(n14880) );
  INV_X1 U14395 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19824) );
  AOI22_X1 U14396 ( .A1(n11400), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11401) );
  OAI21_X1 U14397 ( .B1(n12546), .B2(n19824), .A(n11401), .ZN(n14879) );
  NAND2_X1 U14398 ( .A1(n12547), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14399 ( .A1(n11400), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11403) );
  AND2_X1 U14400 ( .A1(n11404), .A2(n11403), .ZN(n14873) );
  NAND2_X1 U14401 ( .A1(n12547), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14402 ( .A1(n11400), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11405) );
  AND2_X1 U14403 ( .A1(n11406), .A2(n11405), .ZN(n14865) );
  NAND2_X1 U14404 ( .A1(n12547), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14405 ( .A1(n11400), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11407) );
  NAND2_X1 U14406 ( .A1(n11408), .A2(n11407), .ZN(n11409) );
  OAI21_X1 U14407 ( .B1(n14867), .B2(n11409), .A(n12566), .ZN(n14861) );
  INV_X1 U14408 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12561) );
  NAND3_X1 U14409 ( .A1(n12562), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n12561), .ZN(n11410) );
  OAI211_X1 U14410 ( .C1(n16324), .C2(n14861), .A(n11411), .B(n11410), .ZN(
        n11412) );
  AOI211_X1 U14411 ( .C1(n12560), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11413), .B(n11412), .ZN(n11414) );
  NAND2_X1 U14412 ( .A1(n11417), .A2(n11416), .ZN(P2_U3018) );
  NOR2_X2 U14413 ( .A1(n11419), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11425) );
  AND2_X4 U14414 ( .A1(n13261), .A2(n14752), .ZN(n12009) );
  AOI22_X1 U14415 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11424) );
  AND2_X2 U14416 ( .A1(n11420), .A2(n13526), .ZN(n11611) );
  AOI22_X1 U14417 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14418 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11595), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14419 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11421) );
  NAND4_X1 U14420 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11432) );
  AND2_X2 U14421 ( .A1(n11425), .A2(n13261), .ZN(n11870) );
  AOI22_X1 U14422 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11430) );
  BUF_X4 U14423 ( .A(n11479), .Z(n12193) );
  AOI22_X1 U14424 ( .A1(n11479), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11579), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14425 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11473), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14426 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11427) );
  NAND4_X1 U14427 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n11431) );
  AOI22_X1 U14428 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14429 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14430 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14431 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14432 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11595), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14433 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11473), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14434 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14435 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14436 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14437 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11479), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14438 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14439 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14440 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11452) );
  AOI22_X1 U14441 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11595), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14442 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11473), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14443 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14444 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11447) );
  NAND4_X1 U14445 ( .A1(n11450), .A2(n11449), .A3(n11448), .A4(n11447), .ZN(
        n11451) );
  NAND2_X1 U14446 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11456) );
  NAND2_X1 U14447 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11455) );
  NAND2_X1 U14448 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U14449 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11453) );
  NAND2_X1 U14450 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11460) );
  NAND2_X1 U14451 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11459) );
  NAND2_X1 U14452 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11458) );
  NAND2_X1 U14453 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11457) );
  NAND2_X1 U14454 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11464) );
  NAND2_X1 U14455 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11463) );
  NAND2_X1 U14456 ( .A1(n11474), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U14457 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11461) );
  NAND2_X1 U14458 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11468) );
  NAND2_X1 U14459 ( .A1(n11595), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11467) );
  NAND2_X1 U14460 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14461 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11465) );
  AOI22_X1 U14462 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12215), .B1(
        n11595), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14463 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11473), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14464 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11491), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14465 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11475) );
  NAND4_X1 U14466 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11485) );
  AOI22_X1 U14467 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14468 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11501), .B1(
        n11479), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14469 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14470 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11911), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11480) );
  NAND4_X1 U14471 ( .A1(n11483), .A2(n11482), .A3(n11481), .A4(n11480), .ZN(
        n11484) );
  OR2_X2 U14472 ( .A1(n11485), .A2(n11484), .ZN(n11542) );
  INV_X2 U14473 ( .A(n11542), .ZN(n20143) );
  AOI22_X1 U14474 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14475 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14476 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11479), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14477 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11473), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14478 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11497) );
  AOI22_X1 U14479 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14480 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11595), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14481 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14482 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14483 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11496) );
  NAND2_X1 U14484 ( .A1(n20143), .A2(n13580), .ZN(n11543) );
  NAND2_X1 U14485 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11505) );
  NAND2_X1 U14486 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11504) );
  NAND2_X1 U14487 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14488 ( .A1(n12193), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14489 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U14490 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14491 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14492 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11506) );
  NAND2_X1 U14493 ( .A1(n11595), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U14494 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11512) );
  NAND2_X1 U14495 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11511) );
  NAND2_X1 U14496 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11510) );
  NAND2_X1 U14497 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14498 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11516) );
  NAND2_X1 U14499 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11515) );
  NAND2_X1 U14500 ( .A1(n12216), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11514) );
  NAND4_X4 U14501 ( .A1(n11521), .A2(n11520), .A3(n11519), .A4(n11518), .ZN(
        n13402) );
  XNOR2_X1 U14502 ( .A(n20660), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12522) );
  NOR2_X2 U14503 ( .A1(n13278), .A2(n12418), .ZN(n13347) );
  NAND2_X1 U14504 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U14505 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11524) );
  NAND2_X1 U14506 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11523) );
  NAND2_X1 U14507 ( .A1(n12193), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11522) );
  NAND2_X1 U14508 ( .A1(n11579), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14509 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14510 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U14511 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U14512 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11533) );
  NAND2_X1 U14513 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U14514 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U14515 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U14516 ( .A1(n11595), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U14517 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U14518 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11535) );
  NAND2_X1 U14519 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11534) );
  NAND4_X4 U14520 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n13422) );
  NAND3_X1 U14522 ( .A1(n13347), .A2(n14364), .A3(n20139), .ZN(n13245) );
  AOI21_X1 U14523 ( .B1(n13410), .B2(n12522), .A(n13411), .ZN(n11551) );
  INV_X2 U14524 ( .A(n11556), .ZN(n20135) );
  OAI21_X1 U14525 ( .B1(n20139), .B2(n13278), .A(n11672), .ZN(n11544) );
  NAND2_X1 U14526 ( .A1(n13087), .A2(n11544), .ZN(n11547) );
  NAND2_X1 U14527 ( .A1(n11557), .A2(n12418), .ZN(n11546) );
  AND2_X2 U14528 ( .A1(n11547), .A2(n11546), .ZN(n11554) );
  NOR2_X1 U14529 ( .A1(n13088), .A2(n13402), .ZN(n11549) );
  INV_X2 U14530 ( .A(n13422), .ZN(n20124) );
  NAND2_X1 U14531 ( .A1(n11550), .A2(n13422), .ZN(n13273) );
  NAND2_X1 U14532 ( .A1(n11551), .A2(n13397), .ZN(n11552) );
  NAND2_X1 U14533 ( .A1(n13088), .A2(n13278), .ZN(n11553) );
  NAND2_X1 U14534 ( .A1(n11554), .A2(n11553), .ZN(n13248) );
  NAND2_X1 U14535 ( .A1(n13248), .A2(n20107), .ZN(n11559) );
  INV_X1 U14536 ( .A(n13347), .ZN(n11569) );
  NAND2_X1 U14537 ( .A1(n20139), .A2(n13346), .ZN(n11555) );
  NAND2_X1 U14538 ( .A1(n11555), .A2(n13580), .ZN(n12296) );
  NAND2_X1 U14539 ( .A1(n11572), .A2(n12295), .ZN(n11571) );
  NAND2_X1 U14540 ( .A1(n11571), .A2(n11557), .ZN(n11558) );
  NAND2_X1 U14541 ( .A1(n20107), .A2(n13422), .ZN(n13279) );
  NAND4_X1 U14542 ( .A1(n11559), .A2(n11569), .A3(n11558), .A4(n13279), .ZN(
        n11563) );
  NAND2_X1 U14543 ( .A1(n12295), .A2(n13402), .ZN(n11560) );
  NAND2_X1 U14544 ( .A1(n11560), .A2(n20739), .ZN(n11561) );
  NAND2_X1 U14545 ( .A1(n11571), .A2(n11561), .ZN(n13406) );
  INV_X1 U14546 ( .A(n13088), .ZN(n12300) );
  AND2_X1 U14547 ( .A1(n13278), .A2(n13402), .ZN(n11567) );
  AOI21_X1 U14548 ( .B1(n12300), .B2(n14256), .A(n11567), .ZN(n11562) );
  NAND2_X1 U14549 ( .A1(n13406), .A2(n11562), .ZN(n13247) );
  MUX2_X1 U14550 ( .A(n12305), .B(n12294), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11565) );
  INV_X1 U14551 ( .A(n14364), .ZN(n13574) );
  NAND3_X1 U14552 ( .A1(n12295), .A2(n13574), .A3(n12418), .ZN(n11566) );
  NAND2_X1 U14553 ( .A1(n13248), .A2(n11566), .ZN(n11577) );
  INV_X1 U14554 ( .A(n11567), .ZN(n11568) );
  OAI21_X1 U14555 ( .B1(n11569), .B2(n13346), .A(n11568), .ZN(n13404) );
  NAND3_X1 U14556 ( .A1(n13279), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n16083), 
        .ZN(n11570) );
  NOR2_X1 U14557 ( .A1(n13404), .A2(n11570), .ZN(n11576) );
  NAND3_X1 U14558 ( .A1(n11571), .A2(n13422), .A3(n11557), .ZN(n11575) );
  INV_X1 U14559 ( .A(n11572), .ZN(n11573) );
  NAND2_X1 U14560 ( .A1(n11573), .A2(n13319), .ZN(n11574) );
  NAND4_X1 U14561 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11632) );
  INV_X1 U14562 ( .A(n11632), .ZN(n11578) );
  AOI22_X1 U14563 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14564 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14565 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14566 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U14567 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AOI22_X1 U14568 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14569 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14570 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14571 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14572 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  AOI22_X1 U14573 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14574 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14575 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14576 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11591) );
  NAND4_X1 U14577 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(
        n11601) );
  AOI22_X1 U14578 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11599) );
  INV_X2 U14579 ( .A(n11580), .ZN(n12194) );
  AOI22_X1 U14580 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14581 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14582 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11596) );
  NAND4_X1 U14583 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11600) );
  XNOR2_X1 U14584 ( .A(n11606), .B(n12377), .ZN(n11602) );
  NAND2_X1 U14585 ( .A1(n11602), .A2(n11636), .ZN(n11603) );
  INV_X1 U14586 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U14587 ( .A1(n20135), .A2(n12377), .ZN(n11605) );
  OAI211_X1 U14588 ( .C1(n11606), .C2(n13402), .A(n11605), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11607) );
  INV_X1 U14589 ( .A(n11607), .ZN(n11608) );
  NAND2_X1 U14590 ( .A1(n11636), .A2(n12377), .ZN(n11610) );
  INV_X1 U14591 ( .A(n12377), .ZN(n12384) );
  NOR2_X1 U14592 ( .A1(n13402), .A2(n20644), .ZN(n11669) );
  AOI22_X1 U14593 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14594 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14595 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14596 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14597 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11621) );
  AOI22_X1 U14598 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14599 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14600 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14601 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11616) );
  NAND4_X1 U14602 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11620) );
  AOI22_X1 U14603 ( .A1(n11636), .A2(n12384), .B1(n11669), .B2(n12321), .ZN(
        n11623) );
  NAND2_X1 U14604 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U14605 ( .A1(n11623), .A2(n11622), .ZN(n11624) );
  NAND2_X1 U14606 ( .A1(n11625), .A2(n11624), .ZN(n11626) );
  NAND2_X1 U14607 ( .A1(n11643), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11629) );
  NAND2_X1 U14608 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11646) );
  OAI21_X1 U14609 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11646), .ZN(n20415) );
  NAND2_X1 U14610 ( .A1(n15667), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11640) );
  OAI21_X1 U14611 ( .B1(n12305), .B2(n20415), .A(n11640), .ZN(n11627) );
  INV_X1 U14612 ( .A(n11627), .ZN(n11628) );
  XNOR2_X2 U14613 ( .A(n11631), .B(n11630), .ZN(n20216) );
  INV_X1 U14614 ( .A(n20216), .ZN(n11634) );
  INV_X1 U14615 ( .A(n11635), .ZN(n11633) );
  NAND2_X2 U14616 ( .A1(n20216), .A2(n11635), .ZN(n11655) );
  OR2_X2 U14617 ( .A1(n13545), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11638) );
  NAND2_X1 U14618 ( .A1(n11636), .A2(n12321), .ZN(n11637) );
  NAND2_X2 U14619 ( .A1(n11638), .A2(n11637), .ZN(n12314) );
  INV_X1 U14620 ( .A(n11630), .ZN(n11642) );
  NAND2_X1 U14621 ( .A1(n11640), .A2(n9829), .ZN(n11641) );
  NAND2_X1 U14622 ( .A1(n11642), .A2(n11641), .ZN(n11653) );
  NAND2_X1 U14623 ( .A1(n11655), .A2(n11653), .ZN(n11649) );
  NAND2_X1 U14624 ( .A1(n11699), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U14625 ( .A1(n15667), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U14626 ( .A1(n11645), .A2(n11644), .ZN(n11650) );
  INV_X1 U14627 ( .A(n12305), .ZN(n11701) );
  NAND2_X1 U14628 ( .A1(n11646), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11647) );
  NAND3_X1 U14629 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20474), .ZN(n20446) );
  NAND2_X1 U14630 ( .A1(n11647), .A2(n20446), .ZN(n20119) );
  INV_X1 U14631 ( .A(n11650), .ZN(n11654) );
  INV_X1 U14632 ( .A(n11651), .ZN(n11652) );
  NAND4_X1 U14633 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(
        n11656) );
  AOI22_X1 U14634 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11661) );
  INV_X1 U14635 ( .A(n11501), .ZN(n11729) );
  INV_X1 U14636 ( .A(n11729), .ZN(n11657) );
  AOI22_X1 U14637 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14638 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14639 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U14640 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11667) );
  AOI22_X1 U14641 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14642 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14643 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14644 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11662) );
  NAND4_X1 U14645 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11662), .ZN(
        n11666) );
  OAI22_X2 U14646 ( .A1(n13515), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12323), 
        .B2(n12380), .ZN(n11671) );
  AOI22_X1 U14647 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11669), .B2(n11668), .ZN(n11670) );
  NAND2_X1 U14648 ( .A1(n12319), .A2(n11830), .ZN(n11679) );
  AND2_X1 U14649 ( .A1(n11672), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11726) );
  INV_X1 U14650 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11676) );
  NOR2_X2 U14651 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11674) );
  INV_X1 U14652 ( .A(n12240), .ZN(n12209) );
  XNOR2_X1 U14653 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14396) );
  AOI21_X1 U14654 ( .B1(n12209), .B2(n14396), .A(n12241), .ZN(n11675) );
  OAI21_X1 U14655 ( .B1(n12146), .B2(n11676), .A(n11675), .ZN(n11677) );
  AOI21_X1 U14656 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n11726), .A(
        n11677), .ZN(n11678) );
  NAND2_X1 U14657 ( .A1(n11679), .A2(n11678), .ZN(n11680) );
  NAND2_X1 U14658 ( .A1(n12241), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11695) );
  NAND2_X1 U14659 ( .A1(n20185), .A2(n11830), .ZN(n11685) );
  INV_X1 U14660 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11682) );
  INV_X1 U14661 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19988) );
  OAI22_X1 U14662 ( .A1(n12146), .A2(n11682), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n19988), .ZN(n11683) );
  AOI21_X1 U14663 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11726), .A(
        n11683), .ZN(n11684) );
  NAND2_X1 U14664 ( .A1(n11685), .A2(n11684), .ZN(n13361) );
  NAND2_X1 U14665 ( .A1(n20184), .A2(n20143), .ZN(n11687) );
  NAND2_X1 U14666 ( .A1(n11687), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13353) );
  INV_X1 U14667 ( .A(n11726), .ZN(n11744) );
  NAND2_X1 U14668 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14669 ( .A1(n12242), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11690) );
  OAI211_X1 U14670 ( .C1(n11744), .C2(n11419), .A(n11691), .B(n11690), .ZN(
        n11692) );
  AOI21_X1 U14671 ( .B1(n11689), .B2(n11830), .A(n11692), .ZN(n11693) );
  OR2_X1 U14672 ( .A1(n13353), .A2(n11693), .ZN(n13354) );
  INV_X1 U14673 ( .A(n11693), .ZN(n13355) );
  OR2_X1 U14674 ( .A1(n13355), .A2(n12240), .ZN(n11694) );
  NAND2_X1 U14675 ( .A1(n13354), .A2(n11694), .ZN(n13360) );
  INV_X1 U14676 ( .A(n11696), .ZN(n11698) );
  NAND2_X1 U14677 ( .A1(n11699), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11703) );
  NAND3_X1 U14678 ( .A1(n20722), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20335) );
  INV_X1 U14679 ( .A(n20356), .ZN(n11700) );
  NOR3_X1 U14680 ( .A1(n20722), .A2(n20474), .A3(n20412), .ZN(n20591) );
  INV_X1 U14681 ( .A(n20591), .ZN(n20581) );
  AOI21_X1 U14682 ( .B1(n20722), .B2(n11700), .A(n20634), .ZN(n20361) );
  AOI22_X1 U14683 ( .A1(n11701), .A2(n20361), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15667), .ZN(n11702) );
  AOI22_X1 U14684 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14685 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14686 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14687 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U14688 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n11714) );
  AOI22_X1 U14689 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14690 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14691 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14692 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U14693 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11713) );
  AOI22_X1 U14694 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12272), .B2(n12340), .ZN(n11715) );
  INV_X1 U14695 ( .A(n11717), .ZN(n11718) );
  INV_X1 U14696 ( .A(n20108), .ZN(n20250) );
  NAND2_X1 U14697 ( .A1(n11718), .A2(n20250), .ZN(n11719) );
  NAND2_X1 U14698 ( .A1(n11748), .A2(n11719), .ZN(n20710) );
  INV_X1 U14699 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11724) );
  INV_X1 U14700 ( .A(n11720), .ZN(n11722) );
  INV_X1 U14701 ( .A(n11745), .ZN(n11721) );
  OAI21_X1 U14702 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11722), .A(
        n11721), .ZN(n14386) );
  AOI22_X1 U14703 ( .A1(n11674), .A2(n14386), .B1(n12241), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11723) );
  OAI21_X1 U14704 ( .B1(n12146), .B2(n11724), .A(n11723), .ZN(n11725) );
  AOI21_X1 U14705 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11726), .A(
        n11725), .ZN(n11727) );
  NAND2_X1 U14706 ( .A1(n13566), .A2(n13567), .ZN(n13565) );
  INV_X1 U14707 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14708 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11733) );
  INV_X1 U14709 ( .A(n11729), .ZN(n11806) );
  AOI22_X1 U14710 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14711 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14712 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14713 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11739) );
  AOI22_X1 U14714 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14715 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14716 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14717 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14718 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11738) );
  NAND2_X1 U14719 ( .A1(n12272), .A2(n12351), .ZN(n11740) );
  XNOR2_X1 U14720 ( .A(n11748), .B(n11749), .ZN(n12339) );
  NAND2_X1 U14721 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14722 ( .A1(n12242), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11742) );
  OAI211_X1 U14723 ( .C1(n11744), .C2(n16086), .A(n11743), .B(n11742), .ZN(
        n11746) );
  OAI21_X1 U14724 ( .B1(n11745), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11767), .ZN(n14371) );
  MUX2_X1 U14725 ( .A(n11746), .B(n14371), .S(n12209), .Z(n11747) );
  AOI21_X1 U14726 ( .B1(n12339), .B2(n11830), .A(n11747), .ZN(n13670) );
  NOR2_X2 U14727 ( .A1(n13565), .A2(n13670), .ZN(n13671) );
  NAND2_X1 U14728 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11762) );
  AOI22_X1 U14729 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14730 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14731 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14732 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U14733 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n11760) );
  AOI22_X1 U14734 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14735 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14736 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14737 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14738 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11759) );
  NAND2_X1 U14739 ( .A1(n12272), .A2(n12359), .ZN(n11761) );
  NAND2_X1 U14740 ( .A1(n11762), .A2(n11761), .ZN(n11763) );
  INV_X1 U14741 ( .A(n11763), .ZN(n11764) );
  NAND2_X1 U14742 ( .A1(n11765), .A2(n11764), .ZN(n11766) );
  INV_X1 U14743 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11771) );
  INV_X1 U14744 ( .A(n11767), .ZN(n11769) );
  INV_X1 U14745 ( .A(n11786), .ZN(n11768) );
  OAI21_X1 U14746 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11769), .A(
        n11768), .ZN(n19970) );
  AOI22_X1 U14747 ( .A1(n11674), .A2(n19970), .B1(n12241), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11770) );
  OAI21_X1 U14748 ( .B1(n12146), .B2(n11771), .A(n11770), .ZN(n11772) );
  NAND2_X1 U14749 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11784) );
  AOI22_X1 U14750 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14751 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14752 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14753 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11774) );
  NAND4_X1 U14754 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11783) );
  AOI22_X1 U14755 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14756 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14757 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14758 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11778) );
  NAND4_X1 U14759 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11782) );
  NAND2_X1 U14760 ( .A1(n12272), .A2(n12368), .ZN(n11793) );
  AND2_X1 U14761 ( .A1(n11784), .A2(n11793), .ZN(n11785) );
  NAND2_X1 U14762 ( .A1(n11794), .A2(n11785), .ZN(n12358) );
  NAND2_X1 U14763 ( .A1(n12358), .A2(n11830), .ZN(n11792) );
  OAI21_X1 U14764 ( .B1(n11786), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11798), .ZN(n19953) );
  AND2_X1 U14765 ( .A1(n19953), .A2(n12209), .ZN(n11790) );
  INV_X1 U14766 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11788) );
  INV_X1 U14767 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11787) );
  OAI22_X1 U14768 ( .A1(n12146), .A2(n11788), .B1(n11935), .B2(n11787), .ZN(
        n11789) );
  NOR2_X1 U14769 ( .A1(n11790), .A2(n11789), .ZN(n11791) );
  NAND2_X1 U14770 ( .A1(n11792), .A2(n11791), .ZN(n13772) );
  AND2_X2 U14771 ( .A1(n13706), .A2(n13772), .ZN(n13786) );
  INV_X1 U14772 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U14773 ( .A1(n12272), .A2(n12377), .ZN(n11795) );
  OAI21_X1 U14774 ( .B1(n12281), .B2(n11796), .A(n11795), .ZN(n11797) );
  NAND2_X1 U14775 ( .A1(n12372), .A2(n11830), .ZN(n11804) );
  OAI21_X1 U14776 ( .B1(n11799), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11820), .ZN(n19950) );
  INV_X1 U14777 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11801) );
  INV_X1 U14778 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11800) );
  OAI22_X1 U14779 ( .A1(n12146), .A2(n11801), .B1(n11935), .B2(n11800), .ZN(
        n11802) );
  AOI21_X1 U14780 ( .B1(n19950), .B2(n11674), .A(n11802), .ZN(n11803) );
  NAND2_X1 U14781 ( .A1(n11804), .A2(n11803), .ZN(n13785) );
  INV_X1 U14782 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11805) );
  XNOR2_X1 U14783 ( .A(n11820), .B(n11805), .ZN(n13842) );
  NAND2_X1 U14784 ( .A1(n13842), .A2(n11674), .ZN(n11819) );
  AOI22_X1 U14785 ( .A1(n12242), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n12241), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14786 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14787 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14788 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14789 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11807) );
  NAND4_X1 U14790 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11816) );
  AOI22_X1 U14791 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14792 ( .A1(n12193), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14793 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14794 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11811) );
  NAND4_X1 U14795 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11815) );
  OAI21_X1 U14796 ( .B1(n11816), .B2(n11815), .A(n11830), .ZN(n11817) );
  XOR2_X1 U14797 ( .A(n13976), .B(n11839), .Z(n14000) );
  INV_X1 U14798 ( .A(n14000), .ZN(n11837) );
  AOI22_X1 U14799 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14800 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14801 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14802 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11822) );
  NAND4_X1 U14803 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11832) );
  AOI22_X1 U14804 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11500), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14805 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14806 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14807 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U14808 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11831) );
  OAI21_X1 U14809 ( .B1(n11832), .B2(n11831), .A(n11830), .ZN(n11835) );
  NAND2_X1 U14810 ( .A1(n12242), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U14811 ( .A1(n12241), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11833) );
  NAND3_X1 U14812 ( .A1(n11835), .A2(n11834), .A3(n11833), .ZN(n11836) );
  XNOR2_X1 U14813 ( .A(n11856), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14694) );
  NAND2_X1 U14814 ( .A1(n14694), .A2(n11674), .ZN(n11855) );
  INV_X1 U14815 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14033) );
  INV_X1 U14816 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11840) );
  OAI22_X1 U14817 ( .A1(n12146), .A2(n14033), .B1(n11935), .B2(n11840), .ZN(
        n11853) );
  AOI22_X1 U14818 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14819 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14820 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14821 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11841) );
  NAND4_X1 U14822 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11850) );
  AOI22_X1 U14823 ( .A1(n11500), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14824 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14825 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14826 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14827 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11849) );
  NOR2_X1 U14828 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NOR2_X1 U14829 ( .A1(n11939), .A2(n11851), .ZN(n11852) );
  NOR2_X1 U14830 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  INV_X1 U14831 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14054) );
  OAI21_X1 U14832 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11857), .A(
        n11896), .ZN(n15882) );
  AOI22_X1 U14833 ( .A1(n11674), .A2(n15882), .B1(n12241), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11858) );
  OAI21_X1 U14834 ( .B1(n12146), .B2(n14054), .A(n11858), .ZN(n14343) );
  AOI22_X1 U14835 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14836 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14837 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14838 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11859) );
  NAND4_X1 U14839 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11868) );
  AOI22_X1 U14840 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14841 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14842 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14843 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11863) );
  NAND4_X1 U14844 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11867) );
  NOR2_X1 U14845 ( .A1(n11868), .A2(n11867), .ZN(n11869) );
  NOR2_X1 U14846 ( .A1(n11939), .A2(n11869), .ZN(n14043) );
  AOI22_X1 U14847 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14848 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14849 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14850 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11871) );
  NAND4_X1 U14851 ( .A1(n11874), .A2(n11873), .A3(n11872), .A4(n11871), .ZN(
        n11880) );
  AOI22_X1 U14852 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14853 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14854 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14855 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U14856 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n11879) );
  NOR2_X1 U14857 ( .A1(n11880), .A2(n11879), .ZN(n11885) );
  NAND2_X1 U14858 ( .A1(n12242), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11884) );
  INV_X1 U14859 ( .A(n11934), .ZN(n11881) );
  OAI21_X1 U14860 ( .B1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n11882), .A(
        n11881), .ZN(n14673) );
  AOI22_X1 U14861 ( .A1(n11674), .A2(n14673), .B1(n12241), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11883) );
  OAI211_X1 U14862 ( .C1(n11885), .C2(n11939), .A(n11884), .B(n11883), .ZN(
        n14344) );
  OAI21_X1 U14863 ( .B1(n14343), .B2(n14043), .A(n14344), .ZN(n11904) );
  AOI22_X1 U14864 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14865 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14866 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U14867 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11886) );
  NAND4_X1 U14868 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11895) );
  AOI22_X1 U14869 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14870 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14871 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14872 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11890) );
  NAND4_X1 U14873 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11894) );
  NOR2_X1 U14874 ( .A1(n11895), .A2(n11894), .ZN(n11901) );
  NAND2_X1 U14875 ( .A1(n20780), .A2(n11896), .ZN(n11898) );
  AND2_X1 U14876 ( .A1(n11898), .A2(n11897), .ZN(n15870) );
  OAI22_X1 U14877 ( .A1(n15870), .A2(n12240), .B1(n11935), .B2(n20780), .ZN(
        n11899) );
  INV_X1 U14878 ( .A(n11899), .ZN(n11900) );
  OAI21_X1 U14879 ( .B1(n11939), .B2(n11901), .A(n11900), .ZN(n11903) );
  INV_X1 U14880 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14570) );
  NOR2_X1 U14881 ( .A1(n12146), .A2(n14570), .ZN(n11902) );
  NOR2_X1 U14882 ( .A1(n11903), .A2(n11902), .ZN(n14490) );
  AOI22_X1 U14883 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14884 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14885 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12194), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14886 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11907) );
  NAND4_X1 U14887 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11917) );
  AOI22_X1 U14888 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14889 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12223), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14890 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12068), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14891 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12224), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U14892 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  NOR2_X1 U14893 ( .A1(n11917), .A2(n11916), .ZN(n11920) );
  XOR2_X1 U14894 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11934), .Z(
        n15861) );
  INV_X1 U14895 ( .A(n15861), .ZN(n11918) );
  AOI22_X1 U14896 ( .A1(n12241), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11674), .B2(n11918), .ZN(n11919) );
  OAI21_X1 U14897 ( .B1(n11939), .B2(n11920), .A(n11919), .ZN(n11922) );
  INV_X1 U14898 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14050) );
  NOR2_X1 U14899 ( .A1(n12146), .A2(n14050), .ZN(n11921) );
  NOR2_X1 U14900 ( .A1(n11922), .A2(n11921), .ZN(n14035) );
  AOI22_X1 U14901 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14902 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14903 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U14904 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U14905 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11933) );
  AOI22_X1 U14906 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14907 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14908 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U14909 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U14910 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11932) );
  NOR2_X1 U14911 ( .A1(n11933), .A2(n11932), .ZN(n11940) );
  NAND2_X1 U14912 ( .A1(n12242), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11938) );
  XNOR2_X1 U14913 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11956), .ZN(
        n15791) );
  OAI22_X1 U14914 ( .A1(n15791), .A2(n12240), .B1(n11935), .B2(n14669), .ZN(
        n11936) );
  INV_X1 U14915 ( .A(n11936), .ZN(n11937) );
  OAI211_X1 U14916 ( .C1(n11940), .C2(n11939), .A(n11938), .B(n11937), .ZN(
        n14475) );
  AOI22_X1 U14917 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U14918 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U14919 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14920 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U14921 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11951) );
  AOI22_X1 U14922 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U14923 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14924 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U14925 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U14926 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11950) );
  NOR2_X1 U14927 ( .A1(n11951), .A2(n11950), .ZN(n11955) );
  INV_X1 U14928 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14558) );
  NAND2_X1 U14929 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11952) );
  OAI211_X1 U14930 ( .C1(n12146), .C2(n14558), .A(n12240), .B(n11952), .ZN(
        n11953) );
  INV_X1 U14931 ( .A(n11953), .ZN(n11954) );
  OAI21_X1 U14932 ( .B1(n12237), .B2(n11955), .A(n11954), .ZN(n11959) );
  OAI21_X1 U14933 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11957), .A(
        n11989), .ZN(n15854) );
  OR2_X1 U14934 ( .A1(n12240), .A2(n15854), .ZN(n11958) );
  AOI22_X1 U14935 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U14936 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U14937 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U14938 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U14939 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11969) );
  AOI22_X1 U14940 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U14941 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U14942 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U14943 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U14944 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11968) );
  OR2_X1 U14945 ( .A1(n11969), .A2(n11968), .ZN(n11973) );
  INV_X1 U14946 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14553) );
  INV_X1 U14947 ( .A(n11989), .ZN(n11970) );
  XNOR2_X1 U14948 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11970), .ZN(
        n14656) );
  AOI22_X1 U14949 ( .A1(n11674), .A2(n14656), .B1(n12241), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11971) );
  OAI21_X1 U14950 ( .B1(n12146), .B2(n14553), .A(n11971), .ZN(n11972) );
  AOI21_X1 U14951 ( .B1(n12206), .B2(n11973), .A(n11972), .ZN(n14330) );
  AOI22_X1 U14952 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U14953 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U14954 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U14955 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11974) );
  NAND4_X1 U14956 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n11983) );
  AOI22_X1 U14957 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U14958 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U14959 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U14960 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U14961 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n11982) );
  NOR2_X1 U14962 ( .A1(n11983), .A2(n11982), .ZN(n11987) );
  INV_X1 U14963 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U14964 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11984) );
  OAI211_X1 U14965 ( .C1(n12146), .C2(n14549), .A(n12240), .B(n11984), .ZN(
        n11985) );
  INV_X1 U14966 ( .A(n11985), .ZN(n11986) );
  OAI21_X1 U14967 ( .B1(n12237), .B2(n11987), .A(n11986), .ZN(n11992) );
  OAI21_X1 U14968 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11990), .A(
        n12024), .ZN(n15764) );
  OR2_X1 U14969 ( .A1(n12240), .A2(n15764), .ZN(n11991) );
  NAND2_X1 U14970 ( .A1(n11992), .A2(n11991), .ZN(n14453) );
  AOI22_X1 U14971 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U14972 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U14973 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U14974 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11994) );
  NAND4_X1 U14975 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n12003) );
  AOI22_X1 U14976 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U14977 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U14978 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U14979 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U14980 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12002) );
  NOR2_X1 U14981 ( .A1(n12003), .A2(n12002), .ZN(n12006) );
  OAI21_X1 U14982 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14637), .A(n12240), 
        .ZN(n12004) );
  AOI21_X1 U14983 ( .B1(n12242), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12004), .ZN(
        n12005) );
  OAI21_X1 U14984 ( .B1(n12237), .B2(n12006), .A(n12005), .ZN(n12008) );
  XNOR2_X1 U14985 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12024), .ZN(
        n14639) );
  NAND2_X1 U14986 ( .A1(n11674), .A2(n14639), .ZN(n12007) );
  AOI22_X1 U14987 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14988 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U14989 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U14990 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12010) );
  NAND4_X1 U14991 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12019) );
  AOI22_X1 U14992 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U14993 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U14994 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U14995 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U14996 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  NOR2_X1 U14997 ( .A1(n12019), .A2(n12018), .ZN(n12023) );
  INV_X1 U14998 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U14999 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12020) );
  OAI211_X1 U15000 ( .C1(n12146), .C2(n14542), .A(n12240), .B(n12020), .ZN(
        n12021) );
  INV_X1 U15001 ( .A(n12021), .ZN(n12022) );
  OAI21_X1 U15002 ( .B1(n12237), .B2(n12023), .A(n12022), .ZN(n12027) );
  OAI21_X1 U15003 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12025), .A(
        n12058), .ZN(n15750) );
  OR2_X1 U15004 ( .A1(n12240), .A2(n15750), .ZN(n12026) );
  AOI22_X1 U15005 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15006 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15007 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15008 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U15009 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12037) );
  AOI22_X1 U15010 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15011 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15012 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15013 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12032) );
  NAND4_X1 U15014 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12036) );
  NOR2_X1 U15015 ( .A1(n12037), .A2(n12036), .ZN(n12040) );
  OAI21_X1 U15016 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n12057), .A(n12240), 
        .ZN(n12038) );
  AOI21_X1 U15017 ( .B1(n12242), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12038), .ZN(
        n12039) );
  OAI21_X1 U15018 ( .B1(n12237), .B2(n12040), .A(n12039), .ZN(n12042) );
  XNOR2_X1 U15019 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12058), .ZN(
        n15841) );
  NAND2_X1 U15020 ( .A1(n15841), .A2(n11674), .ZN(n12041) );
  NAND2_X1 U15021 ( .A1(n12042), .A2(n12041), .ZN(n14443) );
  AOI22_X1 U15022 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15023 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12068), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15024 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12194), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15025 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15026 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12052) );
  AOI22_X1 U15027 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11806), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15028 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15029 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15030 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12224), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15031 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  NOR2_X1 U15032 ( .A1(n12052), .A2(n12051), .ZN(n12056) );
  INV_X1 U15033 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U15034 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12053) );
  OAI211_X1 U15035 ( .C1(n12146), .C2(n14534), .A(n12240), .B(n12053), .ZN(
        n12054) );
  INV_X1 U15036 ( .A(n12054), .ZN(n12055) );
  OAI21_X1 U15037 ( .B1(n12237), .B2(n12056), .A(n12055), .ZN(n12061) );
  OAI21_X1 U15038 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12059), .A(
        n12109), .ZN(n15840) );
  OR2_X1 U15039 ( .A1(n12240), .A2(n15840), .ZN(n12060) );
  NAND2_X1 U15040 ( .A1(n12061), .A2(n12060), .ZN(n14436) );
  AOI22_X1 U15041 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15042 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15043 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15044 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12064) );
  NAND4_X1 U15045 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12075) );
  AOI22_X1 U15046 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15047 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15048 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15049 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12070) );
  NAND4_X1 U15050 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12074) );
  NOR2_X1 U15051 ( .A1(n12075), .A2(n12074), .ZN(n12094) );
  AOI22_X1 U15052 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15053 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15054 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15055 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15056 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12085) );
  AOI22_X1 U15057 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15058 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15059 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15060 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U15061 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12084) );
  NOR2_X1 U15062 ( .A1(n12085), .A2(n12084), .ZN(n12093) );
  XOR2_X1 U15063 ( .A(n12094), .B(n12093), .Z(n12086) );
  NAND2_X1 U15064 ( .A1(n12086), .A2(n12206), .ZN(n12090) );
  INV_X1 U15065 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14530) );
  INV_X1 U15066 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20535) );
  OAI21_X1 U15067 ( .B1(n20535), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n11673), .ZN(n12087) );
  OAI21_X1 U15068 ( .B1(n12146), .B2(n14530), .A(n12087), .ZN(n12088) );
  INV_X1 U15069 ( .A(n12088), .ZN(n12089) );
  NAND2_X1 U15070 ( .A1(n12090), .A2(n12089), .ZN(n12092) );
  XNOR2_X1 U15071 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12109), .ZN(
        n15719) );
  NAND2_X1 U15072 ( .A1(n11674), .A2(n15719), .ZN(n12091) );
  NAND2_X1 U15073 ( .A1(n12092), .A2(n12091), .ZN(n14430) );
  NOR2_X1 U15074 ( .A1(n12094), .A2(n12093), .ZN(n12115) );
  AOI22_X1 U15075 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15076 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15077 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15078 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15079 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12104) );
  AOI22_X1 U15080 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15081 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15082 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15083 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15084 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  OR2_X1 U15085 ( .A1(n12104), .A2(n12103), .ZN(n12114) );
  INV_X1 U15086 ( .A(n12114), .ZN(n12105) );
  XNOR2_X1 U15087 ( .A(n12115), .B(n12105), .ZN(n12106) );
  NAND2_X1 U15088 ( .A1(n12106), .A2(n12206), .ZN(n12113) );
  INV_X1 U15089 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14525) );
  NAND2_X1 U15090 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12107) );
  OAI211_X1 U15091 ( .C1(n12146), .C2(n14525), .A(n12240), .B(n12107), .ZN(
        n12108) );
  INV_X1 U15092 ( .A(n12108), .ZN(n12112) );
  INV_X1 U15093 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15729) );
  OAI21_X1 U15094 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12110), .A(
        n12149), .ZN(n15833) );
  NOR2_X1 U15095 ( .A1(n15833), .A2(n12240), .ZN(n12111) );
  AOI21_X1 U15096 ( .B1(n12113), .B2(n12112), .A(n12111), .ZN(n14422) );
  NAND2_X1 U15097 ( .A1(n12115), .A2(n12114), .ZN(n12132) );
  AOI22_X1 U15098 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15099 ( .A1(n12193), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15100 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15101 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15102 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12125) );
  AOI22_X1 U15103 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15104 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15105 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15106 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15107 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  NOR2_X1 U15108 ( .A1(n12125), .A2(n12124), .ZN(n12133) );
  XOR2_X1 U15109 ( .A(n12132), .B(n12133), .Z(n12126) );
  NAND2_X1 U15110 ( .A1(n12126), .A2(n12206), .ZN(n12129) );
  INV_X1 U15111 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14620) );
  OAI21_X1 U15112 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14620), .A(n12240), 
        .ZN(n12127) );
  AOI21_X1 U15113 ( .B1(n12242), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12127), .ZN(
        n12128) );
  NAND2_X1 U15114 ( .A1(n12129), .A2(n12128), .ZN(n12131) );
  XNOR2_X1 U15115 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12149), .ZN(
        n14622) );
  NAND2_X1 U15116 ( .A1(n11674), .A2(n14622), .ZN(n12130) );
  NAND2_X1 U15117 ( .A1(n12131), .A2(n12130), .ZN(n14306) );
  NOR2_X1 U15118 ( .A1(n12133), .A2(n12132), .ZN(n12154) );
  AOI22_X1 U15119 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15120 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15121 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15122 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12134) );
  NAND4_X1 U15123 ( .A1(n12137), .A2(n12136), .A3(n12135), .A4(n12134), .ZN(
        n12143) );
  AOI22_X1 U15124 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15125 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15126 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15127 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U15128 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12142) );
  OR2_X1 U15129 ( .A1(n12143), .A2(n12142), .ZN(n12153) );
  INV_X1 U15130 ( .A(n12153), .ZN(n12144) );
  XNOR2_X1 U15131 ( .A(n12154), .B(n12144), .ZN(n12148) );
  INV_X1 U15132 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U15133 ( .A1(n11673), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12145) );
  OAI211_X1 U15134 ( .C1(n12146), .C2(n14517), .A(n12240), .B(n12145), .ZN(
        n12147) );
  AOI21_X1 U15135 ( .B1(n12148), .B2(n12206), .A(n12147), .ZN(n12152) );
  OAI21_X1 U15136 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n12150), .A(
        n12170), .ZN(n15825) );
  NOR2_X1 U15137 ( .A1(n15825), .A2(n12240), .ZN(n12151) );
  NAND2_X1 U15138 ( .A1(n12154), .A2(n12153), .ZN(n12175) );
  AOI22_X1 U15139 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15140 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15141 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15142 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15143 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12165) );
  AOI22_X1 U15144 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15145 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15146 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15147 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U15148 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12164) );
  NOR2_X1 U15149 ( .A1(n12165), .A2(n12164), .ZN(n12176) );
  XOR2_X1 U15150 ( .A(n12175), .B(n12176), .Z(n12166) );
  NAND2_X1 U15151 ( .A1(n12166), .A2(n12206), .ZN(n12169) );
  INV_X1 U15152 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14609) );
  NOR2_X1 U15153 ( .A1(n14609), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12167) );
  AOI211_X1 U15154 ( .C1(n12242), .C2(P1_EAX_REG_27__SCAN_IN), .A(n11674), .B(
        n12167), .ZN(n12168) );
  XNOR2_X1 U15155 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B(n12170), .ZN(
        n14613) );
  AOI22_X1 U15156 ( .A1(n12169), .A2(n12168), .B1(n11674), .B2(n14613), .ZN(
        n14296) );
  INV_X1 U15157 ( .A(n12170), .ZN(n12171) );
  INV_X1 U15158 ( .A(n12172), .ZN(n12173) );
  INV_X1 U15159 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U15160 ( .A1(n12173), .A2(n14287), .ZN(n12174) );
  NAND2_X1 U15161 ( .A1(n12212), .A2(n12174), .ZN(n14602) );
  NOR2_X1 U15162 ( .A1(n12176), .A2(n12175), .ZN(n12192) );
  AOI22_X1 U15163 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15164 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15165 ( .A1(n12222), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15166 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12177) );
  NAND4_X1 U15167 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(
        n12186) );
  AOI22_X1 U15168 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15169 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15170 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15171 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12181) );
  NAND4_X1 U15172 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12185) );
  OR2_X1 U15173 ( .A1(n12186), .A2(n12185), .ZN(n12191) );
  XNOR2_X1 U15174 ( .A(n12192), .B(n12191), .ZN(n12189) );
  AOI21_X1 U15175 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11673), .A(
        n11674), .ZN(n12188) );
  NAND2_X1 U15176 ( .A1(n12242), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12187) );
  OAI211_X1 U15177 ( .C1(n12189), .C2(n12237), .A(n12188), .B(n12187), .ZN(
        n12190) );
  OAI21_X1 U15178 ( .B1(n12240), .B2(n14602), .A(n12190), .ZN(n14286) );
  NAND2_X1 U15179 ( .A1(n12192), .A2(n12191), .ZN(n12231) );
  AOI22_X1 U15180 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12221), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15181 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15182 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12068), .B1(
        n12194), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15183 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12224), .B1(
        n11490), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12195) );
  NAND4_X1 U15184 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12195), .ZN(
        n12205) );
  AOI22_X1 U15185 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9655), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15186 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15187 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15188 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U15189 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12204) );
  NOR2_X1 U15190 ( .A1(n12205), .A2(n12204), .ZN(n12232) );
  XOR2_X1 U15191 ( .A(n12231), .B(n12232), .Z(n12207) );
  NAND2_X1 U15192 ( .A1(n12207), .A2(n12206), .ZN(n12211) );
  INV_X1 U15193 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14583) );
  AOI21_X1 U15194 ( .B1(n14583), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12208) );
  AOI21_X1 U15195 ( .B1(n12242), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12208), .ZN(
        n12210) );
  XNOR2_X1 U15196 ( .A(n12212), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14585) );
  AOI22_X1 U15197 ( .A1(n12211), .A2(n12210), .B1(n12209), .B2(n14585), .ZN(
        n14271) );
  INV_X1 U15198 ( .A(n12212), .ZN(n12213) );
  NAND2_X1 U15199 ( .A1(n12213), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12303) );
  XOR2_X1 U15200 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12303), .Z(
        n14578) );
  AOI22_X1 U15201 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12193), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15202 ( .A1(n9655), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15203 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9658), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15204 ( .A1(n11490), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11474), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15205 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12230) );
  AOI22_X1 U15206 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15207 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12222), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15208 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15209 ( .A1(n12194), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12069), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15210 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  NOR2_X1 U15211 ( .A1(n12230), .A2(n12229), .ZN(n12234) );
  NOR2_X1 U15212 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  XOR2_X1 U15213 ( .A(n12234), .B(n12233), .Z(n12238) );
  AOI21_X1 U15214 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n11673), .A(
        n11674), .ZN(n12236) );
  NAND2_X1 U15215 ( .A1(n12242), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12235) );
  OAI211_X1 U15216 ( .C1(n12238), .C2(n12237), .A(n12236), .B(n12235), .ZN(
        n12239) );
  OAI21_X1 U15217 ( .B1(n12240), .B2(n14578), .A(n12239), .ZN(n14260) );
  AOI22_X1 U15218 ( .A1(n12242), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12241), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12243) );
  NOR2_X2 U15219 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20718) );
  NOR2_X1 U15220 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20643), .ZN(n15673) );
  NAND2_X1 U15221 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n15673), .ZN(n16090) );
  INV_X1 U15222 ( .A(n16090), .ZN(n12244) );
  XNOR2_X1 U15223 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12266) );
  NAND2_X1 U15224 ( .A1(n12267), .A2(n12266), .ZN(n12246) );
  NAND2_X1 U15225 ( .A1(n20412), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12245) );
  NAND2_X1 U15226 ( .A1(n12246), .A2(n12245), .ZN(n12257) );
  XNOR2_X1 U15227 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U15228 ( .A1(n12257), .A2(n12256), .ZN(n12248) );
  NAND2_X1 U15229 ( .A1(n20474), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12247) );
  NAND2_X1 U15230 ( .A1(n12248), .A2(n12247), .ZN(n12255) );
  XNOR2_X1 U15231 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12254) );
  NAND2_X1 U15232 ( .A1(n12255), .A2(n12254), .ZN(n12250) );
  NAND2_X1 U15233 ( .A1(n20722), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12249) );
  NAND2_X1 U15234 ( .A1(n12250), .A2(n12249), .ZN(n12284) );
  NOR2_X1 U15235 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16086), .ZN(
        n12251) );
  NAND2_X1 U15236 ( .A1(n12413), .A2(n12272), .ZN(n12292) );
  XNOR2_X1 U15237 ( .A(n12255), .B(n12254), .ZN(n12410) );
  XNOR2_X1 U15238 ( .A(n12257), .B(n12256), .ZN(n12409) );
  INV_X1 U15239 ( .A(n12409), .ZN(n12258) );
  NAND2_X1 U15240 ( .A1(n20139), .A2(n13402), .ZN(n12259) );
  NAND2_X1 U15241 ( .A1(n12259), .A2(n20124), .ZN(n12279) );
  INV_X1 U15242 ( .A(n12279), .ZN(n12260) );
  AOI211_X1 U15243 ( .C1(n12288), .C2(n12409), .A(n12278), .B(n12260), .ZN(
        n12280) );
  INV_X1 U15244 ( .A(n12272), .ZN(n12268) );
  INV_X1 U15245 ( .A(n12267), .ZN(n12261) );
  OAI21_X1 U15246 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20504), .A(
        n12261), .ZN(n12262) );
  NOR2_X1 U15247 ( .A1(n12268), .A2(n12262), .ZN(n12265) );
  INV_X1 U15248 ( .A(n12262), .ZN(n12263) );
  OAI211_X1 U15249 ( .C1(n20107), .C2(n13088), .A(n12263), .B(n12279), .ZN(
        n12264) );
  OAI21_X1 U15250 ( .B1(n12283), .B2(n12265), .A(n12264), .ZN(n12273) );
  INV_X1 U15251 ( .A(n12273), .ZN(n12277) );
  XNOR2_X1 U15252 ( .A(n12267), .B(n12266), .ZN(n12408) );
  NAND2_X1 U15253 ( .A1(n20139), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12270) );
  OAI21_X1 U15254 ( .B1(n20124), .B2(n12268), .A(n12270), .ZN(n12269) );
  AOI21_X1 U15255 ( .B1(n12288), .B2(n12408), .A(n12269), .ZN(n12274) );
  INV_X1 U15256 ( .A(n12274), .ZN(n12276) );
  NAND2_X1 U15257 ( .A1(n12270), .A2(n13422), .ZN(n12271) );
  AOI22_X1 U15258 ( .A1(n12408), .A2(n12285), .B1(n12274), .B2(n12273), .ZN(
        n12275) );
  NAND2_X1 U15259 ( .A1(n12281), .A2(n12410), .ZN(n12282) );
  INV_X1 U15260 ( .A(n12286), .ZN(n12411) );
  NAND3_X1 U15261 ( .A1(n12288), .A2(n12287), .A3(n12411), .ZN(n12289) );
  AOI21_X1 U15262 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20644), .A(
        n12290), .ZN(n12291) );
  NAND2_X1 U15263 ( .A1(n12294), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19913) );
  OR2_X1 U15264 ( .A1(n12295), .A2(n11556), .ZN(n12298) );
  INV_X1 U15265 ( .A(n12296), .ZN(n12297) );
  AND2_X1 U15266 ( .A1(n12298), .A2(n12297), .ZN(n13403) );
  NAND2_X1 U15267 ( .A1(n11557), .A2(n20107), .ZN(n12299) );
  NAND2_X1 U15268 ( .A1(n13277), .A2(n12300), .ZN(n15658) );
  AND2_X1 U15269 ( .A1(n20590), .A2(n12305), .ZN(n20734) );
  OR2_X1 U15270 ( .A1(n20734), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12301) );
  NAND2_X1 U15271 ( .A1(n20644), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15666) );
  NAND2_X1 U15272 ( .A1(n20535), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U15273 ( .A1(n15666), .A2(n12302), .ZN(n20067) );
  INV_X1 U15274 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14262) );
  NOR2_X1 U15275 ( .A1(n12303), .A2(n14262), .ZN(n12304) );
  XNOR2_X1 U15276 ( .A(n12304), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13840) );
  INV_X2 U15277 ( .A(n16057), .ZN(n20074) );
  NAND2_X1 U15278 ( .A1(n20074), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14712) );
  NAND2_X1 U15279 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12306) );
  OAI211_X1 U15280 ( .C1(n15899), .C2(n13840), .A(n14712), .B(n12306), .ZN(
        n12307) );
  AOI21_X1 U15281 ( .B1(n14216), .B2(n15894), .A(n12307), .ZN(n12406) );
  INV_X1 U15282 ( .A(n12378), .ZN(n13086) );
  NAND2_X1 U15283 ( .A1(n20107), .A2(n12418), .ZN(n12324) );
  OAI21_X1 U15284 ( .B1(n20739), .B2(n12320), .A(n12324), .ZN(n12308) );
  INV_X1 U15285 ( .A(n12308), .ZN(n12309) );
  NAND2_X1 U15286 ( .A1(n20064), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12315) );
  XNOR2_X1 U15287 ( .A(n12321), .B(n12320), .ZN(n12311) );
  OAI211_X1 U15288 ( .C1(n12311), .C2(n20739), .A(n13081), .B(n11548), .ZN(
        n12312) );
  INV_X1 U15289 ( .A(n12312), .ZN(n12313) );
  NAND2_X1 U15290 ( .A1(n13377), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12318) );
  INV_X1 U15291 ( .A(n12315), .ZN(n20065) );
  NAND2_X1 U15292 ( .A1(n20065), .A2(n12316), .ZN(n12317) );
  INV_X1 U15293 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20082) );
  NAND2_X1 U15294 ( .A1(n9672), .A2(n12378), .ZN(n12328) );
  NAND2_X1 U15295 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  NAND2_X1 U15296 ( .A1(n12322), .A2(n12323), .ZN(n12341) );
  OAI21_X1 U15297 ( .B1(n12323), .B2(n12322), .A(n12341), .ZN(n12326) );
  INV_X1 U15298 ( .A(n12324), .ZN(n12325) );
  AOI21_X1 U15299 ( .B1(n12326), .B2(n13319), .A(n12325), .ZN(n12327) );
  NAND2_X1 U15300 ( .A1(n12328), .A2(n12327), .ZN(n13498) );
  NAND2_X1 U15301 ( .A1(n13499), .A2(n13498), .ZN(n12331) );
  NAND2_X1 U15302 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12330) );
  NAND2_X2 U15303 ( .A1(n12331), .A2(n12330), .ZN(n12336) );
  INV_X1 U15304 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13592) );
  OR2_X1 U15305 ( .A1(n20710), .A2(n13086), .ZN(n12335) );
  INV_X1 U15306 ( .A(n12340), .ZN(n12332) );
  XNOR2_X1 U15307 ( .A(n12341), .B(n12332), .ZN(n12333) );
  NAND2_X1 U15308 ( .A1(n12333), .A2(n13319), .ZN(n12334) );
  NAND2_X1 U15309 ( .A1(n12335), .A2(n12334), .ZN(n13589) );
  NAND2_X1 U15310 ( .A1(n13590), .A2(n13589), .ZN(n12338) );
  NAND2_X1 U15311 ( .A1(n12336), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12337) );
  NAND2_X1 U15312 ( .A1(n12338), .A2(n12337), .ZN(n13713) );
  NAND2_X1 U15313 ( .A1(n12339), .A2(n12378), .ZN(n12345) );
  AND2_X1 U15314 ( .A1(n12341), .A2(n12340), .ZN(n12352) );
  INV_X1 U15315 ( .A(n12351), .ZN(n12342) );
  XNOR2_X1 U15316 ( .A(n12352), .B(n12342), .ZN(n12343) );
  NAND2_X1 U15317 ( .A1(n12343), .A2(n13319), .ZN(n12344) );
  NAND2_X1 U15318 ( .A1(n12345), .A2(n12344), .ZN(n12347) );
  INV_X1 U15319 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12346) );
  XNOR2_X1 U15320 ( .A(n12347), .B(n12346), .ZN(n13714) );
  NAND2_X1 U15321 ( .A1(n13713), .A2(n13714), .ZN(n12349) );
  NAND2_X1 U15322 ( .A1(n12347), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12348) );
  NAND2_X2 U15323 ( .A1(n12349), .A2(n12348), .ZN(n15897) );
  NAND2_X1 U15324 ( .A1(n12352), .A2(n12351), .ZN(n12360) );
  XNOR2_X1 U15325 ( .A(n12359), .B(n12360), .ZN(n12353) );
  NAND2_X1 U15326 ( .A1(n13319), .A2(n12353), .ZN(n12354) );
  INV_X1 U15327 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15328 ( .A1(n12356), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12357) );
  NAND3_X1 U15329 ( .A1(n12382), .A2(n12358), .A3(n12378), .ZN(n12365) );
  INV_X1 U15330 ( .A(n12359), .ZN(n12361) );
  NOR2_X1 U15331 ( .A1(n12361), .A2(n12360), .ZN(n12369) );
  INV_X1 U15332 ( .A(n12369), .ZN(n12362) );
  XNOR2_X1 U15333 ( .A(n12368), .B(n12362), .ZN(n12363) );
  NAND2_X1 U15334 ( .A1(n13319), .A2(n12363), .ZN(n12364) );
  AND2_X1 U15335 ( .A1(n12365), .A2(n12364), .ZN(n12366) );
  INV_X1 U15336 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16050) );
  NAND2_X1 U15337 ( .A1(n12366), .A2(n16050), .ZN(n15891) );
  INV_X1 U15338 ( .A(n12366), .ZN(n12367) );
  NAND2_X1 U15339 ( .A1(n12367), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15890) );
  NAND2_X1 U15340 ( .A1(n12369), .A2(n12368), .ZN(n12383) );
  XNOR2_X1 U15341 ( .A(n12384), .B(n12383), .ZN(n12370) );
  NOR2_X1 U15342 ( .A1(n12370), .A2(n20739), .ZN(n12371) );
  AOI21_X1 U15343 ( .B1(n12372), .B2(n12378), .A(n12371), .ZN(n15884) );
  INV_X1 U15344 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15883) );
  NAND2_X1 U15345 ( .A1(n15884), .A2(n15883), .ZN(n12373) );
  NAND2_X1 U15346 ( .A1(n15886), .A2(n12373), .ZN(n12376) );
  INV_X1 U15347 ( .A(n15884), .ZN(n12374) );
  NAND2_X1 U15348 ( .A1(n12374), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12375) );
  NAND2_X2 U15349 ( .A1(n12376), .A2(n12375), .ZN(n13991) );
  NAND2_X1 U15350 ( .A1(n12378), .A2(n12377), .ZN(n12379) );
  NOR2_X1 U15351 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  INV_X4 U15352 ( .A(n12400), .ZN(n15858) );
  NOR2_X1 U15353 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  NAND2_X1 U15354 ( .A1(n12385), .A2(n13319), .ZN(n12386) );
  NAND2_X1 U15355 ( .A1(n15858), .A2(n12386), .ZN(n13989) );
  AND2_X1 U15356 ( .A1(n13989), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12387) );
  INV_X1 U15357 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16056) );
  INV_X1 U15358 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n20884) );
  INV_X1 U15359 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12395) );
  XNOR2_X1 U15360 ( .A(n15858), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14682) );
  INV_X1 U15361 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16021) );
  NAND2_X1 U15362 ( .A1(n15858), .A2(n16021), .ZN(n14681) );
  NAND2_X1 U15363 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12389) );
  NAND2_X1 U15364 ( .A1(n15858), .A2(n12389), .ZN(n14678) );
  AND2_X1 U15365 ( .A1(n14681), .A2(n14678), .ZN(n12390) );
  NAND2_X1 U15366 ( .A1(n14682), .A2(n12390), .ZN(n15855) );
  INV_X1 U15367 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12466) );
  AND2_X1 U15368 ( .A1(n15858), .A2(n12466), .ZN(n12391) );
  OR2_X2 U15369 ( .A1(n15855), .A2(n12391), .ZN(n14662) );
  INV_X1 U15370 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15983) );
  XNOR2_X1 U15371 ( .A(n15858), .B(n15983), .ZN(n15849) );
  INV_X1 U15372 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14690) );
  INV_X1 U15373 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15877) );
  NAND2_X1 U15374 ( .A1(n14690), .A2(n15877), .ZN(n12392) );
  NAND2_X1 U15375 ( .A1(n15874), .A2(n12392), .ZN(n14676) );
  NAND2_X1 U15376 ( .A1(n15874), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14680) );
  AND2_X1 U15377 ( .A1(n14676), .A2(n14680), .ZN(n15856) );
  OAI21_X1 U15378 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n15874), .ZN(n12394) );
  NAND2_X1 U15379 ( .A1(n15856), .A2(n12394), .ZN(n14663) );
  NOR2_X1 U15380 ( .A1(n15858), .A2(n12395), .ZN(n14665) );
  NOR2_X1 U15381 ( .A1(n14663), .A2(n14665), .ZN(n15847) );
  NOR2_X1 U15382 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12396) );
  XNOR2_X1 U15383 ( .A(n12393), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14645) );
  NAND2_X1 U15384 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14713) );
  INV_X1 U15385 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12399) );
  NOR2_X1 U15386 ( .A1(n14713), .A2(n12399), .ZN(n12397) );
  NAND2_X1 U15387 ( .A1(n12398), .A2(n12393), .ZN(n15835) );
  INV_X1 U15388 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15982) );
  INV_X1 U15389 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14066) );
  INV_X1 U15390 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14067) );
  NAND4_X1 U15391 ( .A1(n15982), .A2(n14066), .A3(n14067), .A4(n12399), .ZN(
        n12401) );
  OAI21_X1 U15392 ( .B1(n14644), .B2(n12401), .A(n12400), .ZN(n15834) );
  INV_X1 U15393 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15950) );
  INV_X1 U15394 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15940) );
  INV_X1 U15395 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14617) );
  NAND2_X1 U15396 ( .A1(n15940), .A2(n14617), .ZN(n14594) );
  NAND2_X1 U15397 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15923) );
  NOR2_X1 U15398 ( .A1(n15923), .A2(n14617), .ZN(n14700) );
  NAND2_X1 U15399 ( .A1(n14700), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12402) );
  OAI21_X1 U15400 ( .B1(n14615), .B2(n12402), .A(n12393), .ZN(n14606) );
  NAND2_X1 U15401 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15904) );
  INV_X1 U15402 ( .A(n15904), .ZN(n14729) );
  INV_X1 U15403 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14728) );
  NAND2_X1 U15404 ( .A1(n15874), .A2(n14728), .ZN(n14587) );
  NOR2_X1 U15405 ( .A1(n14587), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12403) );
  NAND2_X1 U15406 ( .A1(n15858), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14586) );
  NAND2_X1 U15407 ( .A1(n12404), .A2(n20070), .ZN(n12405) );
  NAND2_X1 U15408 ( .A1(n12406), .A2(n12405), .ZN(P1_U2968) );
  INV_X1 U15409 ( .A(n13410), .ZN(n12407) );
  NOR4_X1 U15410 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12412) );
  NOR2_X1 U15411 ( .A1(n12413), .A2(n12412), .ZN(n13383) );
  AND2_X1 U15412 ( .A1(n9735), .A2(n13383), .ZN(n13079) );
  NAND2_X1 U15413 ( .A1(n13079), .A2(n13578), .ZN(n13058) );
  NAND2_X1 U15414 ( .A1(n11673), .A2(n20643), .ZN(n16088) );
  INV_X1 U15415 ( .A(n16088), .ZN(n20737) );
  NAND2_X1 U15416 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20737), .ZN(n15669) );
  NAND2_X1 U15417 ( .A1(n11674), .A2(n15673), .ZN(n12414) );
  OAI211_X1 U15418 ( .C1(n15669), .C2(n20644), .A(n16057), .B(n12414), .ZN(
        n12415) );
  NOR2_X1 U15419 ( .A1(n13840), .A2(n20643), .ZN(n12417) );
  NAND2_X1 U15420 ( .A1(n14216), .A2(n19958), .ZN(n12540) );
  INV_X1 U15421 ( .A(n12418), .ZN(n20131) );
  NAND2_X1 U15422 ( .A1(n20131), .A2(n13402), .ZN(n12513) );
  INV_X1 U15423 ( .A(n12513), .ZN(n12419) );
  AND2_X1 U15424 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12420) );
  AOI21_X1 U15425 ( .B1(n13082), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12420), .ZN(
        n14257) );
  INV_X1 U15426 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n19983) );
  NAND2_X1 U15427 ( .A1(n12505), .A2(n19983), .ZN(n12426) );
  INV_X1 U15428 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12422) );
  NAND2_X1 U15429 ( .A1(n12513), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U15430 ( .A1(n13362), .A2(n19983), .ZN(n12423) );
  NAND3_X1 U15431 ( .A1(n12424), .A2(n12421), .A3(n12423), .ZN(n12425) );
  NAND2_X1 U15432 ( .A1(n12513), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12427) );
  OAI21_X1 U15433 ( .B1(n14256), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12427), .ZN(
        n13343) );
  XNOR2_X1 U15434 ( .A(n12428), .B(n13343), .ZN(n19982) );
  NAND2_X1 U15435 ( .A1(n19982), .A2(n13362), .ZN(n13364) );
  NAND2_X1 U15436 ( .A1(n13364), .A2(n12428), .ZN(n13569) );
  MUX2_X1 U15437 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12430) );
  OR2_X1 U15438 ( .A1(n13082), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12429) );
  AND2_X1 U15439 ( .A1(n12430), .A2(n12429), .ZN(n13570) );
  NAND2_X1 U15440 ( .A1(n12513), .A2(n20082), .ZN(n12432) );
  INV_X1 U15441 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n20007) );
  NAND2_X1 U15442 ( .A1(n13362), .A2(n20007), .ZN(n12431) );
  NAND3_X1 U15443 ( .A1(n12432), .A2(n12421), .A3(n12431), .ZN(n12434) );
  NAND2_X1 U15444 ( .A1(n12505), .A2(n20007), .ZN(n12433) );
  NAND2_X1 U15445 ( .A1(n12434), .A2(n12433), .ZN(n14395) );
  NAND2_X1 U15446 ( .A1(n13570), .A2(n14395), .ZN(n12435) );
  NAND2_X1 U15447 ( .A1(n12419), .A2(n13349), .ZN(n12461) );
  NAND2_X1 U15448 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12436) );
  AND2_X1 U15449 ( .A1(n12461), .A2(n12436), .ZN(n12438) );
  MUX2_X1 U15450 ( .A(n12518), .B(n12513), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12437) );
  NAND2_X1 U15451 ( .A1(n12438), .A2(n12437), .ZN(n13709) );
  INV_X1 U15452 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19965) );
  NAND2_X1 U15453 ( .A1(n12471), .A2(n19965), .ZN(n12441) );
  NAND2_X1 U15454 ( .A1(n13362), .A2(n19965), .ZN(n12439) );
  OAI211_X1 U15455 ( .C1(n14256), .C2(n12355), .A(n12513), .B(n12439), .ZN(
        n12440) );
  AND2_X1 U15456 ( .A1(n12441), .A2(n12440), .ZN(n13708) );
  NAND2_X1 U15457 ( .A1(n13709), .A2(n13708), .ZN(n12442) );
  NAND2_X1 U15458 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12443) );
  AND2_X1 U15459 ( .A1(n12461), .A2(n12443), .ZN(n12445) );
  MUX2_X1 U15460 ( .A(n12518), .B(n12513), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12444) );
  NAND2_X1 U15461 ( .A1(n12445), .A2(n12444), .ZN(n13775) );
  INV_X1 U15462 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19938) );
  NAND2_X1 U15463 ( .A1(n12471), .A2(n19938), .ZN(n12448) );
  NAND2_X1 U15464 ( .A1(n13362), .A2(n19938), .ZN(n12446) );
  OAI211_X1 U15465 ( .C1(n14256), .C2(n15883), .A(n12513), .B(n12446), .ZN(
        n12447) );
  NAND2_X1 U15466 ( .A1(n12448), .A2(n12447), .ZN(n13788) );
  MUX2_X1 U15467 ( .A(n12518), .B(n12513), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12450) );
  NAND2_X1 U15468 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12449) );
  INV_X1 U15469 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13984) );
  NAND2_X1 U15470 ( .A1(n12471), .A2(n13984), .ZN(n12453) );
  NAND2_X1 U15471 ( .A1(n13362), .A2(n13984), .ZN(n12451) );
  OAI211_X1 U15472 ( .C1(n14256), .C2(n20884), .A(n12513), .B(n12451), .ZN(
        n12452) );
  NAND2_X1 U15473 ( .A1(n12513), .A2(n14690), .ZN(n12455) );
  INV_X1 U15474 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U15475 ( .A1(n13362), .A2(n14355), .ZN(n12454) );
  NAND3_X1 U15476 ( .A1(n12455), .A2(n12421), .A3(n12454), .ZN(n12457) );
  NAND2_X1 U15477 ( .A1(n12505), .A2(n14355), .ZN(n12456) );
  NAND2_X1 U15478 ( .A1(n12457), .A2(n12456), .ZN(n14026) );
  NAND2_X1 U15479 ( .A1(n15877), .A2(n13345), .ZN(n12459) );
  MUX2_X1 U15480 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12458) );
  NAND2_X1 U15481 ( .A1(n12459), .A2(n12458), .ZN(n14048) );
  MUX2_X1 U15482 ( .A(n12518), .B(n12513), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12462) );
  NAND2_X1 U15483 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12460) );
  MUX2_X1 U15484 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12465) );
  INV_X1 U15485 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12463) );
  NAND2_X1 U15486 ( .A1(n13345), .A2(n12463), .ZN(n12464) );
  NAND2_X1 U15487 ( .A1(n12465), .A2(n12464), .ZN(n14346) );
  NAND2_X1 U15488 ( .A1(n12513), .A2(n12466), .ZN(n12468) );
  INV_X1 U15489 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15795) );
  NAND2_X1 U15490 ( .A1(n13362), .A2(n15795), .ZN(n12467) );
  NAND3_X1 U15491 ( .A1(n12468), .A2(n12421), .A3(n12467), .ZN(n12470) );
  NAND2_X1 U15492 ( .A1(n12505), .A2(n15795), .ZN(n12469) );
  NAND2_X1 U15493 ( .A1(n12470), .A2(n12469), .ZN(n14038) );
  INV_X1 U15494 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14480) );
  NAND2_X1 U15495 ( .A1(n12471), .A2(n14480), .ZN(n12474) );
  NAND2_X1 U15496 ( .A1(n13362), .A2(n14480), .ZN(n12472) );
  OAI211_X1 U15497 ( .C1(n14256), .C2(n12395), .A(n12513), .B(n12472), .ZN(
        n12473) );
  NAND2_X1 U15498 ( .A1(n12474), .A2(n12473), .ZN(n14476) );
  INV_X1 U15499 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14471) );
  NAND2_X1 U15500 ( .A1(n12505), .A2(n14471), .ZN(n12478) );
  NAND2_X1 U15501 ( .A1(n12513), .A2(n15983), .ZN(n12476) );
  NAND2_X1 U15502 ( .A1(n13362), .A2(n14471), .ZN(n12475) );
  NAND3_X1 U15503 ( .A1(n12476), .A2(n12421), .A3(n12475), .ZN(n12477) );
  MUX2_X1 U15504 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12480) );
  INV_X1 U15505 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U15506 ( .A1(n13345), .A2(n14654), .ZN(n12479) );
  INV_X1 U15507 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15760) );
  NAND2_X1 U15508 ( .A1(n12505), .A2(n15760), .ZN(n12484) );
  NAND2_X1 U15509 ( .A1(n12513), .A2(n15982), .ZN(n12482) );
  NAND2_X1 U15510 ( .A1(n13362), .A2(n15760), .ZN(n12481) );
  NAND3_X1 U15511 ( .A1(n12482), .A2(n12421), .A3(n12481), .ZN(n12483) );
  AND2_X1 U15512 ( .A1(n12484), .A2(n12483), .ZN(n14457) );
  MUX2_X1 U15513 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12486) );
  OR2_X1 U15514 ( .A1(n13082), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12485) );
  NAND2_X1 U15515 ( .A1(n12486), .A2(n12485), .ZN(n14318) );
  NAND2_X1 U15516 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12488) );
  MUX2_X1 U15517 ( .A(n12518), .B(n12513), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12487) );
  NAND2_X1 U15518 ( .A1(n12488), .A2(n12487), .ZN(n14071) );
  MUX2_X1 U15519 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12490) );
  NAND2_X1 U15520 ( .A1(n13345), .A2(n12399), .ZN(n12489) );
  INV_X1 U15521 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U15522 ( .A1(n12505), .A2(n12492), .ZN(n12496) );
  INV_X1 U15523 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U15524 ( .A1(n12513), .A2(n12491), .ZN(n12494) );
  NAND2_X1 U15525 ( .A1(n13362), .A2(n12492), .ZN(n12493) );
  NAND3_X1 U15526 ( .A1(n12494), .A2(n12421), .A3(n12493), .ZN(n12495) );
  AND2_X1 U15527 ( .A1(n12496), .A2(n12495), .ZN(n14439) );
  NAND2_X1 U15528 ( .A1(n15950), .A2(n13345), .ZN(n12498) );
  MUX2_X1 U15529 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12497) );
  NAND2_X1 U15530 ( .A1(n12498), .A2(n12497), .ZN(n14432) );
  INV_X1 U15531 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14427) );
  NAND2_X1 U15532 ( .A1(n12505), .A2(n14427), .ZN(n12502) );
  NAND2_X1 U15533 ( .A1(n12513), .A2(n15940), .ZN(n12500) );
  NAND2_X1 U15534 ( .A1(n13362), .A2(n14427), .ZN(n12499) );
  NAND3_X1 U15535 ( .A1(n12500), .A2(n12421), .A3(n12499), .ZN(n12501) );
  NOR2_X2 U15536 ( .A1(n14434), .A2(n14424), .ZN(n14423) );
  MUX2_X1 U15537 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12504) );
  OR2_X1 U15538 ( .A1(n13082), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12503) );
  AND2_X1 U15539 ( .A1(n12504), .A2(n12503), .ZN(n14308) );
  INV_X1 U15540 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U15541 ( .A1(n12505), .A2(n15704), .ZN(n12509) );
  INV_X1 U15542 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U15543 ( .A1(n12513), .A2(n14595), .ZN(n12507) );
  NAND2_X1 U15544 ( .A1(n13362), .A2(n15704), .ZN(n12506) );
  NAND3_X1 U15545 ( .A1(n12507), .A2(n12421), .A3(n12506), .ZN(n12508) );
  AND2_X1 U15546 ( .A1(n12509), .A2(n12508), .ZN(n14414) );
  MUX2_X1 U15547 ( .A(n12510), .B(n12421), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12512) );
  INV_X1 U15548 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15917) );
  NAND2_X1 U15549 ( .A1(n13345), .A2(n15917), .ZN(n12511) );
  NAND2_X1 U15550 ( .A1(n12512), .A2(n12511), .ZN(n14297) );
  NAND2_X1 U15551 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12515) );
  MUX2_X1 U15552 ( .A(n12518), .B(n12513), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12514) );
  NAND2_X1 U15553 ( .A1(n12515), .A2(n12514), .ZN(n14282) );
  OR2_X1 U15554 ( .A1(n13082), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12517) );
  INV_X1 U15555 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U15556 ( .A1(n13362), .A2(n14409), .ZN(n12516) );
  NAND2_X1 U15557 ( .A1(n12517), .A2(n12516), .ZN(n14254) );
  OAI22_X1 U15558 ( .A1(n14254), .A2(n14256), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12518), .ZN(n14275) );
  NAND2_X1 U15559 ( .A1(n14284), .A2(n14275), .ZN(n14277) );
  MUX2_X1 U15560 ( .A(n14257), .B(n12421), .S(n14277), .Z(n12520) );
  AOI22_X1 U15561 ( .A1(n13082), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13349), .ZN(n12519) );
  NOR2_X1 U15562 ( .A1(n14363), .A2(n20107), .ZN(n12533) );
  NAND2_X1 U15563 ( .A1(n13422), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U15564 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20654) );
  AND2_X1 U15565 ( .A1(n20654), .A2(n20535), .ZN(n15663) );
  NOR2_X1 U15566 ( .A1(n12529), .A2(n15663), .ZN(n12521) );
  AND2_X1 U15567 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n12524) );
  INV_X1 U15568 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20657) );
  NAND2_X1 U15569 ( .A1(n12522), .A2(n20657), .ZN(n15689) );
  INV_X1 U15570 ( .A(n15689), .ZN(n13270) );
  OAI21_X1 U15571 ( .B1(n13422), .B2(n13270), .A(n20654), .ZN(n13384) );
  NOR2_X1 U15572 ( .A1(n13384), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12531) );
  INV_X1 U15573 ( .A(n15779), .ZN(n19976) );
  OR2_X1 U15574 ( .A1(n15771), .A2(n19976), .ZN(n19993) );
  NAND2_X1 U15575 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12526) );
  INV_X1 U15576 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15932) );
  INV_X1 U15577 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15948) );
  INV_X1 U15578 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15735) );
  INV_X1 U15579 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20685) );
  INV_X1 U15580 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20681) );
  INV_X1 U15581 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20679) );
  INV_X1 U15582 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20676) );
  INV_X1 U15583 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20671) );
  INV_X1 U15584 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20669) );
  NAND4_X1 U15585 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14366)
         );
  NAND3_X1 U15586 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13849) );
  NOR3_X1 U15587 ( .A1(n20669), .A2(n14366), .A3(n13849), .ZN(n13978) );
  NAND2_X1 U15588 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n13978), .ZN(n14358) );
  NOR2_X1 U15589 ( .A1(n20671), .A2(n14358), .ZN(n14356) );
  NAND3_X1 U15590 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n14356), .ZN(n14348) );
  NOR3_X1 U15591 ( .A1(n20679), .A2(n20676), .A3(n14348), .ZN(n15781) );
  NAND2_X1 U15592 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15781), .ZN(n15769) );
  NOR2_X1 U15593 ( .A1(n20681), .A2(n15769), .ZN(n14328) );
  NAND2_X1 U15594 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14328), .ZN(n14317) );
  NOR2_X1 U15595 ( .A1(n20685), .A2(n14317), .ZN(n14322) );
  NAND2_X1 U15596 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n14322), .ZN(n15747) );
  NAND2_X1 U15597 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15721) );
  NOR4_X1 U15598 ( .A1(n15948), .A2(n15735), .A3(n15747), .A4(n15721), .ZN(
        n15714) );
  NAND2_X1 U15599 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15714), .ZN(n14310) );
  NOR2_X1 U15600 ( .A1(n15932), .A2(n14310), .ZN(n12525) );
  AOI21_X1 U15601 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n12525), .A(n15803), 
        .ZN(n12523) );
  OR2_X1 U15602 ( .A1(n12523), .A2(n19976), .ZN(n15708) );
  AOI21_X1 U15603 ( .B1(n19993), .B2(n12526), .A(n15708), .ZN(n14289) );
  OAI21_X1 U15604 ( .B1(n12524), .B2(n15803), .A(n14289), .ZN(n14266) );
  NAND2_X1 U15605 ( .A1(n15771), .A2(n12525), .ZN(n15702) );
  INV_X1 U15606 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15706) );
  NOR2_X1 U15607 ( .A1(n15702), .A2(n15706), .ZN(n14298) );
  INV_X1 U15608 ( .A(n12526), .ZN(n12527) );
  NAND2_X1 U15609 ( .A1(n14298), .A2(n12527), .ZN(n14274) );
  INV_X1 U15610 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n12528) );
  NAND3_X1 U15611 ( .A1(n12528), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .ZN(n12535) );
  INV_X1 U15612 ( .A(n12529), .ZN(n12530) );
  NOR2_X1 U15613 ( .A1(n12531), .A2(n12530), .ZN(n12532) );
  AOI22_X1 U15614 ( .A1(n19997), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19977), .ZN(n12534) );
  OAI21_X1 U15615 ( .B1(n14274), .B2(n12535), .A(n12534), .ZN(n12536) );
  AOI21_X1 U15616 ( .B1(n14266), .B2(P1_REIP_REG_31__SCAN_IN), .A(n12536), 
        .ZN(n12537) );
  NAND2_X1 U15617 ( .A1(n12540), .A2(n12539), .ZN(P1_U2809) );
  AND2_X1 U15618 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12549) );
  AOI21_X1 U15619 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12549), .A(
        n15241), .ZN(n12542) );
  NOR2_X1 U15620 ( .A1(n15127), .A2(n12542), .ZN(n14247) );
  OAI21_X1 U15621 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15241), .A(
        n14247), .ZN(n12554) );
  INV_X1 U15622 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19832) );
  AOI22_X1 U15623 ( .A1(n11400), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12543) );
  OAI21_X1 U15624 ( .B1(n12546), .B2(n19832), .A(n12543), .ZN(n12544) );
  INV_X1 U15625 ( .A(n12544), .ZN(n12565) );
  INV_X1 U15626 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14235) );
  AOI22_X1 U15627 ( .A1(n11400), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11211), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12545) );
  OAI21_X1 U15628 ( .B1(n12546), .B2(n14235), .A(n12545), .ZN(n12975) );
  AOI222_X1 U15629 ( .A1(n12547), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11400), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11211), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12548) );
  NAND4_X1 U15630 ( .A1(n14242), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n11073), .ZN(n12550) );
  OAI211_X1 U15631 ( .C1(n16324), .C2(n16102), .A(n12551), .B(n12550), .ZN(
        n12552) );
  AOI211_X1 U15632 ( .C1(n12554), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12553), .B(n12552), .ZN(n12556) );
  NAND2_X1 U15633 ( .A1(n9715), .A2(n16313), .ZN(n12555) );
  NOR2_X1 U15634 ( .A1(n11072), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12559) );
  NOR2_X1 U15635 ( .A1(n12558), .A2(n12559), .ZN(n12583) );
  AOI21_X1 U15636 ( .B1(n12562), .B2(n12561), .A(n12560), .ZN(n12571) );
  OAI21_X1 U15637 ( .B1(n12564), .B2(n12563), .A(n12927), .ZN(n14792) );
  INV_X1 U15638 ( .A(n14792), .ZN(n16111) );
  XNOR2_X1 U15639 ( .A(n12566), .B(n12565), .ZN(n14854) );
  NAND2_X1 U15640 ( .A1(n14242), .A2(n12570), .ZN(n12567) );
  NAND2_X1 U15641 ( .A1(n19044), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12578) );
  OAI211_X1 U15642 ( .C1(n16324), .C2(n14854), .A(n12567), .B(n12578), .ZN(
        n12568) );
  AOI21_X1 U15643 ( .B1(n16111), .B2(n16312), .A(n12568), .ZN(n12569) );
  OAI21_X1 U15644 ( .B1(n12571), .B2(n12570), .A(n12569), .ZN(n12572) );
  AOI21_X1 U15645 ( .B1(n12583), .B2(n16313), .A(n12572), .ZN(n12576) );
  NAND2_X1 U15646 ( .A1(n12573), .A2(n14228), .ZN(n12575) );
  XOR2_X1 U15647 ( .A(n12575), .B(n12574), .Z(n12584) );
  NAND2_X1 U15648 ( .A1(n12576), .A2(n10252), .ZN(P2_U3017) );
  AOI21_X1 U15649 ( .B1(n12579), .B2(n11084), .A(n12577), .ZN(n16114) );
  OAI21_X1 U15650 ( .B1(n19229), .B2(n12579), .A(n12578), .ZN(n12580) );
  AOI21_X1 U15651 ( .B1(n19220), .B2(n16114), .A(n12580), .ZN(n12581) );
  OAI21_X1 U15652 ( .B1(n14792), .B2(n16206), .A(n12581), .ZN(n12582) );
  AOI21_X1 U15653 ( .B1(n12583), .B2(n19224), .A(n12582), .ZN(n12585) );
  NAND2_X1 U15654 ( .A1(n12585), .A2(n10260), .ZN(P2_U2985) );
  NAND2_X1 U15655 ( .A1(n12586), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12587) );
  NOR2_X1 U15656 ( .A1(n12599), .A2(n19886), .ZN(n19692) );
  OAI21_X1 U15657 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12598), .A(
        n19864), .ZN(n12588) );
  NOR2_X1 U15658 ( .A1(n12588), .A2(n19745), .ZN(n19584) );
  AOI21_X1 U15659 ( .B1(n12602), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19584), .ZN(n12589) );
  AOI22_X1 U15660 ( .A1(n12602), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19864), .B2(n19896), .ZN(n12591) );
  NAND2_X1 U15661 ( .A1(n12602), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12593) );
  XNOR2_X1 U15662 ( .A(n19886), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19358) );
  NAND2_X1 U15663 ( .A1(n19358), .A2(n19864), .ZN(n19298) );
  INV_X1 U15664 ( .A(n12595), .ZN(n12596) );
  INV_X1 U15665 ( .A(n12598), .ZN(n12601) );
  NAND2_X1 U15666 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19554) );
  NAND2_X1 U15667 ( .A1(n19554), .A2(n12599), .ZN(n12600) );
  NAND2_X1 U15668 ( .A1(n12601), .A2(n12600), .ZN(n19359) );
  NAND2_X1 U15669 ( .A1(n12602), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12603) );
  OAI21_X1 U15670 ( .B1(n19359), .B2(n19652), .A(n12603), .ZN(n12604) );
  NAND2_X1 U15671 ( .A1(n13292), .A2(n13291), .ZN(n12605) );
  NAND2_X1 U15672 ( .A1(n13373), .A2(n13374), .ZN(n12612) );
  INV_X1 U15673 ( .A(n12607), .ZN(n12609) );
  AND2_X1 U15674 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12586), .ZN(
        n12608) );
  AOI21_X1 U15675 ( .B1(n12610), .B2(n12609), .A(n12608), .ZN(n12611) );
  NAND4_X1 U15676 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__5__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12613) );
  NOR3_X1 U15677 ( .A1(n12846), .A2(n13486), .A3(n12613), .ZN(n12614) );
  AOI22_X1 U15678 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15679 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15680 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12618) );
  NAND2_X1 U15681 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12617) );
  AND2_X1 U15682 ( .A1(n12618), .A2(n12617), .ZN(n12620) );
  AOI22_X1 U15683 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12619) );
  NAND4_X1 U15684 ( .A1(n12622), .A2(n12621), .A3(n12620), .A4(n12619), .ZN(
        n12628) );
  AOI22_X1 U15685 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15686 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15687 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U15688 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12623) );
  NAND4_X1 U15689 ( .A1(n12626), .A2(n12625), .A3(n12624), .A4(n12623), .ZN(
        n12627) );
  NOR2_X1 U15690 ( .A1(n12628), .A2(n12627), .ZN(n13832) );
  NAND2_X1 U15691 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12629) );
  OAI21_X1 U15692 ( .B1(n13559), .B2(n12630), .A(n12629), .ZN(n12636) );
  AOI22_X1 U15693 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12634) );
  NAND2_X1 U15694 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12633) );
  NAND2_X1 U15695 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12632) );
  NAND2_X1 U15696 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12631) );
  NAND4_X1 U15697 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n12635) );
  NOR2_X1 U15698 ( .A1(n12636), .A2(n12635), .ZN(n12644) );
  AOI22_X1 U15699 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10613), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15700 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12639) );
  NAND2_X1 U15701 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12638) );
  NAND2_X1 U15702 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12637) );
  AND4_X1 U15703 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12643) );
  AOI22_X1 U15704 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10667), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U15705 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10763), .ZN(n12641) );
  NAND4_X1 U15706 ( .A1(n12644), .A2(n12643), .A3(n12642), .A4(n12641), .ZN(
        n16186) );
  AOI22_X1 U15707 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10667), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15708 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n10763), .ZN(n12649) );
  AOI22_X1 U15709 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12719), .B1(
        n10613), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U15710 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12645) );
  AND2_X1 U15711 ( .A1(n12646), .A2(n12645), .ZN(n12648) );
  AOI22_X1 U15712 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12647) );
  NAND4_X1 U15713 ( .A1(n12650), .A2(n12649), .A3(n12648), .A4(n12647), .ZN(
        n12656) );
  AOI22_X1 U15714 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15715 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15716 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U15717 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12651) );
  NAND4_X1 U15718 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12655) );
  NOR2_X1 U15719 ( .A1(n12656), .A2(n12655), .ZN(n14851) );
  INV_X1 U15720 ( .A(n14851), .ZN(n12657) );
  AOI22_X1 U15721 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10667), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15722 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n10763), .ZN(n12663) );
  AOI22_X1 U15723 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10613), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U15724 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12659) );
  AND2_X1 U15725 ( .A1(n12660), .A2(n12659), .ZN(n12662) );
  AOI22_X1 U15726 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U15727 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12670) );
  AOI22_X1 U15728 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U15729 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U15730 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U15731 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12665) );
  NAND4_X1 U15732 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12669) );
  NOR2_X1 U15733 ( .A1(n12670), .A2(n12669), .ZN(n14935) );
  AOI22_X1 U15734 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15735 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10676), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15736 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U15737 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12671) );
  AND4_X1 U15738 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n12682) );
  AOI22_X1 U15739 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12719), .B1(
        n10613), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12678) );
  NAND2_X1 U15740 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12677) );
  NAND2_X1 U15741 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12676) );
  NAND2_X1 U15742 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12675) );
  AND4_X1 U15743 ( .A1(n12678), .A2(n12677), .A3(n12676), .A4(n12675), .ZN(
        n12681) );
  AOI22_X1 U15744 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10762), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15745 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n10763), .ZN(n12679) );
  NAND4_X1 U15746 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n14840) );
  AOI22_X1 U15747 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15748 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U15749 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15750 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12684) );
  AND2_X1 U15751 ( .A1(n12685), .A2(n12684), .ZN(n12687) );
  AOI22_X1 U15752 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12686) );
  NAND4_X1 U15753 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12696) );
  AOI22_X1 U15754 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15755 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U15756 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U15757 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12691) );
  NAND4_X1 U15758 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12695) );
  NOR2_X1 U15759 ( .A1(n12696), .A2(n12695), .ZN(n14920) );
  AOI22_X1 U15760 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10667), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15761 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10763), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15762 ( .A1(n10613), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12699) );
  NAND2_X1 U15763 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12698) );
  AND2_X1 U15764 ( .A1(n12699), .A2(n12698), .ZN(n12702) );
  AOI22_X1 U15765 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12701) );
  NAND4_X1 U15766 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12711) );
  AOI22_X1 U15767 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15768 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15769 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U15770 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12706) );
  NAND4_X1 U15771 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12710) );
  NOR2_X1 U15772 ( .A1(n12711), .A2(n12710), .ZN(n14836) );
  INV_X1 U15773 ( .A(n14836), .ZN(n12712) );
  INV_X1 U15774 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12713) );
  OR2_X1 U15775 ( .A1(n12714), .A2(n12713), .ZN(n12718) );
  NAND2_X1 U15776 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12717) );
  NAND2_X1 U15777 ( .A1(n10667), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12716) );
  NAND2_X1 U15778 ( .A1(n10763), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12715) );
  AND4_X1 U15779 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12732) );
  AOI22_X1 U15780 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10613), .B1(
        n12719), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15781 ( .A1(n12683), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12722) );
  NAND2_X1 U15782 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12721) );
  NAND2_X1 U15783 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12720) );
  AND4_X1 U15784 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12731) );
  AOI22_X1 U15785 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15786 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10581), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U15787 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12727) );
  NAND2_X1 U15788 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12726) );
  NAND2_X1 U15789 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12725) );
  AND4_X1 U15790 ( .A1(n12728), .A2(n12727), .A3(n12726), .A4(n12725), .ZN(
        n12729) );
  NAND4_X1 U15791 ( .A1(n12732), .A2(n12731), .A3(n12730), .A4(n12729), .ZN(
        n12754) );
  INV_X1 U15792 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U15793 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12736) );
  AND2_X1 U15794 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12735) );
  OR2_X1 U15795 ( .A1(n12735), .A2(n12734), .ZN(n12914) );
  OAI211_X1 U15796 ( .C1(n12882), .C2(n12737), .A(n12736), .B(n12914), .ZN(
        n12738) );
  INV_X1 U15797 ( .A(n12738), .ZN(n12744) );
  INV_X1 U15798 ( .A(n9661), .ZN(n12894) );
  AOI22_X1 U15799 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15800 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15801 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12741) );
  NAND4_X1 U15802 ( .A1(n12744), .A2(n12743), .A3(n12742), .A4(n12741), .ZN(
        n12753) );
  INV_X1 U15803 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15804 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12745) );
  INV_X1 U15805 ( .A(n12914), .ZN(n12836) );
  OAI211_X1 U15806 ( .C1(n12882), .C2(n12746), .A(n12745), .B(n12836), .ZN(
        n12747) );
  INV_X1 U15807 ( .A(n12747), .ZN(n12751) );
  AOI22_X1 U15808 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15809 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15810 ( .A1(n9669), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U15811 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12752) );
  AND2_X1 U15812 ( .A1(n12753), .A2(n12752), .ZN(n12759) );
  NAND2_X1 U15813 ( .A1(n12778), .A2(n11215), .ZN(n12758) );
  INV_X1 U15814 ( .A(n12754), .ZN(n12756) );
  NAND2_X1 U15815 ( .A1(n11215), .A2(n12759), .ZN(n12755) );
  NAND2_X1 U15816 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  NAND2_X1 U15817 ( .A1(n12758), .A2(n12757), .ZN(n12782) );
  INV_X1 U15818 ( .A(n12759), .ZN(n12760) );
  NOR2_X1 U15819 ( .A1(n11215), .A2(n12760), .ZN(n14823) );
  INV_X1 U15820 ( .A(n14835), .ZN(n12761) );
  INV_X1 U15821 ( .A(n12911), .ZN(n12892) );
  NAND2_X1 U15822 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12762) );
  OAI211_X1 U15823 ( .C1(n12892), .C2(n12763), .A(n12762), .B(n12914), .ZN(
        n12764) );
  INV_X1 U15824 ( .A(n12764), .ZN(n12768) );
  AOI22_X1 U15825 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12740), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U15826 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U15827 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12765) );
  NAND4_X1 U15828 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12777) );
  NAND2_X1 U15829 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12769) );
  OAI211_X1 U15830 ( .C1(n12892), .C2(n12770), .A(n12769), .B(n12836), .ZN(
        n12771) );
  INV_X1 U15831 ( .A(n12771), .ZN(n12775) );
  AOI22_X1 U15832 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12740), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15833 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15834 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12772) );
  NAND4_X1 U15835 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  AND2_X1 U15836 ( .A1(n12777), .A2(n12776), .ZN(n14892) );
  INV_X1 U15837 ( .A(n14892), .ZN(n12781) );
  INV_X1 U15838 ( .A(n12778), .ZN(n12779) );
  AOI211_X1 U15839 ( .C1(n12781), .C2(n12779), .A(n12846), .B(n12799), .ZN(
        n14891) );
  INV_X1 U15840 ( .A(n14823), .ZN(n12780) );
  NOR3_X1 U15841 ( .A1(n12782), .A2(n12781), .A3(n12780), .ZN(n12783) );
  INV_X1 U15842 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13948) );
  NAND2_X1 U15843 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12784) );
  OAI211_X1 U15844 ( .C1(n12882), .C2(n13948), .A(n12784), .B(n12914), .ZN(
        n12785) );
  INV_X1 U15845 ( .A(n12785), .ZN(n12789) );
  AOI22_X1 U15846 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U15847 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15848 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U15849 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12798) );
  NAND2_X1 U15850 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12790) );
  OAI211_X1 U15851 ( .C1(n12882), .C2(n12791), .A(n12790), .B(n12836), .ZN(
        n12792) );
  INV_X1 U15852 ( .A(n12792), .ZN(n12796) );
  AOI22_X1 U15853 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U15854 ( .A1(n9671), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U15855 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12793) );
  NAND4_X1 U15856 ( .A1(n12796), .A2(n12795), .A3(n12794), .A4(n12793), .ZN(
        n12797) );
  NAND2_X1 U15857 ( .A1(n12799), .A2(n12800), .ZN(n12824) );
  OAI211_X1 U15858 ( .C1(n12799), .C2(n12800), .A(n13307), .B(n12824), .ZN(
        n12803) );
  INV_X1 U15859 ( .A(n12800), .ZN(n12801) );
  NOR2_X1 U15860 ( .A1(n11215), .A2(n12801), .ZN(n14816) );
  NAND2_X1 U15861 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12807) );
  OAI211_X1 U15862 ( .C1(n12892), .C2(n12808), .A(n12807), .B(n12914), .ZN(
        n12809) );
  INV_X1 U15863 ( .A(n12809), .ZN(n12813) );
  AOI22_X1 U15864 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12740), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15865 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U15866 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12810) );
  NAND4_X1 U15867 ( .A1(n12813), .A2(n12812), .A3(n12811), .A4(n12810), .ZN(
        n12823) );
  NAND2_X1 U15868 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12815) );
  OAI211_X1 U15869 ( .C1(n12882), .C2(n12816), .A(n12815), .B(n12836), .ZN(
        n12817) );
  INV_X1 U15870 ( .A(n12817), .ZN(n12821) );
  AOI22_X1 U15871 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U15872 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15873 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12818) );
  NAND4_X1 U15874 ( .A1(n12821), .A2(n12820), .A3(n12819), .A4(n12818), .ZN(
        n12822) );
  NAND2_X1 U15875 ( .A1(n12823), .A2(n12822), .ZN(n12825) );
  AOI21_X1 U15876 ( .B1(n12824), .B2(n12825), .A(n12846), .ZN(n12827) );
  INV_X1 U15877 ( .A(n12824), .ZN(n12826) );
  INV_X1 U15878 ( .A(n12825), .ZN(n12828) );
  NAND2_X1 U15879 ( .A1(n12826), .A2(n12828), .ZN(n12847) );
  NOR2_X2 U15880 ( .A1(n14812), .A2(n10244), .ZN(n12852) );
  NAND2_X1 U15881 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12830) );
  OAI211_X1 U15882 ( .C1(n12882), .C2(n19249), .A(n12830), .B(n12914), .ZN(
        n12831) );
  INV_X1 U15883 ( .A(n12831), .ZN(n12835) );
  AOI22_X1 U15884 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U15885 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15886 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12832) );
  NAND4_X1 U15887 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12845) );
  INV_X1 U15888 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12838) );
  NAND2_X1 U15889 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12837) );
  OAI211_X1 U15890 ( .C1(n12882), .C2(n12838), .A(n12837), .B(n12836), .ZN(
        n12839) );
  INV_X1 U15891 ( .A(n12839), .ZN(n12843) );
  AOI22_X1 U15892 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15893 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U15894 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12840) );
  NAND4_X1 U15895 ( .A1(n12843), .A2(n12842), .A3(n12841), .A4(n12840), .ZN(
        n12844) );
  NAND2_X1 U15896 ( .A1(n12845), .A2(n12844), .ZN(n12850) );
  AOI21_X1 U15897 ( .B1(n12847), .B2(n12850), .A(n12846), .ZN(n12848) );
  OR2_X1 U15898 ( .A1(n12847), .A2(n12850), .ZN(n12873) );
  NAND2_X1 U15899 ( .A1(n12848), .A2(n12873), .ZN(n12851) );
  INV_X1 U15900 ( .A(n12851), .ZN(n12849) );
  NOR2_X1 U15901 ( .A1(n10294), .A2(n12850), .ZN(n14802) );
  AOI22_X1 U15902 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15903 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U15904 ( .A1(n12854), .A2(n12853), .ZN(n12872) );
  AOI22_X1 U15905 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12856) );
  AOI21_X1 U15906 ( .B1(n12915), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n12914), .ZN(n12855) );
  OAI211_X1 U15907 ( .C1(n9645), .C2(n12857), .A(n12856), .B(n12855), .ZN(
        n12871) );
  OAI22_X1 U15908 ( .A1(n12894), .A2(n12859), .B1(n12892), .B2(n12858), .ZN(
        n12869) );
  NAND2_X1 U15909 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12860) );
  OAI211_X1 U15910 ( .C1(n12882), .C2(n19257), .A(n12860), .B(n12914), .ZN(
        n12868) );
  OAI22_X1 U15911 ( .A1(n9651), .A2(n12863), .B1(n10300), .B2(n12862), .ZN(
        n12867) );
  OAI22_X1 U15912 ( .A1(n13603), .A2(n12865), .B1(n9645), .B2(n12864), .ZN(
        n12866) );
  OR4_X1 U15913 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n12870) );
  INV_X1 U15914 ( .A(n12873), .ZN(n14795) );
  INV_X1 U15915 ( .A(n14797), .ZN(n12874) );
  NAND3_X1 U15916 ( .A1(n14795), .A2(n12874), .A3(n11215), .ZN(n12902) );
  OAI22_X1 U15917 ( .A1(n12894), .A2(n12876), .B1(n12892), .B2(n12875), .ZN(
        n12886) );
  OAI22_X1 U15918 ( .A1(n9651), .A2(n12878), .B1(n13603), .B2(n12877), .ZN(
        n12885) );
  OAI22_X1 U15919 ( .A1(n9664), .A2(n12880), .B1(n9645), .B2(n12879), .ZN(
        n12884) );
  NAND2_X1 U15920 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12881) );
  OAI211_X1 U15921 ( .C1(n12882), .C2(n13474), .A(n12881), .B(n12914), .ZN(
        n12883) );
  NOR4_X1 U15922 ( .A1(n12886), .A2(n12885), .A3(n12884), .A4(n12883), .ZN(
        n12901) );
  AOI22_X1 U15923 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12889) );
  AOI21_X1 U15924 ( .B1(n12915), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n12914), .ZN(n12888) );
  OAI211_X1 U15925 ( .C1(n12733), .C2(n12890), .A(n12889), .B(n12888), .ZN(
        n12899) );
  OAI22_X1 U15926 ( .A1(n12894), .A2(n12893), .B1(n12892), .B2(n12891), .ZN(
        n12898) );
  OAI22_X1 U15927 ( .A1(n9651), .A2(n12896), .B1(n13603), .B2(n12895), .ZN(
        n12897) );
  NOR3_X1 U15928 ( .A1(n12899), .A2(n12898), .A3(n12897), .ZN(n12900) );
  NOR2_X1 U15929 ( .A1(n12901), .A2(n12900), .ZN(n12903) );
  XNOR2_X1 U15930 ( .A(n12902), .B(n12903), .ZN(n14790) );
  INV_X1 U15931 ( .A(n12902), .ZN(n12904) );
  AOI22_X1 U15932 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12910), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U15933 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U15934 ( .A1(n12906), .A2(n12905), .ZN(n12922) );
  AOI22_X1 U15935 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12909) );
  NAND2_X1 U15936 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12908) );
  NAND2_X1 U15937 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12907) );
  NAND4_X1 U15938 ( .A1(n12909), .A2(n12914), .A3(n12908), .A4(n12907), .ZN(
        n12921) );
  AOI22_X1 U15939 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12910), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U15940 ( .A1(n12740), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12912) );
  NAND2_X1 U15941 ( .A1(n12913), .A2(n12912), .ZN(n12920) );
  AOI21_X1 U15942 ( .B1(n12915), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12914), .ZN(n12917) );
  AOI22_X1 U15943 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12916) );
  OAI211_X1 U15944 ( .C1(n12733), .C2(n12918), .A(n12917), .B(n12916), .ZN(
        n12919) );
  OAI22_X1 U15945 ( .A1(n12922), .A2(n12921), .B1(n12920), .B2(n12919), .ZN(
        n12923) );
  INV_X1 U15946 ( .A(n13641), .ZN(n12924) );
  INV_X1 U15947 ( .A(n13554), .ZN(n13637) );
  NAND2_X1 U15948 ( .A1(n12924), .A2(n13637), .ZN(n13154) );
  INV_X1 U15949 ( .A(n11169), .ZN(n12925) );
  INV_X2 U15950 ( .A(n19078), .ZN(n14844) );
  NAND2_X1 U15951 ( .A1(n14250), .A2(n14844), .ZN(n12930) );
  NAND2_X1 U15952 ( .A1(n19078), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12929) );
  OAI21_X1 U15953 ( .B1(n14227), .B2(n16181), .A(n12931), .ZN(P2_U2857) );
  AOI21_X1 U15954 ( .B1(n16123), .B2(n12933), .A(n10973), .ZN(n16122) );
  OR2_X1 U15955 ( .A1(n9769), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12935) );
  NAND2_X1 U15956 ( .A1(n12933), .A2(n12935), .ZN(n14978) );
  INV_X1 U15957 ( .A(n14978), .ZN(n16142) );
  AOI21_X1 U15958 ( .B1(n14988), .B2(n12936), .A(n9769), .ZN(n16154) );
  INV_X1 U15959 ( .A(n12940), .ZN(n12937) );
  NAND2_X1 U15960 ( .A1(n12937), .A2(n10152), .ZN(n12938) );
  AND2_X1 U15961 ( .A1(n12938), .A2(n12936), .ZN(n14997) );
  INV_X1 U15962 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15004) );
  AOI21_X1 U15963 ( .B1(n15004), .B2(n12939), .A(n12940), .ZN(n16165) );
  OAI21_X1 U15964 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9685), .A(
        n12939), .ZN(n15013) );
  INV_X1 U15965 ( .A(n15013), .ZN(n15634) );
  AOI21_X1 U15966 ( .B1(n15031), .B2(n12941), .A(n9685), .ZN(n15034) );
  OAI21_X1 U15967 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12942), .A(
        n12941), .ZN(n15045) );
  INV_X1 U15968 ( .A(n15045), .ZN(n18891) );
  NOR2_X1 U15969 ( .A1(n12943), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12944) );
  NOR2_X1 U15970 ( .A1(n12942), .A2(n12944), .ZN(n18904) );
  AOI21_X1 U15971 ( .B1(n12945), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12946) );
  OR2_X1 U15972 ( .A1(n12943), .A2(n12946), .ZN(n18915) );
  AOI21_X1 U15973 ( .B1(n16198), .B2(n9677), .A(n12945), .ZN(n13951) );
  OAI21_X1 U15974 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12948), .A(
        n12950), .ZN(n16220) );
  INV_X1 U15975 ( .A(n16220), .ZN(n12966) );
  OAI21_X1 U15976 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12951), .A(
        n12952), .ZN(n16238) );
  INV_X1 U15977 ( .A(n16238), .ZN(n18968) );
  OAI21_X1 U15978 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12953), .A(
        n12954), .ZN(n18997) );
  INV_X1 U15979 ( .A(n18997), .ZN(n12964) );
  AOI21_X1 U15980 ( .B1(n16270), .B2(n12955), .A(n12956), .ZN(n16257) );
  AOI21_X1 U15981 ( .B1(n15115), .B2(n12957), .A(n12958), .ZN(n19031) );
  AOI21_X1 U15982 ( .B1(n19228), .B2(n12961), .A(n12962), .ZN(n19219) );
  AOI21_X1 U15983 ( .B1(n19058), .B2(n13824), .A(n12959), .ZN(n13820) );
  AOI22_X1 U15984 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n12960), .ZN(n15333) );
  AOI22_X1 U15985 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19058), .B2(n12960), .ZN(
        n15332) );
  NAND2_X1 U15986 ( .A1(n15333), .A2(n15332), .ZN(n15331) );
  NOR2_X1 U15987 ( .A1(n13820), .A2(n15331), .ZN(n13882) );
  OAI21_X1 U15988 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12959), .A(
        n12961), .ZN(n13883) );
  NAND2_X1 U15989 ( .A1(n13882), .A2(n13883), .ZN(n13808) );
  NOR2_X1 U15990 ( .A1(n19219), .A2(n13808), .ZN(n19046) );
  OAI21_X1 U15991 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12962), .A(
        n12957), .ZN(n19048) );
  NAND2_X1 U15992 ( .A1(n19046), .A2(n19048), .ZN(n19028) );
  NOR2_X1 U15993 ( .A1(n19031), .A2(n19028), .ZN(n19016) );
  OAI21_X1 U15994 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12958), .A(
        n12955), .ZN(n19017) );
  NAND2_X1 U15995 ( .A1(n19016), .A2(n19017), .ZN(n13872) );
  NOR2_X1 U15996 ( .A1(n16257), .A2(n13872), .ZN(n19006) );
  OAI21_X1 U15997 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n12956), .A(
        n12963), .ZN(n19007) );
  NAND2_X1 U15998 ( .A1(n19006), .A2(n19007), .ZN(n18995) );
  NOR2_X1 U15999 ( .A1(n12964), .A2(n18995), .ZN(n18988) );
  AOI21_X1 U16000 ( .B1(n16245), .B2(n12954), .A(n12951), .ZN(n16239) );
  INV_X1 U16001 ( .A(n16239), .ZN(n18991) );
  NAND2_X1 U16002 ( .A1(n18988), .A2(n18991), .ZN(n18967) );
  NOR2_X1 U16003 ( .A1(n18968), .A2(n18967), .ZN(n18964) );
  AOI21_X1 U16004 ( .B1(n12965), .B2(n12952), .A(n12948), .ZN(n18955) );
  INV_X1 U16005 ( .A(n18955), .ZN(n18963) );
  NAND2_X1 U16006 ( .A1(n18964), .A2(n18963), .ZN(n13962) );
  NOR2_X1 U16007 ( .A1(n12966), .A2(n13962), .ZN(n18943) );
  OAI21_X1 U16008 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n12949), .A(
        n9677), .ZN(n18952) );
  NAND2_X1 U16009 ( .A1(n18943), .A2(n18952), .ZN(n18941) );
  NOR2_X1 U16010 ( .A1(n13951), .A2(n18941), .ZN(n18933) );
  XNOR2_X1 U16011 ( .A(n12945), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18932) );
  NAND2_X1 U16012 ( .A1(n18933), .A2(n18932), .ZN(n18931) );
  OAI21_X1 U16013 ( .B1(n19047), .B2(n18915), .A(n18916), .ZN(n18905) );
  NOR2_X1 U16014 ( .A1(n18904), .A2(n18905), .ZN(n18906) );
  NOR2_X1 U16015 ( .A1(n15634), .A2(n15633), .ZN(n15632) );
  NOR2_X1 U16016 ( .A1(n19047), .A2(n15632), .ZN(n16164) );
  NOR2_X1 U16017 ( .A1(n16165), .A2(n16164), .ZN(n16163) );
  NOR2_X1 U16018 ( .A1(n16142), .A2(n16141), .ZN(n16140) );
  NOR2_X1 U16019 ( .A1(n19047), .A2(n14769), .ZN(n16113) );
  NOR2_X1 U16020 ( .A1(n19047), .A2(n16112), .ZN(n12967) );
  XNOR2_X1 U16021 ( .A(n12577), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16104) );
  XNOR2_X1 U16022 ( .A(n12967), .B(n16104), .ZN(n12969) );
  NOR2_X1 U16023 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15691) );
  NAND3_X1 U16024 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15691), .A3(n19470), 
        .ZN(n19759) );
  NAND2_X1 U16025 ( .A1(n12969), .A2(n12968), .ZN(n12998) );
  NAND2_X1 U16026 ( .A1(n13635), .A2(n16343), .ZN(n12970) );
  OR2_X1 U16027 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19778), .ZN(n12985) );
  NOR2_X1 U16028 ( .A1(n12987), .A2(n12985), .ZN(n12971) );
  NAND2_X1 U16029 ( .A1(n19470), .A2(n13158), .ZN(n12980) );
  INV_X1 U16030 ( .A(n12980), .ZN(n13600) );
  NAND2_X1 U16031 ( .A1(n12972), .A2(n13600), .ZN(n12973) );
  NOR2_X2 U16032 ( .A1(n13040), .A2(n12973), .ZN(n18972) );
  OR2_X1 U16033 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  INV_X1 U16034 ( .A(n14245), .ZN(n12978) );
  AOI22_X1 U16035 ( .A1(n14250), .A2(n19067), .B1(n18972), .B2(n12978), .ZN(
        n12996) );
  OR2_X1 U16036 ( .A1(n13599), .A2(n13163), .ZN(n12979) );
  NAND2_X1 U16037 ( .A1(n13147), .A2(n12980), .ZN(n16099) );
  INV_X1 U16038 ( .A(n13052), .ZN(n12982) );
  INV_X1 U16039 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12981) );
  NAND3_X1 U16040 ( .A1(n12982), .A2(n12981), .A3(n12985), .ZN(n12983) );
  INV_X1 U16041 ( .A(n12984), .ZN(n12993) );
  NAND2_X1 U16042 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12985), .ZN(n12986) );
  NOR2_X1 U16043 ( .A1(n12987), .A2(n12986), .ZN(n12988) );
  NOR2_X1 U16044 ( .A1(n19888), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19443) );
  INV_X1 U16045 ( .A(n19443), .ZN(n19755) );
  NOR2_X1 U16046 ( .A1(n19762), .A2(n19755), .ZN(n16340) );
  INV_X1 U16047 ( .A(n16340), .ZN(n12989) );
  NAND2_X1 U16048 ( .A1(n19759), .A2(n12989), .ZN(n12990) );
  NOR2_X1 U16049 ( .A1(n19044), .A2(n12990), .ZN(n12991) );
  NAND2_X1 U16050 ( .A1(n19059), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19057) );
  AOI22_X1 U16051 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19038), .ZN(n12992) );
  OAI21_X1 U16052 ( .B1(n12993), .B2(n19024), .A(n12992), .ZN(n12994) );
  AOI21_X1 U16053 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19055), .A(n12994), .ZN(
        n12995) );
  NAND2_X1 U16054 ( .A1(n12998), .A2(n12997), .ZN(P2_U2825) );
  NOR2_X1 U16055 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13000) );
  NOR4_X1 U16056 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12999) );
  NAND4_X1 U16057 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13000), .A4(n12999), .ZN(n13023) );
  NOR4_X1 U16058 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13004) );
  NOR4_X1 U16059 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13003) );
  NOR4_X1 U16060 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13002) );
  NOR4_X1 U16061 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13001) );
  AND4_X1 U16062 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13010) );
  NOR4_X1 U16063 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_2__SCAN_IN), .ZN(n13008) );
  NOR4_X1 U16064 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13007) );
  NOR4_X1 U16065 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13006) );
  INV_X1 U16066 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13005) );
  AND4_X1 U16067 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  NAND2_X1 U16068 ( .A1(n13010), .A2(n13009), .ZN(n13011) );
  INV_X1 U16069 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20759) );
  NOR3_X1 U16070 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20759), .ZN(n13013) );
  NOR4_X1 U16071 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13012) );
  NAND4_X1 U16072 ( .A1(n20102), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13013), .A4(
        n13012), .ZN(U214) );
  NOR4_X1 U16073 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13017) );
  NOR4_X1 U16074 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13016) );
  NOR4_X1 U16075 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13015) );
  NOR4_X1 U16076 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13014) );
  NAND4_X1 U16077 ( .A1(n13017), .A2(n13016), .A3(n13015), .A4(n13014), .ZN(
        n13022) );
  NOR4_X1 U16078 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_2__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13020) );
  NOR4_X1 U16079 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13019) );
  NOR4_X1 U16080 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13018) );
  INV_X1 U16081 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19790) );
  NAND4_X1 U16082 ( .A1(n13020), .A2(n13019), .A3(n13018), .A4(n19790), .ZN(
        n13021) );
  NOR2_X1 U16083 ( .A1(n14221), .A2(n13023), .ZN(n16422) );
  NAND2_X1 U16084 ( .A1(n16422), .A2(U214), .ZN(U212) );
  AOI211_X1 U16085 ( .C1(n15034), .C2(n10162), .A(n13024), .B(n19759), .ZN(
        n13035) );
  OAI22_X1 U16086 ( .A1(n19816), .A2(n19059), .B1(n15031), .B2(n19057), .ZN(
        n13034) );
  INV_X1 U16087 ( .A(n13025), .ZN(n13026) );
  INV_X1 U16088 ( .A(n19055), .ZN(n19042) );
  OAI22_X1 U16089 ( .A1(n13026), .A2(n19024), .B1(n19042), .B2(n10821), .ZN(
        n13033) );
  NAND2_X1 U16090 ( .A1(n14843), .A2(n13027), .ZN(n13028) );
  NAND2_X1 U16091 ( .A1(n14831), .A2(n13028), .ZN(n16177) );
  OR2_X1 U16092 ( .A1(n14927), .A2(n13029), .ZN(n13030) );
  AND2_X1 U16093 ( .A1(n13030), .A2(n14908), .ZN(n15189) );
  INV_X1 U16094 ( .A(n15189), .ZN(n13031) );
  OAI22_X1 U16095 ( .A1(n16177), .A2(n18958), .B1(n13031), .B2(n19065), .ZN(
        n13032) );
  OR4_X1 U16096 ( .A1(n13035), .A2(n13034), .A3(n13033), .A4(n13032), .ZN(
        P2_U2834) );
  OR2_X1 U16097 ( .A1(n13157), .A2(n13163), .ZN(n19148) );
  NOR2_X1 U16098 ( .A1(n13636), .A2(n19148), .ZN(n19069) );
  INV_X1 U16099 ( .A(n19069), .ZN(n14023) );
  OAI21_X1 U16100 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n19652), .A(n13052), 
        .ZN(n13037) );
  AOI21_X1 U16101 ( .B1(n14023), .B2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n13037), 
        .ZN(n13036) );
  INV_X1 U16102 ( .A(n13036), .ZN(P2_U2814) );
  NOR3_X1 U16103 ( .A1(n13037), .A2(n19069), .A3(P2_READREQUEST_REG_SCAN_IN), 
        .ZN(n13038) );
  AOI21_X1 U16104 ( .B1(n18862), .B2(n13044), .A(n13038), .ZN(P2_U3612) );
  NAND2_X1 U16105 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13758) );
  CLKBUF_X2 U16106 ( .A(n19215), .Z(n19201) );
  NOR2_X1 U16107 ( .A1(n13039), .A2(n19693), .ZN(n13653) );
  OAI21_X1 U16108 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13653), .A(n13040), 
        .ZN(n13041) );
  AOI21_X1 U16109 ( .B1(n19201), .B2(n19764), .A(n13041), .ZN(n13047) );
  INV_X1 U16110 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19774) );
  AOI21_X1 U16111 ( .B1(n19693), .B2(n11027), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16338) );
  AOI21_X1 U16112 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19764), .A(n16338), 
        .ZN(n13042) );
  NOR2_X1 U16113 ( .A1(n13047), .A2(n13042), .ZN(n13046) );
  OAI21_X1 U16114 ( .B1(n10294), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19150), 
        .ZN(n13043) );
  NAND3_X1 U16115 ( .A1(n13044), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13043), 
        .ZN(n13045) );
  AOI22_X1 U16116 ( .A1(n13047), .A2(n19774), .B1(n13046), .B2(n13045), .ZN(
        P2_U3610) );
  INV_X1 U16117 ( .A(n13635), .ZN(n13048) );
  NOR2_X1 U16118 ( .A1(n13636), .A2(n13048), .ZN(n13156) );
  INV_X1 U16119 ( .A(n13156), .ZN(n13050) );
  AND2_X1 U16120 ( .A1(n13049), .A2(n19764), .ZN(n13155) );
  NOR3_X1 U16121 ( .A1(n13050), .A2(n13155), .A3(n13158), .ZN(n13642) );
  NOR2_X1 U16122 ( .A1(n13642), .A2(n13163), .ZN(n19899) );
  OAI21_X1 U16123 ( .B1(n19899), .B2(n15692), .A(n13051), .ZN(P2_U2819) );
  INV_X1 U16124 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13057) );
  NOR2_X1 U16125 ( .A1(n13052), .A2(n19778), .ZN(n13053) );
  INV_X1 U16126 ( .A(n13053), .ZN(n13054) );
  NOR2_X2 U16127 ( .A1(n13054), .A2(n10378), .ZN(n13133) );
  INV_X1 U16128 ( .A(n13133), .ZN(n13056) );
  AOI22_X1 U16129 ( .A1(n14220), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14221), .ZN(n19088) );
  INV_X1 U16130 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13055) );
  OAI222_X1 U16131 ( .A1(n13057), .A2(n13108), .B1(n13056), .B2(n19088), .C1(
        n19147), .C2(n13055), .ZN(P2_U2982) );
  NAND2_X1 U16132 ( .A1(n20718), .A2(n20643), .ZN(n19916) );
  INV_X1 U16133 ( .A(n19916), .ZN(n13846) );
  AOI21_X1 U16134 ( .B1(n13058), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13846), 
        .ZN(n13059) );
  NAND2_X1 U16135 ( .A1(n13059), .A2(n13421), .ZN(P1_U2801) );
  INV_X2 U16136 ( .A(n13108), .ZN(n13075) );
  AOI22_X1 U16137 ( .A1(n13075), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13147), .ZN(n13060) );
  AOI22_X1 U16138 ( .A1(n14220), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14221), .ZN(n13945) );
  INV_X1 U16139 ( .A(n13945), .ZN(n14952) );
  NAND2_X1 U16140 ( .A1(n13133), .A2(n14952), .ZN(n13143) );
  NAND2_X1 U16141 ( .A1(n13060), .A2(n13143), .ZN(P2_U2954) );
  AOI22_X1 U16142 ( .A1(n13075), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13147), .ZN(n13061) );
  AOI22_X1 U16143 ( .A1(n14220), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13132), .ZN(n19246) );
  INV_X1 U16144 ( .A(n19246), .ZN(n14929) );
  NAND2_X1 U16145 ( .A1(n13133), .A2(n14929), .ZN(n13145) );
  NAND2_X1 U16146 ( .A1(n13061), .A2(n13145), .ZN(P2_U2956) );
  AOI22_X1 U16147 ( .A1(n13075), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16148 ( .A1(n14220), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n13132), .ZN(n19102) );
  INV_X1 U16149 ( .A(n19102), .ZN(n13062) );
  NAND2_X1 U16150 ( .A1(n13133), .A2(n13062), .ZN(n13116) );
  NAND2_X1 U16151 ( .A1(n13063), .A2(n13116), .ZN(P2_U2977) );
  AOI22_X1 U16152 ( .A1(n13075), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16153 ( .A1(n14220), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13132), .ZN(n19260) );
  INV_X1 U16154 ( .A(n19260), .ZN(n14913) );
  NAND2_X1 U16155 ( .A1(n13133), .A2(n14913), .ZN(n13125) );
  NAND2_X1 U16156 ( .A1(n13064), .A2(n13125), .ZN(P2_U2973) );
  AOI22_X1 U16157 ( .A1(n13075), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16158 ( .A1(n14220), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13132), .ZN(n19136) );
  INV_X1 U16159 ( .A(n19136), .ZN(n14942) );
  NAND2_X1 U16160 ( .A1(n13133), .A2(n14942), .ZN(n13127) );
  NAND2_X1 U16161 ( .A1(n13065), .A2(n13127), .ZN(P2_U2970) );
  INV_X1 U16162 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19154) );
  NAND2_X1 U16163 ( .A1(n13075), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U16164 ( .A1(n14221), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13068) );
  INV_X1 U16165 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13066) );
  OR2_X1 U16166 ( .A1(n14221), .A2(n13066), .ZN(n13067) );
  NAND2_X1 U16167 ( .A1(n13068), .A2(n13067), .ZN(n19090) );
  NAND2_X1 U16168 ( .A1(n13133), .A2(n19090), .ZN(n13073) );
  OAI211_X1 U16169 ( .C1(n19154), .C2(n19147), .A(n13069), .B(n13073), .ZN(
        P2_U2966) );
  INV_X1 U16170 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19158) );
  NAND2_X1 U16171 ( .A1(n13075), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13072) );
  NAND2_X1 U16172 ( .A1(n14221), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13071) );
  INV_X1 U16173 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16455) );
  OR2_X1 U16174 ( .A1(n14221), .A2(n16455), .ZN(n13070) );
  NAND2_X1 U16175 ( .A1(n13071), .A2(n13070), .ZN(n19097) );
  NAND2_X1 U16176 ( .A1(n13133), .A2(n19097), .ZN(n13076) );
  OAI211_X1 U16177 ( .C1(n19158), .C2(n19147), .A(n13072), .B(n13076), .ZN(
        P2_U2964) );
  INV_X1 U16178 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19187) );
  NAND2_X1 U16179 ( .A1(n13075), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13074) );
  OAI211_X1 U16180 ( .C1(n19187), .C2(n19147), .A(n13074), .B(n13073), .ZN(
        P2_U2981) );
  INV_X1 U16181 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19191) );
  NAND2_X1 U16182 ( .A1(n13075), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13077) );
  OAI211_X1 U16183 ( .C1(n19191), .C2(n19147), .A(n13077), .B(n13076), .ZN(
        P2_U2979) );
  NAND2_X1 U16184 ( .A1(n13391), .A2(n13574), .ZN(n13078) );
  OAI21_X1 U16185 ( .B1(n13079), .B2(n13410), .A(n13078), .ZN(n19914) );
  NAND3_X1 U16186 ( .A1(n13574), .A2(n15689), .A3(n13349), .ZN(n13080) );
  AND2_X1 U16187 ( .A1(n13080), .A2(n20654), .ZN(n20738) );
  NOR2_X1 U16188 ( .A1(n19914), .A2(n20738), .ZN(n15655) );
  OR2_X1 U16189 ( .A1(n15655), .A2(n19913), .ZN(n13096) );
  INV_X1 U16190 ( .A(n13096), .ZN(n19922) );
  INV_X1 U16191 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13098) );
  INV_X1 U16192 ( .A(n13081), .ZN(n13083) );
  NAND2_X1 U16193 ( .A1(n13083), .A2(n13082), .ZN(n13085) );
  INV_X1 U16194 ( .A(n13279), .ZN(n14372) );
  NAND2_X1 U16195 ( .A1(n14372), .A2(n13088), .ZN(n13084) );
  NOR2_X1 U16196 ( .A1(n13087), .A2(n13086), .ZN(n13390) );
  INV_X1 U16197 ( .A(n13401), .ZN(n13259) );
  NAND2_X1 U16198 ( .A1(n20143), .A2(n13402), .ZN(n13090) );
  NAND2_X1 U16199 ( .A1(n13574), .A2(n13088), .ZN(n13089) );
  NAND2_X1 U16200 ( .A1(n13277), .A2(n13089), .ZN(n13396) );
  OAI21_X1 U16201 ( .B1(n13091), .B2(n13090), .A(n13396), .ZN(n13093) );
  INV_X1 U16202 ( .A(n13383), .ZN(n13092) );
  AOI22_X1 U16203 ( .A1(n13093), .A2(n13391), .B1(n9735), .B2(n13092), .ZN(
        n13094) );
  OAI21_X1 U16204 ( .B1(n13391), .B2(n13259), .A(n13094), .ZN(n13095) );
  NAND2_X1 U16205 ( .A1(n13095), .A2(n13580), .ZN(n15656) );
  OR2_X1 U16206 ( .A1(n13096), .A2(n15656), .ZN(n13097) );
  OAI21_X1 U16207 ( .B1(n19922), .B2(n13098), .A(n13097), .ZN(P1_U3484) );
  AOI21_X1 U16208 ( .B1(n15334), .B2(n13100), .A(n13099), .ZN(n13101) );
  INV_X1 U16209 ( .A(n13101), .ZN(n13213) );
  NAND2_X1 U16210 ( .A1(n19044), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13208) );
  OR2_X1 U16211 ( .A1(n19229), .A2(n19058), .ZN(n13102) );
  OAI211_X1 U16212 ( .C1(n13213), .C2(n19234), .A(n13208), .B(n13102), .ZN(
        n13103) );
  AOI21_X1 U16213 ( .B1(n19220), .B2(n19058), .A(n13103), .ZN(n13107) );
  OAI21_X1 U16214 ( .B1(n19056), .B2(n13171), .A(n13104), .ZN(n13105) );
  XOR2_X1 U16215 ( .A(n13105), .B(n15334), .Z(n13205) );
  NAND2_X1 U16216 ( .A1(n13205), .A2(n19222), .ZN(n13106) );
  OAI211_X1 U16217 ( .C1(n10454), .C2(n16206), .A(n13107), .B(n13106), .ZN(
        P2_U3013) );
  AOI22_X1 U16218 ( .A1(n13075), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13147), .ZN(n13110) );
  AOI22_X1 U16219 ( .A1(n14220), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n13132), .ZN(n19100) );
  INV_X1 U16220 ( .A(n19100), .ZN(n13109) );
  NAND2_X1 U16221 ( .A1(n13133), .A2(n13109), .ZN(n13123) );
  NAND2_X1 U16222 ( .A1(n13110), .A2(n13123), .ZN(P2_U2963) );
  AOI22_X1 U16223 ( .A1(n13075), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13147), .ZN(n13111) );
  AOI22_X1 U16224 ( .A1(n14220), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13132), .ZN(n19104) );
  INV_X1 U16225 ( .A(n19104), .ZN(n14884) );
  NAND2_X1 U16226 ( .A1(n13133), .A2(n14884), .ZN(n13141) );
  NAND2_X1 U16227 ( .A1(n13111), .A2(n13141), .ZN(P2_U2961) );
  AOI22_X1 U16228 ( .A1(n13075), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n13147), .ZN(n13113) );
  AOI22_X1 U16229 ( .A1(n14220), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14221), .ZN(n19106) );
  INV_X1 U16230 ( .A(n19106), .ZN(n13112) );
  NAND2_X1 U16231 ( .A1(n13133), .A2(n13112), .ZN(n13137) );
  NAND2_X1 U16232 ( .A1(n13113), .A2(n13137), .ZN(P2_U2960) );
  AOI22_X1 U16233 ( .A1(n13075), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13147), .ZN(n13115) );
  AOI22_X1 U16234 ( .A1(n14220), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13132), .ZN(n19093) );
  INV_X1 U16235 ( .A(n19093), .ZN(n13114) );
  NAND2_X1 U16236 ( .A1(n13133), .A2(n13114), .ZN(n13129) );
  NAND2_X1 U16237 ( .A1(n13115), .A2(n13129), .ZN(P2_U2965) );
  AOI22_X1 U16238 ( .A1(n13075), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n13147), .ZN(n13117) );
  NAND2_X1 U16239 ( .A1(n13117), .A2(n13116), .ZN(P2_U2962) );
  AOI22_X1 U16240 ( .A1(n13075), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16241 ( .A1(n14220), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14221), .ZN(n19250) );
  INV_X1 U16242 ( .A(n19250), .ZN(n13118) );
  NAND2_X1 U16243 ( .A1(n13133), .A2(n13118), .ZN(n13121) );
  NAND2_X1 U16244 ( .A1(n13119), .A2(n13121), .ZN(P2_U2972) );
  AOI22_X1 U16245 ( .A1(n13075), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13120) );
  OAI22_X1 U16246 ( .A1(n13132), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14220), .ZN(n13927) );
  INV_X1 U16247 ( .A(n13927), .ZN(n16189) );
  NAND2_X1 U16248 ( .A1(n13133), .A2(n16189), .ZN(n13135) );
  NAND2_X1 U16249 ( .A1(n13120), .A2(n13135), .ZN(P2_U2953) );
  AOI22_X1 U16250 ( .A1(n13075), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U16251 ( .A1(n13122), .A2(n13121), .ZN(P2_U2957) );
  AOI22_X1 U16252 ( .A1(n13075), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U16253 ( .A1(n13124), .A2(n13123), .ZN(P2_U2978) );
  AOI22_X1 U16254 ( .A1(n13075), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U16255 ( .A1(n13126), .A2(n13125), .ZN(P2_U2958) );
  AOI22_X1 U16256 ( .A1(n13075), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U16257 ( .A1(n13128), .A2(n13127), .ZN(P2_U2955) );
  AOI22_X1 U16258 ( .A1(n13075), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16259 ( .A1(n13130), .A2(n13129), .ZN(P2_U2980) );
  AOI22_X1 U16260 ( .A1(n13075), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16261 ( .A1(n14220), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14221), .ZN(n19108) );
  INV_X1 U16262 ( .A(n19108), .ZN(n14902) );
  NAND2_X1 U16263 ( .A1(n13133), .A2(n14902), .ZN(n13148) );
  NAND2_X1 U16264 ( .A1(n13131), .A2(n13148), .ZN(P2_U2974) );
  AOI22_X1 U16265 ( .A1(n13075), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U16266 ( .A1(n14220), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13132), .ZN(n19146) );
  INV_X1 U16267 ( .A(n19146), .ZN(n14958) );
  NAND2_X1 U16268 ( .A1(n13133), .A2(n14958), .ZN(n13139) );
  NAND2_X1 U16269 ( .A1(n13134), .A2(n13139), .ZN(P2_U2952) );
  AOI22_X1 U16270 ( .A1(n13075), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13136) );
  NAND2_X1 U16271 ( .A1(n13136), .A2(n13135), .ZN(P2_U2968) );
  AOI22_X1 U16272 ( .A1(n13075), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13138) );
  NAND2_X1 U16273 ( .A1(n13138), .A2(n13137), .ZN(P2_U2975) );
  AOI22_X1 U16274 ( .A1(n13075), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U16275 ( .A1(n13140), .A2(n13139), .ZN(P2_U2967) );
  AOI22_X1 U16276 ( .A1(n13075), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U16277 ( .A1(n13142), .A2(n13141), .ZN(P2_U2976) );
  AOI22_X1 U16278 ( .A1(n13075), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13144) );
  NAND2_X1 U16279 ( .A1(n13144), .A2(n13143), .ZN(P2_U2969) );
  AOI22_X1 U16280 ( .A1(n13075), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13146) );
  NAND2_X1 U16281 ( .A1(n13146), .A2(n13145), .ZN(P2_U2971) );
  AOI22_X1 U16282 ( .A1(n13075), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13147), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U16283 ( .A1(n13149), .A2(n13148), .ZN(P2_U2959) );
  NOR2_X1 U16284 ( .A1(n14364), .A2(n14256), .ZN(n13151) );
  OAI21_X1 U16285 ( .B1(n13846), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20733), 
        .ZN(n13150) );
  OAI21_X1 U16286 ( .B1(n20733), .B2(n13151), .A(n13150), .ZN(P1_U3487) );
  INV_X1 U16287 ( .A(n13152), .ZN(n13153) );
  AND2_X1 U16288 ( .A1(n13154), .A2(n13153), .ZN(n13162) );
  AOI22_X1 U16289 ( .A1(n13641), .A2(n13553), .B1(n13156), .B2(n13155), .ZN(
        n13224) );
  INV_X1 U16290 ( .A(n19149), .ZN(n13160) );
  INV_X1 U16291 ( .A(n13157), .ZN(n13159) );
  NAND3_X1 U16292 ( .A1(n13160), .A2(n13159), .A3(n13158), .ZN(n13161) );
  AND3_X1 U16293 ( .A1(n13162), .A2(n13224), .A3(n13161), .ZN(n13647) );
  INV_X1 U16294 ( .A(n13758), .ZN(n19893) );
  NAND2_X1 U16295 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19893), .ZN(n16339) );
  OAI22_X1 U16296 ( .A1(n13647), .A2(n13163), .B1(n15692), .B2(n16339), .ZN(
        n13164) );
  AOI21_X1 U16297 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n12960), .A(n13164), 
        .ZN(n19855) );
  INV_X1 U16298 ( .A(n19855), .ZN(n19857) );
  INV_X1 U16299 ( .A(n13165), .ZN(n13166) );
  NOR2_X1 U16300 ( .A1(n11106), .A2(n13166), .ZN(n13643) );
  NAND4_X1 U16301 ( .A1(n11135), .A2(n19857), .A3(n13643), .A4(n19850), .ZN(
        n13167) );
  OAI21_X1 U16302 ( .B1(n19857), .B2(n13168), .A(n13167), .ZN(P2_U3595) );
  OAI21_X1 U16303 ( .B1(n13170), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13169), .ZN(n19233) );
  OAI21_X1 U16304 ( .B1(n14017), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13171), .ZN(n19235) );
  OAI22_X1 U16305 ( .A1(n16317), .A2(n19235), .B1(n16329), .B2(n14013), .ZN(
        n13172) );
  AOI21_X1 U16306 ( .B1(n13177), .B2(n15264), .A(n13172), .ZN(n13180) );
  NOR2_X1 U16307 ( .A1(n13174), .A2(n13173), .ZN(n13175) );
  NOR2_X1 U16308 ( .A1(n13176), .A2(n13175), .ZN(n19141) );
  NAND2_X1 U16309 ( .A1(n19044), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19232) );
  OAI21_X1 U16310 ( .B1(n13177), .B2(n13209), .A(n19232), .ZN(n13178) );
  AOI21_X1 U16311 ( .B1(n16301), .B2(n19141), .A(n13178), .ZN(n13179) );
  OAI211_X1 U16312 ( .C1(n16330), .C2(n19233), .A(n13180), .B(n13179), .ZN(
        P2_U3046) );
  NAND2_X1 U16313 ( .A1(n13182), .A2(n13181), .ZN(n13184) );
  AND2_X1 U16314 ( .A1(n13184), .A2(n10120), .ZN(n19114) );
  INV_X1 U16315 ( .A(n19114), .ZN(n19874) );
  AOI21_X1 U16316 ( .B1(n13187), .B2(n13186), .A(n13185), .ZN(n13221) );
  NAND2_X1 U16317 ( .A1(n13221), .A2(n16313), .ZN(n13194) );
  INV_X1 U16318 ( .A(n15238), .ZN(n13188) );
  OAI21_X1 U16319 ( .B1(n13737), .B2(n13189), .A(n13188), .ZN(n13193) );
  NAND2_X1 U16320 ( .A1(n19044), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13215) );
  NAND2_X1 U16321 ( .A1(n13191), .A2(n13190), .ZN(n13217) );
  NAND3_X1 U16322 ( .A1(n16334), .A2(n13218), .A3(n13217), .ZN(n13192) );
  NAND4_X1 U16323 ( .A1(n13194), .A2(n13193), .A3(n13215), .A4(n13192), .ZN(
        n13200) );
  AOI21_X1 U16324 ( .B1(n15240), .B2(n13206), .A(n13195), .ZN(n13198) );
  OAI22_X1 U16325 ( .A1(n13198), .A2(n13197), .B1(n13196), .B2(n13206), .ZN(
        n13199) );
  AOI211_X1 U16326 ( .C1(n19874), .C2(n16301), .A(n13200), .B(n13199), .ZN(
        n13201) );
  OAI21_X1 U16327 ( .B1(n10500), .B2(n16329), .A(n13201), .ZN(P2_U3044) );
  AOI21_X1 U16328 ( .B1(n13204), .B2(n13203), .A(n13202), .ZN(n19879) );
  INV_X1 U16329 ( .A(n19879), .ZN(n13239) );
  AOI22_X1 U16330 ( .A1(n16301), .A2(n13239), .B1(n16334), .B2(n13205), .ZN(
        n13212) );
  OAI211_X1 U16331 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15264), .B(n13206), .ZN(n13207) );
  OAI211_X1 U16332 ( .C1(n13209), .C2(n15334), .A(n13208), .B(n13207), .ZN(
        n13210) );
  AOI21_X1 U16333 ( .B1(n19068), .B2(n16312), .A(n13210), .ZN(n13211) );
  OAI211_X1 U16334 ( .C1(n16330), .C2(n13213), .A(n13212), .B(n13211), .ZN(
        P2_U3045) );
  INV_X1 U16335 ( .A(n13820), .ZN(n13216) );
  NAND2_X1 U16336 ( .A1(n19230), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13214) );
  OAI211_X1 U16337 ( .C1(n16256), .C2(n13216), .A(n13215), .B(n13214), .ZN(
        n13220) );
  AND3_X1 U16338 ( .A1(n13218), .A2(n19222), .A3(n13217), .ZN(n13219) );
  AOI211_X1 U16339 ( .C1(n13221), .C2(n19224), .A(n13220), .B(n13219), .ZN(
        n13222) );
  OAI21_X1 U16340 ( .B1(n10500), .B2(n16206), .A(n13222), .ZN(P2_U3012) );
  NAND2_X1 U16341 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  AND2_X1 U16342 ( .A1(n12586), .A2(n13931), .ZN(n13226) );
  NAND2_X1 U16343 ( .A1(n19111), .A2(n13226), .ZN(n14222) );
  INV_X1 U16344 ( .A(n14222), .ZN(n13229) );
  AND2_X1 U16345 ( .A1(n13227), .A2(n13931), .ZN(n13228) );
  OR2_X1 U16346 ( .A1(n13229), .A2(n16190), .ZN(n19096) );
  XNOR2_X1 U16347 ( .A(n19883), .B(n19879), .ZN(n13236) );
  NAND2_X1 U16348 ( .A1(n11215), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13234) );
  AND4_X1 U16349 ( .A1(n9646), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13234), 
        .A4(n19888), .ZN(n13235) );
  NAND2_X1 U16350 ( .A1(n19142), .A2(n19141), .ZN(n19140) );
  NAND2_X1 U16351 ( .A1(n13236), .A2(n19140), .ZN(n13491) );
  OAI21_X1 U16352 ( .B1(n13236), .B2(n19140), .A(n13491), .ZN(n13237) );
  NAND2_X1 U16353 ( .A1(n13237), .A2(n19139), .ZN(n13241) );
  AOI22_X1 U16354 ( .A1(n19138), .A2(n13239), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19137), .ZN(n13240) );
  OAI211_X1 U16355 ( .C1(n19145), .C2(n13927), .A(n13241), .B(n13240), .ZN(
        P2_U2918) );
  INV_X1 U16356 ( .A(n14751), .ZN(n13242) );
  AOI21_X1 U16357 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13242), .A(
        n13258), .ZN(n13243) );
  NAND2_X1 U16358 ( .A1(n11580), .A2(n13243), .ZN(n13269) );
  NAND2_X1 U16359 ( .A1(n13244), .A2(n13245), .ZN(n13246) );
  NOR2_X1 U16360 ( .A1(n13247), .A2(n13246), .ZN(n13256) );
  NAND2_X1 U16361 ( .A1(n13248), .A2(n14364), .ZN(n13254) );
  OAI21_X1 U16362 ( .B1(n13249), .B2(n13346), .A(n13580), .ZN(n13250) );
  OAI21_X1 U16363 ( .B1(n13250), .B2(n13347), .A(n13422), .ZN(n13251) );
  AND2_X1 U16364 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  AND2_X1 U16365 ( .A1(n13254), .A2(n13253), .ZN(n13408) );
  AND3_X1 U16366 ( .A1(n13256), .A2(n13408), .A3(n13255), .ZN(n14757) );
  INV_X1 U16367 ( .A(n14757), .ZN(n13523) );
  NAND2_X1 U16368 ( .A1(n20711), .A2(n13523), .ZN(n13268) );
  NAND2_X1 U16369 ( .A1(n14757), .A2(n13347), .ZN(n13520) );
  INV_X1 U16370 ( .A(n13520), .ZN(n13266) );
  AOI21_X1 U16371 ( .B1(n13261), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13258), .ZN(n13264) );
  NAND2_X1 U16372 ( .A1(n9735), .A2(n13422), .ZN(n13516) );
  NOR2_X1 U16373 ( .A1(n13516), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14753) );
  NAND2_X1 U16374 ( .A1(n14753), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13263) );
  MUX2_X1 U16375 ( .A(n13258), .B(n13257), .S(n14751), .Z(n13260) );
  NAND2_X1 U16376 ( .A1(n13277), .A2(n14364), .ZN(n13272) );
  NAND2_X1 U16377 ( .A1(n13259), .A2(n13272), .ZN(n13518) );
  OAI21_X1 U16378 ( .B1(n13261), .B2(n13260), .A(n13518), .ZN(n13262) );
  OAI211_X1 U16379 ( .C1(n13264), .C2(n13516), .A(n13263), .B(n13262), .ZN(
        n13265) );
  AOI21_X1 U16380 ( .B1(n13266), .B2(n13269), .A(n13265), .ZN(n13267) );
  NAND2_X1 U16381 ( .A1(n13268), .A2(n13267), .ZN(n15641) );
  AOI22_X1 U16382 ( .A1(n15671), .A2(n13269), .B1(n16083), .B2(n15641), .ZN(
        n13290) );
  NAND2_X1 U16383 ( .A1(n13516), .A2(n13244), .ZN(n13271) );
  NAND2_X1 U16384 ( .A1(n13271), .A2(n13270), .ZN(n13315) );
  INV_X1 U16385 ( .A(n20654), .ZN(n20736) );
  OR2_X1 U16386 ( .A1(n13391), .A2(n20736), .ZN(n13284) );
  OAI21_X1 U16387 ( .B1(n13273), .B2(n20736), .A(n13272), .ZN(n13274) );
  NAND2_X1 U16388 ( .A1(n13274), .A2(n13386), .ZN(n13276) );
  INV_X1 U16389 ( .A(n13255), .ZN(n16082) );
  NAND3_X1 U16390 ( .A1(n16082), .A2(n13383), .A3(n20654), .ZN(n13275) );
  OAI21_X1 U16391 ( .B1(n9735), .B2(n13277), .A(n13406), .ZN(n13389) );
  NOR2_X1 U16392 ( .A1(n13279), .A2(n13278), .ZN(n13280) );
  OR2_X1 U16393 ( .A1(n13389), .A2(n13280), .ZN(n13282) );
  NAND2_X1 U16394 ( .A1(n13401), .A2(n13391), .ZN(n13351) );
  INV_X1 U16395 ( .A(n13351), .ZN(n13281) );
  NOR2_X1 U16396 ( .A1(n13282), .A2(n13281), .ZN(n13283) );
  OAI211_X1 U16397 ( .C1(n13315), .C2(n13284), .A(n13577), .B(n13283), .ZN(
        n15646) );
  NAND2_X1 U16398 ( .A1(n15646), .A2(n13578), .ZN(n13287) );
  NAND2_X1 U16399 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16092) );
  INV_X1 U16400 ( .A(n16092), .ZN(n14747) );
  NAND2_X1 U16401 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14747), .ZN(n16096) );
  INV_X1 U16402 ( .A(n16096), .ZN(n13285) );
  NAND2_X1 U16403 ( .A1(n13285), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13286) );
  NAND2_X1 U16404 ( .A1(n13287), .A2(n13286), .ZN(n16081) );
  AND2_X1 U16405 ( .A1(n20644), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13288) );
  OR2_X1 U16406 ( .A1(n16081), .A2(n13288), .ZN(n16087) );
  INV_X1 U16407 ( .A(n16087), .ZN(n13304) );
  NAND2_X1 U16408 ( .A1(n13304), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13289) );
  OAI21_X1 U16409 ( .B1(n13290), .B2(n13304), .A(n13289), .ZN(P1_U3469) );
  MUX2_X1 U16410 ( .A(n13295), .B(n10500), .S(n14844), .Z(n13296) );
  OAI21_X1 U16411 ( .B1(n19872), .B2(n16181), .A(n13296), .ZN(P2_U2885) );
  MUX2_X1 U16412 ( .A(n10643), .B(n14013), .S(n14844), .Z(n13297) );
  OAI21_X1 U16413 ( .B1(n19890), .B2(n16181), .A(n13297), .ZN(P2_U2887) );
  INV_X1 U16414 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n19054) );
  NOR2_X1 U16415 ( .A1(n14844), .A2(n19054), .ZN(n13298) );
  AOI21_X1 U16416 ( .B1(n19068), .B2(n14844), .A(n13298), .ZN(n13299) );
  OAI21_X1 U16417 ( .B1(n19854), .B2(n16181), .A(n13299), .ZN(P2_U2886) );
  NOR2_X1 U16418 ( .A1(n11557), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13300) );
  AOI21_X1 U16419 ( .B1(n11689), .B2(n13523), .A(n13300), .ZN(n15645) );
  INV_X1 U16420 ( .A(n16083), .ZN(n13301) );
  OAI22_X1 U16421 ( .A1(n15645), .A2(n13301), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20643), .ZN(n13302) );
  AOI21_X1 U16422 ( .B1(n15671), .B2(n11419), .A(n13302), .ZN(n13305) );
  NOR2_X1 U16423 ( .A1(n13516), .A2(n11419), .ZN(n15643) );
  AOI22_X1 U16424 ( .A1(n13304), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n16083), .B2(n15643), .ZN(n13303) );
  OAI21_X1 U16425 ( .B1(n13305), .B2(n13304), .A(n13303), .ZN(P1_U3474) );
  AND2_X1 U16426 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13308) );
  NAND2_X1 U16427 ( .A1(n13306), .A2(n13308), .ZN(n13367) );
  OR2_X1 U16428 ( .A1(n13306), .A2(n13308), .ZN(n13309) );
  NAND2_X1 U16429 ( .A1(n13367), .A2(n13309), .ZN(n19125) );
  NOR2_X1 U16430 ( .A1(n13311), .A2(n13310), .ZN(n13312) );
  OR2_X1 U16431 ( .A1(n13469), .A2(n13312), .ZN(n13811) );
  MUX2_X1 U16432 ( .A(n13313), .B(n13811), .S(n14844), .Z(n13314) );
  OAI21_X1 U16433 ( .B1(n19125), .B2(n16181), .A(n13314), .ZN(P2_U2883) );
  INV_X1 U16434 ( .A(n13516), .ZN(n13400) );
  INV_X1 U16435 ( .A(n13315), .ZN(n13318) );
  INV_X1 U16436 ( .A(n13316), .ZN(n13317) );
  INV_X1 U16437 ( .A(n20033), .ZN(n13320) );
  NAND2_X1 U16438 ( .A1(n13320), .A2(n13402), .ZN(n13341) );
  NAND2_X1 U16439 ( .A1(n20644), .A2(n14747), .ZN(n20735) );
  INV_X2 U16440 ( .A(n20735), .ZN(n20031) );
  AOI22_X1 U16441 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13321) );
  OAI21_X1 U16442 ( .B1(n14517), .B2(n13341), .A(n13321), .ZN(P1_U2910) );
  INV_X1 U16443 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16444 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13322) );
  OAI21_X1 U16445 ( .B1(n13323), .B2(n13341), .A(n13322), .ZN(P1_U2908) );
  AOI22_X1 U16446 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13324) );
  OAI21_X1 U16447 ( .B1(n14525), .B2(n13341), .A(n13324), .ZN(P1_U2912) );
  AOI22_X1 U16448 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13325) );
  OAI21_X1 U16449 ( .B1(n14542), .B2(n13341), .A(n13325), .ZN(P1_U2916) );
  AOI22_X1 U16450 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13326) );
  OAI21_X1 U16451 ( .B1(n14549), .B2(n13341), .A(n13326), .ZN(P1_U2918) );
  INV_X1 U16452 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U16453 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13327) );
  OAI21_X1 U16454 ( .B1(n13328), .B2(n13341), .A(n13327), .ZN(P1_U2917) );
  INV_X1 U16455 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13330) );
  AOI22_X1 U16456 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13329) );
  OAI21_X1 U16457 ( .B1(n13330), .B2(n13341), .A(n13329), .ZN(P1_U2915) );
  INV_X1 U16458 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U16459 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13331) );
  OAI21_X1 U16460 ( .B1(n13332), .B2(n13341), .A(n13331), .ZN(P1_U2909) );
  INV_X1 U16461 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20770) );
  AOI22_X1 U16462 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16463 ( .B1(n20770), .B2(n13341), .A(n13333), .ZN(P1_U2906) );
  INV_X1 U16464 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13335) );
  AOI22_X1 U16465 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13334) );
  OAI21_X1 U16466 ( .B1(n13335), .B2(n13341), .A(n13334), .ZN(P1_U2911) );
  AOI22_X1 U16467 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13336) );
  OAI21_X1 U16468 ( .B1(n14534), .B2(n13341), .A(n13336), .ZN(P1_U2914) );
  AOI22_X1 U16469 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13337) );
  OAI21_X1 U16470 ( .B1(n14530), .B2(n13341), .A(n13337), .ZN(P1_U2913) );
  AOI22_X1 U16471 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13338) );
  OAI21_X1 U16472 ( .B1(n14553), .B2(n13341), .A(n13338), .ZN(P1_U2919) );
  AOI22_X1 U16473 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13339) );
  OAI21_X1 U16474 ( .B1(n14558), .B2(n13341), .A(n13339), .ZN(P1_U2920) );
  INV_X1 U16475 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U16476 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13340) );
  OAI21_X1 U16477 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(P1_U2907) );
  INV_X1 U16478 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20094) );
  INV_X1 U16479 ( .A(n13343), .ZN(n13344) );
  AOI21_X1 U16480 ( .B1(n13345), .B2(n20094), .A(n13344), .ZN(n20088) );
  INV_X1 U16481 ( .A(n20088), .ZN(n13358) );
  INV_X1 U16482 ( .A(n13580), .ZN(n20147) );
  NAND4_X1 U16483 ( .A1(n13348), .A2(n13347), .A3(n20147), .A4(n13346), .ZN(
        n13575) );
  OR2_X1 U16484 ( .A1(n13575), .A2(n13349), .ZN(n13350) );
  NAND2_X1 U16485 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  INV_X1 U16486 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13357) );
  INV_X1 U16487 ( .A(n13353), .ZN(n13356) );
  OAI21_X1 U16488 ( .B1(n13356), .B2(n13355), .A(n13354), .ZN(n20072) );
  INV_X2 U16489 ( .A(n20004), .ZN(n14492) );
  OAI222_X1 U16490 ( .A1(n13358), .A2(n14494), .B1(n13357), .B2(n20008), .C1(
        n20072), .C2(n14492), .ZN(P1_U2872) );
  OAI21_X1 U16491 ( .B1(n13361), .B2(n13360), .A(n13359), .ZN(n19992) );
  OR2_X1 U16492 ( .A1(n19982), .A2(n13362), .ZN(n13363) );
  AND2_X1 U16493 ( .A1(n13364), .A2(n13363), .ZN(n13415) );
  INV_X1 U16494 ( .A(n13415), .ZN(n13365) );
  AOI22_X1 U16495 ( .A1(n20003), .A2(n13365), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14483), .ZN(n13366) );
  OAI21_X1 U16496 ( .B1(n19992), .B2(n14492), .A(n13366), .ZN(P1_U2871) );
  INV_X1 U16497 ( .A(n13367), .ZN(n13467) );
  NAND2_X1 U16498 ( .A1(n13467), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13475) );
  XOR2_X1 U16499 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(n13475), .Z(n13372)
         );
  INV_X1 U16500 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U16501 ( .B1(n13368), .B2(n13369), .A(n13478), .ZN(n19032) );
  MUX2_X1 U16502 ( .A(n13370), .B(n19032), .S(n14844), .Z(n13371) );
  OAI21_X1 U16503 ( .B1(n13372), .B2(n16181), .A(n13371), .ZN(P2_U2881) );
  NOR2_X1 U16504 ( .A1(n10490), .A2(n19078), .ZN(n13375) );
  AOI21_X1 U16505 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19078), .A(n13375), .ZN(
        n13376) );
  OAI21_X1 U16506 ( .B1(n19113), .B2(n16181), .A(n13376), .ZN(P2_U2884) );
  XNOR2_X1 U16507 ( .A(n13377), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13419) );
  INV_X1 U16508 ( .A(n19992), .ZN(n13380) );
  AOI22_X1 U16509 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13378) );
  OAI21_X1 U16510 ( .B1(n15899), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13378), .ZN(n13379) );
  AOI21_X1 U16511 ( .B1(n13380), .B2(n15894), .A(n13379), .ZN(n13381) );
  OAI21_X1 U16512 ( .B1(n13419), .B2(n19920), .A(n13381), .ZN(P1_U2998) );
  AOI21_X1 U16513 ( .B1(n13422), .B2(n15689), .A(n20736), .ZN(n13382) );
  NAND2_X1 U16514 ( .A1(n13383), .A2(n13382), .ZN(n13388) );
  OAI211_X1 U16515 ( .C1(n13244), .C2(n13384), .A(n13402), .B(n13584), .ZN(
        n13385) );
  MUX2_X1 U16516 ( .A(n13388), .B(n13387), .S(n13249), .Z(n13394) );
  INV_X1 U16517 ( .A(n13389), .ZN(n13393) );
  NAND2_X1 U16518 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  NAND3_X1 U16519 ( .A1(n13394), .A2(n13393), .A3(n13392), .ZN(n13395) );
  INV_X1 U16520 ( .A(n13411), .ZN(n13398) );
  OAI211_X1 U16521 ( .C1(n20135), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        n13399) );
  NAND2_X1 U16522 ( .A1(n13403), .A2(n13402), .ZN(n13405) );
  AOI21_X1 U16523 ( .B1(n13405), .B2(n14256), .A(n13404), .ZN(n13407) );
  NAND3_X1 U16524 ( .A1(n13408), .A2(n13407), .A3(n13406), .ZN(n13409) );
  AOI21_X1 U16525 ( .B1(n20094), .B2(n14699), .A(n16048), .ZN(n13417) );
  OAI22_X1 U16526 ( .A1(n13414), .A2(n20074), .B1(n20092), .B2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15973) );
  INV_X1 U16527 ( .A(n15973), .ZN(n20078) );
  OAI21_X1 U16528 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20093), .A(
        n20078), .ZN(n20096) );
  NAND2_X1 U16529 ( .A1(n13410), .A2(n20124), .ZN(n15664) );
  NAND2_X1 U16530 ( .A1(n13411), .A2(n20135), .ZN(n13412) );
  NAND2_X1 U16531 ( .A1(n15664), .A2(n13412), .ZN(n13413) );
  INV_X1 U16532 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20724) );
  OAI22_X1 U16533 ( .A1(n13415), .A2(n16079), .B1(n16057), .B2(n20724), .ZN(
        n13416) );
  AOI221_X1 U16534 ( .B1(n13417), .B2(n12422), .C1(n20096), .C2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n13416), .ZN(n13418) );
  OAI21_X1 U16535 ( .B1(n13419), .B2(n16073), .A(n13418), .ZN(P1_U3030) );
  AND2_X1 U16536 ( .A1(n20739), .A2(n20736), .ZN(n13420) );
  AND2_X2 U16537 ( .A1(n13448), .A2(n20124), .ZN(n20061) );
  INV_X2 U16538 ( .A(n13448), .ZN(n20060) );
  AOI22_X1 U16539 ( .A1(n20061), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U16540 ( .A1(n13448), .A2(n13422), .ZN(n13449) );
  INV_X1 U16541 ( .A(n20102), .ZN(n20103) );
  INV_X1 U16542 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13423) );
  NOR2_X1 U16543 ( .A1(n20103), .A2(n13423), .ZN(n13424) );
  AOI21_X1 U16544 ( .B1(DATAI_7_), .B2(n20103), .A(n13424), .ZN(n20152) );
  INV_X1 U16545 ( .A(n20152), .ZN(n13425) );
  NAND2_X1 U16546 ( .A1(n20048), .A2(n13425), .ZN(n13694) );
  NAND2_X1 U16547 ( .A1(n13426), .A2(n13694), .ZN(P1_U2944) );
  AOI22_X1 U16548 ( .A1(n20061), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13430) );
  INV_X1 U16549 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13427) );
  NOR2_X1 U16550 ( .A1(n20103), .A2(n13427), .ZN(n13428) );
  AOI21_X1 U16551 ( .B1(DATAI_0_), .B2(n20103), .A(n13428), .ZN(n20117) );
  INV_X1 U16552 ( .A(n20117), .ZN(n13429) );
  NAND2_X1 U16553 ( .A1(n20048), .A2(n13429), .ZN(n13680) );
  NAND2_X1 U16554 ( .A1(n13430), .A2(n13680), .ZN(P1_U2937) );
  AOI22_X1 U16555 ( .A1(n20061), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U16556 ( .A1(n20103), .A2(DATAI_4_), .ZN(n13432) );
  NAND2_X1 U16557 ( .A1(n20102), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13431) );
  AND2_X1 U16558 ( .A1(n13432), .A2(n13431), .ZN(n20136) );
  INV_X1 U16559 ( .A(n20136), .ZN(n13433) );
  NAND2_X1 U16560 ( .A1(n20048), .A2(n13433), .ZN(n13435) );
  NAND2_X1 U16561 ( .A1(n13434), .A2(n13435), .ZN(P1_U2956) );
  AOI22_X1 U16562 ( .A1(n20061), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U16563 ( .A1(n13436), .A2(n13435), .ZN(P1_U2941) );
  INV_X1 U16564 ( .A(n20061), .ZN(n13450) );
  INV_X1 U16565 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20021) );
  NAND2_X1 U16566 ( .A1(n20060), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13440) );
  INV_X1 U16567 ( .A(DATAI_8_), .ZN(n13438) );
  INV_X1 U16568 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13437) );
  MUX2_X1 U16569 ( .A(n13438), .B(n13437), .S(n20102), .Z(n14526) );
  INV_X1 U16570 ( .A(n14526), .ZN(n13439) );
  NAND2_X1 U16571 ( .A1(n20048), .A2(n13439), .ZN(n13444) );
  OAI211_X1 U16572 ( .C1(n13450), .C2(n20021), .A(n13440), .B(n13444), .ZN(
        P1_U2960) );
  INV_X1 U16573 ( .A(DATAI_14_), .ZN(n13442) );
  NAND2_X1 U16574 ( .A1(n20102), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13441) );
  OAI21_X1 U16575 ( .B1(n20102), .B2(n13442), .A(n13441), .ZN(n14495) );
  NAND2_X1 U16576 ( .A1(n20048), .A2(n14495), .ZN(n20062) );
  NAND2_X1 U16577 ( .A1(n20060), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13443) );
  OAI211_X1 U16578 ( .C1(n13450), .C2(n20770), .A(n20062), .B(n13443), .ZN(
        P1_U2951) );
  NAND2_X1 U16579 ( .A1(n20060), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13445) );
  OAI211_X1 U16580 ( .C1(n13450), .C2(n14525), .A(n13445), .B(n13444), .ZN(
        P1_U2945) );
  INV_X1 U16581 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20011) );
  INV_X1 U16582 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13446) );
  NOR2_X1 U16583 ( .A1(n20103), .A2(n13446), .ZN(n13447) );
  AOI21_X1 U16584 ( .B1(DATAI_15_), .B2(n20103), .A(n13447), .ZN(n14566) );
  INV_X1 U16585 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20012) );
  OAI222_X1 U16586 ( .A1(n13450), .A2(n20011), .B1(n13449), .B2(n14566), .C1(
        n13448), .C2(n20012), .ZN(P1_U2967) );
  INV_X1 U16587 ( .A(n13451), .ZN(n13454) );
  OAI211_X1 U16588 ( .C1(n13454), .C2(n12616), .A(n19079), .B(n13453), .ZN(
        n13458) );
  NOR2_X1 U16589 ( .A1(n13463), .A2(n13483), .ZN(n13462) );
  OR2_X1 U16590 ( .A1(n13455), .A2(n13462), .ZN(n13456) );
  AND2_X1 U16591 ( .A1(n9764), .A2(n13456), .ZN(n18998) );
  NAND2_X1 U16592 ( .A1(n14844), .A2(n18998), .ZN(n13457) );
  OAI211_X1 U16593 ( .C1(n14844), .C2(n10040), .A(n13458), .B(n13457), .ZN(
        P2_U2877) );
  INV_X1 U16594 ( .A(n13459), .ZN(n13461) );
  OAI211_X1 U16595 ( .C1(n13461), .C2(n12615), .A(n19079), .B(n13451), .ZN(
        n13465) );
  AOI21_X1 U16596 ( .B1(n13463), .B2(n13483), .A(n13462), .ZN(n19009) );
  NAND2_X1 U16597 ( .A1(n14844), .A2(n19009), .ZN(n13464) );
  OAI211_X1 U16598 ( .C1(n14844), .C2(n13466), .A(n13465), .B(n13464), .ZN(
        P2_U2878) );
  OAI211_X1 U16599 ( .C1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .C2(n13467), .A(
        n13475), .B(n19079), .ZN(n13473) );
  INV_X1 U16600 ( .A(n13468), .ZN(n13471) );
  INV_X1 U16601 ( .A(n13469), .ZN(n13470) );
  AOI21_X1 U16602 ( .B1(n13471), .B2(n13470), .A(n13368), .ZN(n19050) );
  NAND2_X1 U16603 ( .A1(n19050), .A2(n14844), .ZN(n13472) );
  OAI211_X1 U16604 ( .C1(n14844), .C2(n19041), .A(n13473), .B(n13472), .ZN(
        P2_U2882) );
  NOR2_X1 U16605 ( .A1(n13475), .A2(n13474), .ZN(n13477) );
  INV_X1 U16606 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13935) );
  NOR3_X1 U16607 ( .A1(n13475), .A2(n13935), .A3(n13474), .ZN(n13488) );
  INV_X1 U16608 ( .A(n13488), .ZN(n13476) );
  OAI211_X1 U16609 ( .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n13477), .A(
        n13476), .B(n19079), .ZN(n13481) );
  AOI21_X1 U16610 ( .B1(n13479), .B2(n13478), .A(n13484), .ZN(n19019) );
  NAND2_X1 U16611 ( .A1(n14844), .A2(n19019), .ZN(n13480) );
  OAI211_X1 U16612 ( .C1(n14844), .C2(n13482), .A(n13481), .B(n13480), .ZN(
        P2_U2880) );
  OAI21_X1 U16613 ( .B1(n13485), .B2(n13484), .A(n13483), .ZN(n16328) );
  INV_X1 U16614 ( .A(n13486), .ZN(n13487) );
  OAI211_X1 U16615 ( .C1(n13488), .C2(n13487), .A(n19079), .B(n13459), .ZN(
        n13490) );
  NAND2_X1 U16616 ( .A1(n19078), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13489) );
  OAI211_X1 U16617 ( .C1(n16328), .C2(n19078), .A(n13490), .B(n13489), .ZN(
        P2_U2879) );
  XOR2_X1 U16618 ( .A(n19114), .B(n19872), .Z(n13494) );
  NAND2_X1 U16619 ( .A1(n19854), .A2(n19879), .ZN(n13492) );
  NAND2_X1 U16620 ( .A1(n13492), .A2(n13491), .ZN(n13493) );
  NAND2_X1 U16621 ( .A1(n13494), .A2(n13493), .ZN(n19115) );
  OAI21_X1 U16622 ( .B1(n13494), .B2(n13493), .A(n19115), .ZN(n13495) );
  NAND2_X1 U16623 ( .A1(n13495), .A2(n19139), .ZN(n13497) );
  AOI22_X1 U16624 ( .A1(n19096), .A2(n14952), .B1(n19137), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13496) );
  OAI211_X1 U16625 ( .C1(n19114), .C2(n14962), .A(n13497), .B(n13496), .ZN(
        P2_U2917) );
  XOR2_X1 U16626 ( .A(n13499), .B(n13498), .Z(n20081) );
  INV_X1 U16627 ( .A(n20081), .ZN(n13506) );
  NAND2_X1 U16628 ( .A1(n13500), .A2(n13359), .ZN(n13501) );
  AND2_X1 U16629 ( .A1(n13502), .A2(n13501), .ZN(n20005) );
  AOI22_X1 U16630 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13503) );
  OAI21_X1 U16631 ( .B1(n15899), .B2(n14396), .A(n13503), .ZN(n13504) );
  AOI21_X1 U16632 ( .B1(n20005), .B2(n15894), .A(n13504), .ZN(n13505) );
  OAI21_X1 U16633 ( .B1(n13506), .B2(n19920), .A(n13505), .ZN(P1_U2997) );
  INV_X1 U16634 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13514) );
  INV_X1 U16635 ( .A(n13453), .ZN(n13509) );
  OAI211_X1 U16636 ( .C1(n13509), .C2(n10113), .A(n19079), .B(n13508), .ZN(
        n13513) );
  NAND2_X1 U16637 ( .A1(n9764), .A2(n13510), .ZN(n13511) );
  AND2_X1 U16638 ( .A1(n13659), .A2(n13511), .ZN(n18985) );
  NAND2_X1 U16639 ( .A1(n14844), .A2(n18985), .ZN(n13512) );
  OAI211_X1 U16640 ( .C1(n14844), .C2(n13514), .A(n13513), .B(n13512), .ZN(
        P2_U2876) );
  INV_X1 U16641 ( .A(n13515), .ZN(n20112) );
  NOR2_X1 U16642 ( .A1(n13516), .A2(n9829), .ZN(n13517) );
  MUX2_X1 U16643 ( .A(n13517), .B(n14753), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13522) );
  XNOR2_X1 U16644 ( .A(n14751), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14766) );
  NAND2_X1 U16645 ( .A1(n13518), .A2(n14766), .ZN(n13519) );
  OAI21_X1 U16646 ( .B1(n13520), .B2(n14766), .A(n13519), .ZN(n13521) );
  AOI211_X1 U16647 ( .C1(n20112), .C2(n13523), .A(n13522), .B(n13521), .ZN(
        n13524) );
  INV_X1 U16648 ( .A(n13524), .ZN(n15642) );
  INV_X1 U16649 ( .A(n15646), .ZN(n13536) );
  AOI21_X1 U16650 ( .B1(n15641), .B2(n15642), .A(n13536), .ZN(n13525) );
  INV_X1 U16651 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19921) );
  NAND2_X1 U16652 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n19921), .ZN(n13533) );
  OAI21_X1 U16653 ( .B1(n13525), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n13533), 
        .ZN(n13529) );
  NAND2_X1 U16654 ( .A1(n15646), .A2(n20643), .ZN(n13532) );
  INV_X1 U16655 ( .A(n13526), .ZN(n13527) );
  NAND2_X1 U16656 ( .A1(n13532), .A2(n13527), .ZN(n13528) );
  NAND2_X1 U16657 ( .A1(n13529), .A2(n13528), .ZN(n15659) );
  INV_X1 U16658 ( .A(n20247), .ZN(n20477) );
  OR2_X1 U16659 ( .A1(n13530), .A2(n20477), .ZN(n13531) );
  XNOR2_X1 U16660 ( .A(n13531), .B(n16086), .ZN(n16080) );
  OR3_X1 U16661 ( .A1(n16080), .A2(n13255), .A3(n13532), .ZN(n13538) );
  NOR2_X1 U16662 ( .A1(n16086), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13535) );
  NOR2_X1 U16663 ( .A1(n16086), .A2(n13533), .ZN(n13534) );
  AOI21_X1 U16664 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13537) );
  NAND2_X1 U16665 ( .A1(n13538), .A2(n13537), .ZN(n15661) );
  INV_X1 U16666 ( .A(n15661), .ZN(n13539) );
  OAI21_X1 U16667 ( .B1(n15659), .B2(n14752), .A(n13539), .ZN(n14746) );
  NOR2_X1 U16668 ( .A1(n14746), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13540) );
  OAI21_X1 U16669 ( .B1(n13540), .B2(n16096), .A(n20254), .ZN(n20723) );
  INV_X1 U16670 ( .A(n20723), .ZN(n20720) );
  NAND2_X1 U16671 ( .A1(n20185), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20586) );
  XNOR2_X1 U16672 ( .A(n9672), .B(n20586), .ZN(n13541) );
  NAND2_X1 U16673 ( .A1(n20479), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20712) );
  AOI22_X1 U16674 ( .A1(n13541), .A2(n20718), .B1(n20112), .B2(n20712), .ZN(
        n13543) );
  NAND2_X1 U16675 ( .A1(n20720), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13542) );
  OAI21_X1 U16676 ( .B1(n20720), .B2(n13543), .A(n13542), .ZN(P1_U3476) );
  INV_X1 U16677 ( .A(n20185), .ZN(n13544) );
  AOI21_X1 U16678 ( .B1(n13544), .B2(n20535), .A(n20590), .ZN(n13546) );
  INV_X1 U16679 ( .A(n13545), .ZN(n20538) );
  AOI22_X1 U16680 ( .A1(n13546), .A2(n20586), .B1(n20538), .B2(n20712), .ZN(
        n13548) );
  NAND2_X1 U16681 ( .A1(n20720), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13547) );
  OAI21_X1 U16682 ( .B1(n20720), .B2(n13548), .A(n13547), .ZN(P1_U3477) );
  INV_X1 U16683 ( .A(n19113), .ZN(n19866) );
  INV_X1 U16684 ( .A(n13612), .ZN(n13620) );
  OR2_X1 U16685 ( .A1(n10490), .A2(n13620), .ZN(n13562) );
  OR2_X1 U16686 ( .A1(n11185), .A2(n11169), .ZN(n13608) );
  NAND2_X1 U16687 ( .A1(n13608), .A2(n13603), .ZN(n13552) );
  NAND2_X1 U16688 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13555) );
  INV_X1 U16689 ( .A(n10519), .ZN(n13549) );
  NAND2_X1 U16690 ( .A1(n13549), .A2(n13614), .ZN(n13602) );
  INV_X1 U16691 ( .A(n13602), .ZN(n13550) );
  AOI21_X1 U16692 ( .B1(n13621), .B2(n13555), .A(n13550), .ZN(n13551) );
  AND2_X1 U16693 ( .A1(n13552), .A2(n13551), .ZN(n13558) );
  INV_X1 U16694 ( .A(n13553), .ZN(n13640) );
  NAND2_X1 U16695 ( .A1(n13640), .A2(n13554), .ZN(n13604) );
  INV_X1 U16696 ( .A(n13555), .ZN(n13556) );
  AOI22_X1 U16697 ( .A1(n13604), .A2(n13602), .B1(n13556), .B2(n13621), .ZN(
        n13557) );
  MUX2_X1 U16698 ( .A(n13558), .B(n13557), .S(n10273), .Z(n13560) );
  AND2_X1 U16699 ( .A1(n13560), .A2(n13559), .ZN(n13561) );
  NAND2_X1 U16700 ( .A1(n13562), .A2(n13561), .ZN(n13615) );
  AOI22_X1 U16701 ( .A1(n19866), .A2(n15328), .B1(n19850), .B2(n13615), .ZN(
        n13564) );
  NAND2_X1 U16702 ( .A1(n19855), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13563) );
  OAI21_X1 U16703 ( .B1(n13564), .B2(n19855), .A(n13563), .ZN(P2_U3596) );
  OR2_X1 U16704 ( .A1(n13567), .A2(n13566), .ZN(n13568) );
  NAND2_X1 U16705 ( .A1(n13565), .A2(n13568), .ZN(n14393) );
  INV_X1 U16706 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13573) );
  INV_X1 U16707 ( .A(n13569), .ZN(n13571) );
  AOI21_X1 U16708 ( .B1(n13571), .B2(n14395), .A(n13570), .ZN(n13572) );
  NOR2_X1 U16709 ( .A1(n13572), .A2(n9981), .ZN(n13594) );
  INV_X1 U16710 ( .A(n13594), .ZN(n14389) );
  OAI222_X1 U16711 ( .A1(n14393), .A2(n14492), .B1(n13573), .B2(n20008), .C1(
        n14389), .C2(n14494), .ZN(P1_U2869) );
  AND2_X1 U16712 ( .A1(n20139), .A2(n13580), .ZN(n13583) );
  INV_X1 U16713 ( .A(n13583), .ZN(n13581) );
  AND2_X1 U16714 ( .A1(n13584), .A2(n13581), .ZN(n13582) );
  OR2_X1 U16715 ( .A1(n14567), .A2(n13584), .ZN(n14217) );
  NAND2_X1 U16716 ( .A1(n14559), .A2(n14217), .ZN(n14568) );
  INV_X1 U16717 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20034) );
  OAI222_X1 U16718 ( .A1(n14572), .A2(n20072), .B1(n14571), .B2(n20117), .C1(
        n9648), .C2(n20034), .ZN(P1_U2904) );
  INV_X1 U16719 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13585) );
  NOR2_X1 U16720 ( .A1(n20103), .A2(n13585), .ZN(n13586) );
  AOI21_X1 U16721 ( .B1(DATAI_1_), .B2(n20103), .A(n13586), .ZN(n20125) );
  OAI222_X1 U16722 ( .A1(n14572), .A2(n19992), .B1(n14571), .B2(n20125), .C1(
        n9648), .C2(n11682), .ZN(P1_U2903) );
  INV_X1 U16723 ( .A(n20005), .ZN(n14406) );
  INV_X1 U16724 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13587) );
  NOR2_X1 U16725 ( .A1(n20103), .A2(n13587), .ZN(n13588) );
  AOI21_X1 U16726 ( .B1(DATAI_2_), .B2(n20103), .A(n13588), .ZN(n20128) );
  OAI222_X1 U16727 ( .A1(n14572), .A2(n14406), .B1(n14571), .B2(n20128), .C1(
        n9648), .C2(n11676), .ZN(P1_U2902) );
  XNOR2_X1 U16728 ( .A(n13590), .B(n13589), .ZN(n13669) );
  AOI21_X1 U16729 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20077) );
  INV_X1 U16730 ( .A(n20077), .ZN(n13591) );
  NAND2_X1 U16731 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14058) );
  AOI21_X1 U16732 ( .B1(n14702), .B2(n14058), .A(n15973), .ZN(n14005) );
  OAI21_X1 U16733 ( .B1(n20093), .B2(n13591), .A(n14005), .ZN(n16046) );
  AOI21_X1 U16734 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14706), .A(
        n20097), .ZN(n15938) );
  AOI22_X1 U16735 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16046), .B1(
        n16070), .B2(n13592), .ZN(n13596) );
  INV_X1 U16736 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13593) );
  NOR2_X1 U16737 ( .A1(n16057), .A2(n13593), .ZN(n13664) );
  AOI21_X1 U16738 ( .B1(n20089), .B2(n13594), .A(n13664), .ZN(n13595) );
  OAI211_X1 U16739 ( .C1(n16073), .C2(n13669), .A(n13596), .B(n13595), .ZN(
        P1_U3028) );
  NAND2_X1 U16740 ( .A1(n20103), .A2(DATAI_3_), .ZN(n13598) );
  NAND2_X1 U16741 ( .A1(n20102), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13597) );
  AND2_X1 U16742 ( .A1(n13598), .A2(n13597), .ZN(n20132) );
  OAI222_X1 U16743 ( .A1(n14572), .A2(n14393), .B1(n20132), .B2(n14571), .C1(
        n9648), .C2(n11724), .ZN(P1_U2901) );
  INV_X1 U16744 ( .A(n13599), .ZN(n13601) );
  NAND3_X1 U16745 ( .A1(n13601), .A2(n10378), .A3(n13600), .ZN(n13654) );
  NAND2_X1 U16746 ( .A1(n13603), .A2(n13602), .ZN(n13605) );
  NAND2_X1 U16747 ( .A1(n13604), .A2(n13605), .ZN(n13610) );
  INV_X1 U16748 ( .A(n13605), .ZN(n13607) );
  XNOR2_X1 U16749 ( .A(n13614), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13606) );
  AOI22_X1 U16750 ( .A1(n13608), .A2(n13607), .B1(n13606), .B2(n13621), .ZN(
        n13609) );
  NAND2_X1 U16751 ( .A1(n13610), .A2(n13609), .ZN(n13611) );
  AOI21_X1 U16752 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n15337) );
  INV_X1 U16753 ( .A(n13647), .ZN(n13628) );
  MUX2_X1 U16754 ( .A(n13614), .B(n15337), .S(n13628), .Z(n13651) );
  MUX2_X1 U16755 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13615), .S(
        n13628), .Z(n13633) );
  INV_X1 U16756 ( .A(n13633), .ZN(n13650) );
  NAND2_X1 U16757 ( .A1(n13616), .A2(n11193), .ZN(n13622) );
  OAI21_X1 U16758 ( .B1(n10512), .B2(n13617), .A(n13622), .ZN(n13619) );
  NAND2_X1 U16759 ( .A1(n13621), .A2(n9789), .ZN(n13618) );
  OAI211_X1 U16760 ( .C1(n10454), .C2(n13620), .A(n13619), .B(n13618), .ZN(
        n19851) );
  INV_X1 U16761 ( .A(n19851), .ZN(n13627) );
  OR2_X1 U16762 ( .A1(n14013), .A2(n13620), .ZN(n13625) );
  MUX2_X1 U16763 ( .A(n13622), .B(n13621), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13623) );
  INV_X1 U16764 ( .A(n13623), .ZN(n13624) );
  NAND2_X1 U16765 ( .A1(n13625), .A2(n13624), .ZN(n15324) );
  OAI22_X1 U16766 ( .A1(n19851), .A2(n19886), .B1(n19896), .B2(n15324), .ZN(
        n13626) );
  OAI21_X1 U16767 ( .B1(n13627), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13626), .ZN(n13629) );
  NAND2_X1 U16768 ( .A1(n13629), .A2(n13628), .ZN(n13632) );
  OR2_X1 U16769 ( .A1(n13651), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13631) );
  OAI21_X1 U16770 ( .B1(n19869), .B2(n13633), .A(n12599), .ZN(n13630) );
  AOI222_X1 U16771 ( .A1(n13632), .A2(n13631), .B1(n13632), .B2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C1(n13631), .C2(n13630), .ZN(
        n13634) );
  OAI221_X1 U16772 ( .B1(n13634), .B2(n19869), .C1(n13634), .C2(n13633), .A(
        n15693), .ZN(n13649) );
  NAND2_X1 U16773 ( .A1(n13636), .A2(n13635), .ZN(n13639) );
  NAND2_X1 U16774 ( .A1(n13641), .A2(n13637), .ZN(n13638) );
  OAI211_X1 U16775 ( .C1(n13641), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        n19905) );
  OAI21_X1 U16776 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n13642), .ZN(n13645) );
  AOI22_X1 U16777 ( .A1(n10918), .A2(n13763), .B1(n13643), .B2(n11135), .ZN(
        n13644) );
  NAND2_X1 U16778 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  AOI211_X1 U16779 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n13647), .A(
        n19905), .B(n13646), .ZN(n13648) );
  OAI211_X1 U16780 ( .C1(n13651), .C2(n13650), .A(n13649), .B(n13648), .ZN(
        n16344) );
  OAI21_X1 U16781 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n16344), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13652) );
  OAI21_X1 U16782 ( .B1(n16342), .B2(n12960), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13655) );
  NAND2_X1 U16783 ( .A1(n13655), .A2(n16339), .ZN(P2_U3593) );
  INV_X1 U16784 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13663) );
  INV_X1 U16785 ( .A(n13508), .ZN(n13657) );
  OAI211_X1 U16786 ( .C1(n13657), .C2(n10114), .A(n19076), .B(n19079), .ZN(
        n13662) );
  NAND2_X1 U16787 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  AND2_X1 U16788 ( .A1(n15257), .A2(n13660), .ZN(n18973) );
  NAND2_X1 U16789 ( .A1(n18973), .A2(n14844), .ZN(n13661) );
  OAI211_X1 U16790 ( .C1(n14844), .C2(n13663), .A(n13662), .B(n13661), .ZN(
        P2_U2875) );
  INV_X1 U16791 ( .A(n14393), .ZN(n13667) );
  AOI21_X1 U16792 ( .B1(n20068), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13664), .ZN(n13665) );
  OAI21_X1 U16793 ( .B1(n15899), .B2(n14386), .A(n13665), .ZN(n13666) );
  AOI21_X1 U16794 ( .B1(n13667), .B2(n15894), .A(n13666), .ZN(n13668) );
  OAI21_X1 U16795 ( .B1(n13669), .B2(n19920), .A(n13668), .ZN(P1_U2996) );
  INV_X1 U16796 ( .A(n13565), .ZN(n13673) );
  INV_X1 U16797 ( .A(n13670), .ZN(n13672) );
  INV_X1 U16798 ( .A(n13671), .ZN(n13705) );
  OAI21_X1 U16799 ( .B1(n13673), .B2(n13672), .A(n13705), .ZN(n14380) );
  INV_X1 U16800 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20026) );
  OAI222_X1 U16801 ( .A1(n14572), .A2(n14380), .B1(n20136), .B2(n14571), .C1(
        n9648), .C2(n20026), .ZN(P1_U2900) );
  INV_X1 U16802 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14369) );
  INV_X1 U16803 ( .A(n13709), .ZN(n13674) );
  XNOR2_X1 U16804 ( .A(n13675), .B(n13674), .ZN(n14374) );
  OAI222_X1 U16805 ( .A1(n14492), .A2(n14380), .B1(n20008), .B2(n14369), .C1(
        n14494), .C2(n14374), .ZN(P1_U2868) );
  AOI22_X1 U16806 ( .A1(n20061), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13677) );
  INV_X1 U16807 ( .A(n20128), .ZN(n13676) );
  NAND2_X1 U16808 ( .A1(n20048), .A2(n13676), .ZN(n13702) );
  NAND2_X1 U16809 ( .A1(n13677), .A2(n13702), .ZN(P1_U2939) );
  AOI22_X1 U16810 ( .A1(n20061), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13679) );
  INV_X1 U16811 ( .A(n20132), .ZN(n13678) );
  NAND2_X1 U16812 ( .A1(n20048), .A2(n13678), .ZN(n13700) );
  NAND2_X1 U16813 ( .A1(n13679), .A2(n13700), .ZN(P1_U2940) );
  AOI22_X1 U16814 ( .A1(n20061), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13681) );
  NAND2_X1 U16815 ( .A1(n13681), .A2(n13680), .ZN(P1_U2952) );
  AOI22_X1 U16816 ( .A1(n20061), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13683) );
  INV_X1 U16817 ( .A(n20125), .ZN(n13682) );
  NAND2_X1 U16818 ( .A1(n20048), .A2(n13682), .ZN(n13696) );
  NAND2_X1 U16819 ( .A1(n13683), .A2(n13696), .ZN(P1_U2953) );
  AOI22_X1 U16820 ( .A1(n20061), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13687) );
  INV_X1 U16821 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13684) );
  NOR2_X1 U16822 ( .A1(n20103), .A2(n13684), .ZN(n13685) );
  AOI21_X1 U16823 ( .B1(DATAI_6_), .B2(n20103), .A(n13685), .ZN(n20144) );
  INV_X1 U16824 ( .A(n20144), .ZN(n13686) );
  NAND2_X1 U16825 ( .A1(n20048), .A2(n13686), .ZN(n13692) );
  NAND2_X1 U16826 ( .A1(n13687), .A2(n13692), .ZN(P1_U2943) );
  AOI22_X1 U16827 ( .A1(n20061), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13691) );
  INV_X1 U16828 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13688) );
  NOR2_X1 U16829 ( .A1(n20103), .A2(n13688), .ZN(n13689) );
  AOI21_X1 U16830 ( .B1(DATAI_5_), .B2(n20103), .A(n13689), .ZN(n20140) );
  INV_X1 U16831 ( .A(n20140), .ZN(n13690) );
  NAND2_X1 U16832 ( .A1(n20048), .A2(n13690), .ZN(n13698) );
  NAND2_X1 U16833 ( .A1(n13691), .A2(n13698), .ZN(P1_U2957) );
  AOI22_X1 U16834 ( .A1(n20061), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13693) );
  NAND2_X1 U16835 ( .A1(n13693), .A2(n13692), .ZN(P1_U2958) );
  AOI22_X1 U16836 ( .A1(n20061), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13695) );
  NAND2_X1 U16837 ( .A1(n13695), .A2(n13694), .ZN(P1_U2959) );
  AOI22_X1 U16838 ( .A1(n20061), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13697) );
  NAND2_X1 U16839 ( .A1(n13697), .A2(n13696), .ZN(P1_U2938) );
  AOI22_X1 U16840 ( .A1(n20061), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U16841 ( .A1(n13699), .A2(n13698), .ZN(P1_U2942) );
  AOI22_X1 U16842 ( .A1(n20061), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13701) );
  NAND2_X1 U16843 ( .A1(n13701), .A2(n13700), .ZN(P1_U2955) );
  AOI22_X1 U16844 ( .A1(n20061), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13703) );
  NAND2_X1 U16845 ( .A1(n13703), .A2(n13702), .ZN(P1_U2954) );
  AND2_X1 U16846 ( .A1(n13705), .A2(n13704), .ZN(n13707) );
  OR2_X1 U16847 ( .A1(n13707), .A2(n13706), .ZN(n19971) );
  AOI21_X1 U16848 ( .B1(n9981), .B2(n13709), .A(n13708), .ZN(n13710) );
  OR2_X1 U16849 ( .A1(n13710), .A2(n9763), .ZN(n19966) );
  OAI22_X1 U16850 ( .A1(n19966), .A2(n14494), .B1(n19965), .B2(n20008), .ZN(
        n13711) );
  INV_X1 U16851 ( .A(n13711), .ZN(n13712) );
  OAI21_X1 U16852 ( .B1(n19971), .B2(n14492), .A(n13712), .ZN(P1_U2867) );
  XOR2_X1 U16853 ( .A(n13713), .B(n13714), .Z(n13719) );
  INV_X1 U16854 ( .A(n13719), .ZN(n13718) );
  NAND2_X1 U16855 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16071) );
  OAI211_X1 U16856 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n16070), .B(n16071), .ZN(n13717) );
  INV_X1 U16857 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20663) );
  NOR2_X1 U16858 ( .A1(n16057), .A2(n20663), .ZN(n13721) );
  NOR2_X1 U16859 ( .A1(n16079), .A2(n14374), .ZN(n13715) );
  AOI211_X1 U16860 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n16046), .A(
        n13721), .B(n13715), .ZN(n13716) );
  OAI211_X1 U16861 ( .C1(n13718), .C2(n16073), .A(n13717), .B(n13716), .ZN(
        P1_U3027) );
  OAI222_X1 U16862 ( .A1(n14572), .A2(n19971), .B1(n20140), .B2(n14571), .C1(
        n9648), .C2(n11771), .ZN(P1_U2899) );
  NAND2_X1 U16863 ( .A1(n13719), .A2(n20070), .ZN(n13723) );
  NOR2_X1 U16864 ( .A1(n15899), .A2(n14371), .ZN(n13720) );
  AOI211_X1 U16865 ( .C1(n20068), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13721), .B(n13720), .ZN(n13722) );
  OAI211_X1 U16866 ( .C1(n20104), .C2(n14380), .A(n13723), .B(n13722), .ZN(
        P1_U2995) );
  NAND2_X1 U16867 ( .A1(n13725), .A2(n13724), .ZN(n13727) );
  XNOR2_X1 U16868 ( .A(n13727), .B(n13726), .ZN(n13748) );
  INV_X2 U16869 ( .A(n19044), .ZN(n19023) );
  NOR2_X1 U16870 ( .A1(n19023), .A2(n13729), .ZN(n13741) );
  INV_X1 U16871 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13886) );
  OAI22_X1 U16872 ( .A1(n13886), .A2(n19229), .B1(n16256), .B2(n13883), .ZN(
        n13730) );
  AOI211_X1 U16873 ( .C1(n19239), .C2(n13728), .A(n13741), .B(n13730), .ZN(
        n13735) );
  NAND2_X1 U16874 ( .A1(n13732), .A2(n13733), .ZN(n13745) );
  NAND3_X1 U16875 ( .A1(n13731), .A2(n19224), .A3(n13745), .ZN(n13734) );
  OAI211_X1 U16876 ( .C1(n13748), .C2(n19236), .A(n13735), .B(n13734), .ZN(
        P2_U3011) );
  OAI211_X1 U16877 ( .C1(n13737), .C2(n13736), .A(n10662), .B(n15264), .ZN(
        n13743) );
  OR2_X1 U16878 ( .A1(n13739), .A2(n13738), .ZN(n13740) );
  NAND2_X1 U16879 ( .A1(n13740), .A2(n13801), .ZN(n13892) );
  INV_X1 U16880 ( .A(n13892), .ZN(n19865) );
  AOI21_X1 U16881 ( .B1(n19865), .B2(n16301), .A(n13741), .ZN(n13742) );
  OAI211_X1 U16882 ( .C1(n10490), .C2(n16329), .A(n13743), .B(n13742), .ZN(
        n13744) );
  AOI21_X1 U16883 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13799), .A(
        n13744), .ZN(n13747) );
  NAND3_X1 U16884 ( .A1(n13731), .A2(n13745), .A3(n16313), .ZN(n13746) );
  OAI211_X1 U16885 ( .C1(n13748), .C2(n16317), .A(n13747), .B(n13746), .ZN(
        P2_U3043) );
  INV_X1 U16886 ( .A(n13749), .ZN(n13750) );
  OAI211_X1 U16887 ( .C1(n13752), .C2(n13751), .A(n13750), .B(n19079), .ZN(
        n13756) );
  OR2_X1 U16888 ( .A1(n15258), .A2(n13753), .ZN(n13754) );
  AND2_X1 U16889 ( .A1(n13754), .A2(n13777), .ZN(n16288) );
  NAND2_X1 U16890 ( .A1(n16288), .A2(n14844), .ZN(n13755) );
  OAI211_X1 U16891 ( .C1(n14844), .C2(n11020), .A(n13756), .B(n13755), .ZN(
        P2_U2873) );
  NAND2_X1 U16892 ( .A1(n19113), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19445) );
  OR2_X1 U16893 ( .A1(n19445), .A2(n19624), .ZN(n13757) );
  NAND2_X1 U16894 ( .A1(n13757), .A2(n19864), .ZN(n13768) );
  INV_X1 U16895 ( .A(n13768), .ZN(n13761) );
  NAND3_X1 U16896 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19869), .A3(
        n19886), .ZN(n19362) );
  AOI21_X1 U16897 ( .B1(n13766), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13759) );
  NOR2_X1 U16898 ( .A1(n19896), .A2(n19362), .ZN(n19412) );
  OAI21_X1 U16899 ( .B1(n13759), .B2(n19412), .A(n19702), .ZN(n13760) );
  INV_X1 U16900 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U16901 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19261), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19262), .ZN(n19707) );
  INV_X1 U16902 ( .A(n19707), .ZN(n19649) );
  NOR2_X2 U16903 ( .A1(n19411), .A2(n19624), .ZN(n19405) );
  AOI22_X1 U16904 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19261), .ZN(n19663) );
  NAND2_X1 U16905 ( .A1(n13763), .A2(n19258), .ZN(n19242) );
  INV_X1 U16906 ( .A(n19412), .ZN(n13764) );
  OAI22_X1 U16907 ( .A1(n19663), .A2(n19389), .B1(n19242), .B2(n13764), .ZN(
        n13765) );
  AOI21_X1 U16908 ( .B1(n19649), .B2(n19405), .A(n13765), .ZN(n13770) );
  OAI21_X1 U16909 ( .B1(n10542), .B2(n19412), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13767) );
  OAI21_X1 U16910 ( .B1(n13768), .B2(n19362), .A(n13767), .ZN(n19406) );
  NOR2_X2 U16911 ( .A1(n19146), .A2(n19447), .ZN(n19696) );
  NAND2_X1 U16912 ( .A1(n19406), .A2(n19696), .ZN(n13769) );
  OAI211_X1 U16913 ( .C1(n19410), .C2(n13771), .A(n13770), .B(n13769), .ZN(
        P2_U3088) );
  INV_X1 U16914 ( .A(n13772), .ZN(n13774) );
  INV_X1 U16915 ( .A(n13706), .ZN(n13773) );
  AOI21_X1 U16916 ( .B1(n13774), .B2(n13773), .A(n13786), .ZN(n19957) );
  INV_X1 U16917 ( .A(n19957), .ZN(n13783) );
  XOR2_X1 U16918 ( .A(n13775), .B(n9763), .Z(n19951) );
  AOI22_X1 U16919 ( .A1(n19951), .A2(n20003), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14483), .ZN(n13776) );
  OAI21_X1 U16920 ( .B1(n13783), .B2(n14492), .A(n13776), .ZN(P1_U2866) );
  AOI21_X1 U16921 ( .B1(n13778), .B2(n13777), .A(n13833), .ZN(n18949) );
  INV_X1 U16922 ( .A(n18949), .ZN(n15091) );
  OAI211_X1 U16923 ( .C1(n13749), .C2(n13780), .A(n13831), .B(n19079), .ZN(
        n13782) );
  NAND2_X1 U16924 ( .A1(n19078), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13781) );
  OAI211_X1 U16925 ( .C1(n15091), .C2(n19078), .A(n13782), .B(n13781), .ZN(
        P2_U2872) );
  OAI222_X1 U16926 ( .A1(n14572), .A2(n13783), .B1(n20144), .B2(n14571), .C1(
        n9648), .C2(n11788), .ZN(P1_U2898) );
  OR2_X1 U16927 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  NAND2_X1 U16928 ( .A1(n13784), .A2(n13787), .ZN(n19945) );
  NAND2_X1 U16929 ( .A1(n13789), .A2(n13788), .ZN(n13790) );
  NAND2_X1 U16930 ( .A1(n13843), .A2(n13790), .ZN(n19939) );
  OAI22_X1 U16931 ( .A1(n19939), .A2(n14494), .B1(n19938), .B2(n20008), .ZN(
        n13791) );
  INV_X1 U16932 ( .A(n13791), .ZN(n13792) );
  OAI21_X1 U16933 ( .B1(n19945), .B2(n14492), .A(n13792), .ZN(P1_U2865) );
  XOR2_X1 U16934 ( .A(n13794), .B(n13793), .Z(n19221) );
  INV_X1 U16935 ( .A(n19221), .ZN(n13807) );
  XNOR2_X1 U16936 ( .A(n13795), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13796) );
  XNOR2_X1 U16937 ( .A(n13797), .B(n13796), .ZN(n19225) );
  OR2_X1 U16938 ( .A1(n10662), .A2(n13798), .ZN(n13859) );
  AOI21_X1 U16939 ( .B1(n10662), .B2(n15264), .A(n13799), .ZN(n13864) );
  NAND2_X1 U16940 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19044), .ZN(n13800) );
  OAI221_X1 U16941 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13859), .C1(
        n13860), .C2(n13864), .A(n13800), .ZN(n13805) );
  NAND2_X1 U16942 ( .A1(n13802), .A2(n13801), .ZN(n13803) );
  AND2_X1 U16943 ( .A1(n13803), .A2(n10118), .ZN(n19124) );
  INV_X1 U16944 ( .A(n19124), .ZN(n19117) );
  OAI22_X1 U16945 ( .A1(n13811), .A2(n16329), .B1(n16324), .B2(n19117), .ZN(
        n13804) );
  AOI211_X1 U16946 ( .C1(n19225), .C2(n16313), .A(n13805), .B(n13804), .ZN(
        n13806) );
  OAI21_X1 U16947 ( .B1(n13807), .B2(n16317), .A(n13806), .ZN(P2_U3042) );
  AND2_X1 U16948 ( .A1(n19029), .A2(n13808), .ZN(n13810) );
  AOI21_X1 U16949 ( .B1(n19219), .B2(n13810), .A(n19759), .ZN(n13809) );
  OAI21_X1 U16950 ( .B1(n19219), .B2(n13810), .A(n13809), .ZN(n13818) );
  INV_X1 U16951 ( .A(n13811), .ZN(n19223) );
  AOI22_X1 U16952 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19055), .B1(n18972), .B2(
        n19124), .ZN(n13812) );
  OAI211_X1 U16953 ( .C1(n19057), .C2(n19228), .A(n19023), .B(n13812), .ZN(
        n13813) );
  AOI21_X1 U16954 ( .B1(n19045), .B2(P2_REIP_REG_4__SCAN_IN), .A(n13813), .ZN(
        n13814) );
  OAI21_X1 U16955 ( .B1(n13815), .B2(n19024), .A(n13814), .ZN(n13816) );
  AOI21_X1 U16956 ( .B1(n19223), .B2(n19067), .A(n13816), .ZN(n13817) );
  OAI211_X1 U16957 ( .C1(n19125), .C2(n14023), .A(n13818), .B(n13817), .ZN(
        P2_U2851) );
  OAI222_X1 U16958 ( .A1(n14572), .A2(n19945), .B1(n20152), .B2(n14571), .C1(
        n9648), .C2(n11801), .ZN(P1_U2897) );
  NAND2_X1 U16959 ( .A1(n19029), .A2(n15331), .ZN(n13819) );
  XNOR2_X1 U16960 ( .A(n13820), .B(n13819), .ZN(n13821) );
  NAND2_X1 U16961 ( .A1(n13821), .A2(n12968), .ZN(n13829) );
  AOI22_X1 U16962 ( .A1(n19062), .A2(n13822), .B1(n19045), .B2(
        P2_REIP_REG_2__SCAN_IN), .ZN(n13823) );
  OAI21_X1 U16963 ( .B1(n19042), .B2(n13295), .A(n13823), .ZN(n13826) );
  OAI22_X1 U16964 ( .A1(n19114), .A2(n19065), .B1(n13824), .B2(n19057), .ZN(
        n13825) );
  AOI211_X1 U16965 ( .C1(n19067), .C2(n13613), .A(n13826), .B(n13825), .ZN(
        n13828) );
  OAI211_X1 U16966 ( .C1(n19872), .C2(n14023), .A(n13829), .B(n13828), .ZN(
        P2_U2853) );
  AOI21_X1 U16967 ( .B1(n13832), .B2(n13831), .A(n13830), .ZN(n14964) );
  NAND2_X1 U16968 ( .A1(n14964), .A2(n19079), .ZN(n13837) );
  OR2_X1 U16969 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  NAND2_X1 U16970 ( .A1(n9740), .A2(n13835), .ZN(n16207) );
  INV_X1 U16971 ( .A(n16207), .ZN(n13957) );
  NAND2_X1 U16972 ( .A1(n14844), .A2(n13957), .ZN(n13836) );
  OAI211_X1 U16973 ( .C1(n14844), .C2(n10830), .A(n13837), .B(n13836), .ZN(
        P2_U2871) );
  NAND2_X1 U16974 ( .A1(n13784), .A2(n13838), .ZN(n13839) );
  NAND2_X1 U16975 ( .A1(n9679), .A2(n13839), .ZN(n13995) );
  AND2_X1 U16976 ( .A1(n13840), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13841) );
  INV_X1 U16977 ( .A(n13842), .ZN(n13992) );
  AOI21_X1 U16978 ( .B1(n13844), .B2(n13843), .A(n13973), .ZN(n13845) );
  INV_X1 U16979 ( .A(n13845), .ZN(n16051) );
  NAND2_X1 U16980 ( .A1(n15779), .A2(n13846), .ZN(n19963) );
  AOI21_X1 U16981 ( .B1(n19977), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19955), .ZN(n13848) );
  OAI21_X1 U16982 ( .B1(n15803), .B2(n13978), .A(n15779), .ZN(n13980) );
  AOI22_X1 U16983 ( .A1(n13980), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n19997), .ZN(n13847) );
  OAI211_X1 U16984 ( .C1(n19985), .C2(n16051), .A(n13848), .B(n13847), .ZN(
        n13851) );
  NAND3_X1 U16985 ( .A1(n15771), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n14382) );
  NOR2_X1 U16986 ( .A1(n13593), .A2(n14382), .ZN(n14368) );
  NAND2_X1 U16987 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n14368), .ZN(n19975) );
  NOR3_X1 U16988 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13849), .A3(n19975), .ZN(
        n13850) );
  AOI211_X1 U16989 ( .C1(n19989), .C2(n13992), .A(n13851), .B(n13850), .ZN(
        n13852) );
  OAI21_X1 U16990 ( .B1(n19944), .B2(n13995), .A(n13852), .ZN(P1_U2832) );
  XNOR2_X1 U16991 ( .A(n13853), .B(n13855), .ZN(n13902) );
  NAND2_X1 U16992 ( .A1(n13857), .A2(n13856), .ZN(n13858) );
  AOI221_X1 U16993 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n10739), .C2(n13860), .A(
        n13859), .ZN(n13870) );
  INV_X1 U16994 ( .A(n19050), .ZN(n13868) );
  XNOR2_X1 U16995 ( .A(n13862), .B(n13861), .ZN(n19122) );
  INV_X1 U16996 ( .A(n19122), .ZN(n13866) );
  NOR2_X1 U16997 ( .A1(n19023), .A2(n13863), .ZN(n13898) );
  NOR2_X1 U16998 ( .A1(n10739), .A2(n13864), .ZN(n13865) );
  AOI211_X1 U16999 ( .C1(n16301), .C2(n13866), .A(n13898), .B(n13865), .ZN(
        n13867) );
  OAI21_X1 U17000 ( .B1(n13868), .B2(n16329), .A(n13867), .ZN(n13869) );
  AOI211_X1 U17001 ( .C1(n13899), .C2(n16313), .A(n13870), .B(n13869), .ZN(
        n13871) );
  OAI21_X1 U17002 ( .B1(n13902), .B2(n16317), .A(n13871), .ZN(P2_U3041) );
  NAND2_X1 U17003 ( .A1(n19029), .A2(n13872), .ZN(n13873) );
  XNOR2_X1 U17004 ( .A(n16257), .B(n13873), .ZN(n13875) );
  AOI21_X1 U17005 ( .B1(n13874), .B2(n15301), .A(n15286), .ZN(n16323) );
  AOI22_X1 U17006 ( .A1(n12968), .A2(n13875), .B1(n18972), .B2(n16323), .ZN(
        n13880) );
  INV_X1 U17007 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19796) );
  OAI21_X1 U17008 ( .B1(n19796), .B2(n19059), .A(n19023), .ZN(n13876) );
  AOI21_X1 U17009 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19038), .A(
        n13876), .ZN(n13877) );
  OAI21_X1 U17010 ( .B1(n16328), .B2(n18958), .A(n13877), .ZN(n13878) );
  AOI21_X1 U17011 ( .B1(n19055), .B2(P2_EBX_REG_8__SCAN_IN), .A(n13878), .ZN(
        n13879) );
  OAI211_X1 U17012 ( .C1(n13881), .C2(n19024), .A(n13880), .B(n13879), .ZN(
        P2_U2847) );
  NOR2_X1 U17013 ( .A1(n19047), .A2(n13882), .ZN(n13884) );
  XNOR2_X1 U17014 ( .A(n13884), .B(n13883), .ZN(n13885) );
  NAND2_X1 U17015 ( .A1(n13885), .A2(n12968), .ZN(n13895) );
  OAI22_X1 U17016 ( .A1(n13886), .A2(n19057), .B1(n13729), .B2(n19059), .ZN(
        n13890) );
  NAND2_X1 U17017 ( .A1(n19055), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13887) );
  OAI21_X1 U17018 ( .B1(n19024), .B2(n13888), .A(n13887), .ZN(n13889) );
  NOR2_X1 U17019 ( .A1(n13890), .A2(n13889), .ZN(n13891) );
  OAI21_X1 U17020 ( .B1(n13892), .B2(n19065), .A(n13891), .ZN(n13893) );
  AOI21_X1 U17021 ( .B1(n13728), .B2(n19067), .A(n13893), .ZN(n13894) );
  OAI211_X1 U17022 ( .C1(n19113), .C2(n14023), .A(n13895), .B(n13894), .ZN(
        P2_U2852) );
  INV_X1 U17023 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13896) );
  OAI22_X1 U17024 ( .A1(n19229), .A2(n13896), .B1(n16256), .B2(n19048), .ZN(
        n13897) );
  AOI211_X1 U17025 ( .C1(n19050), .C2(n19239), .A(n13898), .B(n13897), .ZN(
        n13901) );
  NAND2_X1 U17026 ( .A1(n13899), .A2(n19224), .ZN(n13900) );
  OAI211_X1 U17027 ( .C1(n13902), .C2(n19236), .A(n13901), .B(n13900), .ZN(
        P2_U3009) );
  OAI222_X1 U17028 ( .A1(n13995), .A2(n14572), .B1(n14526), .B2(n14571), .C1(
        n20021), .C2(n9648), .ZN(P1_U2896) );
  INV_X1 U17029 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13903) );
  OAI222_X1 U17030 ( .A1(n13995), .A2(n14492), .B1(n20008), .B2(n13903), .C1(
        n16051), .C2(n14494), .ZN(P1_U2864) );
  OAI21_X1 U17031 ( .B1(n19547), .B2(n19579), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13904) );
  NAND2_X1 U17032 ( .A1(n13904), .A2(n19864), .ZN(n13914) );
  INV_X1 U17033 ( .A(n13914), .ZN(n13907) );
  NAND2_X1 U17034 ( .A1(n12599), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19553) );
  INV_X1 U17035 ( .A(n19553), .ZN(n19557) );
  NAND2_X1 U17036 ( .A1(n19358), .A2(n19557), .ZN(n13913) );
  AOI21_X1 U17037 ( .B1(n10541), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13905) );
  NAND2_X1 U17038 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19896), .ZN(
        n19296) );
  NOR2_X1 U17039 ( .A1(n19296), .A2(n19553), .ZN(n19546) );
  OAI21_X1 U17040 ( .B1(n13905), .B2(n19546), .A(n19702), .ZN(n13906) );
  INV_X1 U17041 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13917) );
  INV_X1 U17042 ( .A(n19546), .ZN(n13908) );
  OAI22_X1 U17043 ( .A1(n19663), .A2(n13909), .B1(n19242), .B2(n13908), .ZN(
        n13910) );
  AOI21_X1 U17044 ( .B1(n19547), .B2(n19649), .A(n13910), .ZN(n13916) );
  INV_X1 U17045 ( .A(n10541), .ZN(n13911) );
  OAI21_X1 U17046 ( .B1(n13911), .B2(n19546), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13912) );
  NAND2_X1 U17047 ( .A1(n19548), .A2(n19696), .ZN(n13915) );
  OAI211_X1 U17048 ( .C1(n19552), .C2(n13917), .A(n13916), .B(n13915), .ZN(
        P2_U3128) );
  NOR2_X2 U17049 ( .A1(n19502), .A2(n19411), .ZN(n19292) );
  OAI21_X1 U17050 ( .B1(n19749), .B2(n19292), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13918) );
  NAND2_X1 U17051 ( .A1(n13918), .A2(n19864), .ZN(n13926) );
  INV_X1 U17052 ( .A(n13926), .ZN(n13921) );
  NAND2_X1 U17053 ( .A1(n19869), .A2(n12599), .ZN(n19328) );
  OR2_X1 U17054 ( .A1(n19328), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19269) );
  NOR2_X1 U17055 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19269), .ZN(
        n19259) );
  NOR2_X1 U17056 ( .A1(n19745), .A2(n19259), .ZN(n13925) );
  AOI21_X1 U17057 ( .B1(n10695), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13919) );
  OAI21_X1 U17058 ( .B1(n13919), .B2(n19259), .A(n19702), .ZN(n13920) );
  AOI22_X1 U17059 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19261), .ZN(n19713) );
  INV_X1 U17060 ( .A(n19713), .ZN(n19594) );
  AOI22_X1 U17061 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19261), .ZN(n19597) );
  INV_X1 U17062 ( .A(n19292), .ZN(n13943) );
  INV_X1 U17063 ( .A(n19259), .ZN(n13942) );
  NAND2_X1 U17064 ( .A1(n10294), .A2(n19258), .ZN(n19274) );
  OAI22_X1 U17065 ( .A1(n19597), .A2(n13943), .B1(n13942), .B2(n19274), .ZN(
        n13922) );
  AOI21_X1 U17066 ( .B1(n19749), .B2(n19594), .A(n13922), .ZN(n13929) );
  INV_X1 U17067 ( .A(n10695), .ZN(n13923) );
  OAI21_X1 U17068 ( .B1(n13923), .B2(n19259), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13924) );
  NOR2_X2 U17069 ( .A1(n13927), .A2(n19447), .ZN(n19709) );
  NAND2_X1 U17070 ( .A1(n19263), .A2(n19709), .ZN(n13928) );
  OAI211_X1 U17071 ( .C1(n19266), .C2(n13930), .A(n13929), .B(n13928), .ZN(
        P2_U3049) );
  INV_X1 U17072 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16423) );
  INV_X1 U17073 ( .A(n19262), .ZN(n19253) );
  INV_X1 U17074 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18236) );
  INV_X1 U17075 ( .A(n19261), .ZN(n19251) );
  OAI22_X2 U17076 ( .A1(n16423), .A2(n19253), .B1(n18236), .B2(n19251), .ZN(
        n19684) );
  AOI22_X1 U17077 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19261), .ZN(n19689) );
  NAND2_X1 U17078 ( .A1(n13931), .A2(n19258), .ZN(n19289) );
  OAI22_X1 U17079 ( .A1(n19689), .A2(n13943), .B1(n13942), .B2(n19289), .ZN(
        n13932) );
  AOI21_X1 U17080 ( .B1(n19749), .B2(n19684), .A(n13932), .ZN(n13934) );
  NOR2_X2 U17081 ( .A1(n19108), .A2(n19447), .ZN(n19746) );
  NAND2_X1 U17082 ( .A1(n19263), .A2(n19746), .ZN(n13933) );
  OAI211_X1 U17083 ( .C1(n19266), .C2(n13935), .A(n13934), .B(n13933), .ZN(
        P2_U3055) );
  AOI22_X1 U17084 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19261), .ZN(n19725) );
  AOI22_X1 U17085 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19261), .ZN(n19673) );
  NAND2_X1 U17086 ( .A1(n13936), .A2(n19258), .ZN(n19280) );
  OAI22_X1 U17087 ( .A1(n19673), .A2(n13943), .B1(n13942), .B2(n19280), .ZN(
        n13937) );
  AOI21_X1 U17088 ( .B1(n19749), .B2(n19670), .A(n13937), .ZN(n13939) );
  NOR2_X2 U17089 ( .A1(n19136), .A2(n19447), .ZN(n19721) );
  NAND2_X1 U17090 ( .A1(n19263), .A2(n19721), .ZN(n13938) );
  OAI211_X1 U17091 ( .C1(n19266), .C2(n13940), .A(n13939), .B(n13938), .ZN(
        P2_U3051) );
  AOI22_X1 U17092 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19261), .ZN(n19719) );
  INV_X1 U17093 ( .A(n19719), .ZN(n19666) );
  AOI22_X1 U17094 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19261), .ZN(n19669) );
  NAND2_X1 U17095 ( .A1(n13941), .A2(n19258), .ZN(n19277) );
  OAI22_X1 U17096 ( .A1(n19669), .A2(n13943), .B1(n13942), .B2(n19277), .ZN(
        n13944) );
  AOI21_X1 U17097 ( .B1(n19749), .B2(n19666), .A(n13944), .ZN(n13947) );
  NOR2_X2 U17098 ( .A1(n13945), .A2(n19447), .ZN(n19715) );
  NAND2_X1 U17099 ( .A1(n19263), .A2(n19715), .ZN(n13946) );
  OAI211_X1 U17100 ( .C1(n19266), .C2(n13948), .A(n13947), .B(n13946), .ZN(
        P2_U3050) );
  INV_X1 U17101 ( .A(n16273), .ZN(n13949) );
  XNOR2_X1 U17102 ( .A(n13950), .B(n13949), .ZN(n15622) );
  INV_X1 U17103 ( .A(n13951), .ZN(n16196) );
  NAND2_X1 U17104 ( .A1(n19029), .A2(n18941), .ZN(n13952) );
  XOR2_X1 U17105 ( .A(n16196), .B(n13952), .Z(n13953) );
  AOI22_X1 U17106 ( .A1(n15622), .A2(n18972), .B1(n12968), .B2(n13953), .ZN(
        n13959) );
  INV_X1 U17107 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19808) );
  OAI21_X1 U17108 ( .B1(n19808), .B2(n19059), .A(n19023), .ZN(n13954) );
  AOI21_X1 U17109 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19038), .A(
        n13954), .ZN(n13955) );
  OAI21_X1 U17110 ( .B1(n19042), .B2(n10830), .A(n13955), .ZN(n13956) );
  AOI21_X1 U17111 ( .B1(n19067), .B2(n13957), .A(n13956), .ZN(n13958) );
  OAI211_X1 U17112 ( .C1(n13960), .C2(n19024), .A(n13959), .B(n13958), .ZN(
        P2_U2839) );
  AOI21_X1 U17113 ( .B1(n13961), .B2(n15254), .A(n16271), .ZN(n16285) );
  NAND2_X1 U17114 ( .A1(n19029), .A2(n13962), .ZN(n18961) );
  XOR2_X1 U17115 ( .A(n16220), .B(n18961), .Z(n13963) );
  AOI22_X1 U17116 ( .A1(n16285), .A2(n18972), .B1(n12968), .B2(n13963), .ZN(
        n13968) );
  INV_X1 U17117 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U17118 ( .B1(n19805), .B2(n19059), .A(n19023), .ZN(n13964) );
  AOI21_X1 U17119 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19038), .A(
        n13964), .ZN(n13965) );
  OAI21_X1 U17120 ( .B1(n19042), .B2(n11020), .A(n13965), .ZN(n13966) );
  AOI21_X1 U17121 ( .B1(n16288), .B2(n19067), .A(n13966), .ZN(n13967) );
  OAI211_X1 U17122 ( .C1(n13969), .C2(n19024), .A(n13968), .B(n13967), .ZN(
        P2_U2841) );
  AOI21_X1 U17123 ( .B1(n13971), .B2(n9679), .A(n13970), .ZN(n14003) );
  INV_X1 U17124 ( .A(n14003), .ZN(n13988) );
  NOR2_X1 U17125 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15803), .ZN(n13979) );
  NOR2_X1 U17126 ( .A1(n13973), .A2(n13972), .ZN(n13974) );
  OR2_X1 U17127 ( .A1(n14027), .A2(n13974), .ZN(n13983) );
  INV_X1 U17128 ( .A(n13983), .ZN(n14009) );
  AOI22_X1 U17129 ( .A1(n14009), .A2(n19994), .B1(n19997), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n13975) );
  OAI211_X1 U17130 ( .C1(n19996), .C2(n13976), .A(n13975), .B(n19963), .ZN(
        n13977) );
  AOI21_X1 U17131 ( .B1(n13979), .B2(n13978), .A(n13977), .ZN(n13982) );
  AOI22_X1 U17132 ( .A1(n13980), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n19989), 
        .B2(n14000), .ZN(n13981) );
  OAI211_X1 U17133 ( .C1(n13988), .C2(n19944), .A(n13982), .B(n13981), .ZN(
        P1_U2831) );
  OAI222_X1 U17134 ( .A1(n13988), .A2(n14492), .B1(n13984), .B2(n20008), .C1(
        n13983), .C2(n14494), .ZN(P1_U2863) );
  INV_X1 U17135 ( .A(DATAI_9_), .ZN(n13986) );
  INV_X1 U17136 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13985) );
  MUX2_X1 U17137 ( .A(n13986), .B(n13985), .S(n20102), .Z(n20035) );
  INV_X1 U17138 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13987) );
  OAI222_X1 U17139 ( .A1(n13988), .A2(n14572), .B1(n20035), .B2(n14571), .C1(
        n13987), .C2(n9648), .ZN(P1_U2895) );
  XNOR2_X1 U17140 ( .A(n13989), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13990) );
  XNOR2_X1 U17141 ( .A(n13991), .B(n13990), .ZN(n16054) );
  AOI22_X1 U17142 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13994) );
  NAND2_X1 U17143 ( .A1(n15871), .A2(n13992), .ZN(n13993) );
  OAI211_X1 U17144 ( .C1(n13995), .C2(n20104), .A(n13994), .B(n13993), .ZN(
        n13996) );
  AOI21_X1 U17145 ( .B1(n16054), .B2(n20070), .A(n13996), .ZN(n13997) );
  INV_X1 U17146 ( .A(n13997), .ZN(P1_U2991) );
  XNOR2_X1 U17147 ( .A(n12393), .B(n20884), .ZN(n13998) );
  XNOR2_X1 U17148 ( .A(n13999), .B(n13998), .ZN(n14012) );
  NAND2_X1 U17149 ( .A1(n15871), .A2(n14000), .ZN(n14001) );
  NAND2_X1 U17150 ( .A1(n20074), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14007) );
  OAI211_X1 U17151 ( .C1(n15902), .C2(n13976), .A(n14001), .B(n14007), .ZN(
        n14002) );
  AOI21_X1 U17152 ( .B1(n14003), .B2(n15894), .A(n14002), .ZN(n14004) );
  OAI21_X1 U17153 ( .B1(n14012), .B2(n19920), .A(n14004), .ZN(P1_U2990) );
  NOR2_X1 U17154 ( .A1(n12355), .A2(n16071), .ZN(n16064) );
  NAND4_X1 U17155 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16064), .ZN(n14057) );
  NOR2_X1 U17156 ( .A1(n20077), .A2(n14057), .ZN(n16037) );
  AOI22_X1 U17157 ( .A1(n16048), .A2(n20078), .B1(n16037), .B2(n14005), .ZN(
        n16040) );
  AND2_X1 U17158 ( .A1(n16037), .A2(n16036), .ZN(n14006) );
  AOI22_X1 U17159 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16040), .B1(
        n14006), .B2(n20884), .ZN(n14011) );
  INV_X1 U17160 ( .A(n14007), .ZN(n14008) );
  AOI21_X1 U17161 ( .B1(n14009), .B2(n20089), .A(n14008), .ZN(n14010) );
  OAI211_X1 U17162 ( .C1(n14012), .C2(n16073), .A(n14011), .B(n14010), .ZN(
        P1_U3022) );
  NAND2_X1 U17163 ( .A1(n19055), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n14020) );
  INV_X1 U17164 ( .A(n15333), .ZN(n15323) );
  NOR2_X1 U17165 ( .A1(n19047), .A2(n19759), .ZN(n18942) );
  NAND2_X1 U17166 ( .A1(n15323), .A2(n18942), .ZN(n14015) );
  NOR2_X1 U17167 ( .A1(n19759), .A2(n19029), .ZN(n18956) );
  OAI21_X1 U17168 ( .B1(n19038), .B2(n18956), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U17169 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  AOI21_X1 U17170 ( .B1(n19062), .B2(n14017), .A(n14016), .ZN(n14019) );
  AOI22_X1 U17171 ( .A1(n18972), .A2(n19141), .B1(n19045), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n14018) );
  NAND3_X1 U17172 ( .A1(n14020), .A2(n14019), .A3(n14018), .ZN(n14021) );
  AOI21_X1 U17173 ( .B1(n10461), .B2(n19067), .A(n14021), .ZN(n14022) );
  OAI21_X1 U17174 ( .B1(n19890), .B2(n14023), .A(n14022), .ZN(P2_U2855) );
  INV_X1 U17175 ( .A(n13970), .ZN(n14025) );
  AOI21_X1 U17176 ( .B1(n9772), .B2(n14025), .A(n11906), .ZN(n14696) );
  INV_X1 U17177 ( .A(n14696), .ZN(n14362) );
  OR2_X1 U17178 ( .A1(n14027), .A2(n14026), .ZN(n14028) );
  NAND2_X1 U17179 ( .A1(n14047), .A2(n14028), .ZN(n16038) );
  OAI22_X1 U17180 ( .A1(n16038), .A2(n14494), .B1(n14355), .B2(n20008), .ZN(
        n14029) );
  INV_X1 U17181 ( .A(n14029), .ZN(n14030) );
  OAI21_X1 U17182 ( .B1(n14362), .B2(n14492), .A(n14030), .ZN(P1_U2862) );
  INV_X1 U17183 ( .A(DATAI_10_), .ZN(n14032) );
  INV_X1 U17184 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14031) );
  MUX2_X1 U17185 ( .A(n14032), .B(n14031), .S(n20102), .Z(n20038) );
  OAI222_X1 U17186 ( .A1(n14572), .A2(n14362), .B1(n20038), .B2(n14571), .C1(
        n14033), .C2(n9648), .ZN(P1_U2894) );
  AND2_X1 U17187 ( .A1(n14034), .A2(n14035), .ZN(n14037) );
  OR2_X1 U17188 ( .A1(n14037), .A2(n14036), .ZN(n15797) );
  OR2_X1 U17189 ( .A1(n14345), .A2(n14038), .ZN(n14039) );
  NAND2_X1 U17190 ( .A1(n14477), .A2(n14039), .ZN(n16006) );
  OAI22_X1 U17191 ( .A1(n16006), .A2(n14494), .B1(n15795), .B2(n20008), .ZN(
        n14040) );
  INV_X1 U17192 ( .A(n14040), .ZN(n14041) );
  OAI21_X1 U17193 ( .B1(n15797), .B2(n14492), .A(n14041), .ZN(P1_U2858) );
  XOR2_X1 U17194 ( .A(n14343), .B(n14042), .Z(n14045) );
  INV_X1 U17195 ( .A(n14043), .ZN(n14044) );
  NOR2_X1 U17196 ( .A1(n14045), .A2(n14044), .ZN(n14342) );
  AOI21_X1 U17197 ( .B1(n14045), .B2(n14044), .A(n14342), .ZN(n15879) );
  INV_X1 U17198 ( .A(n15879), .ZN(n14055) );
  INV_X1 U17199 ( .A(n14486), .ZN(n14046) );
  AOI21_X1 U17200 ( .B1(n14048), .B2(n14047), .A(n14046), .ZN(n16029) );
  AOI22_X1 U17201 ( .A1(n16029), .A2(n20003), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14483), .ZN(n14049) );
  OAI21_X1 U17202 ( .B1(n14055), .B2(n14492), .A(n14049), .ZN(P1_U2861) );
  INV_X1 U17203 ( .A(n14495), .ZN(n14051) );
  OAI222_X1 U17204 ( .A1(n15797), .A2(n14572), .B1(n14051), .B2(n14571), .C1(
        n14050), .C2(n9648), .ZN(P1_U2890) );
  INV_X1 U17205 ( .A(DATAI_11_), .ZN(n14053) );
  INV_X1 U17206 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14052) );
  MUX2_X1 U17207 ( .A(n14053), .B(n14052), .S(n20102), .Z(n20041) );
  OAI222_X1 U17208 ( .A1(n14055), .A2(n14572), .B1(n20041), .B2(n14571), .C1(
        n14054), .C2(n9648), .ZN(P1_U2893) );
  NOR2_X1 U17209 ( .A1(n14690), .A2(n20884), .ZN(n16045) );
  NAND2_X1 U17210 ( .A1(n16045), .A2(n16037), .ZN(n16035) );
  NOR3_X1 U17211 ( .A1(n16021), .A2(n15877), .A3(n16035), .ZN(n15971) );
  INV_X1 U17212 ( .A(n16045), .ZN(n14056) );
  NOR3_X1 U17213 ( .A1(n14058), .A2(n14057), .A3(n14056), .ZN(n16020) );
  NAND3_X1 U17214 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n16020), .ZN(n14076) );
  NOR3_X1 U17215 ( .A1(n20094), .A2(n20092), .A3(n14076), .ZN(n14059) );
  AOI21_X1 U17216 ( .B1(n15971), .B2(n20075), .A(n14059), .ZN(n14075) );
  NAND2_X1 U17217 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14060) );
  NAND3_X1 U17218 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15975) );
  NOR3_X1 U17219 ( .A1(n15982), .A2(n14060), .A3(n15975), .ZN(n14061) );
  NAND2_X1 U17220 ( .A1(n14061), .A2(n15971), .ZN(n14701) );
  INV_X1 U17221 ( .A(n14701), .ZN(n14063) );
  INV_X1 U17222 ( .A(n14076), .ZN(n15972) );
  NAND2_X1 U17223 ( .A1(n15972), .A2(n14061), .ZN(n14703) );
  OAI21_X1 U17224 ( .B1(n14066), .B2(n14703), .A(n14702), .ZN(n14062) );
  OAI211_X1 U17225 ( .C1(n20093), .C2(n14063), .A(n14062), .B(n20078), .ZN(
        n15965) );
  INV_X1 U17226 ( .A(n15965), .ZN(n14064) );
  OAI21_X1 U17227 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14075), .A(
        n14064), .ZN(n14074) );
  INV_X1 U17228 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20689) );
  NOR2_X1 U17229 ( .A1(n16057), .A2(n20689), .ZN(n14631) );
  INV_X1 U17230 ( .A(n14065), .ZN(n14643) );
  OAI21_X1 U17231 ( .B1(n15858), .B2(n15982), .A(n14643), .ZN(n14634) );
  NAND2_X1 U17232 ( .A1(n15874), .A2(n14066), .ZN(n14633) );
  NAND2_X1 U17233 ( .A1(n15858), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14737) );
  OAI22_X1 U17234 ( .A1(n14634), .A2(n14633), .B1(n14643), .B2(n14737), .ZN(
        n14068) );
  INV_X1 U17235 ( .A(n14068), .ZN(n14070) );
  NAND2_X1 U17236 ( .A1(n14068), .A2(n14067), .ZN(n14740) );
  INV_X1 U17237 ( .A(n14740), .ZN(n14069) );
  NOR2_X1 U17238 ( .A1(n14320), .A2(n14071), .ZN(n14072) );
  OR2_X1 U17239 ( .A1(n14446), .A2(n14072), .ZN(n15758) );
  OAI22_X1 U17240 ( .A1(n14629), .A2(n16073), .B1(n16079), .B2(n15758), .ZN(
        n14073) );
  AOI211_X1 U17241 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n14074), .A(
        n14631), .B(n14073), .ZN(n14079) );
  OAI21_X1 U17242 ( .B1(n14699), .B2(n14076), .A(n14075), .ZN(n16012) );
  NAND3_X1 U17243 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n16012), .ZN(n15995) );
  NOR2_X1 U17244 ( .A1(n15975), .A2(n15995), .ZN(n15980) );
  NAND2_X1 U17245 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15980), .ZN(
        n15970) );
  INV_X1 U17246 ( .A(n15970), .ZN(n14077) );
  NAND3_X1 U17247 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14067), .A3(
        n14077), .ZN(n14078) );
  NAND2_X1 U17248 ( .A1(n14079), .A2(n14078), .ZN(P1_U3011) );
  INV_X1 U17249 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18801) );
  NAND2_X1 U17250 ( .A1(n18801), .A2(n18791), .ZN(n18851) );
  NOR2_X2 U17251 ( .A1(n14089), .A2(n14086), .ZN(n15482) );
  AOI22_X1 U17252 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17253 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17254 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17255 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14080) );
  NAND4_X1 U17256 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14095) );
  INV_X2 U17257 ( .A(n15479), .ZN(n15423) );
  AOI22_X1 U17258 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U17259 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14092) );
  NOR2_X2 U17260 ( .A1(n14087), .A2(n14086), .ZN(n15486) );
  CLKBUF_X3 U17261 ( .A(n15486), .Z(n17186) );
  NOR2_X2 U17262 ( .A1(n14087), .A2(n18661), .ZN(n14106) );
  AOI22_X1 U17263 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17264 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14090) );
  NAND4_X1 U17265 ( .A1(n14093), .A2(n14092), .A3(n14091), .A4(n14090), .ZN(
        n14094) );
  AOI22_X1 U17266 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U17267 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17268 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U17269 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14096) );
  NAND4_X1 U17270 ( .A1(n14099), .A2(n14098), .A3(n14097), .A4(n14096), .ZN(
        n14105) );
  AOI22_X1 U17271 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U17272 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U17273 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14101) );
  AOI22_X1 U17274 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14100) );
  NAND4_X1 U17275 ( .A1(n14103), .A2(n14102), .A3(n14101), .A4(n14100), .ZN(
        n14104) );
  AOI22_X1 U17276 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n9647), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17188), .ZN(n14110) );
  AOI22_X1 U17277 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U17278 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17279 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n15518), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14107) );
  NAND4_X1 U17280 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        n14117) );
  AOI22_X1 U17281 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U17282 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17283 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9654), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17284 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n9653), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17097), .ZN(n14112) );
  NAND4_X1 U17285 ( .A1(n14115), .A2(n14114), .A3(n14113), .A4(n14112), .ZN(
        n14116) );
  INV_X2 U17286 ( .A(n17342), .ZN(n18234) );
  AOI22_X1 U17287 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17288 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17289 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14118) );
  OAI21_X1 U17290 ( .B1(n9694), .B2(n20869), .A(n14118), .ZN(n14124) );
  AOI22_X1 U17291 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17292 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17293 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U17294 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14119) );
  NAND4_X1 U17295 ( .A1(n14122), .A2(n14121), .A3(n14120), .A4(n14119), .ZN(
        n14123) );
  NAND3_X2 U17296 ( .A1(n14127), .A2(n14126), .A3(n14125), .ZN(n18195) );
  NAND2_X1 U17297 ( .A1(n18234), .A2(n15695), .ZN(n14174) );
  INV_X1 U17298 ( .A(n14174), .ZN(n14175) );
  AOI22_X1 U17299 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U17300 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U17301 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14129) );
  AOI22_X1 U17302 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14128) );
  NAND4_X1 U17303 ( .A1(n14131), .A2(n14130), .A3(n14129), .A4(n14128), .ZN(
        n14137) );
  AOI22_X1 U17304 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U17305 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14134) );
  AOI22_X1 U17306 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14133) );
  AOI22_X1 U17307 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14132) );
  NAND4_X1 U17308 ( .A1(n14135), .A2(n14134), .A3(n14133), .A4(n14132), .ZN(
        n14136) );
  AOI22_X1 U17309 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17310 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U17311 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U17312 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14138) );
  NAND4_X1 U17313 ( .A1(n14141), .A2(n14140), .A3(n14139), .A4(n14138), .ZN(
        n14147) );
  AOI22_X1 U17314 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U17315 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U17316 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9642), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17317 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14142) );
  NAND4_X1 U17318 ( .A1(n14145), .A2(n14144), .A3(n14143), .A4(n14142), .ZN(
        n14146) );
  NOR2_X1 U17319 ( .A1(n17239), .A2(n14168), .ZN(n15558) );
  NAND4_X1 U17320 ( .A1(n15415), .A2(n18213), .A3(n14175), .A4(n15558), .ZN(
        n14177) );
  AOI22_X1 U17321 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17322 ( .A1(n15518), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U17323 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U17324 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14148) );
  NAND4_X1 U17325 ( .A1(n14151), .A2(n14150), .A3(n14149), .A4(n14148), .ZN(
        n14157) );
  AOI22_X1 U17326 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U17327 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15344), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17328 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17329 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14152) );
  NAND4_X1 U17330 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14156) );
  NAND2_X1 U17331 ( .A1(n15559), .A2(n18224), .ZN(n15562) );
  INV_X1 U17332 ( .A(n15415), .ZN(n18219) );
  NAND2_X1 U17333 ( .A1(n17239), .A2(n18219), .ZN(n18635) );
  INV_X1 U17334 ( .A(n17239), .ZN(n18229) );
  NAND2_X1 U17335 ( .A1(n14168), .A2(n18229), .ZN(n14193) );
  NAND3_X1 U17336 ( .A1(n15559), .A2(n18635), .A3(n14193), .ZN(n14169) );
  NAND2_X1 U17337 ( .A1(n15562), .A2(n14169), .ZN(n14176) );
  AOI22_X1 U17338 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U17339 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U17340 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U17341 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14158) );
  NAND4_X1 U17342 ( .A1(n14161), .A2(n14160), .A3(n14159), .A4(n14158), .ZN(
        n14167) );
  AOI22_X1 U17343 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14165) );
  AOI22_X1 U17344 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14164) );
  AOI22_X1 U17345 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14163) );
  AOI22_X1 U17346 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14162) );
  NAND4_X1 U17347 ( .A1(n14165), .A2(n14164), .A3(n14163), .A4(n14162), .ZN(
        n14166) );
  NOR2_X1 U17348 ( .A1(n15695), .A2(n18203), .ZN(n15602) );
  NOR2_X1 U17349 ( .A1(n18229), .A2(n14168), .ZN(n14194) );
  NAND2_X1 U17350 ( .A1(n18234), .A2(n18645), .ZN(n15698) );
  NAND2_X1 U17351 ( .A1(n15602), .A2(n15698), .ZN(n14198) );
  NOR2_X1 U17352 ( .A1(n18195), .A2(n14169), .ZN(n14173) );
  NOR2_X1 U17353 ( .A1(n17342), .A2(n15558), .ZN(n14171) );
  INV_X1 U17354 ( .A(n15603), .ZN(n14178) );
  NAND2_X1 U17355 ( .A1(n15559), .A2(n14178), .ZN(n14196) );
  AOI21_X1 U17356 ( .B1(n15415), .B2(n18224), .A(n14196), .ZN(n14170) );
  OAI22_X1 U17357 ( .A1(n15415), .A2(n14171), .B1(n15558), .B2(n14170), .ZN(
        n14172) );
  AOI211_X1 U17358 ( .C1(n18213), .C2(n14174), .A(n14173), .B(n14172), .ZN(
        n14197) );
  OAI211_X1 U17359 ( .C1(n18213), .C2(n14176), .A(n14198), .B(n14197), .ZN(
        n15607) );
  NOR2_X1 U17360 ( .A1(n14177), .A2(n15607), .ZN(n15601) );
  NAND2_X1 U17361 ( .A1(n15559), .A2(n18213), .ZN(n18634) );
  NOR2_X1 U17362 ( .A1(n14193), .A2(n18634), .ZN(n15414) );
  NAND3_X1 U17363 ( .A1(n14175), .A2(n15414), .A3(n18841), .ZN(n14179) );
  INV_X1 U17364 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16865) );
  NAND2_X1 U17365 ( .A1(n14180), .A2(n16865), .ZN(n14211) );
  NAND2_X1 U17366 ( .A1(n18660), .A2(n14211), .ZN(n18674) );
  NOR2_X1 U17367 ( .A1(n18851), .A2(n18674), .ZN(n14210) );
  NOR2_X1 U17368 ( .A1(n18203), .A2(n17429), .ZN(n18681) );
  NOR2_X2 U17369 ( .A1(n20897), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18777) );
  AND2_X1 U17370 ( .A1(n18832), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18724) );
  NOR2_X1 U17371 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18702) );
  NOR3_X1 U17372 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18724), .A3(n18702), 
        .ZN(n16542) );
  OAI21_X1 U17373 ( .B1(n14181), .B2(n18681), .A(n16542), .ZN(n17389) );
  NAND2_X1 U17374 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18842) );
  INV_X1 U17375 ( .A(n18842), .ZN(n18708) );
  AOI22_X1 U17376 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18651), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18815), .ZN(n14203) );
  XNOR2_X1 U17377 ( .A(n14203), .B(n14201), .ZN(n14192) );
  OAI22_X1 U17378 ( .A1(n18808), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18192), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14187) );
  OAI22_X1 U17379 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18191), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14184), .ZN(n14189) );
  NOR2_X1 U17380 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18191), .ZN(
        n14185) );
  NAND2_X1 U17381 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14184), .ZN(
        n14190) );
  AOI22_X1 U17382 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14189), .B1(
        n14185), .B2(n14190), .ZN(n14202) );
  NAND2_X1 U17383 ( .A1(n14188), .A2(n14187), .ZN(n14186) );
  OAI211_X1 U17384 ( .C1(n14188), .C2(n14187), .A(n14202), .B(n14186), .ZN(
        n15566) );
  AOI21_X1 U17385 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14190), .A(
        n14189), .ZN(n14191) );
  AOI211_X1 U17386 ( .C1(n15697), .C2(n17389), .A(n18708), .B(n16522), .ZN(
        n14208) );
  OAI211_X1 U17387 ( .C1(n15415), .C2(n14194), .A(n15606), .B(n14193), .ZN(
        n14195) );
  NOR2_X1 U17388 ( .A1(n14196), .A2(n14195), .ZN(n15557) );
  NAND2_X1 U17389 ( .A1(n15557), .A2(n14197), .ZN(n14200) );
  INV_X1 U17390 ( .A(n14198), .ZN(n14199) );
  AOI21_X1 U17391 ( .B1(n14200), .B2(n16524), .A(n14199), .ZN(n15564) );
  AOI21_X1 U17392 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20913), .A(
        n14201), .ZN(n15567) );
  NAND3_X1 U17393 ( .A1(n14203), .A2(n14202), .A3(n15567), .ZN(n14204) );
  NAND3_X1 U17394 ( .A1(n14205), .A2(n15566), .A3(n14204), .ZN(n16349) );
  INV_X1 U17395 ( .A(n16349), .ZN(n18630) );
  NAND2_X1 U17396 ( .A1(n18630), .A2(n15604), .ZN(n15417) );
  NAND2_X1 U17397 ( .A1(n15564), .A2(n15417), .ZN(n14207) );
  NAND2_X1 U17398 ( .A1(n18788), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18193) );
  INV_X1 U17399 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16526) );
  NAND3_X1 U17400 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18790)
         );
  OR2_X1 U17401 ( .A1(n16526), .A2(n18790), .ZN(n14209) );
  OAI211_X1 U17402 ( .C1(n18688), .C2(n18678), .A(n18193), .B(n14209), .ZN(
        n18820) );
  INV_X1 U17403 ( .A(n18820), .ZN(n18822) );
  MUX2_X1 U17404 ( .A(n14210), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18822), .Z(P3_U3284) );
  NOR2_X1 U17405 ( .A1(n15518), .A2(n14211), .ZN(n18183) );
  NOR2_X1 U17406 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18844) );
  AOI21_X1 U17407 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18844), .ZN(n18697) );
  OAI221_X1 U17408 ( .B1(n18790), .B2(n18183), .C1(n18790), .C2(n16526), .A(
        n18265), .ZN(n18190) );
  INV_X1 U17409 ( .A(n18190), .ZN(n18186) );
  INV_X1 U17410 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18840) );
  NOR2_X1 U17411 ( .A1(n18801), .A2(n18840), .ZN(n17831) );
  INV_X1 U17412 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18682) );
  NAND2_X1 U17413 ( .A1(n18682), .A2(n18791), .ZN(n16520) );
  NAND2_X1 U17414 ( .A1(n18851), .A2(n16520), .ZN(n18184) );
  INV_X1 U17415 ( .A(n18184), .ZN(n18835) );
  NOR2_X1 U17416 ( .A1(n17831), .A2(n18835), .ZN(n15438) );
  AOI21_X1 U17417 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15438), .ZN(n15439) );
  NOR2_X1 U17418 ( .A1(n18186), .A2(n15439), .ZN(n14213) );
  NAND3_X1 U17419 ( .A1(n18682), .A2(n18791), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18540) );
  INV_X1 U17420 ( .A(n18540), .ZN(n18447) );
  NAND2_X1 U17421 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18650), .ZN(n18243) );
  NAND2_X1 U17422 ( .A1(n18243), .A2(n18190), .ZN(n15437) );
  OR2_X1 U17423 ( .A1(n18447), .A2(n15437), .ZN(n14212) );
  MUX2_X1 U17424 ( .A(n14213), .B(n14212), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17425 ( .A(n14217), .ZN(n14214) );
  NAND2_X1 U17426 ( .A1(n14214), .A2(n20102), .ZN(n14508) );
  AND2_X1 U17427 ( .A1(n9648), .A2(n20147), .ZN(n14215) );
  NAND2_X1 U17428 ( .A1(n14216), .A2(n14215), .ZN(n14219) );
  AOI22_X1 U17429 ( .A1(n14562), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14567), .ZN(n14218) );
  OAI211_X1 U17430 ( .C1(n14508), .C2(n16423), .A(n14219), .B(n14218), .ZN(
        P1_U2873) );
  NOR2_X2 U17431 ( .A1(n14222), .A2(n14220), .ZN(n19084) );
  NOR2_X2 U17432 ( .A1(n14222), .A2(n14221), .ZN(n19085) );
  AOI22_X1 U17433 ( .A1(n19084), .A2(BUF2_REG_30__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U17434 ( .A1(n16190), .A2(n19090), .B1(n19137), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14223) );
  OAI211_X1 U17435 ( .C1(n14245), .C2(n14962), .A(n14224), .B(n14223), .ZN(
        n14225) );
  INV_X1 U17436 ( .A(n14225), .ZN(n14226) );
  OAI21_X1 U17437 ( .B1(n14227), .B2(n14947), .A(n14226), .ZN(P2_U2889) );
  XNOR2_X1 U17438 ( .A(n12558), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14253) );
  NAND2_X1 U17439 ( .A1(n14229), .A2(n14228), .ZN(n14234) );
  INV_X1 U17440 ( .A(n14230), .ZN(n14232) );
  NAND2_X1 U17441 ( .A1(n14232), .A2(n14231), .ZN(n14233) );
  NAND2_X1 U17442 ( .A1(n14240), .A2(n19222), .ZN(n14239) );
  NOR2_X1 U17443 ( .A1(n19023), .A2(n14235), .ZN(n14241) );
  AOI21_X1 U17444 ( .B1(n19230), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14241), .ZN(n14236) );
  OAI21_X1 U17445 ( .B1(n16256), .B2(n16104), .A(n14236), .ZN(n14237) );
  AOI21_X1 U17446 ( .B1(n14250), .B2(n19239), .A(n14237), .ZN(n14238) );
  NAND2_X1 U17447 ( .A1(n14240), .A2(n16334), .ZN(n14252) );
  INV_X1 U17448 ( .A(n14241), .ZN(n14244) );
  INV_X1 U17449 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14246) );
  NAND3_X1 U17450 ( .A1(n14242), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14246), .ZN(n14243) );
  OAI211_X1 U17451 ( .C1(n16324), .C2(n14245), .A(n14244), .B(n14243), .ZN(
        n14249) );
  NOR2_X1 U17452 ( .A1(n14247), .A2(n14246), .ZN(n14248) );
  AOI211_X1 U17453 ( .C1(n16312), .C2(n14250), .A(n14249), .B(n14248), .ZN(
        n14251) );
  OAI211_X1 U17454 ( .C1(n14253), .C2(n16330), .A(n14252), .B(n14251), .ZN(
        P2_U3016) );
  INV_X1 U17455 ( .A(n14254), .ZN(n14255) );
  AOI22_X1 U17456 ( .A1(n14277), .A2(n14256), .B1(n14255), .B2(n14284), .ZN(
        n14258) );
  XNOR2_X1 U17457 ( .A(n14258), .B(n14257), .ZN(n14720) );
  NAND2_X1 U17458 ( .A1(n14580), .A2(n19958), .ZN(n14268) );
  INV_X1 U17459 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14582) );
  INV_X1 U17460 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14261) );
  OAI21_X1 U17461 ( .B1(n14274), .B2(n14582), .A(n14261), .ZN(n14265) );
  INV_X1 U17462 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14408) );
  NOR2_X1 U17463 ( .A1(n19984), .A2(n14408), .ZN(n14264) );
  OAI22_X1 U17464 ( .A1(n14262), .A2(n19996), .B1(n19995), .B2(n14578), .ZN(
        n14263) );
  AOI211_X1 U17465 ( .C1(n14266), .C2(n14265), .A(n14264), .B(n14263), .ZN(
        n14267) );
  OAI211_X1 U17466 ( .C1(n19985), .C2(n14720), .A(n14268), .B(n14267), .ZN(
        P1_U2810) );
  OAI21_X1 U17467 ( .B1(n14269), .B2(n14271), .A(n14270), .ZN(n14592) );
  INV_X1 U17468 ( .A(n14289), .ZN(n14280) );
  AOI22_X1 U17469 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19977), .B1(
        n19989), .B2(n14585), .ZN(n14273) );
  NAND2_X1 U17470 ( .A1(n19997), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14272) );
  OAI211_X1 U17471 ( .C1(n14274), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14273), 
        .B(n14272), .ZN(n14279) );
  OR2_X1 U17472 ( .A1(n14284), .A2(n14275), .ZN(n14276) );
  NAND2_X1 U17473 ( .A1(n14277), .A2(n14276), .ZN(n14732) );
  NOR2_X1 U17474 ( .A1(n14732), .A2(n19985), .ZN(n14278) );
  AOI211_X1 U17475 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14280), .A(n14279), 
        .B(n14278), .ZN(n14281) );
  OAI21_X1 U17476 ( .B1(n14592), .B2(n19944), .A(n14281), .ZN(P1_U2811) );
  NOR2_X1 U17477 ( .A1(n9732), .A2(n14282), .ZN(n14283) );
  AOI21_X1 U17478 ( .B1(n14286), .B2(n14295), .A(n14269), .ZN(n14604) );
  NAND2_X1 U17479 ( .A1(n14604), .A2(n19958), .ZN(n14293) );
  OAI22_X1 U17480 ( .A1(n14287), .A2(n19996), .B1(n19995), .B2(n14602), .ZN(
        n14291) );
  AOI21_X1 U17481 ( .B1(n14298), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14288) );
  NOR2_X1 U17482 ( .A1(n14289), .A2(n14288), .ZN(n14290) );
  AOI211_X1 U17483 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n19997), .A(n14291), .B(
        n14290), .ZN(n14292) );
  OAI211_X1 U17484 ( .C1(n15911), .C2(n19985), .A(n14293), .B(n14292), .ZN(
        P1_U2812) );
  OAI21_X2 U17485 ( .B1(n14294), .B2(n14296), .A(n14295), .ZN(n14610) );
  AOI21_X1 U17486 ( .B1(n14297), .B2(n14417), .A(n9732), .ZN(n15913) );
  INV_X1 U17487 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15915) );
  AOI22_X1 U17488 ( .A1(n14613), .A2(n19989), .B1(n14298), .B2(n15915), .ZN(
        n14300) );
  AOI22_X1 U17489 ( .A1(n15708), .A2(P1_REIP_REG_27__SCAN_IN), .B1(n19997), 
        .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n14299) );
  OAI211_X1 U17490 ( .C1(n14609), .C2(n19996), .A(n14300), .B(n14299), .ZN(
        n14301) );
  AOI21_X1 U17491 ( .B1(n15913), .B2(n19994), .A(n14301), .ZN(n14302) );
  OAI21_X1 U17492 ( .B1(n14610), .B2(n19944), .A(n14302), .ZN(P1_U2813) );
  INV_X1 U17493 ( .A(n14304), .ZN(n14305) );
  AOI21_X1 U17494 ( .B1(n14306), .B2(n14303), .A(n14305), .ZN(n14619) );
  INV_X1 U17495 ( .A(n14619), .ZN(n14524) );
  NOR2_X1 U17496 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15803), .ZN(n15713) );
  OR2_X1 U17497 ( .A1(n15714), .A2(n15803), .ZN(n14307) );
  NAND2_X1 U17498 ( .A1(n14307), .A2(n15779), .ZN(n15722) );
  OAI21_X1 U17499 ( .B1(n15713), .B2(n15722), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14315) );
  OR2_X1 U17500 ( .A1(n14423), .A2(n14308), .ZN(n14309) );
  AND2_X1 U17501 ( .A1(n14309), .A2(n14415), .ZN(n15930) );
  NOR3_X1 U17502 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15803), .A3(n14310), 
        .ZN(n14313) );
  AOI22_X1 U17503 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(n19997), .B1(n19989), 
        .B2(n14622), .ZN(n14311) );
  OAI21_X1 U17504 ( .B1(n14620), .B2(n19996), .A(n14311), .ZN(n14312) );
  AOI211_X1 U17505 ( .C1(n15930), .C2(n19994), .A(n14313), .B(n14312), .ZN(
        n14314) );
  OAI211_X1 U17506 ( .C1(n14524), .C2(n19944), .A(n14315), .B(n14314), .ZN(
        P1_U2815) );
  XNOR2_X1 U17507 ( .A(n14455), .B(n14316), .ZN(n14642) );
  NOR3_X1 U17508 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15803), .A3(n14317), 
        .ZN(n15762) );
  AOI21_X1 U17509 ( .B1(n14317), .B2(n15771), .A(n19976), .ZN(n14340) );
  INV_X1 U17510 ( .A(n14340), .ZN(n15763) );
  OAI21_X1 U17511 ( .B1(n15762), .B2(n15763), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14327) );
  AND2_X1 U17512 ( .A1(n14460), .A2(n14318), .ZN(n14319) );
  NOR2_X1 U17513 ( .A1(n14320), .A2(n14319), .ZN(n15966) );
  AOI22_X1 U17514 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19997), .B1(n19989), 
        .B2(n14639), .ZN(n14321) );
  OAI211_X1 U17515 ( .C1(n19996), .C2(n14637), .A(n14321), .B(n19963), .ZN(
        n14325) );
  INV_X1 U17516 ( .A(n14322), .ZN(n14323) );
  NOR3_X1 U17517 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15803), .A3(n14323), 
        .ZN(n14324) );
  AOI211_X1 U17518 ( .C1(n15966), .C2(n19994), .A(n14325), .B(n14324), .ZN(
        n14326) );
  OAI211_X1 U17519 ( .C1(n14642), .C2(n19944), .A(n14327), .B(n14326), .ZN(
        P1_U2821) );
  AOI21_X1 U17520 ( .B1(n15771), .B2(n14328), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14341) );
  INV_X1 U17521 ( .A(n14329), .ZN(n14454) );
  AOI21_X1 U17522 ( .B1(n14330), .B2(n14467), .A(n14329), .ZN(n14658) );
  NAND2_X1 U17523 ( .A1(n14658), .A2(n19958), .ZN(n14339) );
  OR2_X1 U17524 ( .A1(n14469), .A2(n14331), .ZN(n14332) );
  AND2_X1 U17525 ( .A1(n14458), .A2(n14332), .ZN(n15986) );
  NAND2_X1 U17526 ( .A1(n19997), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14336) );
  INV_X1 U17527 ( .A(n14656), .ZN(n14333) );
  NAND2_X1 U17528 ( .A1(n19989), .A2(n14333), .ZN(n14335) );
  NAND2_X1 U17529 ( .A1(n19977), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14334) );
  NAND4_X1 U17530 ( .A1(n14336), .A2(n14335), .A3(n14334), .A4(n19963), .ZN(
        n14337) );
  AOI21_X1 U17531 ( .B1(n15986), .B2(n19994), .A(n14337), .ZN(n14338) );
  OAI211_X1 U17532 ( .C1(n14341), .C2(n14340), .A(n14339), .B(n14338), .ZN(
        P1_U2823) );
  AOI21_X1 U17533 ( .B1(n11906), .B2(n14343), .A(n14342), .ZN(n14491) );
  NOR2_X1 U17534 ( .A1(n14491), .A2(n14490), .ZN(n14489) );
  OAI21_X1 U17535 ( .B1(n14489), .B2(n14344), .A(n14034), .ZN(n14686) );
  NOR2_X1 U17536 ( .A1(n15803), .A2(n14348), .ZN(n15793) );
  AOI21_X1 U17537 ( .B1(n14346), .B2(n14488), .A(n14345), .ZN(n16013) );
  INV_X1 U17538 ( .A(n16013), .ZN(n14347) );
  OAI22_X1 U17539 ( .A1(n14347), .A2(n19985), .B1(n14673), .B2(n19995), .ZN(
        n14351) );
  AOI21_X1 U17540 ( .B1(n15771), .B2(n14348), .A(n19976), .ZN(n15808) );
  AOI22_X1 U17541 ( .A1(n19997), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19977), .ZN(n14349) );
  OAI211_X1 U17542 ( .C1(n20676), .C2(n15808), .A(n14349), .B(n19963), .ZN(
        n14350) );
  AOI211_X1 U17543 ( .C1(n15793), .C2(n20676), .A(n14351), .B(n14350), .ZN(
        n14352) );
  OAI21_X1 U17544 ( .B1(n14686), .B2(n19944), .A(n14352), .ZN(P1_U2827) );
  OAI21_X1 U17545 ( .B1(n15803), .B2(n14356), .A(n15779), .ZN(n15811) );
  NOR2_X1 U17546 ( .A1(n19995), .A2(n14694), .ZN(n14353) );
  AOI211_X1 U17547 ( .C1(n19977), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19955), .B(n14353), .ZN(n14354) );
  OAI21_X1 U17548 ( .B1(n14355), .B2(n19984), .A(n14354), .ZN(n14360) );
  INV_X1 U17549 ( .A(n14356), .ZN(n15802) );
  NAND2_X1 U17550 ( .A1(n15771), .A2(n15802), .ZN(n14357) );
  OAI22_X1 U17551 ( .A1(n19985), .A2(n16038), .B1(n14358), .B2(n14357), .ZN(
        n14359) );
  AOI211_X1 U17552 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15811), .A(n14360), 
        .B(n14359), .ZN(n14361) );
  OAI21_X1 U17553 ( .B1(n14362), .B2(n19944), .A(n14361), .ZN(P1_U2830) );
  INV_X1 U17554 ( .A(n14363), .ZN(n14373) );
  NAND2_X1 U17555 ( .A1(n14373), .A2(n14364), .ZN(n14365) );
  AOI21_X1 U17556 ( .B1(n14366), .B2(n15771), .A(n19976), .ZN(n14367) );
  INV_X1 U17557 ( .A(n14367), .ZN(n19969) );
  OAI21_X1 U17558 ( .B1(n14368), .B2(P1_REIP_REG_4__SCAN_IN), .A(n19969), .ZN(
        n14379) );
  NOR2_X1 U17559 ( .A1(n19984), .A2(n14369), .ZN(n14377) );
  INV_X1 U17560 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14370) );
  OAI22_X1 U17561 ( .A1(n14371), .A2(n19995), .B1(n19996), .B2(n14370), .ZN(
        n14376) );
  NAND2_X1 U17562 ( .A1(n14373), .A2(n14372), .ZN(n19980) );
  OAI22_X1 U17563 ( .A1(n19985), .A2(n14374), .B1(n16080), .B2(n19980), .ZN(
        n14375) );
  NOR4_X1 U17564 ( .A1(n14377), .A2(n14376), .A3(n19955), .A4(n14375), .ZN(
        n14378) );
  OAI211_X1 U17565 ( .C1(n20002), .C2(n14380), .A(n14379), .B(n14378), .ZN(
        P1_U2836) );
  NAND3_X1 U17566 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14381) );
  AND2_X1 U17567 ( .A1(n15771), .A2(n14381), .ZN(n14384) );
  NAND2_X1 U17568 ( .A1(n13593), .A2(n14382), .ZN(n14383) );
  OAI21_X1 U17569 ( .B1(n19976), .B2(n14384), .A(n14383), .ZN(n14392) );
  INV_X1 U17570 ( .A(n19980), .ZN(n19998) );
  OAI22_X1 U17571 ( .A1(n14386), .A2(n19995), .B1(n19996), .B2(n14385), .ZN(
        n14387) );
  AOI21_X1 U17572 ( .B1(n19997), .B2(P1_EBX_REG_3__SCAN_IN), .A(n14387), .ZN(
        n14388) );
  OAI21_X1 U17573 ( .B1(n19985), .B2(n14389), .A(n14388), .ZN(n14390) );
  AOI21_X1 U17574 ( .B1(n20711), .B2(n19998), .A(n14390), .ZN(n14391) );
  OAI211_X1 U17575 ( .C1(n20002), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P1_U2837) );
  NAND2_X1 U17576 ( .A1(n15771), .A2(n20724), .ZN(n19978) );
  INV_X1 U17577 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14394) );
  AOI21_X1 U17578 ( .B1(n19978), .B2(n15779), .A(n14394), .ZN(n14404) );
  XNOR2_X1 U17579 ( .A(n13569), .B(n14395), .ZN(n20073) );
  INV_X1 U17580 ( .A(n20073), .ZN(n14402) );
  NOR2_X1 U17581 ( .A1(n19995), .A2(n14396), .ZN(n14400) );
  INV_X1 U17582 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14398) );
  NAND2_X1 U17583 ( .A1(n15771), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14397) );
  OAI22_X1 U17584 ( .A1(n19996), .A2(n14398), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n14397), .ZN(n14399) );
  AOI211_X1 U17585 ( .C1(P1_EBX_REG_2__SCAN_IN), .C2(n19997), .A(n14400), .B(
        n14399), .ZN(n14401) );
  OAI21_X1 U17586 ( .B1(n14402), .B2(n19985), .A(n14401), .ZN(n14403) );
  AOI211_X1 U17587 ( .C1(n19998), .C2(n20112), .A(n14404), .B(n14403), .ZN(
        n14405) );
  OAI21_X1 U17588 ( .B1(n14406), .B2(n20002), .A(n14405), .ZN(P1_U2838) );
  INV_X1 U17589 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14407) );
  OAI22_X1 U17590 ( .A1(n14711), .A2(n14494), .B1(n20008), .B2(n14407), .ZN(
        P1_U2841) );
  OAI222_X1 U17591 ( .A1(n14492), .A2(n14500), .B1(n14408), .B2(n20008), .C1(
        n14720), .C2(n14494), .ZN(P1_U2842) );
  OAI222_X1 U17592 ( .A1(n14492), .A2(n14592), .B1(n14409), .B2(n20008), .C1(
        n14732), .C2(n14494), .ZN(P1_U2843) );
  INV_X1 U17593 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14410) );
  INV_X1 U17594 ( .A(n14604), .ZN(n14513) );
  OAI222_X1 U17595 ( .A1(n15911), .A2(n14494), .B1(n14410), .B2(n20008), .C1(
        n14513), .C2(n14492), .ZN(P1_U2844) );
  AOI22_X1 U17596 ( .A1(n15913), .A2(n20003), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14483), .ZN(n14411) );
  OAI21_X1 U17597 ( .B1(n14610), .B2(n14492), .A(n14411), .ZN(P1_U2845) );
  AND2_X1 U17598 ( .A1(n14304), .A2(n14412), .ZN(n14413) );
  NAND2_X1 U17599 ( .A1(n14415), .A2(n14414), .ZN(n14416) );
  NAND2_X1 U17600 ( .A1(n14417), .A2(n14416), .ZN(n15928) );
  OAI22_X1 U17601 ( .A1(n15928), .A2(n14494), .B1(n15704), .B2(n20008), .ZN(
        n14418) );
  INV_X1 U17602 ( .A(n14418), .ZN(n14419) );
  OAI21_X1 U17603 ( .B1(n15817), .B2(n14492), .A(n14419), .ZN(P1_U2846) );
  AOI22_X1 U17604 ( .A1(n15930), .A2(n20003), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14483), .ZN(n14420) );
  OAI21_X1 U17605 ( .B1(n14524), .B2(n14492), .A(n14420), .ZN(P1_U2847) );
  OAI21_X1 U17606 ( .B1(n14421), .B2(n14422), .A(n14303), .ZN(n15712) );
  INV_X1 U17607 ( .A(n14423), .ZN(n14426) );
  NAND2_X1 U17608 ( .A1(n14434), .A2(n14424), .ZN(n14425) );
  NAND2_X1 U17609 ( .A1(n14426), .A2(n14425), .ZN(n15947) );
  OAI22_X1 U17610 ( .A1(n15947), .A2(n14494), .B1(n14427), .B2(n20008), .ZN(
        n14428) );
  INV_X1 U17611 ( .A(n14428), .ZN(n14429) );
  OAI21_X1 U17612 ( .B1(n15712), .B2(n14492), .A(n14429), .ZN(P1_U2848) );
  AOI21_X1 U17613 ( .B1(n14430), .B2(n14438), .A(n14421), .ZN(n14431) );
  INV_X1 U17614 ( .A(n14431), .ZN(n15725) );
  INV_X1 U17615 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14435) );
  NAND2_X1 U17616 ( .A1(n9697), .A2(n14432), .ZN(n14433) );
  NAND2_X1 U17617 ( .A1(n14434), .A2(n14433), .ZN(n15720) );
  OAI222_X1 U17618 ( .A1(n14492), .A2(n15725), .B1(n14435), .B2(n20008), .C1(
        n15720), .C2(n14494), .ZN(P1_U2849) );
  NAND2_X1 U17619 ( .A1(n9700), .A2(n14436), .ZN(n14437) );
  AND2_X1 U17620 ( .A1(n14438), .A2(n14437), .ZN(n15837) );
  NAND2_X1 U17621 ( .A1(n9746), .A2(n14439), .ZN(n14440) );
  NAND2_X1 U17622 ( .A1(n9697), .A2(n14440), .ZN(n15731) );
  INV_X1 U17623 ( .A(n15731), .ZN(n15958) );
  AOI22_X1 U17624 ( .A1(n15958), .A2(n20003), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14483), .ZN(n14441) );
  OAI21_X1 U17625 ( .B1(n15732), .B2(n14492), .A(n14441), .ZN(P1_U2850) );
  NAND2_X1 U17626 ( .A1(n14442), .A2(n14443), .ZN(n14444) );
  AND2_X1 U17627 ( .A1(n9700), .A2(n14444), .ZN(n15842) );
  INV_X1 U17628 ( .A(n15842), .ZN(n14541) );
  INV_X1 U17629 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14448) );
  OR2_X1 U17630 ( .A1(n14446), .A2(n14445), .ZN(n14447) );
  NAND2_X1 U17631 ( .A1(n9746), .A2(n14447), .ZN(n15741) );
  OAI222_X1 U17632 ( .A1(n14541), .A2(n14492), .B1(n14448), .B2(n20008), .C1(
        n15741), .C2(n14494), .ZN(P1_U2851) );
  OAI21_X1 U17633 ( .B1(n14450), .B2(n14449), .A(n14442), .ZN(n15755) );
  INV_X1 U17634 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14451) );
  OAI222_X1 U17635 ( .A1(n15755), .A2(n14492), .B1(n20008), .B2(n14451), .C1(
        n15758), .C2(n14494), .ZN(P1_U2852) );
  AOI22_X1 U17636 ( .A1(n15966), .A2(n20003), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14483), .ZN(n14452) );
  OAI21_X1 U17637 ( .B1(n14642), .B2(n14492), .A(n14452), .ZN(P1_U2853) );
  AND2_X1 U17638 ( .A1(n14454), .A2(n14453), .ZN(n14456) );
  OR2_X1 U17639 ( .A1(n14456), .A2(n14455), .ZN(n15765) );
  NAND2_X1 U17640 ( .A1(n14458), .A2(n14457), .ZN(n14459) );
  NAND2_X1 U17641 ( .A1(n14460), .A2(n14459), .ZN(n15976) );
  OAI22_X1 U17642 ( .A1(n15976), .A2(n14494), .B1(n15760), .B2(n20008), .ZN(
        n14461) );
  INV_X1 U17643 ( .A(n14461), .ZN(n14462) );
  OAI21_X1 U17644 ( .B1(n15765), .B2(n14492), .A(n14462), .ZN(P1_U2854) );
  INV_X1 U17645 ( .A(n14658), .ZN(n14557) );
  AOI22_X1 U17646 ( .A1(n15986), .A2(n20003), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14483), .ZN(n14463) );
  OAI21_X1 U17647 ( .B1(n14557), .B2(n14492), .A(n14463), .ZN(P1_U2855) );
  OR2_X1 U17648 ( .A1(n14464), .A2(n14465), .ZN(n14466) );
  AND2_X1 U17649 ( .A1(n14467), .A2(n14466), .ZN(n15851) );
  INV_X1 U17650 ( .A(n15851), .ZN(n14565) );
  AND2_X1 U17651 ( .A1(n14479), .A2(n14468), .ZN(n14470) );
  OR2_X1 U17652 ( .A1(n14470), .A2(n14469), .ZN(n15998) );
  OAI22_X1 U17653 ( .A1(n15998), .A2(n14494), .B1(n14471), .B2(n20008), .ZN(
        n14472) );
  INV_X1 U17654 ( .A(n14472), .ZN(n14473) );
  OAI21_X1 U17655 ( .B1(n14565), .B2(n14492), .A(n14473), .ZN(P1_U2856) );
  INV_X1 U17656 ( .A(n14464), .ZN(n14474) );
  OAI21_X1 U17657 ( .B1(n14036), .B2(n14475), .A(n14474), .ZN(n15789) );
  NAND2_X1 U17658 ( .A1(n14477), .A2(n14476), .ZN(n14478) );
  NAND2_X1 U17659 ( .A1(n14479), .A2(n14478), .ZN(n16004) );
  OAI22_X1 U17660 ( .A1(n16004), .A2(n14494), .B1(n14480), .B2(n20008), .ZN(
        n14481) );
  INV_X1 U17661 ( .A(n14481), .ZN(n14482) );
  OAI21_X1 U17662 ( .B1(n15789), .B2(n14492), .A(n14482), .ZN(P1_U2857) );
  AOI22_X1 U17663 ( .A1(n16013), .A2(n20003), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14483), .ZN(n14484) );
  OAI21_X1 U17664 ( .B1(n14686), .B2(n14492), .A(n14484), .ZN(P1_U2859) );
  NAND2_X1 U17665 ( .A1(n14486), .A2(n14485), .ZN(n14487) );
  NAND2_X1 U17666 ( .A1(n14488), .A2(n14487), .ZN(n16028) );
  INV_X1 U17667 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14493) );
  AOI21_X1 U17668 ( .B1(n14491), .B2(n14490), .A(n14489), .ZN(n15869) );
  INV_X1 U17669 ( .A(n15869), .ZN(n14573) );
  OAI222_X1 U17670 ( .A1(n16028), .A2(n14494), .B1(n14493), .B2(n20008), .C1(
        n14573), .C2(n14492), .ZN(P1_U2860) );
  INV_X1 U17671 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U17672 ( .A1(n14503), .A2(n14495), .B1(n14567), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14496) );
  OAI21_X1 U17673 ( .B1(n14508), .B2(n14497), .A(n14496), .ZN(n14498) );
  AOI21_X1 U17674 ( .B1(n14562), .B2(DATAI_30_), .A(n14498), .ZN(n14499) );
  OAI21_X1 U17675 ( .B1(n14500), .B2(n14572), .A(n14499), .ZN(P1_U2874) );
  INV_X1 U17676 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14505) );
  INV_X1 U17677 ( .A(DATAI_13_), .ZN(n14502) );
  NAND2_X1 U17678 ( .A1(n20102), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14501) );
  OAI21_X1 U17679 ( .B1(n20102), .B2(n14502), .A(n14501), .ZN(n20047) );
  AOI22_X1 U17680 ( .A1(n14503), .A2(n20047), .B1(n14567), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14504) );
  OAI21_X1 U17681 ( .B1(n14508), .B2(n14505), .A(n14504), .ZN(n14506) );
  AOI21_X1 U17682 ( .B1(n14562), .B2(DATAI_29_), .A(n14506), .ZN(n14507) );
  OAI21_X1 U17683 ( .B1(n14592), .B2(n14572), .A(n14507), .ZN(P1_U2875) );
  INV_X1 U17684 ( .A(DATAI_12_), .ZN(n14509) );
  MUX2_X1 U17685 ( .A(n14509), .B(n16455), .S(n20102), .Z(n20044) );
  OAI22_X1 U17686 ( .A1(n14559), .A2(n20044), .B1(n9648), .B2(n13323), .ZN(
        n14510) );
  AOI21_X1 U17687 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14561), .A(n14510), .ZN(
        n14512) );
  NAND2_X1 U17688 ( .A1(n14562), .A2(DATAI_28_), .ZN(n14511) );
  OAI211_X1 U17689 ( .C1(n14513), .C2(n14572), .A(n14512), .B(n14511), .ZN(
        P1_U2876) );
  OAI22_X1 U17690 ( .A1(n14559), .A2(n20041), .B1(n9648), .B2(n13332), .ZN(
        n14514) );
  AOI21_X1 U17691 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14561), .A(n14514), .ZN(
        n14516) );
  NAND2_X1 U17692 ( .A1(n14562), .A2(DATAI_27_), .ZN(n14515) );
  OAI211_X1 U17693 ( .C1(n14610), .C2(n14572), .A(n14516), .B(n14515), .ZN(
        P1_U2877) );
  OAI22_X1 U17694 ( .A1(n14559), .A2(n20038), .B1(n9648), .B2(n14517), .ZN(
        n14518) );
  AOI21_X1 U17695 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14561), .A(n14518), .ZN(
        n14520) );
  NAND2_X1 U17696 ( .A1(n14562), .A2(DATAI_26_), .ZN(n14519) );
  OAI211_X1 U17697 ( .C1(n15817), .C2(n14572), .A(n14520), .B(n14519), .ZN(
        P1_U2878) );
  OAI22_X1 U17698 ( .A1(n14559), .A2(n20035), .B1(n9648), .B2(n13335), .ZN(
        n14521) );
  AOI21_X1 U17699 ( .B1(n14561), .B2(BUF1_REG_25__SCAN_IN), .A(n14521), .ZN(
        n14523) );
  NAND2_X1 U17700 ( .A1(n14562), .A2(DATAI_25_), .ZN(n14522) );
  OAI211_X1 U17701 ( .C1(n14524), .C2(n14572), .A(n14523), .B(n14522), .ZN(
        P1_U2879) );
  OAI22_X1 U17702 ( .A1(n14559), .A2(n14526), .B1(n9648), .B2(n14525), .ZN(
        n14527) );
  AOI21_X1 U17703 ( .B1(n14561), .B2(BUF1_REG_24__SCAN_IN), .A(n14527), .ZN(
        n14529) );
  NAND2_X1 U17704 ( .A1(n14562), .A2(DATAI_24_), .ZN(n14528) );
  OAI211_X1 U17705 ( .C1(n15712), .C2(n14572), .A(n14529), .B(n14528), .ZN(
        P1_U2880) );
  OAI22_X1 U17706 ( .A1(n14559), .A2(n20152), .B1(n9648), .B2(n14530), .ZN(
        n14531) );
  AOI21_X1 U17707 ( .B1(n14561), .B2(BUF1_REG_23__SCAN_IN), .A(n14531), .ZN(
        n14533) );
  NAND2_X1 U17708 ( .A1(n14562), .A2(DATAI_23_), .ZN(n14532) );
  OAI211_X1 U17709 ( .C1(n15725), .C2(n14572), .A(n14533), .B(n14532), .ZN(
        P1_U2881) );
  OAI22_X1 U17710 ( .A1(n14559), .A2(n20144), .B1(n9648), .B2(n14534), .ZN(
        n14535) );
  AOI21_X1 U17711 ( .B1(n14561), .B2(BUF1_REG_22__SCAN_IN), .A(n14535), .ZN(
        n14537) );
  NAND2_X1 U17712 ( .A1(n14562), .A2(DATAI_22_), .ZN(n14536) );
  OAI211_X1 U17713 ( .C1(n15732), .C2(n14572), .A(n14537), .B(n14536), .ZN(
        P1_U2882) );
  OAI22_X1 U17714 ( .A1(n14559), .A2(n20140), .B1(n9648), .B2(n13330), .ZN(
        n14538) );
  AOI21_X1 U17715 ( .B1(n14561), .B2(BUF1_REG_21__SCAN_IN), .A(n14538), .ZN(
        n14540) );
  NAND2_X1 U17716 ( .A1(n14562), .A2(DATAI_21_), .ZN(n14539) );
  OAI211_X1 U17717 ( .C1(n14541), .C2(n14572), .A(n14540), .B(n14539), .ZN(
        P1_U2883) );
  OAI22_X1 U17718 ( .A1(n14559), .A2(n20136), .B1(n9648), .B2(n14542), .ZN(
        n14543) );
  AOI21_X1 U17719 ( .B1(n14561), .B2(BUF1_REG_20__SCAN_IN), .A(n14543), .ZN(
        n14545) );
  NAND2_X1 U17720 ( .A1(n14562), .A2(DATAI_20_), .ZN(n14544) );
  OAI211_X1 U17721 ( .C1(n15755), .C2(n14572), .A(n14545), .B(n14544), .ZN(
        P1_U2884) );
  OAI22_X1 U17722 ( .A1(n14559), .A2(n20132), .B1(n9648), .B2(n13328), .ZN(
        n14546) );
  AOI21_X1 U17723 ( .B1(n14561), .B2(BUF1_REG_19__SCAN_IN), .A(n14546), .ZN(
        n14548) );
  NAND2_X1 U17724 ( .A1(n14562), .A2(DATAI_19_), .ZN(n14547) );
  OAI211_X1 U17725 ( .C1(n14642), .C2(n14572), .A(n14548), .B(n14547), .ZN(
        P1_U2885) );
  OAI22_X1 U17726 ( .A1(n14559), .A2(n20128), .B1(n9648), .B2(n14549), .ZN(
        n14550) );
  AOI21_X1 U17727 ( .B1(n14561), .B2(BUF1_REG_18__SCAN_IN), .A(n14550), .ZN(
        n14552) );
  NAND2_X1 U17728 ( .A1(n14562), .A2(DATAI_18_), .ZN(n14551) );
  OAI211_X1 U17729 ( .C1(n15765), .C2(n14572), .A(n14552), .B(n14551), .ZN(
        P1_U2886) );
  OAI22_X1 U17730 ( .A1(n14559), .A2(n20125), .B1(n9648), .B2(n14553), .ZN(
        n14554) );
  AOI21_X1 U17731 ( .B1(n14561), .B2(BUF1_REG_17__SCAN_IN), .A(n14554), .ZN(
        n14556) );
  NAND2_X1 U17732 ( .A1(n14562), .A2(DATAI_17_), .ZN(n14555) );
  OAI211_X1 U17733 ( .C1(n14557), .C2(n14572), .A(n14556), .B(n14555), .ZN(
        P1_U2887) );
  OAI22_X1 U17734 ( .A1(n14559), .A2(n20117), .B1(n9648), .B2(n14558), .ZN(
        n14560) );
  AOI21_X1 U17735 ( .B1(n14561), .B2(BUF1_REG_16__SCAN_IN), .A(n14560), .ZN(
        n14564) );
  NAND2_X1 U17736 ( .A1(n14562), .A2(DATAI_16_), .ZN(n14563) );
  OAI211_X1 U17737 ( .C1(n14565), .C2(n14572), .A(n14564), .B(n14563), .ZN(
        P1_U2888) );
  OAI222_X1 U17738 ( .A1(n15789), .A2(n14572), .B1(n9648), .B2(n20011), .C1(
        n14571), .C2(n14566), .ZN(P1_U2889) );
  AOI22_X1 U17739 ( .A1(n14568), .A2(n20047), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14567), .ZN(n14569) );
  OAI21_X1 U17740 ( .B1(n14686), .B2(n14572), .A(n14569), .ZN(P1_U2891) );
  OAI222_X1 U17741 ( .A1(n14573), .A2(n14572), .B1(n20044), .B2(n14571), .C1(
        n14570), .C2(n9648), .ZN(P1_U2892) );
  NOR2_X1 U17742 ( .A1(n14587), .A2(n9784), .ZN(n14575) );
  AOI21_X1 U17743 ( .B1(n14607), .B2(n14575), .A(n14574), .ZN(n14576) );
  XOR2_X1 U17744 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14576), .Z(
        n14725) );
  NAND2_X1 U17745 ( .A1(n20074), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U17746 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14577) );
  OAI211_X1 U17747 ( .C1(n15899), .C2(n14578), .A(n14719), .B(n14577), .ZN(
        n14579) );
  AOI21_X1 U17748 ( .B1(n14580), .B2(n15894), .A(n14579), .ZN(n14581) );
  OAI21_X1 U17749 ( .B1(n14725), .B2(n19920), .A(n14581), .ZN(P1_U2969) );
  NOR2_X1 U17750 ( .A1(n16057), .A2(n14582), .ZN(n14727) );
  NOR2_X1 U17751 ( .A1(n15902), .A2(n14583), .ZN(n14584) );
  AOI211_X1 U17752 ( .C1(n15871), .C2(n14585), .A(n14727), .B(n14584), .ZN(
        n14591) );
  NAND2_X1 U17753 ( .A1(n14587), .A2(n14586), .ZN(n14588) );
  XNOR2_X1 U17754 ( .A(n14589), .B(n14588), .ZN(n14726) );
  NAND2_X1 U17755 ( .A1(n14726), .A2(n20070), .ZN(n14590) );
  OAI211_X1 U17756 ( .C1(n14592), .C2(n20104), .A(n14591), .B(n14590), .ZN(
        P1_U2970) );
  INV_X1 U17757 ( .A(n14700), .ZN(n15818) );
  NOR2_X1 U17758 ( .A1(n15858), .A2(n14594), .ZN(n15820) );
  NAND3_X1 U17759 ( .A1(n15858), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U17760 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_28__SCAN_IN), .ZN(n14601) );
  OAI21_X1 U17761 ( .B1(n15899), .B2(n14602), .A(n14601), .ZN(n14603) );
  AOI21_X1 U17762 ( .B1(n14604), .B2(n15894), .A(n14603), .ZN(n14605) );
  OAI21_X1 U17763 ( .B1(n15907), .B2(n19920), .A(n14605), .ZN(P1_U2971) );
  OAI21_X1 U17764 ( .B1(n14607), .B2(n12393), .A(n14606), .ZN(n14608) );
  XNOR2_X1 U17765 ( .A(n14608), .B(n15917), .ZN(n15912) );
  OAI22_X1 U17766 ( .A1(n15902), .A2(n14609), .B1(n16057), .B2(n15915), .ZN(
        n14612) );
  NOR2_X1 U17767 ( .A1(n14610), .A2(n20104), .ZN(n14611) );
  OAI21_X1 U17768 ( .B1(n19920), .B2(n15912), .A(n14614), .ZN(P1_U2972) );
  AOI21_X1 U17769 ( .B1(n14615), .B2(n12393), .A(n15950), .ZN(n15828) );
  MUX2_X1 U17770 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n9723), .S(
        n15874), .Z(n14616) );
  OAI21_X1 U17771 ( .B1(n15828), .B2(n15940), .A(n14616), .ZN(n14618) );
  XNOR2_X1 U17772 ( .A(n14618), .B(n14617), .ZN(n15929) );
  NAND2_X1 U17773 ( .A1(n14619), .A2(n15894), .ZN(n14624) );
  OAI22_X1 U17774 ( .A1(n15902), .A2(n14620), .B1(n16057), .B2(n15932), .ZN(
        n14621) );
  AOI21_X1 U17775 ( .B1(n15871), .B2(n14622), .A(n14621), .ZN(n14623) );
  OAI211_X1 U17776 ( .C1(n15929), .C2(n19920), .A(n14624), .B(n14623), .ZN(
        P1_U2974) );
  XNOR2_X1 U17777 ( .A(n12393), .B(n15950), .ZN(n14625) );
  XNOR2_X1 U17778 ( .A(n14593), .B(n14625), .ZN(n15952) );
  OAI22_X1 U17779 ( .A1(n15902), .A2(n15729), .B1(n16057), .B2(n15948), .ZN(
        n14627) );
  NOR2_X1 U17780 ( .A1(n15725), .A2(n20104), .ZN(n14626) );
  AOI211_X1 U17781 ( .C1(n15871), .C2(n15719), .A(n14627), .B(n14626), .ZN(
        n14628) );
  OAI21_X1 U17782 ( .B1(n15952), .B2(n19920), .A(n14628), .ZN(P1_U2976) );
  OAI22_X1 U17783 ( .A1(n14629), .A2(n19920), .B1(n15899), .B2(n15750), .ZN(
        n14630) );
  OAI21_X1 U17784 ( .B1(n15755), .B2(n20104), .A(n14632), .ZN(P1_U2979) );
  NAND2_X1 U17785 ( .A1(n14633), .A2(n14737), .ZN(n14635) );
  XOR2_X1 U17786 ( .A(n14635), .B(n14634), .Z(n15967) );
  NAND2_X1 U17787 ( .A1(n15967), .A2(n20070), .ZN(n14641) );
  INV_X1 U17788 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14636) );
  OAI22_X1 U17789 ( .A1(n15902), .A2(n14637), .B1(n16057), .B2(n14636), .ZN(
        n14638) );
  AOI21_X1 U17790 ( .B1(n15871), .B2(n14639), .A(n14638), .ZN(n14640) );
  OAI211_X1 U17791 ( .C1(n20104), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        P1_U2980) );
  OAI21_X1 U17792 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n15977) );
  INV_X1 U17793 ( .A(n15765), .ZN(n14648) );
  AOI22_X1 U17794 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14646) );
  OAI21_X1 U17795 ( .B1(n15899), .B2(n15764), .A(n14646), .ZN(n14647) );
  AOI21_X1 U17796 ( .B1(n14648), .B2(n15894), .A(n14647), .ZN(n14649) );
  OAI21_X1 U17797 ( .B1(n19920), .B2(n15977), .A(n14649), .ZN(P1_U2981) );
  NAND2_X1 U17798 ( .A1(n14650), .A2(n15847), .ZN(n14652) );
  NOR3_X1 U17799 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n12393), .ZN(n14651) );
  AOI21_X1 U17800 ( .B1(n15858), .B2(n14652), .A(n14651), .ZN(n14653) );
  XOR2_X1 U17801 ( .A(n14654), .B(n14653), .Z(n15987) );
  INV_X1 U17802 ( .A(n15987), .ZN(n14660) );
  AOI22_X1 U17803 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14655) );
  OAI21_X1 U17804 ( .B1(n15899), .B2(n14656), .A(n14655), .ZN(n14657) );
  AOI21_X1 U17805 ( .B1(n14658), .B2(n15894), .A(n14657), .ZN(n14659) );
  OAI21_X1 U17806 ( .B1(n14660), .B2(n19920), .A(n14659), .ZN(P1_U2982) );
  OR2_X1 U17807 ( .A1(n14661), .A2(n14662), .ZN(n15848) );
  INV_X1 U17808 ( .A(n15848), .ZN(n14664) );
  NOR2_X1 U17809 ( .A1(n14664), .A2(n14663), .ZN(n14667) );
  NOR2_X1 U17810 ( .A1(n14665), .A2(n15846), .ZN(n14666) );
  XNOR2_X1 U17811 ( .A(n14667), .B(n14666), .ZN(n16001) );
  NAND2_X1 U17812 ( .A1(n16001), .A2(n20070), .ZN(n14672) );
  INV_X1 U17813 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14668) );
  OAI22_X1 U17814 ( .A1(n15902), .A2(n14669), .B1(n16057), .B2(n14668), .ZN(
        n14670) );
  AOI21_X1 U17815 ( .B1(n15871), .B2(n15791), .A(n14670), .ZN(n14671) );
  OAI211_X1 U17816 ( .C1(n20104), .C2(n15789), .A(n14672), .B(n14671), .ZN(
        P1_U2984) );
  INV_X1 U17817 ( .A(n14673), .ZN(n14675) );
  OAI22_X1 U17818 ( .A1(n15902), .A2(n20886), .B1(n16057), .B2(n20676), .ZN(
        n14674) );
  AOI21_X1 U17819 ( .B1(n14675), .B2(n15871), .A(n14674), .ZN(n14685) );
  INV_X1 U17820 ( .A(n14661), .ZN(n14679) );
  INV_X1 U17821 ( .A(n14676), .ZN(n14677) );
  AOI21_X1 U17822 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n15867) );
  AND2_X1 U17823 ( .A1(n14680), .A2(n14681), .ZN(n15866) );
  NAND2_X1 U17824 ( .A1(n15867), .A2(n15866), .ZN(n15865) );
  NAND2_X1 U17825 ( .A1(n15865), .A2(n14681), .ZN(n14683) );
  XNOR2_X1 U17826 ( .A(n14683), .B(n14682), .ZN(n16014) );
  NAND2_X1 U17827 ( .A1(n16014), .A2(n20070), .ZN(n14684) );
  OAI211_X1 U17828 ( .C1(n14686), .C2(n20104), .A(n14685), .B(n14684), .ZN(
        P1_U2986) );
  NAND2_X1 U17829 ( .A1(n14689), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14688) );
  XNOR2_X1 U17830 ( .A(n14661), .B(n14690), .ZN(n14687) );
  MUX2_X1 U17831 ( .A(n14688), .B(n14687), .S(n15858), .Z(n14692) );
  INV_X1 U17832 ( .A(n14689), .ZN(n14691) );
  NAND3_X1 U17833 ( .A1(n14691), .A2(n15874), .A3(n14690), .ZN(n15876) );
  NAND2_X1 U17834 ( .A1(n14692), .A2(n15876), .ZN(n16041) );
  INV_X1 U17835 ( .A(n16041), .ZN(n14698) );
  AOI22_X1 U17836 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14693) );
  OAI21_X1 U17837 ( .B1(n15899), .B2(n14694), .A(n14693), .ZN(n14695) );
  AOI21_X1 U17838 ( .B1(n14696), .B2(n15894), .A(n14695), .ZN(n14697) );
  OAI21_X1 U17839 ( .B1(n14698), .B2(n19920), .A(n14697), .ZN(P1_U2989) );
  INV_X1 U17840 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14718) );
  OAI22_X1 U17841 ( .A1(n14700), .A2(n14699), .B1(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n20093), .ZN(n14705) );
  NAND2_X1 U17842 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15960) );
  AOI211_X1 U17843 ( .C1(n14703), .C2(n14702), .A(n14701), .B(n14713), .ZN(
        n14704) );
  OAI21_X1 U17844 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20093), .A(
        n15949), .ZN(n15939) );
  AOI211_X1 U17845 ( .C1(n14706), .C2(n15923), .A(n14705), .B(n15939), .ZN(
        n14707) );
  NAND2_X1 U17846 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14707), .ZN(
        n15924) );
  INV_X1 U17847 ( .A(n15924), .ZN(n14708) );
  OAI21_X1 U17848 ( .B1(n14729), .B2(n14710), .A(n14709), .ZN(n14734) );
  AOI211_X1 U17849 ( .C1(n14728), .C2(n16049), .A(n14718), .B(n14734), .ZN(
        n14716) );
  INV_X1 U17850 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14758) );
  NOR3_X1 U17851 ( .A1(n14716), .A2(n14710), .A3(n14758), .ZN(n14715) );
  NAND3_X1 U17852 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15961), .ZN(n15957) );
  NOR2_X1 U17853 ( .A1(n15818), .A2(n15957), .ZN(n15925) );
  NAND3_X1 U17854 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14729), .ZN(n14717) );
  NOR3_X1 U17855 ( .A1(n14717), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14718), .ZN(n14714) );
  INV_X1 U17856 ( .A(n14716), .ZN(n14723) );
  NAND2_X1 U17857 ( .A1(n14718), .A2(n14717), .ZN(n14722) );
  OAI21_X1 U17858 ( .B1(n14720), .B2(n16079), .A(n14719), .ZN(n14721) );
  AOI21_X1 U17859 ( .B1(n14723), .B2(n14722), .A(n14721), .ZN(n14724) );
  OAI21_X1 U17860 ( .B1(n14725), .B2(n16073), .A(n14724), .ZN(P1_U3001) );
  INV_X1 U17861 ( .A(n14726), .ZN(n14736) );
  INV_X1 U17862 ( .A(n14727), .ZN(n14731) );
  NAND3_X1 U17863 ( .A1(n15918), .A2(n14729), .A3(n14728), .ZN(n14730) );
  OAI211_X1 U17864 ( .C1(n14732), .C2(n16079), .A(n14731), .B(n14730), .ZN(
        n14733) );
  AOI21_X1 U17865 ( .B1(n14734), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14733), .ZN(n14735) );
  OAI21_X1 U17866 ( .B1(n14736), .B2(n16073), .A(n14735), .ZN(P1_U3002) );
  INV_X1 U17867 ( .A(n14737), .ZN(n14738) );
  NAND3_X1 U17868 ( .A1(n14065), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n14738), .ZN(n14739) );
  OAI21_X1 U17869 ( .B1(n14740), .B2(n12393), .A(n14739), .ZN(n14741) );
  XNOR2_X1 U17870 ( .A(n14741), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15845) );
  INV_X1 U17871 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14742) );
  OAI22_X1 U17872 ( .A1(n15741), .A2(n16079), .B1(n16057), .B2(n14742), .ZN(
        n14743) );
  NAND2_X1 U17873 ( .A1(n15961), .A2(n12399), .ZN(n14744) );
  OAI211_X1 U17874 ( .C1(n15845), .C2(n16073), .A(n14745), .B(n14744), .ZN(
        P1_U3010) );
  INV_X1 U17875 ( .A(n14746), .ZN(n14748) );
  NAND2_X1 U17876 ( .A1(n14748), .A2(n14747), .ZN(n15670) );
  AOI22_X1 U17877 ( .A1(n20109), .A2(n20718), .B1(n11689), .B2(n20712), .ZN(
        n14749) );
  NAND2_X1 U17878 ( .A1(n15670), .A2(n14749), .ZN(n14750) );
  MUX2_X1 U17879 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14750), .S(
        n20723), .Z(P1_U3478) );
  INV_X1 U17880 ( .A(n15671), .ZN(n14767) );
  NOR2_X1 U17881 ( .A1(n14752), .A2(n14751), .ZN(n14754) );
  INV_X1 U17882 ( .A(n14754), .ZN(n14760) );
  AOI21_X1 U17883 ( .B1(n14755), .B2(n14754), .A(n14753), .ZN(n14756) );
  OAI21_X1 U17884 ( .B1(n13545), .B2(n14757), .A(n14756), .ZN(n15647) );
  NOR2_X1 U17885 ( .A1(n20643), .A2(n20094), .ZN(n14764) );
  OAI22_X1 U17886 ( .A1(n14758), .A2(n12422), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14762) );
  AOI22_X1 U17887 ( .A1(n15647), .A2(n16083), .B1(n14764), .B2(n14762), .ZN(
        n14759) );
  OAI21_X1 U17888 ( .B1(n14767), .B2(n14760), .A(n14759), .ZN(n14761) );
  MUX2_X1 U17889 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14761), .S(
        n16087), .Z(P1_U3473) );
  INV_X1 U17890 ( .A(n14762), .ZN(n14763) );
  AOI22_X1 U17891 ( .A1(n15642), .A2(n16083), .B1(n14764), .B2(n14763), .ZN(
        n14765) );
  OAI21_X1 U17892 ( .B1(n14767), .B2(n14766), .A(n14765), .ZN(n14768) );
  MUX2_X1 U17893 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14768), .S(
        n16087), .Z(P1_U3472) );
  AOI211_X1 U17894 ( .C1(n14771), .C2(n14770), .A(n14769), .B(n19759), .ZN(
        n14772) );
  INV_X1 U17895 ( .A(n14772), .ZN(n14778) );
  AOI22_X1 U17896 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19038), .ZN(n14773) );
  OAI21_X1 U17897 ( .B1(n19065), .B2(n14861), .A(n14773), .ZN(n14776) );
  NOR2_X1 U17898 ( .A1(n14774), .A2(n19024), .ZN(n14775) );
  AOI211_X1 U17899 ( .C1(P2_EBX_REG_28__SCAN_IN), .C2(n19055), .A(n14776), .B(
        n14775), .ZN(n14777) );
  OAI211_X1 U17900 ( .C1(n14799), .C2(n18958), .A(n14778), .B(n14777), .ZN(
        P2_U2827) );
  OR2_X1 U17901 ( .A1(n14827), .A2(n14779), .ZN(n14780) );
  NAND2_X1 U17902 ( .A1(n9744), .A2(n14780), .ZN(n15152) );
  XNOR2_X1 U17903 ( .A(n14880), .B(n14899), .ZN(n15157) );
  AOI22_X1 U17904 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19038), .ZN(n14784) );
  INV_X1 U17905 ( .A(n14781), .ZN(n14782) );
  AOI22_X1 U17906 ( .A1(n14782), .A2(n19062), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19055), .ZN(n14783) );
  OAI211_X1 U17907 ( .C1(n15157), .C2(n19065), .A(n14784), .B(n14783), .ZN(
        n14788) );
  AOI211_X1 U17908 ( .C1(n14997), .C2(n14786), .A(n14785), .B(n19759), .ZN(
        n14787) );
  NOR2_X1 U17909 ( .A1(n14788), .A2(n14787), .ZN(n14789) );
  OAI21_X1 U17910 ( .B1(n18958), .B2(n15152), .A(n14789), .ZN(P2_U2831) );
  XNOR2_X1 U17911 ( .A(n14791), .B(n14790), .ZN(n14858) );
  NOR2_X1 U17912 ( .A1(n14792), .A2(n19078), .ZN(n14793) );
  AOI21_X1 U17913 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n19078), .A(n14793), .ZN(
        n14794) );
  OAI21_X1 U17914 ( .B1(n14858), .B2(n16181), .A(n14794), .ZN(P2_U2858) );
  NOR2_X1 U17915 ( .A1(n14796), .A2(n14795), .ZN(n14798) );
  XNOR2_X1 U17916 ( .A(n14798), .B(n14797), .ZN(n14864) );
  NOR2_X1 U17917 ( .A1(n14799), .A2(n19078), .ZN(n14800) );
  AOI21_X1 U17918 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19078), .A(n14800), .ZN(
        n14801) );
  OAI21_X1 U17919 ( .B1(n14864), .B2(n16181), .A(n14801), .ZN(P2_U2859) );
  XNOR2_X1 U17920 ( .A(n14803), .B(n14802), .ZN(n14871) );
  OR2_X1 U17921 ( .A1(n14810), .A2(n14804), .ZN(n14805) );
  NAND2_X1 U17922 ( .A1(n14806), .A2(n14805), .ZN(n16130) );
  NOR2_X1 U17923 ( .A1(n16130), .A2(n19078), .ZN(n14807) );
  AOI21_X1 U17924 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19078), .A(n14807), .ZN(
        n14808) );
  OAI21_X1 U17925 ( .B1(n14871), .B2(n16181), .A(n14808), .ZN(P2_U2860) );
  AND2_X1 U17926 ( .A1(n9696), .A2(n14809), .ZN(n14811) );
  OR2_X1 U17927 ( .A1(n14811), .A2(n14810), .ZN(n16138) );
  NAND2_X1 U17928 ( .A1(n14872), .A2(n19079), .ZN(n14814) );
  NAND2_X1 U17929 ( .A1(n19078), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14813) );
  OAI211_X1 U17930 ( .C1(n16138), .C2(n19078), .A(n14814), .B(n14813), .ZN(
        P2_U2861) );
  OAI21_X1 U17931 ( .B1(n14817), .B2(n14816), .A(n14815), .ZN(n14889) );
  NAND2_X1 U17932 ( .A1(n19078), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14821) );
  INV_X1 U17933 ( .A(n9696), .ZN(n14818) );
  AOI21_X1 U17934 ( .B1(n14819), .B2(n9744), .A(n14818), .ZN(n16151) );
  NAND2_X1 U17935 ( .A1(n16151), .A2(n14844), .ZN(n14820) );
  OAI211_X1 U17936 ( .C1(n14889), .C2(n16181), .A(n14821), .B(n14820), .ZN(
        P2_U2862) );
  OAI21_X1 U17937 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14907) );
  NOR2_X1 U17938 ( .A1(n14832), .A2(n14825), .ZN(n14826) );
  OR2_X1 U17939 ( .A1(n14827), .A2(n14826), .ZN(n16161) );
  NOR2_X1 U17940 ( .A1(n16161), .A2(n19078), .ZN(n14828) );
  AOI21_X1 U17941 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n19078), .A(n14828), .ZN(
        n14829) );
  OAI21_X1 U17942 ( .B1(n14907), .B2(n16181), .A(n14829), .ZN(P2_U2864) );
  AND2_X1 U17943 ( .A1(n14831), .A2(n14830), .ZN(n14833) );
  OR2_X1 U17944 ( .A1(n14833), .A2(n14832), .ZN(n15630) );
  AOI21_X1 U17945 ( .B1(n14836), .B2(n14919), .A(n14835), .ZN(n14917) );
  NAND2_X1 U17946 ( .A1(n14917), .A2(n19079), .ZN(n14838) );
  NAND2_X1 U17947 ( .A1(n19078), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14837) );
  OAI211_X1 U17948 ( .C1(n15630), .C2(n19078), .A(n14838), .B(n14837), .ZN(
        P2_U2865) );
  OAI21_X1 U17949 ( .B1(n14938), .B2(n14840), .A(n14839), .ZN(n14934) );
  NAND2_X1 U17950 ( .A1(n19078), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U17951 ( .A1(n15059), .A2(n14841), .ZN(n14842) );
  AND2_X1 U17952 ( .A1(n14843), .A2(n14842), .ZN(n18888) );
  NAND2_X1 U17953 ( .A1(n18888), .A2(n14844), .ZN(n14845) );
  OAI211_X1 U17954 ( .C1(n14934), .C2(n16181), .A(n14846), .B(n14845), .ZN(
        P2_U2867) );
  AND2_X1 U17955 ( .A1(n9753), .A2(n14847), .ZN(n14848) );
  OR2_X1 U17956 ( .A1(n15057), .A2(n14848), .ZN(n18922) );
  INV_X1 U17957 ( .A(n14936), .ZN(n14850) );
  AOI21_X1 U17958 ( .B1(n14851), .B2(n16185), .A(n14850), .ZN(n14956) );
  NAND2_X1 U17959 ( .A1(n14956), .A2(n19079), .ZN(n14853) );
  NAND2_X1 U17960 ( .A1(n19078), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14852) );
  OAI211_X1 U17961 ( .C1(n18922), .C2(n19078), .A(n14853), .B(n14852), .ZN(
        P2_U2869) );
  INV_X1 U17962 ( .A(n14854), .ZN(n16110) );
  INV_X1 U17963 ( .A(n16190), .ZN(n14921) );
  INV_X1 U17964 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19156) );
  OAI22_X1 U17965 ( .A1(n14921), .A2(n19093), .B1(n19111), .B2(n19156), .ZN(
        n14855) );
  AOI21_X1 U17966 ( .B1(n19138), .B2(n16110), .A(n14855), .ZN(n14857) );
  AOI22_X1 U17967 ( .A1(n19084), .A2(BUF2_REG_29__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U17968 ( .A1(n19084), .A2(BUF2_REG_28__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14860) );
  AOI22_X1 U17969 ( .A1(n16190), .A2(n19097), .B1(n19137), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n14859) );
  OAI211_X1 U17970 ( .C1(n14962), .C2(n14861), .A(n14860), .B(n14859), .ZN(
        n14862) );
  INV_X1 U17971 ( .A(n14862), .ZN(n14863) );
  OAI21_X1 U17972 ( .B1(n14864), .B2(n14947), .A(n14863), .ZN(P2_U2891) );
  AND2_X1 U17973 ( .A1(n9693), .A2(n14865), .ZN(n14866) );
  NOR2_X1 U17974 ( .A1(n14867), .A2(n14866), .ZN(n16133) );
  INV_X1 U17975 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19160) );
  OAI22_X1 U17976 ( .A1(n14921), .A2(n19100), .B1(n19111), .B2(n19160), .ZN(
        n14868) );
  AOI21_X1 U17977 ( .B1(n19138), .B2(n16133), .A(n14868), .ZN(n14870) );
  AOI22_X1 U17978 ( .A1(n19084), .A2(BUF2_REG_27__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14869) );
  OAI211_X1 U17979 ( .C1(n14871), .C2(n14947), .A(n14870), .B(n14869), .ZN(
        P2_U2892) );
  INV_X1 U17980 ( .A(n14872), .ZN(n14878) );
  NAND2_X1 U17981 ( .A1(n9706), .A2(n14873), .ZN(n14874) );
  AND2_X1 U17982 ( .A1(n9693), .A2(n14874), .ZN(n16136) );
  INV_X1 U17983 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19162) );
  OAI22_X1 U17984 ( .A1(n14921), .A2(n19102), .B1(n19111), .B2(n19162), .ZN(
        n14875) );
  AOI21_X1 U17985 ( .B1(n19138), .B2(n16136), .A(n14875), .ZN(n14877) );
  AOI22_X1 U17986 ( .A1(n19084), .A2(BUF2_REG_26__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14876) );
  OAI211_X1 U17987 ( .C1(n14878), .C2(n14947), .A(n14877), .B(n14876), .ZN(
        P2_U2893) );
  INV_X1 U17988 ( .A(n14879), .ZN(n14882) );
  NAND2_X1 U17989 ( .A1(n14880), .A2(n14899), .ZN(n14881) );
  NAND2_X1 U17990 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  NAND2_X1 U17991 ( .A1(n14883), .A2(n9706), .ZN(n16149) );
  AOI22_X1 U17992 ( .A1(n19084), .A2(BUF2_REG_25__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U17993 ( .A1(n16190), .A2(n14884), .B1(n19137), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n14885) );
  OAI211_X1 U17994 ( .C1(n14962), .C2(n16149), .A(n14886), .B(n14885), .ZN(
        n14887) );
  INV_X1 U17995 ( .A(n14887), .ZN(n14888) );
  OAI21_X1 U17996 ( .B1(n14889), .B2(n14947), .A(n14888), .ZN(P2_U2894) );
  AOI21_X1 U17997 ( .B1(n10378), .B2(n14892), .A(n14891), .ZN(n14893) );
  XNOR2_X1 U17998 ( .A(n14890), .B(n14893), .ZN(n16174) );
  INV_X1 U17999 ( .A(n16174), .ZN(n14898) );
  INV_X1 U18000 ( .A(n15157), .ZN(n14895) );
  INV_X1 U18001 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19166) );
  OAI22_X1 U18002 ( .A1(n14921), .A2(n19106), .B1(n19111), .B2(n19166), .ZN(
        n14894) );
  AOI21_X1 U18003 ( .B1(n19138), .B2(n14895), .A(n14894), .ZN(n14897) );
  AOI22_X1 U18004 ( .A1(n19084), .A2(BUF2_REG_24__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14896) );
  OAI211_X1 U18005 ( .C1(n14898), .C2(n14947), .A(n14897), .B(n14896), .ZN(
        P2_U2895) );
  INV_X1 U18006 ( .A(n14899), .ZN(n14900) );
  OAI21_X1 U18007 ( .B1(n14901), .B2(n14910), .A(n14900), .ZN(n16160) );
  AOI22_X1 U18008 ( .A1(n19084), .A2(BUF2_REG_23__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14904) );
  AOI22_X1 U18009 ( .A1(n16190), .A2(n14902), .B1(n19137), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n14903) );
  OAI211_X1 U18010 ( .C1(n14962), .C2(n16160), .A(n14904), .B(n14903), .ZN(
        n14905) );
  INV_X1 U18011 ( .A(n14905), .ZN(n14906) );
  OAI21_X1 U18012 ( .B1(n14907), .B2(n14947), .A(n14906), .ZN(P2_U2896) );
  NAND2_X1 U18013 ( .A1(n14909), .A2(n14908), .ZN(n14912) );
  INV_X1 U18014 ( .A(n14910), .ZN(n14911) );
  NAND2_X1 U18015 ( .A1(n14912), .A2(n14911), .ZN(n15629) );
  AOI22_X1 U18016 ( .A1(n19084), .A2(BUF2_REG_22__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14915) );
  AOI22_X1 U18017 ( .A1(n16190), .A2(n14913), .B1(n19137), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n14914) );
  OAI211_X1 U18018 ( .C1(n14962), .C2(n15629), .A(n14915), .B(n14914), .ZN(
        n14916) );
  AOI21_X1 U18019 ( .B1(n14917), .B2(n19139), .A(n14916), .ZN(n14918) );
  INV_X1 U18020 ( .A(n14918), .ZN(P2_U2897) );
  AOI21_X1 U18021 ( .B1(n14920), .B2(n14839), .A(n14834), .ZN(n16179) );
  INV_X1 U18022 ( .A(n16179), .ZN(n14925) );
  INV_X1 U18023 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19172) );
  OAI22_X1 U18024 ( .A1(n14921), .A2(n19250), .B1(n19111), .B2(n19172), .ZN(
        n14922) );
  AOI21_X1 U18025 ( .B1(n19138), .B2(n15189), .A(n14922), .ZN(n14924) );
  AOI22_X1 U18026 ( .A1(n19084), .A2(BUF2_REG_21__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14923) );
  OAI211_X1 U18027 ( .C1(n14925), .C2(n14947), .A(n14924), .B(n14923), .ZN(
        P2_U2898) );
  AND2_X1 U18028 ( .A1(n14941), .A2(n14926), .ZN(n14928) );
  OR2_X1 U18029 ( .A1(n14928), .A2(n14927), .ZN(n18886) );
  AOI22_X1 U18030 ( .A1(n19084), .A2(BUF2_REG_20__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U18031 ( .A1(n16190), .A2(n14929), .B1(n19137), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n14930) );
  OAI211_X1 U18032 ( .C1(n14962), .C2(n18886), .A(n14931), .B(n14930), .ZN(
        n14932) );
  INV_X1 U18033 ( .A(n14932), .ZN(n14933) );
  OAI21_X1 U18034 ( .B1(n14934), .B2(n14947), .A(n14933), .ZN(P2_U2899) );
  AND2_X1 U18035 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  OR2_X1 U18036 ( .A1(n14938), .A2(n14937), .ZN(n16182) );
  NAND2_X1 U18037 ( .A1(n14951), .A2(n14939), .ZN(n14940) );
  NAND2_X1 U18038 ( .A1(n14941), .A2(n14940), .ZN(n18914) );
  AOI22_X1 U18039 ( .A1(n19084), .A2(BUF2_REG_19__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U18040 ( .A1(n16190), .A2(n14942), .B1(n19137), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14943) );
  OAI211_X1 U18041 ( .C1(n14962), .C2(n18914), .A(n14944), .B(n14943), .ZN(
        n14945) );
  INV_X1 U18042 ( .A(n14945), .ZN(n14946) );
  OAI21_X1 U18043 ( .B1(n16182), .B2(n14947), .A(n14946), .ZN(P2_U2900) );
  NAND2_X1 U18044 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  AND2_X1 U18045 ( .A1(n14951), .A2(n14950), .ZN(n15229) );
  INV_X1 U18046 ( .A(n15229), .ZN(n18921) );
  AOI22_X1 U18047 ( .A1(n19084), .A2(BUF2_REG_18__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U18048 ( .A1(n16190), .A2(n14952), .B1(n19137), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n14953) );
  OAI211_X1 U18049 ( .C1(n14962), .C2(n18921), .A(n14954), .B(n14953), .ZN(
        n14955) );
  AOI21_X1 U18050 ( .B1(n14956), .B2(n19139), .A(n14955), .ZN(n14957) );
  INV_X1 U18051 ( .A(n14957), .ZN(P2_U2901) );
  INV_X1 U18052 ( .A(n15622), .ZN(n14961) );
  AOI22_X1 U18053 ( .A1(n19084), .A2(BUF2_REG_16__SCAN_IN), .B1(n19085), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U18054 ( .A1(n16190), .A2(n14958), .B1(n19137), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14959) );
  OAI211_X1 U18055 ( .C1(n14962), .C2(n14961), .A(n14960), .B(n14959), .ZN(
        n14963) );
  AOI21_X1 U18056 ( .B1(n14964), .B2(n19139), .A(n14963), .ZN(n14965) );
  INV_X1 U18057 ( .A(n14965), .ZN(P2_U2903) );
  INV_X1 U18058 ( .A(n14966), .ZN(n14967) );
  OAI21_X1 U18059 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n9698), .A(
        n14967), .ZN(n15130) );
  NAND3_X1 U18060 ( .A1(n15121), .A2(n15120), .A3(n19222), .ZN(n14972) );
  NAND2_X1 U18061 ( .A1(n19044), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15122) );
  OAI21_X1 U18062 ( .B1(n19229), .B2(n16123), .A(n15122), .ZN(n14970) );
  NOR2_X1 U18063 ( .A1(n16130), .A2(n16206), .ZN(n14969) );
  AOI211_X1 U18064 ( .C1(n19220), .C2(n16122), .A(n14970), .B(n14969), .ZN(
        n14971) );
  OAI211_X1 U18065 ( .C1(n19234), .C2(n15130), .A(n14972), .B(n14971), .ZN(
        P2_U2987) );
  INV_X1 U18066 ( .A(n14973), .ZN(n14983) );
  NOR2_X1 U18067 ( .A1(n14974), .A2(n14983), .ZN(n14975) );
  XOR2_X1 U18068 ( .A(n14976), .B(n14975), .Z(n15140) );
  AOI21_X1 U18069 ( .B1(n15132), .B2(n14977), .A(n9698), .ZN(n15138) );
  INV_X1 U18070 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19826) );
  NOR2_X1 U18071 ( .A1(n19023), .A2(n19826), .ZN(n15134) );
  NOR2_X1 U18072 ( .A1(n16256), .A2(n14978), .ZN(n14979) );
  AOI211_X1 U18073 ( .C1(n19230), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15134), .B(n14979), .ZN(n14980) );
  OAI21_X1 U18074 ( .B1(n16138), .B2(n16206), .A(n14980), .ZN(n14981) );
  AOI21_X1 U18075 ( .B1(n15138), .B2(n19224), .A(n14981), .ZN(n14982) );
  OAI21_X1 U18076 ( .B1(n15140), .B2(n19236), .A(n14982), .ZN(P2_U2988) );
  NOR2_X1 U18077 ( .A1(n14984), .A2(n14983), .ZN(n14986) );
  XOR2_X1 U18078 ( .A(n14986), .B(n14985), .Z(n15151) );
  NAND2_X1 U18079 ( .A1(n19220), .A2(n16154), .ZN(n14987) );
  NAND2_X1 U18080 ( .A1(n19044), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15141) );
  OAI211_X1 U18081 ( .C1(n19229), .C2(n14988), .A(n14987), .B(n15141), .ZN(
        n14989) );
  AOI21_X1 U18082 ( .B1(n16151), .B2(n19239), .A(n14989), .ZN(n14993) );
  INV_X1 U18083 ( .A(n14977), .ZN(n14991) );
  AOI21_X1 U18084 ( .B1(n15146), .B2(n14990), .A(n14991), .ZN(n15149) );
  NAND2_X1 U18085 ( .A1(n15149), .A2(n19224), .ZN(n14992) );
  OAI211_X1 U18086 ( .C1(n15151), .C2(n19236), .A(n14993), .B(n14992), .ZN(
        P2_U2989) );
  XNOR2_X1 U18087 ( .A(n14995), .B(n15154), .ZN(n14996) );
  XNOR2_X1 U18088 ( .A(n14994), .B(n14996), .ZN(n15161) );
  INV_X1 U18089 ( .A(n15161), .ZN(n15001) );
  INV_X1 U18090 ( .A(n15152), .ZN(n16173) );
  NAND2_X1 U18091 ( .A1(n19220), .A2(n14997), .ZN(n14998) );
  NAND2_X1 U18092 ( .A1(n19044), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15156) );
  OAI211_X1 U18093 ( .C1(n19229), .C2(n10152), .A(n14998), .B(n15156), .ZN(
        n15000) );
  XNOR2_X1 U18094 ( .A(n15003), .B(n15002), .ZN(n15176) );
  AOI21_X1 U18095 ( .B1(n15172), .B2(n9678), .A(n9641), .ZN(n15174) );
  OAI22_X1 U18096 ( .A1(n19229), .A2(n15004), .B1(n19820), .B2(n19023), .ZN(
        n15005) );
  AOI21_X1 U18097 ( .B1(n19220), .B2(n16165), .A(n15005), .ZN(n15006) );
  OAI21_X1 U18098 ( .B1(n16161), .B2(n16206), .A(n15006), .ZN(n15007) );
  AOI21_X1 U18099 ( .B1(n15174), .B2(n19224), .A(n15007), .ZN(n15008) );
  OAI21_X1 U18100 ( .B1(n19236), .B2(n15176), .A(n15008), .ZN(P2_U2991) );
  OAI21_X1 U18101 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n9970), .A(
        n9678), .ZN(n15185) );
  OAI21_X1 U18102 ( .B1(n15012), .B2(n15011), .A(n15010), .ZN(n15183) );
  INV_X1 U18103 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19818) );
  OAI22_X1 U18104 ( .A1(n19818), .A2(n19023), .B1(n16256), .B2(n15013), .ZN(
        n15015) );
  OAI22_X1 U18105 ( .A1(n15630), .A2(n16206), .B1(n10153), .B2(n19229), .ZN(
        n15014) );
  AOI211_X1 U18106 ( .C1(n15183), .C2(n19222), .A(n15015), .B(n15014), .ZN(
        n15016) );
  OAI21_X1 U18107 ( .B1(n15185), .B2(n19234), .A(n15016), .ZN(P2_U2992) );
  AND2_X1 U18108 ( .A1(n15019), .A2(n15018), .ZN(n15252) );
  NAND2_X1 U18109 ( .A1(n15017), .A2(n15252), .ZN(n15251) );
  INV_X1 U18110 ( .A(n15075), .ZN(n15024) );
  INV_X1 U18111 ( .A(n15022), .ZN(n15023) );
  AOI21_X2 U18112 ( .B1(n15024), .B2(n15076), .A(n15023), .ZN(n15067) );
  INV_X1 U18113 ( .A(n15026), .ZN(n15040) );
  NAND2_X1 U18114 ( .A1(n15029), .A2(n15028), .ZN(n15030) );
  NAND2_X1 U18115 ( .A1(n19044), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15191) );
  OAI21_X1 U18116 ( .B1(n19229), .B2(n15031), .A(n15191), .ZN(n15033) );
  NOR2_X1 U18117 ( .A1(n16177), .A2(n16206), .ZN(n15032) );
  AOI211_X1 U18118 ( .C1(n19220), .C2(n15034), .A(n15033), .B(n15032), .ZN(
        n15037) );
  NAND2_X1 U18119 ( .A1(n15036), .A2(n15196), .ZN(n15186) );
  NOR2_X1 U18120 ( .A1(n9705), .A2(n15038), .ZN(n15042) );
  NOR2_X1 U18121 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  XNOR2_X1 U18122 ( .A(n15042), .B(n15041), .ZN(n15214) );
  NOR2_X1 U18123 ( .A1(n19023), .A2(n15043), .ZN(n15207) );
  AOI21_X1 U18124 ( .B1(n19230), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15207), .ZN(n15044) );
  OAI21_X1 U18125 ( .B1(n16256), .B2(n15045), .A(n15044), .ZN(n15048) );
  OAI21_X1 U18126 ( .B1(n15046), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15036), .ZN(n15201) );
  NOR2_X1 U18127 ( .A1(n15201), .A2(n19234), .ZN(n15047) );
  AOI211_X1 U18128 ( .C1(n19239), .C2(n18888), .A(n15048), .B(n15047), .ZN(
        n15049) );
  OAI21_X1 U18129 ( .B1(n15214), .B2(n19236), .A(n15049), .ZN(P2_U2994) );
  NAND2_X1 U18130 ( .A1(n15051), .A2(n15050), .ZN(n15054) );
  INV_X1 U18131 ( .A(n15064), .ZN(n15052) );
  OAI21_X1 U18132 ( .B1(n15067), .B2(n15052), .A(n15065), .ZN(n15053) );
  XOR2_X1 U18133 ( .A(n15054), .B(n15053), .Z(n15225) );
  AOI21_X1 U18134 ( .B1(n15220), .B2(n15055), .A(n15046), .ZN(n15223) );
  OR2_X1 U18135 ( .A1(n15057), .A2(n15056), .ZN(n15058) );
  NAND2_X1 U18136 ( .A1(n15059), .A2(n15058), .ZN(n18911) );
  NAND2_X1 U18137 ( .A1(n18904), .A2(n19220), .ZN(n15061) );
  NOR2_X1 U18138 ( .A1(n19023), .A2(n19813), .ZN(n15216) );
  AOI21_X1 U18139 ( .B1(n19230), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15216), .ZN(n15060) );
  OAI211_X1 U18140 ( .C1(n16206), .C2(n18911), .A(n15061), .B(n15060), .ZN(
        n15062) );
  AOI21_X1 U18141 ( .B1(n15223), .B2(n19224), .A(n15062), .ZN(n15063) );
  OAI21_X1 U18142 ( .B1(n15225), .B2(n19236), .A(n15063), .ZN(P2_U2995) );
  NAND2_X1 U18143 ( .A1(n15065), .A2(n15064), .ZN(n15066) );
  XNOR2_X1 U18144 ( .A(n15067), .B(n15066), .ZN(n15236) );
  INV_X1 U18145 ( .A(n15055), .ZN(n15069) );
  AOI21_X1 U18146 ( .B1(n15203), .B2(n15068), .A(n15069), .ZN(n15234) );
  NOR2_X1 U18147 ( .A1(n19023), .A2(n15070), .ZN(n15228) );
  NOR2_X1 U18148 ( .A1(n18922), .A2(n16206), .ZN(n15071) );
  AOI211_X1 U18149 ( .C1(n19230), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15228), .B(n15071), .ZN(n15072) );
  OAI21_X1 U18150 ( .B1(n16256), .B2(n18915), .A(n15072), .ZN(n15073) );
  AOI21_X1 U18151 ( .B1(n15234), .B2(n19224), .A(n15073), .ZN(n15074) );
  OAI21_X1 U18152 ( .B1(n15236), .B2(n19236), .A(n15074), .ZN(P2_U2996) );
  XOR2_X1 U18153 ( .A(n15076), .B(n15075), .Z(n15250) );
  INV_X1 U18154 ( .A(n9753), .ZN(n15077) );
  AOI21_X1 U18155 ( .B1(n15078), .B2(n9740), .A(n15077), .ZN(n18930) );
  NOR2_X1 U18156 ( .A1(n19810), .A2(n19023), .ZN(n15081) );
  INV_X1 U18157 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15079) );
  OAI22_X1 U18158 ( .A1(n19229), .A2(n15079), .B1(n16256), .B2(n18932), .ZN(
        n15080) );
  AOI211_X1 U18159 ( .C1(n18930), .C2(n19239), .A(n15081), .B(n15080), .ZN(
        n15084) );
  INV_X1 U18160 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16277) );
  OAI211_X1 U18161 ( .C1(n15237), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19224), .B(n15068), .ZN(n15083) );
  OAI211_X1 U18162 ( .C1(n15250), .C2(n19236), .A(n15084), .B(n15083), .ZN(
        P2_U2997) );
  NAND2_X1 U18163 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  XNOR2_X1 U18164 ( .A(n15088), .B(n15087), .ZN(n16282) );
  AOI21_X1 U18165 ( .B1(n16277), .B2(n16209), .A(n16203), .ZN(n16279) );
  INV_X1 U18166 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15089) );
  OAI22_X1 U18167 ( .A1(n19229), .A2(n15089), .B1(n16256), .B2(n18952), .ZN(
        n15093) );
  OAI22_X1 U18168 ( .A1(n16206), .A2(n15091), .B1(n19023), .B2(n15090), .ZN(
        n15092) );
  AOI211_X1 U18169 ( .C1(n16279), .C2(n19224), .A(n15093), .B(n15092), .ZN(
        n15094) );
  OAI21_X1 U18170 ( .B1(n16282), .B2(n19236), .A(n15094), .ZN(P2_U2999) );
  NAND2_X1 U18171 ( .A1(n16246), .A2(n15095), .ZN(n15097) );
  XOR2_X1 U18172 ( .A(n15097), .B(n15096), .Z(n15298) );
  NAND2_X1 U18173 ( .A1(n15098), .A2(n15292), .ZN(n15285) );
  NAND3_X1 U18174 ( .A1(n15285), .A2(n19224), .A3(n16251), .ZN(n15101) );
  AND2_X1 U18175 ( .A1(n19044), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n15289) );
  INV_X1 U18176 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19004) );
  OAI22_X1 U18177 ( .A1(n19229), .A2(n19004), .B1(n16256), .B2(n19007), .ZN(
        n15099) );
  AOI211_X1 U18178 ( .C1(n19239), .C2(n19009), .A(n15289), .B(n15099), .ZN(
        n15100) );
  OAI211_X1 U18179 ( .C1(n19236), .C2(n15298), .A(n15101), .B(n15100), .ZN(
        P2_U3005) );
  XNOR2_X1 U18180 ( .A(n15102), .B(n15103), .ZN(n15310) );
  NAND2_X1 U18181 ( .A1(n16260), .A2(n16262), .ZN(n15105) );
  XNOR2_X1 U18182 ( .A(n15104), .B(n15105), .ZN(n15308) );
  INV_X1 U18183 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15106) );
  OAI22_X1 U18184 ( .A1(n19229), .A2(n15106), .B1(n16256), .B2(n19017), .ZN(
        n15109) );
  INV_X1 U18185 ( .A(n19019), .ZN(n15107) );
  OAI22_X1 U18186 ( .A1(n16206), .A2(n15107), .B1(n19023), .B2(n19794), .ZN(
        n15108) );
  AOI211_X1 U18187 ( .C1(n15308), .C2(n19222), .A(n15109), .B(n15108), .ZN(
        n15110) );
  OAI21_X1 U18188 ( .B1(n15310), .B2(n19234), .A(n15110), .ZN(P2_U3007) );
  CLKBUF_X1 U18189 ( .A(n15112), .Z(n15113) );
  XNOR2_X1 U18190 ( .A(n15111), .B(n15113), .ZN(n15322) );
  XNOR2_X1 U18191 ( .A(n15114), .B(n15313), .ZN(n15320) );
  OAI22_X1 U18192 ( .A1(n19229), .A2(n15115), .B1(n19792), .B2(n19023), .ZN(
        n15116) );
  AOI21_X1 U18193 ( .B1(n19220), .B2(n19031), .A(n15116), .ZN(n15117) );
  OAI21_X1 U18194 ( .B1(n19032), .B2(n16206), .A(n15117), .ZN(n15118) );
  AOI21_X1 U18195 ( .B1(n15320), .B2(n19224), .A(n15118), .ZN(n15119) );
  OAI21_X1 U18196 ( .B1(n19236), .B2(n15322), .A(n15119), .ZN(P2_U3008) );
  NAND3_X1 U18197 ( .A1(n15121), .A2(n15120), .A3(n16334), .ZN(n15129) );
  NOR2_X1 U18198 ( .A1(n16130), .A2(n16329), .ZN(n15126) );
  INV_X1 U18199 ( .A(n16133), .ZN(n15124) );
  OAI211_X1 U18200 ( .C1(n16324), .C2(n15124), .A(n15123), .B(n15122), .ZN(
        n15125) );
  AOI211_X1 U18201 ( .C1(n15127), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15126), .B(n15125), .ZN(n15128) );
  OAI211_X1 U18202 ( .C1(n15130), .C2(n16330), .A(n15129), .B(n15128), .ZN(
        P2_U3019) );
  NOR2_X1 U18203 ( .A1(n15147), .A2(n15132), .ZN(n15137) );
  NAND2_X1 U18204 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15153), .ZN(
        n15142) );
  AOI211_X1 U18205 ( .C1(n15132), .C2(n15146), .A(n15131), .B(n15142), .ZN(
        n15133) );
  AOI211_X1 U18206 ( .C1(n16301), .C2(n16136), .A(n15134), .B(n15133), .ZN(
        n15135) );
  OAI21_X1 U18207 ( .B1(n16138), .B2(n16329), .A(n15135), .ZN(n15136) );
  AOI211_X1 U18208 ( .C1(n15138), .C2(n16313), .A(n15137), .B(n15136), .ZN(
        n15139) );
  OAI21_X1 U18209 ( .B1(n15140), .B2(n16317), .A(n15139), .ZN(P2_U3020) );
  NOR2_X1 U18210 ( .A1(n16324), .A2(n16149), .ZN(n15144) );
  OAI21_X1 U18211 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15142), .A(
        n15141), .ZN(n15143) );
  AOI211_X1 U18212 ( .C1(n16151), .C2(n16312), .A(n15144), .B(n15143), .ZN(
        n15145) );
  OAI21_X1 U18213 ( .B1(n15147), .B2(n15146), .A(n15145), .ZN(n15148) );
  AOI21_X1 U18214 ( .B1(n15149), .B2(n16313), .A(n15148), .ZN(n15150) );
  OAI21_X1 U18215 ( .B1(n15151), .B2(n16317), .A(n15150), .ZN(P2_U3021) );
  NOR2_X1 U18216 ( .A1(n15152), .A2(n16329), .ZN(n15159) );
  NAND2_X1 U18217 ( .A1(n15154), .A2(n15153), .ZN(n15155) );
  OAI211_X1 U18218 ( .C1(n16324), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        n15158) );
  AOI211_X1 U18219 ( .C1(n15160), .C2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15159), .B(n15158), .ZN(n15163) );
  NAND2_X1 U18220 ( .A1(n15161), .A2(n16334), .ZN(n15162) );
  OAI211_X1 U18221 ( .C1(n15164), .C2(n16330), .A(n15163), .B(n15162), .ZN(
        P2_U3022) );
  INV_X1 U18222 ( .A(n16161), .ZN(n15170) );
  AOI21_X1 U18223 ( .B1(n15172), .B2(n15179), .A(n15165), .ZN(n15167) );
  NOR2_X1 U18224 ( .A1(n19820), .A2(n19023), .ZN(n15166) );
  AOI21_X1 U18225 ( .B1(n15177), .B2(n15167), .A(n15166), .ZN(n15168) );
  OAI21_X1 U18226 ( .B1(n16324), .B2(n16160), .A(n15168), .ZN(n15169) );
  AOI21_X1 U18227 ( .B1(n15170), .B2(n16312), .A(n15169), .ZN(n15171) );
  OAI21_X1 U18228 ( .B1(n15197), .B2(n15172), .A(n15171), .ZN(n15173) );
  AOI21_X1 U18229 ( .B1(n15174), .B2(n16313), .A(n15173), .ZN(n15175) );
  OAI21_X1 U18230 ( .B1(n16317), .B2(n15176), .A(n15175), .ZN(P2_U3023) );
  INV_X1 U18231 ( .A(n15177), .ZN(n15180) );
  NAND2_X1 U18232 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19044), .ZN(n15178) );
  OAI221_X1 U18233 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15180), 
        .C1(n15179), .C2(n15197), .A(n15178), .ZN(n15182) );
  OAI22_X1 U18234 ( .A1(n15630), .A2(n16329), .B1(n16324), .B2(n15629), .ZN(
        n15181) );
  AOI211_X1 U18235 ( .C1(n15183), .C2(n16334), .A(n15182), .B(n15181), .ZN(
        n15184) );
  OAI21_X1 U18236 ( .B1(n15185), .B2(n16330), .A(n15184), .ZN(P2_U3024) );
  NAND3_X1 U18237 ( .A1(n15187), .A2(n16313), .A3(n15186), .ZN(n15195) );
  AND2_X1 U18238 ( .A1(n15188), .A2(n15196), .ZN(n15193) );
  NAND2_X1 U18239 ( .A1(n16301), .A2(n15189), .ZN(n15190) );
  OAI211_X1 U18240 ( .C1(n16177), .C2(n16329), .A(n15191), .B(n15190), .ZN(
        n15192) );
  AOI21_X1 U18241 ( .B1(n15273), .B2(n15193), .A(n15192), .ZN(n15194) );
  OAI211_X1 U18242 ( .C1(n15197), .C2(n15196), .A(n15195), .B(n15194), .ZN(
        n15198) );
  INV_X1 U18243 ( .A(n15198), .ZN(n15199) );
  OAI21_X1 U18244 ( .B1(n15200), .B2(n16317), .A(n15199), .ZN(P2_U3025) );
  INV_X1 U18245 ( .A(n15201), .ZN(n15212) );
  OAI21_X1 U18246 ( .B1(n15202), .B2(n15241), .A(n15293), .ZN(n15226) );
  AOI21_X1 U18247 ( .B1(n15203), .B2(n15264), .A(n15226), .ZN(n15221) );
  INV_X1 U18248 ( .A(n15232), .ZN(n15206) );
  NAND3_X1 U18249 ( .A1(n15206), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15220), .ZN(n15218) );
  AOI21_X1 U18250 ( .B1(n15221), .B2(n15218), .A(n15204), .ZN(n15211) );
  NAND3_X1 U18251 ( .A1(n15206), .A2(n15205), .A3(n15204), .ZN(n15209) );
  AOI21_X1 U18252 ( .B1(n18888), .B2(n16312), .A(n15207), .ZN(n15208) );
  OAI211_X1 U18253 ( .C1(n16324), .C2(n18886), .A(n15209), .B(n15208), .ZN(
        n15210) );
  AOI211_X1 U18254 ( .C1(n15212), .C2(n16313), .A(n15211), .B(n15210), .ZN(
        n15213) );
  OAI21_X1 U18255 ( .B1(n15214), .B2(n16317), .A(n15213), .ZN(P2_U3026) );
  INV_X1 U18256 ( .A(n18911), .ZN(n15217) );
  NOR2_X1 U18257 ( .A1(n16324), .A2(n18914), .ZN(n15215) );
  AOI211_X1 U18258 ( .C1(n15217), .C2(n16312), .A(n15216), .B(n15215), .ZN(
        n15219) );
  OAI211_X1 U18259 ( .C1(n15221), .C2(n15220), .A(n15219), .B(n15218), .ZN(
        n15222) );
  AOI21_X1 U18260 ( .B1(n15223), .B2(n16313), .A(n15222), .ZN(n15224) );
  OAI21_X1 U18261 ( .B1(n15225), .B2(n16317), .A(n15224), .ZN(P2_U3027) );
  NAND2_X1 U18262 ( .A1(n15226), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15231) );
  NOR2_X1 U18263 ( .A1(n16329), .A2(n18922), .ZN(n15227) );
  AOI211_X1 U18264 ( .C1(n16301), .C2(n15229), .A(n15228), .B(n15227), .ZN(
        n15230) );
  OAI211_X1 U18265 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15232), .A(
        n15231), .B(n15230), .ZN(n15233) );
  AOI21_X1 U18266 ( .B1(n15234), .B2(n16313), .A(n15233), .ZN(n15235) );
  OAI21_X1 U18267 ( .B1(n15236), .B2(n16317), .A(n15235), .ZN(P2_U3028) );
  OAI21_X1 U18268 ( .B1(n15239), .B2(n15241), .A(n15293), .ZN(n16276) );
  OAI211_X1 U18269 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15241), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15626), .ZN(n15248) );
  NAND2_X1 U18270 ( .A1(n15242), .A2(n15273), .ZN(n16299) );
  NOR2_X1 U18271 ( .A1(n15243), .A2(n16299), .ZN(n16278) );
  AOI22_X1 U18272 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16278), .B1(
        n16313), .B2(n16203), .ZN(n15628) );
  INV_X1 U18273 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15627) );
  OAI21_X1 U18274 ( .B1(n15628), .B2(n15627), .A(n10841), .ZN(n15247) );
  XNOR2_X1 U18275 ( .A(n15244), .B(n9738), .ZN(n16191) );
  AOI22_X1 U18276 ( .A1(n16312), .A2(n18930), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n19044), .ZN(n15245) );
  OAI21_X1 U18277 ( .B1(n16191), .B2(n16324), .A(n15245), .ZN(n15246) );
  AOI21_X1 U18278 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(n15249) );
  OAI21_X1 U18279 ( .B1(n15250), .B2(n16317), .A(n15249), .ZN(P2_U3029) );
  OAI21_X1 U18280 ( .B1(n15017), .B2(n15252), .A(n15251), .ZN(n16222) );
  INV_X1 U18281 ( .A(n16222), .ZN(n15268) );
  NOR2_X1 U18282 ( .A1(n10813), .A2(n16299), .ZN(n15262) );
  OR2_X1 U18283 ( .A1(n15253), .A2(n16294), .ZN(n15255) );
  NAND2_X1 U18284 ( .A1(n15255), .A2(n15254), .ZN(n19094) );
  AND2_X1 U18285 ( .A1(n15257), .A2(n15256), .ZN(n15259) );
  OR2_X1 U18286 ( .A1(n15259), .A2(n15258), .ZN(n19082) );
  INV_X1 U18287 ( .A(n19082), .ZN(n16221) );
  NAND2_X1 U18288 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16228), .ZN(
        n16229) );
  NAND2_X1 U18289 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16284) );
  INV_X1 U18290 ( .A(n16284), .ZN(n15260) );
  AND2_X1 U18291 ( .A1(n16228), .A2(n15260), .ZN(n16208) );
  AOI21_X1 U18292 ( .B1(n15261), .B2(n16229), .A(n16208), .ZN(n16223) );
  NAND2_X1 U18293 ( .A1(n19044), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16224) );
  AOI21_X1 U18294 ( .B1(n15265), .B2(n15264), .A(n15263), .ZN(n16298) );
  OAI21_X1 U18295 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16299), .A(
        n16298), .ZN(n15266) );
  NAND2_X1 U18296 ( .A1(n15266), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15267) );
  INV_X1 U18297 ( .A(n16228), .ZN(n15269) );
  XNOR2_X1 U18298 ( .A(n15271), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15272) );
  XNOR2_X1 U18299 ( .A(n15270), .B(n15272), .ZN(n16240) );
  NAND2_X1 U18300 ( .A1(n15273), .A2(n15292), .ZN(n15291) );
  NAND2_X1 U18301 ( .A1(n15293), .A2(n15291), .ZN(n16311) );
  NOR2_X1 U18302 ( .A1(n11310), .A2(n19023), .ZN(n15276) );
  NAND2_X1 U18303 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15273), .ZN(
        n16308) );
  AOI221_X1 U18304 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n16252), .C2(n15274), .A(
        n16308), .ZN(n15275) );
  AOI211_X1 U18305 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16311), .A(
        n15276), .B(n15275), .ZN(n15282) );
  OR2_X1 U18306 ( .A1(n15278), .A2(n15277), .ZN(n15279) );
  NAND2_X1 U18307 ( .A1(n15279), .A2(n16295), .ZN(n19101) );
  INV_X1 U18308 ( .A(n19101), .ZN(n15280) );
  AOI22_X1 U18309 ( .A1(n16301), .A2(n15280), .B1(n16312), .B2(n18985), .ZN(
        n15281) );
  OAI211_X1 U18310 ( .C1(n16240), .C2(n16317), .A(n15282), .B(n15281), .ZN(
        n15283) );
  INV_X1 U18311 ( .A(n15283), .ZN(n15284) );
  OAI21_X1 U18312 ( .B1(n16241), .B2(n16330), .A(n15284), .ZN(P2_U3035) );
  NAND3_X1 U18313 ( .A1(n15285), .A2(n16313), .A3(n16251), .ZN(n15297) );
  OR2_X1 U18314 ( .A1(n15287), .A2(n15286), .ZN(n15288) );
  NAND2_X1 U18315 ( .A1(n15288), .A2(n16306), .ZN(n19105) );
  INV_X1 U18316 ( .A(n15289), .ZN(n15290) );
  OAI211_X1 U18317 ( .C1(n16324), .C2(n19105), .A(n15291), .B(n15290), .ZN(
        n15295) );
  NOR2_X1 U18318 ( .A1(n15293), .A2(n15292), .ZN(n15294) );
  AOI211_X1 U18319 ( .C1(n19009), .C2(n16312), .A(n15295), .B(n15294), .ZN(
        n15296) );
  OAI211_X1 U18320 ( .C1(n15298), .C2(n16317), .A(n15297), .B(n15296), .ZN(
        P2_U3037) );
  NAND2_X1 U18321 ( .A1(n15312), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15306) );
  NOR2_X1 U18322 ( .A1(n19794), .A2(n19023), .ZN(n15304) );
  OR2_X1 U18323 ( .A1(n15300), .A2(n15299), .ZN(n15302) );
  NAND2_X1 U18324 ( .A1(n15302), .A2(n15301), .ZN(n19109) );
  NOR2_X1 U18325 ( .A1(n16324), .A2(n19109), .ZN(n15303) );
  AOI211_X1 U18326 ( .C1(n19019), .C2(n16312), .A(n15304), .B(n15303), .ZN(
        n15305) );
  OAI211_X1 U18327 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16320), .A(
        n15306), .B(n15305), .ZN(n15307) );
  AOI21_X1 U18328 ( .B1(n15308), .B2(n16334), .A(n15307), .ZN(n15309) );
  OAI21_X1 U18329 ( .B1(n15310), .B2(n16330), .A(n15309), .ZN(P2_U3039) );
  NOR2_X1 U18330 ( .A1(n19792), .A2(n19023), .ZN(n15311) );
  AOI221_X1 U18331 ( .B1(n15314), .B2(n15313), .C1(n15312), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n15311), .ZN(n15315) );
  INV_X1 U18332 ( .A(n15315), .ZN(n15319) );
  XNOR2_X1 U18333 ( .A(n15317), .B(n15316), .ZN(n19110) );
  OAI22_X1 U18334 ( .A1(n19032), .A2(n16329), .B1(n16324), .B2(n19110), .ZN(
        n15318) );
  AOI211_X1 U18335 ( .C1(n15320), .C2(n16313), .A(n15319), .B(n15318), .ZN(
        n15321) );
  OAI21_X1 U18336 ( .B1(n16317), .B2(n15322), .A(n15321), .ZN(P2_U3040) );
  INV_X1 U18337 ( .A(n15328), .ZN(n19853) );
  AOI22_X1 U18338 ( .A1(n19047), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15323), .B2(n19029), .ZN(n15330) );
  NAND2_X1 U18339 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15330), .ZN(n15326) );
  NAND2_X1 U18340 ( .A1(n15324), .A2(n19850), .ZN(n15325) );
  OAI211_X1 U18341 ( .C1(n12594), .C2(n19853), .A(n15326), .B(n15325), .ZN(
        n15327) );
  MUX2_X1 U18342 ( .A(n15327), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n19855), .Z(P2_U3601) );
  INV_X1 U18343 ( .A(n19872), .ZN(n15329) );
  NAND2_X1 U18344 ( .A1(n15329), .A2(n15328), .ZN(n15336) );
  NOR2_X1 U18345 ( .A1(n15330), .A2(n11027), .ZN(n19846) );
  OAI211_X1 U18346 ( .C1(n15333), .C2(n15332), .A(n19029), .B(n15331), .ZN(
        n19072) );
  OAI21_X1 U18347 ( .B1(n19029), .B2(n15334), .A(n19072), .ZN(n19848) );
  NAND2_X1 U18348 ( .A1(n19846), .A2(n19848), .ZN(n15335) );
  OAI211_X1 U18349 ( .C1(n19861), .C2(n15337), .A(n15336), .B(n15335), .ZN(
        n15338) );
  MUX2_X1 U18350 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15338), .S(
        n19857), .Z(P2_U3599) );
  AOI22_X1 U18351 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15343) );
  AOI22_X1 U18352 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15482), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U18353 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15341) );
  INV_X2 U18354 ( .A(n9694), .ZN(n17138) );
  AOI22_X1 U18355 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15340) );
  NAND4_X1 U18356 ( .A1(n15343), .A2(n15342), .A3(n15341), .A4(n15340), .ZN(
        n15350) );
  AOI22_X1 U18357 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15348) );
  AOI22_X1 U18358 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15347) );
  AOI22_X1 U18359 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16937), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U18360 ( .A1(n9654), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15345) );
  NAND4_X1 U18361 ( .A1(n15348), .A2(n15347), .A3(n15346), .A4(n15345), .ZN(
        n15349) );
  NOR2_X1 U18362 ( .A1(n15350), .A2(n15349), .ZN(n16966) );
  AOI22_X1 U18363 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U18364 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15353) );
  AOI22_X1 U18365 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U18366 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15351) );
  NAND4_X1 U18367 ( .A1(n15354), .A2(n15353), .A3(n15352), .A4(n15351), .ZN(
        n15361) );
  AOI22_X1 U18368 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15359) );
  AOI22_X1 U18369 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15358) );
  AOI22_X1 U18370 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15357) );
  AOI22_X1 U18371 ( .A1(n15518), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15356) );
  NAND4_X1 U18372 ( .A1(n15359), .A2(n15358), .A3(n15357), .A4(n15356), .ZN(
        n15360) );
  NOR2_X1 U18373 ( .A1(n15361), .A2(n15360), .ZN(n16978) );
  AOI22_X1 U18374 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U18375 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U18376 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15363) );
  AOI22_X1 U18377 ( .A1(n17098), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15362) );
  NAND4_X1 U18378 ( .A1(n15365), .A2(n15364), .A3(n15363), .A4(n15362), .ZN(
        n15371) );
  AOI22_X1 U18379 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U18380 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U18381 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15367) );
  AOI22_X1 U18382 ( .A1(n14111), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15366) );
  NAND4_X1 U18383 ( .A1(n15369), .A2(n15368), .A3(n15367), .A4(n15366), .ZN(
        n15370) );
  NOR2_X1 U18384 ( .A1(n15371), .A2(n15370), .ZN(n16988) );
  AOI22_X1 U18385 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17098), .B1(
        n17099), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U18386 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17097), .ZN(n15374) );
  AOI22_X1 U18387 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U18388 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17188), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15372) );
  NAND4_X1 U18389 ( .A1(n15375), .A2(n15374), .A3(n15373), .A4(n15372), .ZN(
        n15381) );
  AOI22_X1 U18390 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n9654), .B1(
        n16937), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15379) );
  AOI22_X1 U18391 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15378) );
  AOI22_X1 U18392 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17138), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n15518), .ZN(n15377) );
  AOI22_X1 U18393 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15376) );
  NAND4_X1 U18394 ( .A1(n15379), .A2(n15378), .A3(n15377), .A4(n15376), .ZN(
        n15380) );
  NOR2_X1 U18395 ( .A1(n15381), .A2(n15380), .ZN(n16989) );
  NOR2_X1 U18396 ( .A1(n16988), .A2(n16989), .ZN(n16987) );
  AOI22_X1 U18397 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U18398 ( .A1(n15518), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U18399 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15382) );
  OAI21_X1 U18400 ( .B1(n9694), .B2(n20889), .A(n15382), .ZN(n15388) );
  AOI22_X1 U18401 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16937), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U18402 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U18403 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U18404 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15383) );
  NAND4_X1 U18405 ( .A1(n15386), .A2(n15385), .A3(n15384), .A4(n15383), .ZN(
        n15387) );
  AOI211_X1 U18406 ( .C1(n17110), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n15388), .B(n15387), .ZN(n15389) );
  NAND3_X1 U18407 ( .A1(n15391), .A2(n15390), .A3(n15389), .ZN(n16983) );
  NAND2_X1 U18408 ( .A1(n16987), .A2(n16983), .ZN(n16982) );
  NOR2_X1 U18409 ( .A1(n16978), .A2(n16982), .ZN(n16977) );
  AOI22_X1 U18410 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U18411 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15401) );
  INV_X1 U18412 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U18413 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15392) );
  OAI21_X1 U18414 ( .B1(n15393), .B2(n17218), .A(n15392), .ZN(n15399) );
  AOI22_X1 U18415 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U18416 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U18417 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15395) );
  AOI22_X1 U18418 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15394) );
  NAND4_X1 U18419 ( .A1(n15397), .A2(n15396), .A3(n15395), .A4(n15394), .ZN(
        n15398) );
  AOI211_X1 U18420 ( .C1(n17115), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n15399), .B(n15398), .ZN(n15400) );
  NAND3_X1 U18421 ( .A1(n15402), .A2(n15401), .A3(n15400), .ZN(n16972) );
  NAND2_X1 U18422 ( .A1(n16977), .A2(n16972), .ZN(n16971) );
  NOR2_X1 U18423 ( .A1(n16966), .A2(n16971), .ZN(n16965) );
  AOI22_X1 U18424 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U18425 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15411) );
  INV_X1 U18426 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U18427 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15403) );
  OAI21_X1 U18428 ( .B1(n9699), .B2(n20772), .A(n15403), .ZN(n15409) );
  AOI22_X1 U18429 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U18430 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16937), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15406) );
  AOI22_X1 U18431 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15405) );
  AOI22_X1 U18432 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15404) );
  NAND4_X1 U18433 ( .A1(n15407), .A2(n15406), .A3(n15405), .A4(n15404), .ZN(
        n15408) );
  AOI211_X1 U18434 ( .C1(n15482), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15409), .B(n15408), .ZN(n15410) );
  NAND3_X1 U18435 ( .A1(n15412), .A2(n15411), .A3(n15410), .ZN(n15413) );
  NAND2_X1 U18436 ( .A1(n16965), .A2(n15413), .ZN(n16960) );
  OAI21_X1 U18437 ( .B1(n16965), .B2(n15413), .A(n16960), .ZN(n17255) );
  NAND3_X1 U18438 ( .A1(n15415), .A2(n17342), .A3(n15414), .ZN(n15416) );
  INV_X1 U18439 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16969) );
  INV_X1 U18440 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17060) );
  INV_X1 U18441 ( .A(n17232), .ZN(n17229) );
  INV_X1 U18442 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16743) );
  INV_X1 U18443 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16758) );
  NAND4_X1 U18444 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n15419)
         );
  INV_X1 U18445 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16882) );
  NAND3_X1 U18446 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17216) );
  NOR2_X1 U18447 ( .A1(n16882), .A2(n17216), .ZN(n17213) );
  NAND2_X1 U18448 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17213), .ZN(n17212) );
  NAND3_X1 U18449 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n15435) );
  NOR2_X1 U18450 ( .A1(n17212), .A2(n15435), .ZN(n17197) );
  NAND4_X1 U18451 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n17197), .ZN(n15418) );
  NOR4_X1 U18452 ( .A1(n16743), .A2(n16758), .A3(n15419), .A4(n15418), .ZN(
        n17073) );
  NAND3_X1 U18453 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17229), .A3(n17073), 
        .ZN(n17048) );
  NOR2_X1 U18454 ( .A1(n17060), .A2(n17048), .ZN(n17046) );
  NAND2_X1 U18455 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17046), .ZN(n17045) );
  NOR2_X1 U18456 ( .A1(n18234), .A2(n17045), .ZN(n17033) );
  NAND2_X1 U18457 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17033), .ZN(n16975) );
  INV_X1 U18458 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16624) );
  INV_X1 U18459 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16647) );
  NOR2_X1 U18460 ( .A1(n16624), .A2(n16647), .ZN(n15420) );
  NAND4_X1 U18461 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n15420), .ZN(n16926) );
  NOR2_X1 U18462 ( .A1(n16975), .A2(n16926), .ZN(n16981) );
  NAND2_X1 U18463 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16981), .ZN(n16970) );
  INV_X1 U18464 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16589) );
  OAI21_X1 U18465 ( .B1(n16969), .B2(n16970), .A(n16589), .ZN(n15421) );
  NOR2_X1 U18466 ( .A1(n16589), .A2(n16969), .ZN(n16958) );
  NOR2_X1 U18467 ( .A1(n18234), .A2(n17232), .ZN(n17223) );
  INV_X1 U18468 ( .A(n17223), .ZN(n17235) );
  NAND2_X1 U18469 ( .A1(n17219), .A2(n16970), .ZN(n16968) );
  OAI21_X1 U18470 ( .B1(n16958), .B2(n17235), .A(n16968), .ZN(n16962) );
  NAND2_X1 U18471 ( .A1(n15421), .A2(n16962), .ZN(n15422) );
  OAI21_X1 U18472 ( .B1(n17255), .B2(n17219), .A(n15422), .ZN(P3_U2675) );
  AOI22_X1 U18473 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16937), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18474 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18475 ( .A1(n14111), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U18476 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15425) );
  NAND4_X1 U18477 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n15434) );
  AOI22_X1 U18478 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18479 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U18480 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U18481 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15429) );
  NAND4_X1 U18482 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15433) );
  NOR2_X1 U18483 ( .A1(n15434), .A2(n15433), .ZN(n17326) );
  INV_X1 U18484 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17124) );
  NOR2_X1 U18485 ( .A1(n17232), .A2(n17212), .ZN(n17208) );
  INV_X1 U18486 ( .A(n17208), .ZN(n17203) );
  NOR2_X1 U18487 ( .A1(n15435), .A2(n17203), .ZN(n17195) );
  NAND3_X1 U18488 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17195), .ZN(n17179) );
  INV_X1 U18489 ( .A(n17179), .ZN(n17153) );
  AND2_X1 U18490 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17153), .ZN(n17168) );
  NAND2_X1 U18491 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17168), .ZN(n17150) );
  NOR2_X1 U18492 ( .A1(n17124), .A2(n17150), .ZN(n17137) );
  NAND2_X1 U18493 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17137), .ZN(n17078) );
  OAI21_X1 U18494 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17137), .A(n17078), .ZN(
        n15436) );
  AOI22_X1 U18495 ( .A1(n17233), .A2(n17326), .B1(n15436), .B2(n17219), .ZN(
        P3_U2690) );
  NAND2_X1 U18496 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18378) );
  AOI221_X1 U18497 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18378), .C1(n15438), 
        .C2(n18378), .A(n15437), .ZN(n18189) );
  NOR2_X1 U18498 ( .A1(n15439), .A2(n18651), .ZN(n15440) );
  OAI21_X1 U18499 ( .B1(n15440), .B2(n18447), .A(n18190), .ZN(n18187) );
  AOI22_X1 U18500 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18189), .B1(
        n18187), .B2(n18192), .ZN(P3_U2865) );
  AOI22_X1 U18501 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15444) );
  AOI22_X1 U18502 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15443) );
  AOI22_X1 U18503 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15442) );
  AOI22_X1 U18504 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15441) );
  NAND4_X1 U18505 ( .A1(n15444), .A2(n15443), .A3(n15442), .A4(n15441), .ZN(
        n15450) );
  AOI22_X1 U18506 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9654), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18507 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15447) );
  AOI22_X1 U18508 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15446) );
  AOI22_X1 U18509 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15445) );
  NAND4_X1 U18510 ( .A1(n15448), .A2(n15447), .A3(n15446), .A4(n15445), .ZN(
        n15449) );
  AOI22_X1 U18511 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U18512 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9656), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U18513 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U18514 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15451) );
  NAND4_X1 U18515 ( .A1(n15454), .A2(n15453), .A3(n15452), .A4(n15451), .ZN(
        n15460) );
  AOI22_X1 U18516 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U18517 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18518 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18519 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15455) );
  NAND4_X1 U18520 ( .A1(n15458), .A2(n15457), .A3(n15456), .A4(n15455), .ZN(
        n15459) );
  AOI22_X1 U18521 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18522 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15463) );
  AOI22_X1 U18523 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15462) );
  AOI22_X1 U18524 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15461) );
  NAND4_X1 U18525 ( .A1(n15464), .A2(n15463), .A3(n15462), .A4(n15461), .ZN(
        n15470) );
  AOI22_X1 U18526 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15468) );
  AOI22_X1 U18527 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18528 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18529 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15465) );
  NAND4_X1 U18530 ( .A1(n15468), .A2(n15467), .A3(n15466), .A4(n15465), .ZN(
        n15469) );
  AOI22_X1 U18531 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18532 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15473) );
  AOI22_X1 U18533 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18534 ( .A1(n14111), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18535 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18536 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18537 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15478) );
  OAI21_X1 U18538 ( .B1(n15479), .B2(n20889), .A(n15478), .ZN(n15480) );
  NAND3_X1 U18539 ( .A1(n10248), .A2(n10250), .A3(n15481), .ZN(n17380) );
  AOI22_X1 U18540 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15494) );
  AOI22_X1 U18541 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15493) );
  INV_X1 U18542 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U18543 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15483) );
  OAI21_X1 U18544 ( .B1(n17140), .B2(n17155), .A(n15483), .ZN(n15492) );
  AOI22_X1 U18545 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14106), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18546 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U18547 ( .A1(n15344), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15485), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15488) );
  NAND4_X1 U18548 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15491) );
  NAND2_X1 U18549 ( .A1(n17380), .A2(n15576), .ZN(n15532) );
  NOR2_X1 U18550 ( .A1(n17371), .A2(n15532), .ZN(n15534) );
  AOI22_X1 U18551 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U18552 ( .A1(n9656), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15504) );
  INV_X1 U18553 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U18554 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15495) );
  OAI21_X1 U18555 ( .B1(n9694), .B2(n15496), .A(n15495), .ZN(n15502) );
  AOI22_X1 U18556 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18557 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18558 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U18559 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15497) );
  NAND4_X1 U18560 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15501) );
  AOI211_X1 U18561 ( .C1(n15517), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15502), .B(n15501), .ZN(n15503) );
  NAND3_X1 U18562 ( .A1(n15505), .A2(n15504), .A3(n15503), .ZN(n17366) );
  NAND2_X1 U18563 ( .A1(n15534), .A2(n17366), .ZN(n15516) );
  AOI22_X1 U18564 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U18565 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U18566 ( .A1(n9654), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U18567 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15506) );
  NAND4_X1 U18568 ( .A1(n15509), .A2(n15508), .A3(n15507), .A4(n15506), .ZN(
        n15515) );
  AOI22_X1 U18569 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17099), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U18570 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15512) );
  AOI22_X1 U18571 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U18572 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15510) );
  NAND4_X1 U18573 ( .A1(n15513), .A2(n15512), .A3(n15511), .A4(n15510), .ZN(
        n15514) );
  INV_X1 U18574 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17898) );
  INV_X1 U18575 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18090) );
  INV_X1 U18576 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18104) );
  XNOR2_X1 U18577 ( .A(n15516), .B(n17363), .ZN(n17812) );
  INV_X1 U18578 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18802) );
  AOI22_X1 U18579 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U18580 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18581 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15519) );
  OAI21_X1 U18582 ( .B1(n17140), .B2(n20869), .A(n15519), .ZN(n15525) );
  AOI22_X1 U18583 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18584 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15344), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18585 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15521) );
  AOI22_X1 U18586 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15520) );
  NAND4_X1 U18587 ( .A1(n15523), .A2(n15522), .A3(n15521), .A4(n15520), .ZN(
        n15524) );
  AOI211_X1 U18588 ( .C1(n17098), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n15525), .B(n15524), .ZN(n15526) );
  NAND3_X1 U18589 ( .A1(n15528), .A2(n15527), .A3(n15526), .ZN(n17867) );
  NAND2_X1 U18590 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17867), .ZN(
        n17866) );
  INV_X1 U18591 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18154) );
  NOR2_X1 U18592 ( .A1(n18154), .A2(n15529), .ZN(n15530) );
  INV_X1 U18593 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18128) );
  NOR2_X1 U18594 ( .A1(n15531), .A2(n18128), .ZN(n15533) );
  NOR2_X2 U18595 ( .A1(n15533), .A2(n17837), .ZN(n17821) );
  XNOR2_X1 U18596 ( .A(n15534), .B(n17366), .ZN(n17822) );
  INV_X1 U18597 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18105) );
  XOR2_X1 U18598 ( .A(n18105), .B(n15538), .Z(n17802) );
  OAI21_X1 U18599 ( .B1(n15540), .B2(n17354), .A(n17770), .ZN(n15541) );
  NOR2_X1 U18600 ( .A1(n15542), .A2(n15541), .ZN(n15543) );
  NOR4_X1 U18601 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15544) );
  AOI21_X1 U18602 ( .B1(n17710), .B2(n15544), .A(n17758), .ZN(n17658) );
  NAND2_X1 U18603 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18058) );
  INV_X1 U18604 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17744) );
  NOR2_X1 U18605 ( .A1(n18058), .A2(n17744), .ZN(n18060) );
  INV_X1 U18606 ( .A(n18060), .ZN(n18036) );
  NOR2_X1 U18607 ( .A1(n18036), .A2(n17718), .ZN(n18021) );
  INV_X1 U18608 ( .A(n18021), .ZN(n17708) );
  NAND2_X1 U18609 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17677) );
  NOR2_X1 U18610 ( .A1(n17708), .A2(n17677), .ZN(n17999) );
  INV_X1 U18611 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18004) );
  NAND2_X1 U18612 ( .A1(n17758), .A2(n18004), .ZN(n15546) );
  INV_X1 U18613 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17987) );
  NAND2_X1 U18614 ( .A1(n17654), .A2(n17987), .ZN(n17653) );
  INV_X1 U18615 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17924) );
  NOR2_X1 U18616 ( .A1(n18004), .A2(n17987), .ZN(n17979) );
  INV_X1 U18617 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17637) );
  NAND2_X1 U18618 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17938) );
  INV_X1 U18619 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17937) );
  NOR3_X1 U18620 ( .A1(n17637), .A2(n17938), .A3(n17937), .ZN(n17584) );
  AND2_X1 U18621 ( .A1(n17584), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15552) );
  NAND2_X1 U18622 ( .A1(n17979), .A2(n15552), .ZN(n17574) );
  NOR2_X1 U18623 ( .A1(n17924), .A2(n17574), .ZN(n17920) );
  INV_X1 U18624 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17621) );
  NAND2_X1 U18625 ( .A1(n17643), .A2(n17621), .ZN(n15549) );
  NOR2_X1 U18626 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15549), .ZN(
        n17605) );
  NAND2_X1 U18627 ( .A1(n17605), .A2(n17937), .ZN(n17592) );
  NAND2_X1 U18628 ( .A1(n17979), .A2(n17593), .ZN(n17603) );
  NOR2_X1 U18629 ( .A1(n17546), .A2(n17770), .ZN(n15553) );
  NAND2_X1 U18630 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17879) );
  INV_X1 U18631 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U18632 ( .A1(n17758), .A2(n17500), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17770), .ZN(n17504) );
  NOR2_X1 U18633 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15556), .ZN(
        n15678) );
  AOI21_X1 U18634 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15556), .A(
        n15678), .ZN(n16390) );
  NAND2_X1 U18635 ( .A1(n15559), .A2(n18203), .ZN(n15560) );
  NOR2_X1 U18636 ( .A1(n17239), .A2(n15560), .ZN(n15569) );
  NAND2_X1 U18637 ( .A1(n15569), .A2(n15557), .ZN(n16407) );
  INV_X1 U18638 ( .A(n16407), .ZN(n18627) );
  AOI21_X1 U18639 ( .B1(n15559), .B2(n15558), .A(n18219), .ZN(n15565) );
  INV_X1 U18640 ( .A(n15559), .ZN(n18208) );
  AOI21_X1 U18641 ( .B1(n18841), .B2(n18208), .A(n16542), .ZN(n15561) );
  AOI21_X1 U18642 ( .B1(n15561), .B2(n15560), .A(n18708), .ZN(n16523) );
  NAND3_X1 U18643 ( .A1(n18622), .A2(n16523), .A3(n15562), .ZN(n15563) );
  OAI211_X1 U18644 ( .C1(n15565), .C2(n16349), .A(n15564), .B(n15563), .ZN(
        n15570) );
  INV_X1 U18645 ( .A(n15566), .ZN(n15568) );
  AOI21_X1 U18646 ( .B1(n15568), .B2(n15567), .A(n16522), .ZN(n16348) );
  INV_X1 U18647 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17524) );
  INV_X1 U18648 ( .A(n17879), .ZN(n15611) );
  INV_X1 U18649 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17919) );
  INV_X1 U18650 ( .A(n17371), .ZN(n15574) );
  INV_X1 U18651 ( .A(n15576), .ZN(n17375) );
  NAND2_X1 U18652 ( .A1(n17380), .A2(n17867), .ZN(n15575) );
  NAND2_X1 U18653 ( .A1(n17375), .A2(n15575), .ZN(n15573) );
  INV_X1 U18654 ( .A(n17363), .ZN(n15572) );
  NAND2_X1 U18655 ( .A1(n15571), .A2(n15572), .ZN(n15589) );
  NOR2_X1 U18656 ( .A1(n17360), .A2(n15589), .ZN(n15593) );
  NAND2_X1 U18657 ( .A1(n15593), .A2(n17354), .ZN(n15594) );
  XOR2_X1 U18658 ( .A(n15572), .B(n15571), .Z(n15587) );
  AND2_X1 U18659 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15587), .ZN(
        n15588) );
  XNOR2_X1 U18660 ( .A(n15574), .B(n15573), .ZN(n15583) );
  NOR2_X1 U18661 ( .A1(n18128), .A2(n15583), .ZN(n15584) );
  XNOR2_X1 U18662 ( .A(n15576), .B(n15575), .ZN(n15577) );
  NOR2_X1 U18663 ( .A1(n15577), .A2(n18154), .ZN(n15582) );
  XOR2_X1 U18664 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15577), .Z(
        n17850) );
  INV_X1 U18665 ( .A(n17380), .ZN(n15579) );
  INV_X1 U18666 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18819) );
  NOR2_X1 U18667 ( .A1(n15579), .A2(n18819), .ZN(n15580) );
  INV_X1 U18668 ( .A(n17867), .ZN(n15701) );
  NAND3_X1 U18669 ( .A1(n15701), .A2(n15579), .A3(n18819), .ZN(n15578) );
  OAI221_X1 U18670 ( .B1(n15580), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15701), .C2(n15579), .A(n15578), .ZN(n17849) );
  NOR2_X1 U18671 ( .A1(n17850), .A2(n17849), .ZN(n15581) );
  NOR2_X1 U18672 ( .A1(n15582), .A2(n15581), .ZN(n17840) );
  XOR2_X1 U18673 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15583), .Z(
        n17839) );
  NOR2_X1 U18674 ( .A1(n17840), .A2(n17839), .ZN(n17838) );
  NOR2_X1 U18675 ( .A1(n15584), .A2(n17838), .ZN(n17825) );
  XNOR2_X1 U18676 ( .A(n17366), .B(n15585), .ZN(n17826) );
  NOR2_X1 U18677 ( .A1(n17825), .A2(n17826), .ZN(n15586) );
  NAND2_X1 U18678 ( .A1(n17825), .A2(n17826), .ZN(n17824) );
  OAI21_X1 U18679 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15586), .A(
        n17824), .ZN(n17810) );
  XOR2_X1 U18680 ( .A(n10148), .B(n15587), .Z(n17809) );
  NOR2_X1 U18681 ( .A1(n17810), .A2(n17809), .ZN(n17808) );
  XNOR2_X1 U18682 ( .A(n17360), .B(n15589), .ZN(n15591) );
  NOR2_X1 U18683 ( .A1(n15590), .A2(n15591), .ZN(n15592) );
  XNOR2_X1 U18684 ( .A(n15591), .B(n15590), .ZN(n17798) );
  NOR2_X1 U18685 ( .A1(n15592), .A2(n17797), .ZN(n15595) );
  XOR2_X1 U18686 ( .A(n16409), .B(n15593), .Z(n15596) );
  NAND2_X1 U18687 ( .A1(n15595), .A2(n15596), .ZN(n17784) );
  NAND2_X1 U18688 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17784), .ZN(
        n15598) );
  NOR2_X1 U18689 ( .A1(n15594), .A2(n15598), .ZN(n15600) );
  INV_X1 U18690 ( .A(n15594), .ZN(n15599) );
  OR2_X1 U18691 ( .A1(n15596), .A2(n15595), .ZN(n17785) );
  OAI21_X1 U18692 ( .B1(n15599), .B2(n15598), .A(n17785), .ZN(n15597) );
  AOI21_X1 U18693 ( .B1(n15599), .B2(n15598), .A(n15597), .ZN(n17779) );
  NOR2_X2 U18694 ( .A1(n15600), .A2(n17778), .ZN(n18053) );
  NAND2_X1 U18695 ( .A1(n15611), .A2(n17538), .ZN(n17875) );
  NOR3_X1 U18696 ( .A1(n17524), .A2(n17500), .A3(n17875), .ZN(n16384) );
  INV_X1 U18697 ( .A(n16384), .ZN(n16411) );
  NOR2_X2 U18698 ( .A1(n15601), .A2(n15609), .ZN(n18639) );
  NOR2_X1 U18699 ( .A1(n15603), .A2(n15602), .ZN(n18852) );
  NOR3_X1 U18700 ( .A1(n15606), .A2(n18841), .A3(n15605), .ZN(n15608) );
  NOR2_X1 U18701 ( .A1(n15608), .A2(n15607), .ZN(n18633) );
  NAND2_X1 U18702 ( .A1(n18054), .A2(n18175), .ZN(n18172) );
  NAND3_X1 U18703 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18006) );
  INV_X1 U18704 ( .A(n18006), .ZN(n18101) );
  OAI21_X1 U18705 ( .B1(n18802), .B2(n18819), .A(n18154), .ZN(n18145) );
  NAND2_X1 U18706 ( .A1(n18101), .A2(n18145), .ZN(n18085) );
  NAND3_X1 U18707 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18007) );
  NOR2_X1 U18708 ( .A1(n18085), .A2(n18007), .ZN(n17995) );
  NAND2_X1 U18709 ( .A1(n17975), .A2(n17995), .ZN(n17933) );
  INV_X1 U18710 ( .A(n17933), .ZN(n17978) );
  OAI21_X1 U18711 ( .B1(n18657), .B2(n18819), .A(n18639), .ZN(n18155) );
  NOR2_X1 U18712 ( .A1(n18154), .A2(n18802), .ZN(n18125) );
  NAND2_X1 U18713 ( .A1(n18101), .A2(n18125), .ZN(n18084) );
  NOR2_X1 U18714 ( .A1(n18007), .A2(n18084), .ZN(n17994) );
  NAND2_X1 U18715 ( .A1(n17975), .A2(n17994), .ZN(n15612) );
  INV_X1 U18716 ( .A(n15612), .ZN(n17976) );
  AOI22_X1 U18717 ( .A1(n18148), .A2(n17978), .B1(n18155), .B2(n17976), .ZN(
        n16403) );
  NOR2_X1 U18718 ( .A1(n16403), .A2(n17574), .ZN(n17901) );
  NOR2_X1 U18719 ( .A1(n17924), .A2(n17919), .ZN(n17900) );
  NAND2_X1 U18720 ( .A1(n15611), .A2(n17900), .ZN(n17874) );
  INV_X1 U18721 ( .A(n17874), .ZN(n15615) );
  NAND2_X1 U18722 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15615), .ZN(
        n15610) );
  NOR2_X1 U18723 ( .A1(n18167), .A2(n15610), .ZN(n16406) );
  NAND2_X1 U18724 ( .A1(n17901), .A2(n16406), .ZN(n16392) );
  INV_X1 U18725 ( .A(n17759), .ZN(n17739) );
  NOR3_X1 U18726 ( .A1(n17883), .A2(n17524), .A3(n17500), .ZN(n16387) );
  INV_X1 U18727 ( .A(n16387), .ZN(n16410) );
  NAND2_X1 U18728 ( .A1(n18627), .A2(n18175), .ZN(n18182) );
  NOR2_X1 U18729 ( .A1(n17354), .A2(n18182), .ZN(n18093) );
  OAI222_X1 U18730 ( .A1(n16411), .A2(n18172), .B1(n16392), .B2(n17500), .C1(
        n16410), .C2(n17974), .ZN(n15685) );
  INV_X1 U18731 ( .A(n15685), .ZN(n15618) );
  NAND3_X1 U18732 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16371) );
  NOR2_X1 U18733 ( .A1(n16371), .A2(n17875), .ZN(n16373) );
  OAI22_X1 U18734 ( .A1(n16373), .A2(n18172), .B1(n16372), .B2(n17974), .ZN(
        n15683) );
  OR3_X2 U18735 ( .A1(n18851), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18132) );
  INV_X2 U18736 ( .A(n18132), .ZN(n18174) );
  INV_X1 U18737 ( .A(n18061), .ZN(n18067) );
  NOR2_X1 U18738 ( .A1(n17574), .A2(n15612), .ZN(n17876) );
  NAND4_X1 U18739 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n15615), .A4(n17876), .ZN(
        n15613) );
  NOR2_X1 U18740 ( .A1(n17574), .A2(n17933), .ZN(n17915) );
  AOI21_X1 U18741 ( .B1(n15615), .B2(n17915), .A(n18665), .ZN(n17878) );
  AOI211_X1 U18742 ( .C1(n17997), .C2(n15613), .A(n17878), .B(n18167), .ZN(
        n15614) );
  OAI221_X1 U18743 ( .B1(n18639), .B2(n15615), .C1(n18639), .C2(n17876), .A(
        n15614), .ZN(n15681) );
  AOI21_X1 U18744 ( .B1(n18067), .B2(n17524), .A(n15681), .ZN(n16413) );
  NAND2_X1 U18745 ( .A1(n18175), .A2(n18087), .ZN(n18162) );
  OAI22_X1 U18746 ( .A1(n18174), .A2(n16413), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18162), .ZN(n15616) );
  NOR2_X1 U18747 ( .A1(n15683), .A2(n15616), .ZN(n15617) );
  MUX2_X1 U18748 ( .A(n15618), .B(n15617), .S(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(n15619) );
  NAND2_X1 U18749 ( .A1(n18174), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16381) );
  OAI211_X1 U18750 ( .C1(n16390), .C2(n18098), .A(n15619), .B(n16381), .ZN(
        P3_U2833) );
  XOR2_X1 U18751 ( .A(n15621), .B(n15620), .Z(n16201) );
  NAND2_X1 U18752 ( .A1(n19044), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16197) );
  NAND2_X1 U18753 ( .A1(n16301), .A2(n15622), .ZN(n15623) );
  OAI211_X1 U18754 ( .C1(n16329), .C2(n16207), .A(n16197), .B(n15623), .ZN(
        n15624) );
  AOI21_X1 U18755 ( .B1(n16201), .B2(n16334), .A(n15624), .ZN(n15625) );
  OAI221_X1 U18756 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15628), 
        .C1(n15627), .C2(n15626), .A(n15625), .ZN(P2_U3030) );
  OAI22_X1 U18757 ( .A1(n15630), .A2(n18958), .B1(n19065), .B2(n15629), .ZN(
        n15631) );
  INV_X1 U18758 ( .A(n15631), .ZN(n15640) );
  AOI211_X1 U18759 ( .C1(n15634), .C2(n15633), .A(n15632), .B(n19759), .ZN(
        n15638) );
  OAI222_X1 U18760 ( .A1(n19024), .A2(n15636), .B1(n15635), .B2(n19042), .C1(
        n19818), .C2(n19059), .ZN(n15637) );
  AOI211_X1 U18761 ( .C1(n19038), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15638), .B(n15637), .ZN(n15639) );
  NAND2_X1 U18762 ( .A1(n15640), .A2(n15639), .ZN(P2_U2833) );
  NAND2_X1 U18763 ( .A1(n15646), .A2(n15641), .ZN(n15654) );
  AND2_X1 U18764 ( .A1(n15646), .A2(n15642), .ZN(n15652) );
  NOR2_X1 U18765 ( .A1(n15643), .A2(n20504), .ZN(n15644) );
  AND2_X1 U18766 ( .A1(n15645), .A2(n15644), .ZN(n15650) );
  INV_X1 U18767 ( .A(n15650), .ZN(n15648) );
  OAI211_X1 U18768 ( .C1(n15648), .C2(n20412), .A(n15647), .B(n15646), .ZN(
        n15649) );
  OAI21_X1 U18769 ( .B1(n15650), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15649), .ZN(n15651) );
  AOI222_X1 U18770 ( .A1(n15652), .A2(n20474), .B1(n15652), .B2(n15651), .C1(
        n20474), .C2(n15651), .ZN(n15653) );
  AOI222_X1 U18771 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15654), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15653), .C1(n15654), 
        .C2(n15653), .ZN(n15662) );
  OAI21_X1 U18772 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15655), .ZN(n15657) );
  NAND4_X1 U18773 ( .A1(n15659), .A2(n15658), .A3(n15657), .A4(n15656), .ZN(
        n15660) );
  AOI211_X1 U18774 ( .C1(n15662), .C2(n20101), .A(n15661), .B(n15660), .ZN(
        n15677) );
  INV_X1 U18775 ( .A(n15663), .ZN(n15665) );
  NOR3_X1 U18776 ( .A1(n15665), .A2(n15664), .A3(n15689), .ZN(n15668) );
  OAI22_X1 U18777 ( .A1(n15668), .A2(n15667), .B1(n20654), .B2(n15666), .ZN(
        n16091) );
  AOI21_X1 U18778 ( .B1(n15677), .B2(n16091), .A(n20644), .ZN(n16097) );
  INV_X1 U18779 ( .A(n16097), .ZN(n16095) );
  OAI211_X1 U18780 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20654), .A(n15670), 
        .B(n15669), .ZN(n15675) );
  AND2_X1 U18781 ( .A1(n20644), .A2(n15671), .ZN(n15672) );
  AOI22_X1 U18782 ( .A1(n15673), .A2(n16091), .B1(n20737), .B2(n15672), .ZN(
        n15674) );
  OAI21_X1 U18783 ( .B1(n16095), .B2(n15675), .A(n15674), .ZN(n15676) );
  OAI21_X1 U18784 ( .B1(n15677), .B2(n19913), .A(n15676), .ZN(P1_U3161) );
  NAND3_X1 U18785 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n16408), .ZN(n16358) );
  NAND2_X1 U18786 ( .A1(n17758), .A2(n16358), .ZN(n16357) );
  NOR2_X1 U18787 ( .A1(n17758), .A2(n15678), .ZN(n16360) );
  INV_X1 U18788 ( .A(n16360), .ZN(n15679) );
  NAND2_X1 U18789 ( .A1(n16357), .A2(n15679), .ZN(n15680) );
  XOR2_X1 U18790 ( .A(n15680), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16376) );
  INV_X1 U18791 ( .A(n18162), .ZN(n15682) );
  AOI22_X1 U18792 ( .A1(n15682), .A2(n16371), .B1(n18132), .B2(n15681), .ZN(
        n16391) );
  INV_X1 U18793 ( .A(n16391), .ZN(n15684) );
  INV_X1 U18794 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18779) );
  NOR2_X1 U18795 ( .A1(n18132), .A2(n18779), .ZN(n16370) );
  AOI221_X1 U18796 ( .B1(n15684), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), 
        .C1(n15683), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n16370), .ZN(
        n15687) );
  INV_X1 U18797 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16393) );
  NAND3_X1 U18798 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16393), .A3(
        n15685), .ZN(n15686) );
  OAI211_X1 U18799 ( .C1(n16376), .C2(n18098), .A(n15687), .B(n15686), .ZN(
        P3_U2832) );
  INV_X1 U18800 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19911) );
  INV_X1 U18801 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20743) );
  NOR2_X1 U18802 ( .A1(n20657), .A2(n20743), .ZN(n20652) );
  INV_X1 U18803 ( .A(HOLD), .ZN(n20648) );
  NOR2_X1 U18804 ( .A1(n19911), .A2(n20648), .ZN(n20650) );
  OAI22_X1 U18805 ( .A1(n20652), .A2(n20650), .B1(n20660), .B2(n20648), .ZN(
        n15688) );
  OAI211_X1 U18806 ( .C1(n20654), .C2(n19911), .A(n15689), .B(n15688), .ZN(
        P1_U3195) );
  INV_X1 U18807 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16510) );
  NOR2_X1 U18808 ( .A1(n20010), .A2(n16510), .ZN(P1_U2905) );
  NOR3_X1 U18809 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12960), .A3(n19764), 
        .ZN(n19757) );
  OAI21_X1 U18810 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n16339), .ZN(n15690) );
  AOI211_X1 U18811 ( .C1(n15691), .C2(n19470), .A(n19757), .B(n15690), .ZN(
        P2_U3178) );
  OAI221_X1 U18812 ( .B1(n15692), .B2(n16339), .C1(n19900), .C2(n16339), .A(
        n19447), .ZN(n19894) );
  NOR2_X1 U18813 ( .A1(n15693), .A2(n19894), .ZN(P2_U3047) );
  NAND3_X1 U18814 ( .A1(n18622), .A2(n18836), .A3(n18842), .ZN(n17428) );
  NAND3_X1 U18815 ( .A1(n18841), .A2(n15695), .A3(n15694), .ZN(n15696) );
  AOI22_X1 U18816 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17382), .B1(n15699), .B2(
        P3_EAX_REG_0__SCAN_IN), .ZN(n15700) );
  INV_X1 U18817 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17462) );
  NAND2_X1 U18818 ( .A1(n17462), .A2(n17356), .ZN(n17383) );
  OAI211_X1 U18819 ( .C1(n15701), .C2(n17376), .A(n15700), .B(n17383), .ZN(
        P3_U2735) );
  INV_X1 U18820 ( .A(n15702), .ZN(n15707) );
  INV_X1 U18821 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15703) );
  OAI22_X1 U18822 ( .A1(n19984), .A2(n15704), .B1(n15703), .B2(n19996), .ZN(
        n15705) );
  AOI221_X1 U18823 ( .B1(n15708), .B2(P1_REIP_REG_26__SCAN_IN), .C1(n15707), 
        .C2(n15706), .A(n15705), .ZN(n15711) );
  OAI22_X1 U18824 ( .A1(n15817), .A2(n19944), .B1(n15825), .B2(n19995), .ZN(
        n15709) );
  INV_X1 U18825 ( .A(n15709), .ZN(n15710) );
  OAI211_X1 U18826 ( .C1(n19985), .C2(n15928), .A(n15711), .B(n15710), .ZN(
        P1_U2814) );
  INV_X1 U18827 ( .A(n15712), .ZN(n15830) );
  AOI22_X1 U18828 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15722), .B1(n15714), 
        .B2(n15713), .ZN(n15716) );
  AOI22_X1 U18829 ( .A1(n19997), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19977), .ZN(n15715) );
  OAI211_X1 U18830 ( .C1(n15947), .C2(n19985), .A(n15716), .B(n15715), .ZN(
        n15717) );
  AOI21_X1 U18831 ( .B1(n15830), .B2(n19958), .A(n15717), .ZN(n15718) );
  OAI21_X1 U18832 ( .B1(n15833), .B2(n19995), .A(n15718), .ZN(P1_U2816) );
  AOI22_X1 U18833 ( .A1(n19997), .A2(P1_EBX_REG_23__SCAN_IN), .B1(n19989), 
        .B2(n15719), .ZN(n15728) );
  INV_X1 U18834 ( .A(n15720), .ZN(n15953) );
  NOR3_X1 U18835 ( .A1(n15803), .A2(n15747), .A3(n15721), .ZN(n15736) );
  AOI21_X1 U18836 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15736), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15724) );
  INV_X1 U18837 ( .A(n15722), .ZN(n15723) );
  OAI22_X1 U18838 ( .A1(n15725), .A2(n19944), .B1(n15724), .B2(n15723), .ZN(
        n15726) );
  AOI21_X1 U18839 ( .B1(n19994), .B2(n15953), .A(n15726), .ZN(n15727) );
  OAI211_X1 U18840 ( .C1(n15729), .C2(n19996), .A(n15728), .B(n15727), .ZN(
        P1_U2817) );
  AOI22_X1 U18841 ( .A1(n19997), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19977), .ZN(n15730) );
  INV_X1 U18842 ( .A(n15730), .ZN(n15734) );
  OAI22_X1 U18843 ( .A1(n15732), .A2(n19944), .B1(n19985), .B2(n15731), .ZN(
        n15733) );
  AOI211_X1 U18844 ( .C1(n15736), .C2(n15735), .A(n15734), .B(n15733), .ZN(
        n15738) );
  NOR2_X1 U18845 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15803), .ZN(n15739) );
  NOR2_X1 U18846 ( .A1(n15747), .A2(n20689), .ZN(n15740) );
  OAI21_X1 U18847 ( .B1(n15740), .B2(n15803), .A(n15779), .ZN(n15748) );
  OAI21_X1 U18848 ( .B1(n15739), .B2(n15748), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15737) );
  OAI211_X1 U18849 ( .C1(n19995), .C2(n15840), .A(n15738), .B(n15737), .ZN(
        P1_U2818) );
  AOI22_X1 U18850 ( .A1(n19997), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19977), .ZN(n15746) );
  AOI22_X1 U18851 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15748), .B1(n15740), 
        .B2(n15739), .ZN(n15745) );
  NOR2_X1 U18852 ( .A1(n15741), .A2(n19985), .ZN(n15742) );
  AOI21_X1 U18853 ( .B1(n15842), .B2(n19958), .A(n15742), .ZN(n15744) );
  NAND2_X1 U18854 ( .A1(n15841), .A2(n19989), .ZN(n15743) );
  NAND4_X1 U18855 ( .A1(n15746), .A2(n15745), .A3(n15744), .A4(n15743), .ZN(
        P1_U2819) );
  NOR2_X1 U18856 ( .A1(n15803), .A2(n15747), .ZN(n15749) );
  OAI21_X1 U18857 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n15749), .A(n15748), 
        .ZN(n15754) );
  INV_X1 U18858 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15751) );
  OAI22_X1 U18859 ( .A1(n15751), .A2(n19996), .B1(n19995), .B2(n15750), .ZN(
        n15752) );
  AOI21_X1 U18860 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n19997), .A(n15752), .ZN(
        n15753) );
  OAI211_X1 U18861 ( .C1(n15755), .C2(n19944), .A(n15754), .B(n15753), .ZN(
        n15756) );
  INV_X1 U18862 ( .A(n15756), .ZN(n15757) );
  OAI21_X1 U18863 ( .B1(n19985), .B2(n15758), .A(n15757), .ZN(P1_U2820) );
  AOI21_X1 U18864 ( .B1(n19977), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19955), .ZN(n15759) );
  OAI21_X1 U18865 ( .B1(n19984), .B2(n15760), .A(n15759), .ZN(n15761) );
  AOI211_X1 U18866 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15763), .A(n15762), 
        .B(n15761), .ZN(n15768) );
  OAI22_X1 U18867 ( .A1(n15765), .A2(n19944), .B1(n15764), .B2(n19995), .ZN(
        n15766) );
  INV_X1 U18868 ( .A(n15766), .ZN(n15767) );
  OAI211_X1 U18869 ( .C1(n19985), .C2(n15976), .A(n15768), .B(n15767), .ZN(
        P1_U2822) );
  NOR2_X1 U18870 ( .A1(n15769), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15770) );
  NAND2_X1 U18871 ( .A1(n15771), .A2(n15770), .ZN(n15777) );
  NAND2_X1 U18872 ( .A1(n19997), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15776) );
  NAND2_X1 U18873 ( .A1(n19977), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15772) );
  AND2_X1 U18874 ( .A1(n15772), .A2(n19963), .ZN(n15775) );
  INV_X1 U18875 ( .A(n15854), .ZN(n15773) );
  NAND2_X1 U18876 ( .A1(n19989), .A2(n15773), .ZN(n15774) );
  NAND4_X1 U18877 ( .A1(n15777), .A2(n15776), .A3(n15775), .A4(n15774), .ZN(
        n15778) );
  AOI21_X1 U18878 ( .B1(n15851), .B2(n19958), .A(n15778), .ZN(n15784) );
  NAND2_X1 U18879 ( .A1(n15779), .A2(n15781), .ZN(n15780) );
  AND2_X1 U18880 ( .A1(n19993), .A2(n15780), .ZN(n15794) );
  INV_X1 U18881 ( .A(n15781), .ZN(n15782) );
  NOR3_X1 U18882 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15803), .A3(n15782), 
        .ZN(n15785) );
  OAI21_X1 U18883 ( .B1(n15794), .B2(n15785), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15783) );
  OAI211_X1 U18884 ( .C1(n15998), .C2(n19985), .A(n15784), .B(n15783), .ZN(
        P1_U2824) );
  AOI211_X1 U18885 ( .C1(n19977), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15785), .B(n19955), .ZN(n15786) );
  OAI21_X1 U18886 ( .B1(n19984), .B2(n14480), .A(n15786), .ZN(n15787) );
  AOI21_X1 U18887 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15794), .A(n15787), 
        .ZN(n15788) );
  OAI21_X1 U18888 ( .B1(n15789), .B2(n19944), .A(n15788), .ZN(n15790) );
  AOI21_X1 U18889 ( .B1(n15791), .B2(n19989), .A(n15790), .ZN(n15792) );
  OAI21_X1 U18890 ( .B1(n19985), .B2(n16004), .A(n15792), .ZN(P1_U2825) );
  AOI21_X1 U18891 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15793), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15801) );
  INV_X1 U18892 ( .A(n15794), .ZN(n15800) );
  OAI22_X1 U18893 ( .A1(n16006), .A2(n19985), .B1(n15795), .B2(n19984), .ZN(
        n15796) );
  AOI211_X1 U18894 ( .C1(n19977), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19955), .B(n15796), .ZN(n15799) );
  INV_X1 U18895 ( .A(n15797), .ZN(n15862) );
  AOI22_X1 U18896 ( .A1(n15862), .A2(n19958), .B1(n19989), .B2(n15861), .ZN(
        n15798) );
  OAI211_X1 U18897 ( .C1(n15801), .C2(n15800), .A(n15799), .B(n15798), .ZN(
        P1_U2826) );
  NOR2_X1 U18898 ( .A1(n15803), .A2(n15802), .ZN(n15810) );
  AOI21_X1 U18899 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15810), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15809) );
  OAI21_X1 U18900 ( .B1(n19996), .B2(n20780), .A(n19963), .ZN(n15805) );
  NOR2_X1 U18901 ( .A1(n16028), .A2(n19985), .ZN(n15804) );
  AOI211_X1 U18902 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n19997), .A(n15805), .B(
        n15804), .ZN(n15807) );
  AOI22_X1 U18903 ( .A1(n15870), .A2(n19989), .B1(n19958), .B2(n15869), .ZN(
        n15806) );
  OAI211_X1 U18904 ( .C1(n15809), .C2(n15808), .A(n15807), .B(n15806), .ZN(
        P1_U2828) );
  INV_X1 U18905 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U18906 ( .A1(n19994), .A2(n16029), .B1(n15810), .B2(n20674), .ZN(
        n15816) );
  INV_X1 U18907 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U18908 ( .A1(n15811), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n19997), 
        .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n15812) );
  OAI211_X1 U18909 ( .C1(n19996), .C2(n15813), .A(n15812), .B(n19963), .ZN(
        n15814) );
  AOI21_X1 U18910 ( .B1(n19958), .B2(n15879), .A(n15814), .ZN(n15815) );
  OAI211_X1 U18911 ( .C1(n15882), .C2(n19995), .A(n15816), .B(n15815), .ZN(
        P1_U2829) );
  AOI22_X1 U18912 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n15824) );
  INV_X1 U18913 ( .A(n15817), .ZN(n15822) );
  NOR3_X1 U18914 ( .A1(n14593), .A2(n15874), .A3(n15818), .ZN(n15819) );
  AOI21_X1 U18915 ( .B1(n9723), .B2(n15820), .A(n15819), .ZN(n15821) );
  XNOR2_X1 U18916 ( .A(n15821), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15922) );
  AOI22_X1 U18917 ( .A1(n15822), .A2(n15894), .B1(n20070), .B2(n15922), .ZN(
        n15823) );
  OAI211_X1 U18918 ( .C1(n15899), .C2(n15825), .A(n15824), .B(n15823), .ZN(
        P1_U2973) );
  AOI22_X1 U18919 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15832) );
  INV_X1 U18920 ( .A(n14593), .ZN(n15826) );
  NOR2_X1 U18921 ( .A1(n15826), .A2(n15828), .ZN(n15827) );
  MUX2_X1 U18922 ( .A(n15828), .B(n15827), .S(n15874), .Z(n15829) );
  XNOR2_X1 U18923 ( .A(n15829), .B(n15940), .ZN(n15945) );
  AOI22_X1 U18924 ( .A1(n15945), .A2(n20070), .B1(n15830), .B2(n15894), .ZN(
        n15831) );
  OAI211_X1 U18925 ( .C1(n15899), .C2(n15833), .A(n15832), .B(n15831), .ZN(
        P1_U2975) );
  AOI22_X1 U18926 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15839) );
  NAND2_X1 U18927 ( .A1(n15835), .A2(n15834), .ZN(n15836) );
  XNOR2_X1 U18928 ( .A(n15836), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15959) );
  AOI22_X1 U18929 ( .A1(n15837), .A2(n15894), .B1(n20070), .B2(n15959), .ZN(
        n15838) );
  OAI211_X1 U18930 ( .C1(n15899), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        P1_U2977) );
  AOI22_X1 U18931 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15844) );
  AOI22_X1 U18932 ( .A1(n15842), .A2(n15894), .B1(n15871), .B2(n15841), .ZN(
        n15843) );
  OAI211_X1 U18933 ( .C1(n15845), .C2(n19920), .A(n15844), .B(n15843), .ZN(
        P1_U2978) );
  AOI22_X1 U18934 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15853) );
  AOI21_X1 U18935 ( .B1(n15848), .B2(n15847), .A(n15846), .ZN(n15850) );
  XNOR2_X1 U18936 ( .A(n15850), .B(n15849), .ZN(n15994) );
  AOI22_X1 U18937 ( .A1(n15994), .A2(n20070), .B1(n15894), .B2(n15851), .ZN(
        n15852) );
  OAI211_X1 U18938 ( .C1(n15899), .C2(n15854), .A(n15853), .B(n15852), .ZN(
        P1_U2983) );
  AOI21_X1 U18939 ( .B1(n14661), .B2(n15856), .A(n15855), .ZN(n15857) );
  AOI21_X1 U18940 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15874), .A(
        n15857), .ZN(n15860) );
  MUX2_X1 U18941 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n12466), .S(
        n15858), .Z(n15859) );
  XNOR2_X1 U18942 ( .A(n15860), .B(n15859), .ZN(n16007) );
  AOI22_X1 U18943 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15864) );
  AOI22_X1 U18944 ( .A1(n15862), .A2(n15894), .B1(n15871), .B2(n15861), .ZN(
        n15863) );
  OAI211_X1 U18945 ( .C1(n16007), .C2(n19920), .A(n15864), .B(n15863), .ZN(
        P1_U2985) );
  OAI21_X1 U18946 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(n15868) );
  INV_X1 U18947 ( .A(n15868), .ZN(n16023) );
  AOI22_X1 U18948 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15873) );
  AOI22_X1 U18949 ( .A1(n15871), .A2(n15870), .B1(n15894), .B2(n15869), .ZN(
        n15872) );
  OAI211_X1 U18950 ( .C1(n16023), .C2(n19920), .A(n15873), .B(n15872), .ZN(
        P1_U2987) );
  AOI22_X1 U18951 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15881) );
  OR3_X1 U18952 ( .A1(n14661), .A2(n15874), .A3(n14690), .ZN(n15875) );
  NAND2_X1 U18953 ( .A1(n15876), .A2(n15875), .ZN(n15878) );
  XNOR2_X1 U18954 ( .A(n15878), .B(n15877), .ZN(n16031) );
  AOI22_X1 U18955 ( .A1(n20070), .A2(n16031), .B1(n15894), .B2(n15879), .ZN(
        n15880) );
  OAI211_X1 U18956 ( .C1(n15899), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        P1_U2988) );
  AOI22_X1 U18957 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15889) );
  XNOR2_X1 U18958 ( .A(n15884), .B(n15883), .ZN(n15885) );
  XNOR2_X1 U18959 ( .A(n15886), .B(n15885), .ZN(n16060) );
  INV_X1 U18960 ( .A(n19945), .ZN(n15887) );
  AOI22_X1 U18961 ( .A1(n16060), .A2(n20070), .B1(n15894), .B2(n15887), .ZN(
        n15888) );
  OAI211_X1 U18962 ( .C1(n15899), .C2(n19950), .A(n15889), .B(n15888), .ZN(
        P1_U2992) );
  AOI22_X1 U18963 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20074), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15896) );
  NAND2_X1 U18964 ( .A1(n15891), .A2(n15890), .ZN(n15892) );
  XNOR2_X1 U18965 ( .A(n15893), .B(n15892), .ZN(n16065) );
  AOI22_X1 U18966 ( .A1(n16065), .A2(n20070), .B1(n19957), .B2(n15894), .ZN(
        n15895) );
  OAI211_X1 U18967 ( .C1(n15899), .C2(n19953), .A(n15896), .B(n15895), .ZN(
        P1_U2993) );
  XOR2_X1 U18968 ( .A(n15898), .B(n15897), .Z(n16069) );
  OAI22_X1 U18969 ( .A1(n19971), .A2(n20104), .B1(n19970), .B2(n15899), .ZN(
        n15900) );
  AOI21_X1 U18970 ( .B1(n16069), .B2(n20070), .A(n15900), .ZN(n15901) );
  NAND2_X1 U18971 ( .A1(n20074), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16077) );
  OAI211_X1 U18972 ( .C1(n19964), .C2(n15902), .A(n15901), .B(n16077), .ZN(
        P1_U2994) );
  OAI21_X1 U18973 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n15918), .ZN(n15903) );
  INV_X1 U18974 ( .A(n15903), .ZN(n15905) );
  AOI22_X1 U18975 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20074), .B1(n15905), 
        .B2(n15904), .ZN(n15910) );
  INV_X1 U18976 ( .A(n15908), .ZN(n15909) );
  OAI211_X1 U18977 ( .C1(n16079), .C2(n15911), .A(n15910), .B(n15909), .ZN(
        P1_U3003) );
  INV_X1 U18978 ( .A(n15912), .ZN(n15914) );
  AOI22_X1 U18979 ( .A1(n15914), .A2(n20090), .B1(n20089), .B2(n15913), .ZN(
        n15921) );
  NOR2_X1 U18980 ( .A1(n16057), .A2(n15915), .ZN(n15916) );
  AOI221_X1 U18981 ( .B1(n15919), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n15918), .C2(n15917), .A(n15916), .ZN(n15920) );
  NAND2_X1 U18982 ( .A1(n15921), .A2(n15920), .ZN(P1_U3004) );
  AOI22_X1 U18983 ( .A1(n15922), .A2(n20090), .B1(n20074), .B2(
        P1_REIP_REG_26__SCAN_IN), .ZN(n15927) );
  NOR3_X1 U18984 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15923), .A3(
        n15957), .ZN(n15933) );
  OAI22_X1 U18985 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15925), .B1(
        n15933), .B2(n15924), .ZN(n15926) );
  OAI211_X1 U18986 ( .C1(n16079), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P1_U3005) );
  INV_X1 U18987 ( .A(n15929), .ZN(n15931) );
  NOR2_X1 U18988 ( .A1(n16057), .A2(n15932), .ZN(n15934) );
  AOI211_X1 U18989 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15935), .A(
        n15934), .B(n15933), .ZN(n15936) );
  NAND2_X1 U18990 ( .A1(n15937), .A2(n15936), .ZN(P1_U3006) );
  NOR3_X1 U18991 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15950), .A3(
        n15957), .ZN(n15944) );
  INV_X1 U18992 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15942) );
  INV_X1 U18993 ( .A(n15938), .ZN(n20083) );
  AOI21_X1 U18994 ( .B1(n20083), .B2(n15950), .A(n15939), .ZN(n15941) );
  OAI22_X1 U18995 ( .A1(n16057), .A2(n15942), .B1(n15941), .B2(n15940), .ZN(
        n15943) );
  AOI211_X1 U18996 ( .C1(n15945), .C2(n20090), .A(n15944), .B(n15943), .ZN(
        n15946) );
  OAI21_X1 U18997 ( .B1(n16079), .B2(n15947), .A(n15946), .ZN(P1_U3007) );
  OAI22_X1 U18998 ( .A1(n15950), .A2(n15949), .B1(n16057), .B2(n15948), .ZN(
        n15951) );
  INV_X1 U18999 ( .A(n15951), .ZN(n15956) );
  INV_X1 U19000 ( .A(n15952), .ZN(n15954) );
  AOI22_X1 U19001 ( .A1(n15954), .A2(n20090), .B1(n20089), .B2(n15953), .ZN(
        n15955) );
  OAI211_X1 U19002 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15957), .A(
        n15956), .B(n15955), .ZN(P1_U3008) );
  AOI22_X1 U19003 ( .A1(n15959), .A2(n20090), .B1(n20089), .B2(n15958), .ZN(
        n15963) );
  OAI211_X1 U19004 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15961), .B(n15960), .ZN(
        n15962) );
  NAND3_X1 U19005 ( .A1(n15964), .A2(n15963), .A3(n15962), .ZN(P1_U3009) );
  AOI22_X1 U19006 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15965), .B1(
        n20074), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19007 ( .A1(n15967), .A2(n20090), .B1(n20089), .B2(n15966), .ZN(
        n15968) );
  OAI211_X1 U19008 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15970), .A(
        n15969), .B(n15968), .ZN(P1_U3012) );
  NAND2_X1 U19009 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15971), .ZN(
        n16005) );
  AOI21_X1 U19010 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15972), .A(
        n20079), .ZN(n15974) );
  AOI211_X1 U19011 ( .C1(n20075), .C2(n16005), .A(n15974), .B(n15973), .ZN(
        n16018) );
  OAI21_X1 U19012 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16048), .A(
        n16018), .ZN(n16000) );
  AOI21_X1 U19013 ( .B1(n16049), .B2(n15975), .A(n16000), .ZN(n15991) );
  NOR2_X1 U19014 ( .A1(n16057), .A2(n20685), .ZN(n15979) );
  OAI22_X1 U19015 ( .A1(n15977), .A2(n16073), .B1(n16079), .B2(n15976), .ZN(
        n15978) );
  AOI211_X1 U19016 ( .C1(n15980), .C2(n15982), .A(n15979), .B(n15978), .ZN(
        n15981) );
  OAI21_X1 U19017 ( .B1(n15991), .B2(n15982), .A(n15981), .ZN(P1_U3013) );
  NOR2_X1 U19018 ( .A1(n12395), .A2(n15983), .ZN(n15985) );
  INV_X1 U19019 ( .A(n15995), .ZN(n15984) );
  AOI21_X1 U19020 ( .B1(n15985), .B2(n15984), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15990) );
  AOI22_X1 U19021 ( .A1(n15987), .A2(n20090), .B1(n20089), .B2(n15986), .ZN(
        n15989) );
  NAND2_X1 U19022 ( .A1(n20074), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15988) );
  OAI211_X1 U19023 ( .C1(n15991), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        P1_U3014) );
  NOR3_X1 U19024 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n12395), .A3(
        n15995), .ZN(n15993) );
  NOR2_X1 U19025 ( .A1(n16057), .A2(n20681), .ZN(n15992) );
  AOI211_X1 U19026 ( .C1(n15994), .C2(n20090), .A(n15993), .B(n15992), .ZN(
        n15997) );
  NOR2_X1 U19027 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15995), .ZN(
        n15999) );
  OAI21_X1 U19028 ( .B1(n15999), .B2(n16000), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15996) );
  OAI211_X1 U19029 ( .C1(n16079), .C2(n15998), .A(n15997), .B(n15996), .ZN(
        P1_U3015) );
  AOI21_X1 U19030 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n20074), .A(n15999), 
        .ZN(n16003) );
  AOI22_X1 U19031 ( .A1(n16001), .A2(n20090), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16000), .ZN(n16002) );
  OAI211_X1 U19032 ( .C1(n16079), .C2(n16004), .A(n16003), .B(n16002), .ZN(
        P1_U3016) );
  NOR2_X1 U19033 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16005), .ZN(
        n16009) );
  OAI22_X1 U19034 ( .A1(n16007), .A2(n16073), .B1(n16079), .B2(n16006), .ZN(
        n16008) );
  AOI21_X1 U19035 ( .B1(n16009), .B2(n16036), .A(n16008), .ZN(n16011) );
  NAND2_X1 U19036 ( .A1(n20074), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16010) );
  OAI211_X1 U19037 ( .C1(n16018), .C2(n12466), .A(n16011), .B(n16010), .ZN(
        P1_U3017) );
  NOR2_X1 U19038 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16012), .ZN(
        n16017) );
  AOI22_X1 U19039 ( .A1(n16014), .A2(n20090), .B1(n20089), .B2(n16013), .ZN(
        n16016) );
  NAND2_X1 U19040 ( .A1(n20074), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16015) );
  OAI211_X1 U19041 ( .C1(n16018), .C2(n16017), .A(n16016), .B(n16015), .ZN(
        P1_U3018) );
  NOR3_X1 U19042 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15877), .A3(
        n16035), .ZN(n16025) );
  OAI21_X1 U19043 ( .B1(n15877), .B2(n16035), .A(n20075), .ZN(n16019) );
  OAI211_X1 U19044 ( .C1(n20079), .C2(n16020), .A(n20078), .B(n16019), .ZN(
        n16030) );
  AOI21_X1 U19045 ( .B1(n20083), .B2(n15877), .A(n16030), .ZN(n16022) );
  OAI22_X1 U19046 ( .A1(n16023), .A2(n16073), .B1(n16022), .B2(n16021), .ZN(
        n16024) );
  AOI21_X1 U19047 ( .B1(n16025), .B2(n16036), .A(n16024), .ZN(n16027) );
  NAND2_X1 U19048 ( .A1(n20074), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16026) );
  OAI211_X1 U19049 ( .C1(n16079), .C2(n16028), .A(n16027), .B(n16026), .ZN(
        P1_U3019) );
  NAND2_X1 U19050 ( .A1(n15877), .A2(n16036), .ZN(n16034) );
  AOI22_X1 U19051 ( .A1(n20074), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20089), 
        .B2(n16029), .ZN(n16033) );
  AOI22_X1 U19052 ( .A1(n16031), .A2(n20090), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16030), .ZN(n16032) );
  OAI211_X1 U19053 ( .C1(n16035), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        P1_U3020) );
  OAI211_X1 U19054 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16037), .B(n16036), .ZN(n16044) );
  OAI22_X1 U19055 ( .A1(n16057), .A2(n20671), .B1(n16079), .B2(n16038), .ZN(
        n16039) );
  INV_X1 U19056 ( .A(n16039), .ZN(n16043) );
  AOI22_X1 U19057 ( .A1(n16041), .A2(n20090), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16040), .ZN(n16042) );
  OAI211_X1 U19058 ( .C1(n16045), .C2(n16044), .A(n16043), .B(n16042), .ZN(
        P1_U3021) );
  INV_X1 U19059 ( .A(n16046), .ZN(n16047) );
  OAI21_X1 U19060 ( .B1(n16048), .B2(n16064), .A(n16047), .ZN(n16076) );
  AOI21_X1 U19061 ( .B1(n16050), .B2(n16049), .A(n16076), .ZN(n16062) );
  OAI22_X1 U19062 ( .A1(n16051), .A2(n16079), .B1(n20669), .B2(n16057), .ZN(
        n16053) );
  NAND3_X1 U19063 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16064), .A3(
        n16070), .ZN(n16063) );
  AOI221_X1 U19064 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16056), .C2(n15883), .A(
        n16063), .ZN(n16052) );
  AOI211_X1 U19065 ( .C1(n16054), .C2(n20090), .A(n16053), .B(n16052), .ZN(
        n16055) );
  OAI21_X1 U19066 ( .B1(n16062), .B2(n16056), .A(n16055), .ZN(P1_U3023) );
  INV_X1 U19067 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n16058) );
  OAI22_X1 U19068 ( .A1(n16079), .A2(n19939), .B1(n16058), .B2(n16057), .ZN(
        n16059) );
  AOI21_X1 U19069 ( .B1(n16060), .B2(n20090), .A(n16059), .ZN(n16061) );
  OAI221_X1 U19070 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16063), .C1(
        n15883), .C2(n16062), .A(n16061), .ZN(P1_U3024) );
  NAND2_X1 U19071 ( .A1(n16064), .A2(n16070), .ZN(n16068) );
  AOI22_X1 U19072 ( .A1(n20074), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20089), 
        .B2(n19951), .ZN(n16067) );
  AOI22_X1 U19073 ( .A1(n16065), .A2(n20090), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16076), .ZN(n16066) );
  OAI211_X1 U19074 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16068), .A(
        n16067), .B(n16066), .ZN(P1_U3025) );
  INV_X1 U19075 ( .A(n16069), .ZN(n16074) );
  NAND2_X1 U19076 ( .A1(n16070), .A2(n12355), .ZN(n16072) );
  OAI22_X1 U19077 ( .A1(n16074), .A2(n16073), .B1(n16072), .B2(n16071), .ZN(
        n16075) );
  AOI21_X1 U19078 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16076), .A(
        n16075), .ZN(n16078) );
  OAI211_X1 U19079 ( .C1(n16079), .C2(n19966), .A(n16078), .B(n16077), .ZN(
        P1_U3026) );
  INV_X1 U19080 ( .A(n16080), .ZN(n16084) );
  NAND4_X1 U19081 ( .A1(n16084), .A2(n16083), .A3(n16082), .A4(n16081), .ZN(
        n16085) );
  OAI21_X1 U19082 ( .B1(n16087), .B2(n16086), .A(n16085), .ZN(P1_U3468) );
  AOI21_X1 U19083 ( .B1(n20479), .B2(n20654), .A(n16088), .ZN(n16094) );
  NAND4_X1 U19084 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n11673), .A4(n20654), .ZN(n16089) );
  AND2_X1 U19085 ( .A1(n16090), .A2(n16089), .ZN(n20645) );
  AOI21_X1 U19086 ( .B1(n20645), .B2(n16092), .A(n16091), .ZN(n16093) );
  AOI211_X1 U19087 ( .C1(n20643), .C2(n16095), .A(n16094), .B(n16093), .ZN(
        P1_U3162) );
  OAI21_X1 U19088 ( .B1(n16097), .B2(n20479), .A(n16096), .ZN(P1_U3466) );
  INV_X1 U19089 ( .A(n16098), .ZN(n16101) );
  INV_X1 U19090 ( .A(n16099), .ZN(n16100) );
  AOI22_X1 U19091 ( .A1(n16101), .A2(n19062), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n16100), .ZN(n16108) );
  AOI22_X1 U19092 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19038), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19045), .ZN(n16107) );
  INV_X1 U19093 ( .A(n16102), .ZN(n19083) );
  AOI22_X1 U19094 ( .A1(n16103), .A2(n19067), .B1(n18972), .B2(n19083), .ZN(
        n16106) );
  NAND4_X1 U19095 ( .A1(n12968), .A2(n16112), .A3(n16104), .A4(n19029), .ZN(
        n16105) );
  NAND4_X1 U19096 ( .A1(n16108), .A2(n16107), .A3(n16106), .A4(n16105), .ZN(
        P2_U2824) );
  AOI22_X1 U19097 ( .A1(n16109), .A2(n19062), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19038), .ZN(n16119) );
  AOI22_X1 U19098 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19045), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19055), .ZN(n16118) );
  AOI22_X1 U19099 ( .A1(n16111), .A2(n19067), .B1(n18972), .B2(n16110), .ZN(
        n16117) );
  AOI21_X1 U19100 ( .B1(n16114), .B2(n16113), .A(n16112), .ZN(n16115) );
  NAND2_X1 U19101 ( .A1(n12968), .A2(n16115), .ZN(n16116) );
  NAND4_X1 U19102 ( .A1(n16119), .A2(n16118), .A3(n16117), .A4(n16116), .ZN(
        P2_U2826) );
  AOI211_X1 U19103 ( .C1(n16122), .C2(n16121), .A(n16120), .B(n19759), .ZN(
        n16132) );
  INV_X1 U19104 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19829) );
  OAI22_X1 U19105 ( .A1(n19059), .A2(n19829), .B1(n19057), .B2(n16123), .ZN(
        n16124) );
  AOI21_X1 U19106 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19055), .A(n16124), .ZN(
        n16129) );
  OAI211_X1 U19107 ( .C1(n16127), .C2(n16126), .A(n16125), .B(n19062), .ZN(
        n16128) );
  OAI211_X1 U19108 ( .C1(n16130), .C2(n18958), .A(n16129), .B(n16128), .ZN(
        n16131) );
  AOI211_X1 U19109 ( .C1(n18972), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16134) );
  INV_X1 U19110 ( .A(n16134), .ZN(P2_U2828) );
  AOI22_X1 U19111 ( .A1(n16135), .A2(n19062), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n19045), .ZN(n16147) );
  AOI22_X1 U19112 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19055), .ZN(n16146) );
  INV_X1 U19113 ( .A(n16136), .ZN(n16137) );
  OAI22_X1 U19114 ( .A1(n16138), .A2(n18958), .B1(n16137), .B2(n19065), .ZN(
        n16139) );
  INV_X1 U19115 ( .A(n16139), .ZN(n16145) );
  AOI21_X1 U19116 ( .B1(n16142), .B2(n16141), .A(n16140), .ZN(n16143) );
  NAND2_X1 U19117 ( .A1(n12968), .A2(n16143), .ZN(n16144) );
  NAND4_X1 U19118 ( .A1(n16147), .A2(n16146), .A3(n16145), .A4(n16144), .ZN(
        P2_U2829) );
  AOI22_X1 U19119 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19038), .ZN(n16159) );
  AOI22_X1 U19120 ( .A1(n16148), .A2(n19062), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19055), .ZN(n16158) );
  INV_X1 U19121 ( .A(n16149), .ZN(n16150) );
  AOI22_X1 U19122 ( .A1(n16151), .A2(n19067), .B1(n16150), .B2(n18972), .ZN(
        n16157) );
  AOI21_X1 U19123 ( .B1(n16154), .B2(n16153), .A(n16152), .ZN(n16155) );
  NAND2_X1 U19124 ( .A1(n12968), .A2(n16155), .ZN(n16156) );
  NAND4_X1 U19125 ( .A1(n16159), .A2(n16158), .A3(n16157), .A4(n16156), .ZN(
        P2_U2830) );
  OAI22_X1 U19126 ( .A1(n16161), .A2(n18958), .B1(n19065), .B2(n16160), .ZN(
        n16162) );
  INV_X1 U19127 ( .A(n16162), .ZN(n16171) );
  AOI211_X1 U19128 ( .C1(n16165), .C2(n16164), .A(n16163), .B(n19759), .ZN(
        n16169) );
  AOI22_X1 U19129 ( .A1(n19055), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19038), .ZN(n16166) );
  OAI21_X1 U19130 ( .B1(n16167), .B2(n19024), .A(n16166), .ZN(n16168) );
  AOI211_X1 U19131 ( .C1(n19045), .C2(P2_REIP_REG_23__SCAN_IN), .A(n16169), 
        .B(n16168), .ZN(n16170) );
  NAND2_X1 U19132 ( .A1(n16171), .A2(n16170), .ZN(P2_U2832) );
  AOI22_X1 U19133 ( .A1(n14844), .A2(n16172), .B1(n12981), .B2(n19078), .ZN(
        P2_U2856) );
  INV_X1 U19134 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16176) );
  AOI22_X1 U19135 ( .A1(n16174), .A2(n19079), .B1(n14844), .B2(n16173), .ZN(
        n16175) );
  OAI21_X1 U19136 ( .B1(n14844), .B2(n16176), .A(n16175), .ZN(P2_U2863) );
  INV_X1 U19137 ( .A(n16177), .ZN(n16178) );
  AOI22_X1 U19138 ( .A1(n16179), .A2(n19079), .B1(n14844), .B2(n16178), .ZN(
        n16180) );
  OAI21_X1 U19139 ( .B1(n14844), .B2(n10821), .A(n16180), .ZN(P2_U2866) );
  INV_X1 U19140 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n18898) );
  OAI22_X1 U19141 ( .A1(n16182), .A2(n16181), .B1(n19078), .B2(n18911), .ZN(
        n16183) );
  INV_X1 U19142 ( .A(n16183), .ZN(n16184) );
  OAI21_X1 U19143 ( .B1(n14844), .B2(n18898), .A(n16184), .ZN(P2_U2868) );
  OAI21_X1 U19144 ( .B1(n13830), .B2(n16186), .A(n16185), .ZN(n16187) );
  INV_X1 U19145 ( .A(n16187), .ZN(n16192) );
  AOI22_X1 U19146 ( .A1(n16192), .A2(n19079), .B1(n14844), .B2(n18930), .ZN(
        n16188) );
  OAI21_X1 U19147 ( .B1(n14844), .B2(n10817), .A(n16188), .ZN(P2_U2870) );
  AOI22_X1 U19148 ( .A1(n16190), .A2(n16189), .B1(n19137), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16195) );
  AOI22_X1 U19149 ( .A1(n19085), .A2(BUF1_REG_17__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n16194) );
  INV_X1 U19150 ( .A(n16191), .ZN(n18929) );
  AOI22_X1 U19151 ( .A1(n16192), .A2(n19139), .B1(n19138), .B2(n18929), .ZN(
        n16193) );
  NAND3_X1 U19152 ( .A1(n16195), .A2(n16194), .A3(n16193), .ZN(P2_U2902) );
  NOR2_X1 U19153 ( .A1(n16196), .A2(n16256), .ZN(n16200) );
  OAI21_X1 U19154 ( .B1(n19229), .B2(n16198), .A(n16197), .ZN(n16199) );
  AOI211_X1 U19155 ( .C1(n16201), .C2(n19222), .A(n16200), .B(n16199), .ZN(
        n16205) );
  OAI211_X1 U19156 ( .C1(n16203), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16202), .B(n19224), .ZN(n16204) );
  OAI211_X1 U19157 ( .C1(n16207), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        P2_U2998) );
  AOI22_X1 U19158 ( .A1(n19230), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19044), .ZN(n16219) );
  NAND2_X1 U19159 ( .A1(n16288), .A2(n19239), .ZN(n16216) );
  INV_X1 U19160 ( .A(n16210), .ZN(n16211) );
  OR2_X1 U19161 ( .A1(n16212), .A2(n16211), .ZN(n16213) );
  XNOR2_X1 U19162 ( .A(n16214), .B(n16213), .ZN(n16291) );
  NAND2_X1 U19163 ( .A1(n16291), .A2(n19222), .ZN(n16215) );
  OAI211_X1 U19164 ( .C1(n16290), .C2(n19234), .A(n16216), .B(n16215), .ZN(
        n16217) );
  INV_X1 U19165 ( .A(n16217), .ZN(n16218) );
  OAI211_X1 U19166 ( .C1(n16256), .C2(n16220), .A(n16219), .B(n16218), .ZN(
        P2_U3000) );
  AOI22_X1 U19167 ( .A1(n19230), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19220), .B2(n18955), .ZN(n16227) );
  AOI22_X1 U19168 ( .A1(n16222), .A2(n19222), .B1(n19239), .B2(n16221), .ZN(
        n16226) );
  NAND2_X1 U19169 ( .A1(n19224), .A2(n16223), .ZN(n16225) );
  NAND4_X1 U19170 ( .A1(n16227), .A2(n16226), .A3(n16225), .A4(n16224), .ZN(
        P2_U3001) );
  AOI22_X1 U19171 ( .A1(n19230), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19044), .ZN(n16237) );
  OR2_X1 U19172 ( .A1(n16228), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16230) );
  NAND2_X1 U19173 ( .A1(n16230), .A2(n16229), .ZN(n16305) );
  INV_X1 U19174 ( .A(n16305), .ZN(n16235) );
  AND2_X1 U19175 ( .A1(n16233), .A2(n16232), .ZN(n16234) );
  XNOR2_X1 U19176 ( .A(n16231), .B(n16234), .ZN(n16302) );
  AOI222_X1 U19177 ( .A1(n16235), .A2(n19224), .B1(n19222), .B2(n16302), .C1(
        n19239), .C2(n18973), .ZN(n16236) );
  OAI211_X1 U19178 ( .C1(n16256), .C2(n16238), .A(n16237), .B(n16236), .ZN(
        P2_U3002) );
  AOI22_X1 U19179 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19044), .B1(n19220), 
        .B2(n16239), .ZN(n16244) );
  OAI22_X1 U19180 ( .A1(n16241), .A2(n19234), .B1(n16240), .B2(n19236), .ZN(
        n16242) );
  AOI21_X1 U19181 ( .B1(n19239), .B2(n18985), .A(n16242), .ZN(n16243) );
  OAI211_X1 U19182 ( .C1(n19229), .C2(n16245), .A(n16244), .B(n16243), .ZN(
        P2_U3003) );
  AOI22_X1 U19183 ( .A1(n19230), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19044), .ZN(n16255) );
  NAND2_X1 U19184 ( .A1(n16247), .A2(n16246), .ZN(n16250) );
  NOR2_X1 U19185 ( .A1(n16248), .A2(n9766), .ZN(n16249) );
  XNOR2_X1 U19186 ( .A(n16250), .B(n16249), .ZN(n16318) );
  INV_X1 U19187 ( .A(n16318), .ZN(n16253) );
  AOI222_X1 U19188 ( .A1(n16253), .A2(n19222), .B1(n19239), .B2(n18998), .C1(
        n19224), .C2(n16314), .ZN(n16254) );
  OAI211_X1 U19189 ( .C1(n16256), .C2(n18997), .A(n16255), .B(n16254), .ZN(
        P2_U3004) );
  AOI22_X1 U19190 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19044), .B1(n19220), 
        .B2(n16257), .ZN(n16269) );
  NAND2_X1 U19191 ( .A1(n16259), .A2(n16258), .ZN(n16264) );
  INV_X1 U19192 ( .A(n16260), .ZN(n16261) );
  AOI21_X1 U19193 ( .B1(n15104), .B2(n16262), .A(n16261), .ZN(n16263) );
  XOR2_X1 U19194 ( .A(n16264), .B(n16263), .Z(n16333) );
  INV_X1 U19195 ( .A(n16328), .ZN(n16267) );
  XOR2_X1 U19196 ( .A(n16265), .B(n16266), .Z(n16327) );
  AOI222_X1 U19197 ( .A1(n16333), .A2(n19222), .B1(n19239), .B2(n16267), .C1(
        n16327), .C2(n19224), .ZN(n16268) );
  OAI211_X1 U19198 ( .C1(n19229), .C2(n16270), .A(n16269), .B(n16268), .ZN(
        P2_U3006) );
  OR2_X1 U19199 ( .A1(n16272), .A2(n16271), .ZN(n16274) );
  NAND2_X1 U19200 ( .A1(n16274), .A2(n16273), .ZN(n19089) );
  OAI22_X1 U19201 ( .A1(n16324), .A2(n19089), .B1(n15090), .B2(n19023), .ZN(
        n16275) );
  AOI221_X1 U19202 ( .B1(n16278), .B2(n16277), .C1(n16276), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16275), .ZN(n16281) );
  AOI22_X1 U19203 ( .A1(n16279), .A2(n16313), .B1(n16312), .B2(n18949), .ZN(
        n16280) );
  OAI211_X1 U19204 ( .C1(n16282), .C2(n16317), .A(n16281), .B(n16280), .ZN(
        P2_U3031) );
  AOI211_X1 U19205 ( .C1(n10847), .C2(n16284), .A(n16283), .B(n16299), .ZN(
        n16287) );
  INV_X1 U19206 ( .A(n16285), .ZN(n19092) );
  OAI22_X1 U19207 ( .A1(n16324), .A2(n19092), .B1(n19805), .B2(n19023), .ZN(
        n16286) );
  NOR2_X1 U19208 ( .A1(n16287), .A2(n16286), .ZN(n16293) );
  INV_X1 U19209 ( .A(n16288), .ZN(n16289) );
  OAI211_X1 U19210 ( .C1(n16298), .C2(n10847), .A(n16293), .B(n16292), .ZN(
        P2_U3032) );
  AOI21_X1 U19211 ( .B1(n16296), .B2(n16295), .A(n16294), .ZN(n19095) );
  NAND2_X1 U19212 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19044), .ZN(n16297) );
  OAI221_X1 U19213 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16299), 
        .C1(n10813), .C2(n16298), .A(n16297), .ZN(n16300) );
  AOI21_X1 U19214 ( .B1(n16301), .B2(n19095), .A(n16300), .ZN(n16304) );
  AOI22_X1 U19215 ( .A1(n16302), .A2(n16334), .B1(n16312), .B2(n18973), .ZN(
        n16303) );
  OAI211_X1 U19216 ( .C1(n16330), .C2(n16305), .A(n16304), .B(n16303), .ZN(
        P2_U3034) );
  INV_X1 U19217 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19799) );
  NOR2_X1 U19218 ( .A1(n19799), .A2(n19023), .ZN(n16310) );
  XNOR2_X1 U19219 ( .A(n16307), .B(n16306), .ZN(n19103) );
  OAI22_X1 U19220 ( .A1(n16324), .A2(n19103), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16308), .ZN(n16309) );
  AOI211_X1 U19221 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16311), .A(
        n16310), .B(n16309), .ZN(n16316) );
  AOI22_X1 U19222 ( .A1(n16314), .A2(n16313), .B1(n16312), .B2(n18998), .ZN(
        n16315) );
  OAI211_X1 U19223 ( .C1(n16318), .C2(n16317), .A(n16316), .B(n16315), .ZN(
        P2_U3036) );
  INV_X1 U19224 ( .A(n16319), .ZN(n16321) );
  AOI211_X1 U19225 ( .C1(n10962), .C2(n16322), .A(n16321), .B(n16320), .ZN(
        n16326) );
  INV_X1 U19226 ( .A(n16323), .ZN(n19107) );
  OAI22_X1 U19227 ( .A1(n16324), .A2(n19107), .B1(n19796), .B2(n19023), .ZN(
        n16325) );
  NOR2_X1 U19228 ( .A1(n16326), .A2(n16325), .ZN(n16336) );
  INV_X1 U19229 ( .A(n16327), .ZN(n16331) );
  OAI22_X1 U19230 ( .A1(n16331), .A2(n16330), .B1(n16329), .B2(n16328), .ZN(
        n16332) );
  AOI21_X1 U19231 ( .B1(n16334), .B2(n16333), .A(n16332), .ZN(n16335) );
  OAI211_X1 U19232 ( .C1(n16337), .C2(n10962), .A(n16336), .B(n16335), .ZN(
        P2_U3038) );
  INV_X1 U19233 ( .A(n16342), .ZN(n19756) );
  NOR2_X1 U19234 ( .A1(n19756), .A2(n19764), .ZN(n19758) );
  AOI21_X1 U19235 ( .B1(n12960), .B2(n19853), .A(n16338), .ZN(n16347) );
  INV_X1 U19236 ( .A(n16339), .ZN(n16341) );
  AOI211_X1 U19237 ( .C1(n19900), .C2(n16341), .A(n19757), .B(n16340), .ZN(
        n16346) );
  AOI22_X1 U19238 ( .A1(n16344), .A2(n16343), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n16342), .ZN(n16345) );
  OAI211_X1 U19239 ( .C1(n19758), .C2(n16347), .A(n16346), .B(n16345), .ZN(
        P2_U3176) );
  INV_X1 U19240 ( .A(n16348), .ZN(n18625) );
  INV_X1 U19241 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18803) );
  NAND2_X1 U19242 ( .A1(n16372), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16350) );
  XNOR2_X1 U19243 ( .A(n18803), .B(n16350), .ZN(n16401) );
  INV_X1 U19244 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16567) );
  INV_X1 U19245 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17864) );
  NAND2_X1 U19246 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17772) );
  INV_X1 U19247 ( .A(n17772), .ZN(n16351) );
  NAND4_X1 U19248 ( .A1(n16351), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16746) );
  NOR2_X1 U19249 ( .A1(n17716), .A2(n17721), .ZN(n17702) );
  NAND2_X1 U19250 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17663) );
  NAND2_X1 U19251 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17629) );
  NAND2_X1 U19252 ( .A1(n17610), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17585) );
  NAND2_X1 U19253 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17586) );
  NAND2_X1 U19254 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17568), .ZN(
        n17540) );
  NAND2_X1 U19255 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17541) );
  NAND2_X1 U19256 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17530), .ZN(
        n17508) );
  NAND2_X1 U19257 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17509) );
  INV_X1 U19258 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18776) );
  NOR2_X1 U19259 ( .A1(n18776), .A2(n18132), .ZN(n16395) );
  NAND2_X1 U19260 ( .A1(n18788), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18700) );
  OR2_X1 U19261 ( .A1(n16353), .A2(n17700), .ZN(n16367) );
  XNOR2_X1 U19262 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16355) );
  NOR2_X1 U19263 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17617), .ZN(
        n16377) );
  AND2_X1 U19264 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16379), .ZN(
        n16548) );
  NAND2_X1 U19265 ( .A1(n18570), .A2(n16353), .ZN(n16354) );
  OAI211_X1 U19266 ( .C1(n16548), .C2(n18700), .A(n17868), .B(n16354), .ZN(
        n16378) );
  NOR2_X1 U19267 ( .A1(n16377), .A2(n16378), .ZN(n16368) );
  OAI22_X1 U19268 ( .A1(n16367), .A2(n16355), .B1(n16368), .B2(n16567), .ZN(
        n16356) );
  AOI211_X1 U19269 ( .C1(n17730), .C2(n16909), .A(n16395), .B(n16356), .ZN(
        n16366) );
  AOI22_X1 U19270 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17770), .B1(
        n17758), .B2(n18803), .ZN(n16362) );
  OAI21_X1 U19271 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16393), .A(
        n16358), .ZN(n16359) );
  OAI22_X1 U19272 ( .A1(n16360), .A2(n16359), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18803), .ZN(n16361) );
  NAND2_X1 U19273 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16373), .ZN(
        n16363) );
  XOR2_X1 U19274 ( .A(n18803), .B(n16363), .Z(n16399) );
  NOR2_X2 U19275 ( .A1(n18203), .A2(n16525), .ZN(n17842) );
  OAI211_X1 U19276 ( .C1(n17733), .C2(n16401), .A(n16366), .B(n16365), .ZN(
        P3_U2799) );
  XNOR2_X1 U19277 ( .A(n9887), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16570) );
  AOI22_X1 U19278 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16368), .B1(
        n16367), .B2(n9886), .ZN(n16369) );
  AOI211_X1 U19279 ( .C1(n17730), .C2(n16570), .A(n16370), .B(n16369), .ZN(
        n16375) );
  OAI22_X2 U19280 ( .A1(n17733), .A2(n18051), .B1(n17872), .B2(n18053), .ZN(
        n17766) );
  NAND2_X1 U19281 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n9707), .ZN(
        n17523) );
  NOR2_X1 U19282 ( .A1(n16372), .A2(n17733), .ZN(n16386) );
  NOR2_X1 U19283 ( .A1(n16373), .A2(n17872), .ZN(n16385) );
  NOR2_X1 U19284 ( .A1(n16386), .A2(n16385), .ZN(n16374) );
  NOR2_X1 U19285 ( .A1(n17730), .A2(n16377), .ZN(n16382) );
  OAI21_X1 U19286 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16548), .A(
        n9887), .ZN(n16584) );
  OAI221_X1 U19287 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16379), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18570), .A(n16378), .ZN(
        n16380) );
  OAI211_X1 U19288 ( .C1(n16382), .C2(n16584), .A(n16381), .B(n16380), .ZN(
        n16383) );
  AOI221_X1 U19289 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16385), 
        .C1(n16384), .C2(n16385), .A(n16383), .ZN(n16389) );
  OAI21_X1 U19290 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16387), .A(
        n16386), .ZN(n16388) );
  OAI211_X1 U19291 ( .C1(n16390), .C2(n17783), .A(n16389), .B(n16388), .ZN(
        P3_U2801) );
  OAI21_X1 U19292 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18162), .A(
        n16391), .ZN(n16397) );
  NAND2_X1 U19293 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16394) );
  NOR4_X1 U19294 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16394), .A3(
        n16393), .A4(n16392), .ZN(n16396) );
  AOI211_X1 U19295 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16397), .A(
        n16396), .B(n16395), .ZN(n16400) );
  INV_X1 U19296 ( .A(n17574), .ZN(n16404) );
  NOR2_X1 U19297 ( .A1(n17354), .A2(n16407), .ZN(n18052) );
  AOI22_X1 U19298 ( .A1(n18054), .A2(n18014), .B1(n17591), .B2(n18052), .ZN(
        n16402) );
  NAND2_X1 U19299 ( .A1(n16403), .A2(n16402), .ZN(n17942) );
  NAND2_X1 U19300 ( .A1(n16404), .A2(n17942), .ZN(n17925) );
  NOR2_X1 U19301 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17925), .ZN(
        n16405) );
  AOI22_X1 U19302 ( .A1(n18174), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n16406), 
        .B2(n16405), .ZN(n16419) );
  AOI21_X1 U19303 ( .B1(n17758), .B2(n17516), .A(n17514), .ZN(n17503) );
  NOR2_X1 U19304 ( .A1(n17504), .A2(n17503), .ZN(n17502) );
  NOR4_X1 U19305 ( .A1(n16409), .A2(n16408), .A3(n17502), .A4(n16407), .ZN(
        n16415) );
  AOI22_X1 U19306 ( .A1(n18054), .A2(n16411), .B1(n18052), .B2(n16410), .ZN(
        n16412) );
  NAND2_X1 U19307 ( .A1(n16413), .A2(n16412), .ZN(n16414) );
  OAI211_X1 U19308 ( .C1(n16415), .C2(n16414), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18132), .ZN(n16418) );
  INV_X1 U19309 ( .A(n18182), .ZN(n18165) );
  NAND4_X1 U19310 ( .A1(n17758), .A2(n18165), .A3(n17503), .A4(n17500), .ZN(
        n16417) );
  NAND3_X1 U19311 ( .A1(n17504), .A2(n17514), .A3(n18076), .ZN(n16416) );
  NAND4_X1 U19312 ( .A1(n16419), .A2(n16418), .A3(n16417), .A4(n16416), .ZN(
        P3_U2834) );
  NOR3_X1 U19313 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16421) );
  NOR4_X1 U19314 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16420) );
  NAND4_X1 U19315 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16421), .A3(n16420), .A4(
        U215), .ZN(U213) );
  INV_X1 U19316 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16509) );
  INV_X2 U19317 ( .A(U214), .ZN(n16470) );
  NOR2_X2 U19318 ( .A1(n16470), .A2(n16422), .ZN(n16473) );
  OAI222_X1 U19319 ( .A1(U212), .A2(n16509), .B1(n16472), .B2(n16423), .C1(
        U214), .C2(n16510), .ZN(U216) );
  AOI22_X1 U19320 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16469), .ZN(n16424) );
  OAI21_X1 U19321 ( .B1(n14497), .B2(n16472), .A(n16424), .ZN(U217) );
  AOI22_X1 U19322 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16469), .ZN(n16425) );
  OAI21_X1 U19323 ( .B1(n14505), .B2(n16472), .A(n16425), .ZN(U218) );
  INV_X1 U19324 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U19325 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16469), .ZN(n16426) );
  OAI21_X1 U19326 ( .B1(n16427), .B2(n16472), .A(n16426), .ZN(U219) );
  INV_X1 U19327 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20750) );
  AOI22_X1 U19328 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16469), .ZN(n16428) );
  OAI21_X1 U19329 ( .B1(n20750), .B2(n16472), .A(n16428), .ZN(U220) );
  INV_X1 U19330 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16430) );
  AOI22_X1 U19331 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16469), .ZN(n16429) );
  OAI21_X1 U19332 ( .B1(n16430), .B2(n16472), .A(n16429), .ZN(U221) );
  INV_X1 U19333 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16432) );
  AOI22_X1 U19334 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16469), .ZN(n16431) );
  OAI21_X1 U19335 ( .B1(n16432), .B2(n16472), .A(n16431), .ZN(U222) );
  INV_X1 U19336 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19337 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16469), .ZN(n16433) );
  OAI21_X1 U19338 ( .B1(n16434), .B2(n16472), .A(n16433), .ZN(U223) );
  INV_X1 U19339 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U19340 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16469), .ZN(n16435) );
  OAI21_X1 U19341 ( .B1(n16436), .B2(n16472), .A(n16435), .ZN(U224) );
  INV_X1 U19342 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16438) );
  AOI22_X1 U19343 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16469), .ZN(n16437) );
  OAI21_X1 U19344 ( .B1(n16438), .B2(n16472), .A(n16437), .ZN(U225) );
  INV_X1 U19345 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19254) );
  AOI22_X1 U19346 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16469), .ZN(n16439) );
  OAI21_X1 U19347 ( .B1(n19254), .B2(n16472), .A(n16439), .ZN(U226) );
  INV_X1 U19348 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16441) );
  AOI22_X1 U19349 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16469), .ZN(n16440) );
  OAI21_X1 U19350 ( .B1(n16441), .B2(n16472), .A(n16440), .ZN(U227) );
  INV_X1 U19351 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16443) );
  AOI22_X1 U19352 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16469), .ZN(n16442) );
  OAI21_X1 U19353 ( .B1(n16443), .B2(n16472), .A(n16442), .ZN(U228) );
  INV_X1 U19354 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U19355 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16469), .ZN(n16444) );
  OAI21_X1 U19356 ( .B1(n16445), .B2(n16472), .A(n16444), .ZN(U229) );
  INV_X1 U19357 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16447) );
  AOI22_X1 U19358 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16469), .ZN(n16446) );
  OAI21_X1 U19359 ( .B1(n16447), .B2(n16472), .A(n16446), .ZN(U230) );
  INV_X1 U19360 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16449) );
  AOI22_X1 U19361 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16469), .ZN(n16448) );
  OAI21_X1 U19362 ( .B1(n16449), .B2(n16472), .A(n16448), .ZN(U231) );
  INV_X1 U19363 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n20009) );
  AOI22_X1 U19364 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16469), .ZN(n16450) );
  OAI21_X1 U19365 ( .B1(n20009), .B2(U214), .A(n16450), .ZN(U232) );
  INV_X1 U19366 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16452) );
  AOI22_X1 U19367 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16470), .ZN(n16451) );
  OAI21_X1 U19368 ( .B1(n16452), .B2(U212), .A(n16451), .ZN(U233) );
  INV_X1 U19369 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16488) );
  AOI22_X1 U19370 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16470), .ZN(n16453) );
  OAI21_X1 U19371 ( .B1(n16488), .B2(U212), .A(n16453), .ZN(U234) );
  AOI22_X1 U19372 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16469), .ZN(n16454) );
  OAI21_X1 U19373 ( .B1(n16455), .B2(n16472), .A(n16454), .ZN(U235) );
  INV_X1 U19374 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16457) );
  AOI22_X1 U19375 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16470), .ZN(n16456) );
  OAI21_X1 U19376 ( .B1(n16457), .B2(U212), .A(n16456), .ZN(U236) );
  INV_X1 U19377 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16459) );
  AOI22_X1 U19378 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16470), .ZN(n16458) );
  OAI21_X1 U19379 ( .B1(n16459), .B2(U212), .A(n16458), .ZN(U237) );
  INV_X1 U19380 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16484) );
  AOI22_X1 U19381 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16470), .ZN(n16460) );
  OAI21_X1 U19382 ( .B1(n16484), .B2(U212), .A(n16460), .ZN(U238) );
  INV_X1 U19383 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19384 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16470), .ZN(n16461) );
  OAI21_X1 U19385 ( .B1(n16462), .B2(U212), .A(n16461), .ZN(U239) );
  INV_X1 U19386 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19387 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16470), .ZN(n16463) );
  OAI21_X1 U19388 ( .B1(n16482), .B2(U212), .A(n16463), .ZN(U240) );
  INV_X1 U19389 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16481) );
  AOI22_X1 U19390 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16470), .ZN(n16464) );
  OAI21_X1 U19391 ( .B1(n16481), .B2(U212), .A(n16464), .ZN(U241) );
  INV_X1 U19392 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19393 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16470), .ZN(n16465) );
  OAI21_X1 U19394 ( .B1(n16480), .B2(U212), .A(n16465), .ZN(U242) );
  INV_X1 U19395 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U19396 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16470), .ZN(n16466) );
  OAI21_X1 U19397 ( .B1(n16479), .B2(U212), .A(n16466), .ZN(U243) );
  INV_X1 U19398 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U19399 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16470), .ZN(n16467) );
  OAI21_X1 U19400 ( .B1(n16478), .B2(U212), .A(n16467), .ZN(U244) );
  INV_X1 U19401 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16477) );
  AOI22_X1 U19402 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16470), .ZN(n16468) );
  OAI21_X1 U19403 ( .B1(n16477), .B2(U212), .A(n16468), .ZN(U245) );
  AOI22_X1 U19404 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16469), .ZN(n16471) );
  OAI21_X1 U19405 ( .B1(n13585), .B2(n16472), .A(n16471), .ZN(U246) );
  INV_X1 U19406 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19407 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16470), .ZN(n16474) );
  OAI21_X1 U19408 ( .B1(n16475), .B2(U212), .A(n16474), .ZN(U247) );
  INV_X1 U19409 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18196) );
  AOI22_X1 U19410 ( .A1(n16507), .A2(n16475), .B1(n18196), .B2(U215), .ZN(U251) );
  OAI22_X1 U19411 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16507), .ZN(n16476) );
  INV_X1 U19412 ( .A(n16476), .ZN(U252) );
  INV_X1 U19413 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U19414 ( .A1(n16507), .A2(n16477), .B1(n18210), .B2(U215), .ZN(U253) );
  INV_X1 U19415 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U19416 ( .A1(n16507), .A2(n16478), .B1(n18215), .B2(U215), .ZN(U254) );
  INV_X1 U19417 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18221) );
  AOI22_X1 U19418 ( .A1(n16507), .A2(n16479), .B1(n18221), .B2(U215), .ZN(U255) );
  INV_X1 U19419 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18226) );
  AOI22_X1 U19420 ( .A1(n16507), .A2(n16480), .B1(n18226), .B2(U215), .ZN(U256) );
  INV_X1 U19421 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18231) );
  AOI22_X1 U19422 ( .A1(n16507), .A2(n16481), .B1(n18231), .B2(U215), .ZN(U257) );
  INV_X1 U19423 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U19424 ( .A1(n16507), .A2(n16482), .B1(n18237), .B2(U215), .ZN(U258) );
  OAI22_X1 U19425 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16496), .ZN(n16483) );
  INV_X1 U19426 ( .A(n16483), .ZN(U259) );
  INV_X1 U19427 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U19428 ( .A1(n16507), .A2(n16484), .B1(n17346), .B2(U215), .ZN(U260) );
  OAI22_X1 U19429 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16496), .ZN(n16485) );
  INV_X1 U19430 ( .A(n16485), .ZN(U261) );
  OAI22_X1 U19431 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16496), .ZN(n16486) );
  INV_X1 U19432 ( .A(n16486), .ZN(U262) );
  OAI22_X1 U19433 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16496), .ZN(n16487) );
  INV_X1 U19434 ( .A(n16487), .ZN(U263) );
  INV_X1 U19435 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U19436 ( .A1(n16507), .A2(n16488), .B1(n17329), .B2(U215), .ZN(U264) );
  OAI22_X1 U19437 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16496), .ZN(n16489) );
  INV_X1 U19438 ( .A(n16489), .ZN(U265) );
  OAI22_X1 U19439 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16496), .ZN(n16490) );
  INV_X1 U19440 ( .A(n16490), .ZN(U266) );
  OAI22_X1 U19441 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16496), .ZN(n16491) );
  INV_X1 U19442 ( .A(n16491), .ZN(U267) );
  OAI22_X1 U19443 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16507), .ZN(n16492) );
  INV_X1 U19444 ( .A(n16492), .ZN(U268) );
  OAI22_X1 U19445 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16496), .ZN(n16493) );
  INV_X1 U19446 ( .A(n16493), .ZN(U269) );
  OAI22_X1 U19447 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16507), .ZN(n16494) );
  INV_X1 U19448 ( .A(n16494), .ZN(U270) );
  OAI22_X1 U19449 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16496), .ZN(n16495) );
  INV_X1 U19450 ( .A(n16495), .ZN(U271) );
  OAI22_X1 U19451 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16496), .ZN(n16497) );
  INV_X1 U19452 ( .A(n16497), .ZN(U272) );
  OAI22_X1 U19453 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16507), .ZN(n16498) );
  INV_X1 U19454 ( .A(n16498), .ZN(U273) );
  OAI22_X1 U19455 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16507), .ZN(n16499) );
  INV_X1 U19456 ( .A(n16499), .ZN(U274) );
  OAI22_X1 U19457 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16507), .ZN(n16500) );
  INV_X1 U19458 ( .A(n16500), .ZN(U275) );
  OAI22_X1 U19459 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16507), .ZN(n16501) );
  INV_X1 U19460 ( .A(n16501), .ZN(U276) );
  OAI22_X1 U19461 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16507), .ZN(n16502) );
  INV_X1 U19462 ( .A(n16502), .ZN(U277) );
  OAI22_X1 U19463 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16507), .ZN(n16503) );
  INV_X1 U19464 ( .A(n16503), .ZN(U278) );
  OAI22_X1 U19465 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16507), .ZN(n16504) );
  INV_X1 U19466 ( .A(n16504), .ZN(U279) );
  OAI22_X1 U19467 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16507), .ZN(n16505) );
  INV_X1 U19468 ( .A(n16505), .ZN(U280) );
  OAI22_X1 U19469 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16507), .ZN(n16506) );
  INV_X1 U19470 ( .A(n16506), .ZN(U281) );
  AOI22_X1 U19471 ( .A1(n16507), .A2(n16509), .B1(n18236), .B2(U215), .ZN(U282) );
  INV_X1 U19472 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16508) );
  AOI222_X1 U19473 ( .A1(n16510), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16509), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16508), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16511) );
  INV_X2 U19474 ( .A(n16513), .ZN(n16512) );
  INV_X1 U19475 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18737) );
  INV_X1 U19476 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U19477 ( .A1(n16512), .A2(n18737), .B1(n19800), .B2(n16513), .ZN(
        U347) );
  INV_X1 U19478 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18735) );
  INV_X1 U19479 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U19480 ( .A1(n16512), .A2(n18735), .B1(n19798), .B2(n16513), .ZN(
        U348) );
  INV_X1 U19481 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18732) );
  INV_X1 U19482 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19797) );
  AOI22_X1 U19483 ( .A1(n16512), .A2(n18732), .B1(n19797), .B2(n16513), .ZN(
        U349) );
  INV_X1 U19484 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18731) );
  INV_X1 U19485 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19795) );
  AOI22_X1 U19486 ( .A1(n16512), .A2(n18731), .B1(n19795), .B2(n16513), .ZN(
        U350) );
  INV_X1 U19487 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18729) );
  INV_X1 U19488 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19793) );
  AOI22_X1 U19489 ( .A1(n16512), .A2(n18729), .B1(n19793), .B2(n16513), .ZN(
        U351) );
  INV_X1 U19490 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18726) );
  INV_X1 U19491 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19492 ( .A1(n16512), .A2(n18726), .B1(n19791), .B2(n16513), .ZN(
        U352) );
  INV_X1 U19493 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20898) );
  AOI22_X1 U19494 ( .A1(n16512), .A2(n20898), .B1(n19790), .B2(n16513), .ZN(
        U353) );
  INV_X1 U19495 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18723) );
  INV_X1 U19496 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19497 ( .A1(n16512), .A2(n18723), .B1(n19788), .B2(n16513), .ZN(
        U354) );
  INV_X1 U19498 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18778) );
  INV_X1 U19499 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19836) );
  AOI22_X1 U19500 ( .A1(n16512), .A2(n18778), .B1(n19836), .B2(n16513), .ZN(
        U355) );
  INV_X1 U19501 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18774) );
  INV_X1 U19502 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19833) );
  AOI22_X1 U19503 ( .A1(n16512), .A2(n18774), .B1(n19833), .B2(n16513), .ZN(
        U356) );
  INV_X1 U19504 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18771) );
  INV_X1 U19505 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U19506 ( .A1(n16512), .A2(n18771), .B1(n19831), .B2(n16513), .ZN(
        U357) );
  INV_X1 U19507 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18770) );
  INV_X1 U19508 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19828) );
  AOI22_X1 U19509 ( .A1(n16512), .A2(n18770), .B1(n19828), .B2(n16513), .ZN(
        U358) );
  INV_X1 U19510 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18768) );
  INV_X1 U19511 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19827) );
  AOI22_X1 U19512 ( .A1(n16512), .A2(n18768), .B1(n19827), .B2(n16513), .ZN(
        U359) );
  INV_X1 U19513 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18766) );
  INV_X1 U19514 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U19515 ( .A1(n16512), .A2(n18766), .B1(n19825), .B2(n16513), .ZN(
        U360) );
  INV_X1 U19516 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18764) );
  INV_X1 U19517 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U19518 ( .A1(n16512), .A2(n18764), .B1(n19823), .B2(n16513), .ZN(
        U361) );
  INV_X1 U19519 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18762) );
  INV_X1 U19520 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U19521 ( .A1(n16512), .A2(n18762), .B1(n19821), .B2(n16513), .ZN(
        U362) );
  INV_X1 U19522 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18760) );
  INV_X1 U19523 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U19524 ( .A1(n16512), .A2(n18760), .B1(n19819), .B2(n16513), .ZN(
        U363) );
  INV_X1 U19525 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20900) );
  INV_X1 U19526 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19817) );
  AOI22_X1 U19527 ( .A1(n16512), .A2(n20900), .B1(n19817), .B2(n16513), .ZN(
        U364) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18721) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U19530 ( .A1(n16512), .A2(n18721), .B1(n19787), .B2(n16513), .ZN(
        U365) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18756) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U19533 ( .A1(n16512), .A2(n18756), .B1(n19815), .B2(n16513), .ZN(
        U366) );
  INV_X1 U19534 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18755) );
  INV_X1 U19535 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U19536 ( .A1(n16512), .A2(n18755), .B1(n19814), .B2(n16513), .ZN(
        U367) );
  INV_X1 U19537 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18753) );
  INV_X1 U19538 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19812) );
  AOI22_X1 U19539 ( .A1(n16512), .A2(n18753), .B1(n19812), .B2(n16513), .ZN(
        U368) );
  INV_X1 U19540 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18750) );
  INV_X1 U19541 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U19542 ( .A1(n16512), .A2(n18750), .B1(n19811), .B2(n16513), .ZN(
        U369) );
  INV_X1 U19543 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18749) );
  INV_X1 U19544 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19545 ( .A1(n16512), .A2(n18749), .B1(n19809), .B2(n16513), .ZN(
        U370) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18747) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U19548 ( .A1(n16512), .A2(n18747), .B1(n19807), .B2(n16513), .ZN(
        U371) );
  INV_X1 U19549 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18744) );
  INV_X1 U19550 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U19551 ( .A1(n16512), .A2(n18744), .B1(n19806), .B2(n16513), .ZN(
        U372) );
  INV_X1 U19552 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18743) );
  INV_X1 U19553 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U19554 ( .A1(n16512), .A2(n18743), .B1(n19804), .B2(n16513), .ZN(
        U373) );
  INV_X1 U19555 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18741) );
  INV_X1 U19556 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19803) );
  AOI22_X1 U19557 ( .A1(n16512), .A2(n18741), .B1(n19803), .B2(n16513), .ZN(
        U374) );
  INV_X1 U19558 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18739) );
  INV_X1 U19559 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19801) );
  AOI22_X1 U19560 ( .A1(n16512), .A2(n18739), .B1(n19801), .B2(n16513), .ZN(
        U375) );
  INV_X1 U19561 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18719) );
  INV_X1 U19562 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19563 ( .A1(n16512), .A2(n18719), .B1(n19785), .B2(n16513), .ZN(
        U376) );
  INV_X1 U19564 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18718) );
  NAND2_X1 U19565 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18718), .ZN(n18705) );
  INV_X1 U19566 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18716) );
  AOI22_X1 U19567 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18705), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18716), .ZN(n18787) );
  AOI21_X1 U19568 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18787), .ZN(n16514) );
  INV_X1 U19569 ( .A(n16514), .ZN(P3_U2633) );
  INV_X1 U19570 ( .A(n18692), .ZN(n16519) );
  NOR2_X1 U19571 ( .A1(n16516), .A2(n16515), .ZN(n16517) );
  OAI21_X1 U19572 ( .B1(n16517), .B2(n17427), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16518) );
  OAI21_X1 U19573 ( .B1(n16520), .B2(n16519), .A(n16518), .ZN(P3_U2634) );
  AOI21_X1 U19574 ( .B1(n18716), .B2(n18718), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16521) );
  AOI22_X1 U19575 ( .A1(n18832), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16521), 
        .B2(n18849), .ZN(P3_U2635) );
  OAI21_X1 U19576 ( .B1(n18702), .B2(BS16), .A(n18787), .ZN(n18785) );
  OAI21_X1 U19577 ( .B1(n18787), .B2(n18840), .A(n18785), .ZN(P3_U2636) );
  AOI211_X1 U19578 ( .C1(n17429), .C2(n16524), .A(n16523), .B(n16522), .ZN(
        n18632) );
  NOR2_X1 U19579 ( .A1(n18632), .A2(n18688), .ZN(n18833) );
  OAI21_X1 U19580 ( .B1(n18833), .B2(n16526), .A(n16525), .ZN(P3_U2637) );
  NOR4_X1 U19581 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16530) );
  NOR4_X1 U19582 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16529) );
  NOR4_X1 U19583 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16528) );
  NOR4_X1 U19584 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16527) );
  NAND4_X1 U19585 ( .A1(n16530), .A2(n16529), .A3(n16528), .A4(n16527), .ZN(
        n16536) );
  NOR4_X1 U19586 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16534) );
  AOI211_X1 U19587 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16533) );
  NOR4_X1 U19588 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16532) );
  NOR4_X1 U19589 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16531) );
  NAND4_X1 U19590 ( .A1(n16534), .A2(n16533), .A3(n16532), .A4(n16531), .ZN(
        n16535) );
  NOR2_X1 U19591 ( .A1(n16536), .A2(n16535), .ZN(n18830) );
  INV_X1 U19592 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16538) );
  NOR3_X1 U19593 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16539) );
  OAI21_X1 U19594 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16539), .A(n18830), .ZN(
        n16537) );
  OAI21_X1 U19595 ( .B1(n18830), .B2(n16538), .A(n16537), .ZN(P3_U2638) );
  INV_X1 U19596 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18823) );
  INV_X1 U19597 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18786) );
  AOI21_X1 U19598 ( .B1(n18823), .B2(n18786), .A(n16539), .ZN(n16540) );
  INV_X1 U19599 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18780) );
  INV_X1 U19600 ( .A(n18830), .ZN(n18825) );
  AOI22_X1 U19601 ( .A1(n18830), .A2(n16540), .B1(n18780), .B2(n18825), .ZN(
        P3_U2639) );
  NAND2_X1 U19602 ( .A1(n18682), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18690) );
  INV_X1 U19603 ( .A(n18690), .ZN(n18538) );
  NAND2_X1 U19604 ( .A1(n18538), .A2(n18801), .ZN(n18684) );
  NAND4_X1 U19605 ( .A1(n18682), .A2(n18788), .A3(n18840), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18696) );
  NOR2_X1 U19606 ( .A1(n18174), .A2(n16908), .ZN(n16541) );
  AOI21_X1 U19607 ( .B1(n18624), .B2(n18623), .A(n17427), .ZN(n16543) );
  INV_X1 U19608 ( .A(n16543), .ZN(n18853) );
  INV_X1 U19609 ( .A(n16542), .ZN(n18839) );
  AOI211_X1 U19610 ( .C1(n18839), .C2(n18841), .A(n18708), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18680) );
  NAND2_X1 U19611 ( .A1(n16543), .A2(n18195), .ZN(n16547) );
  AOI211_X4 U19612 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18203), .A(n18680), .B(
        n16547), .ZN(n16886) );
  INV_X1 U19613 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18769) );
  INV_X1 U19614 ( .A(n18680), .ZN(n16544) );
  INV_X1 U19615 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18767) );
  INV_X1 U19616 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18763) );
  INV_X1 U19617 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18757) );
  INV_X1 U19618 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18745) );
  INV_X1 U19619 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18740) );
  INV_X1 U19620 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18727) );
  INV_X1 U19621 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18725) );
  INV_X1 U19622 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18722) );
  NAND2_X1 U19623 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16899) );
  OR2_X1 U19624 ( .A1(n18722), .A2(n16899), .ZN(n16874) );
  OR3_X1 U19625 ( .A1(n18727), .A2(n18725), .A3(n16874), .ZN(n16828) );
  NAND3_X1 U19626 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16780) );
  NOR2_X1 U19627 ( .A1(n16828), .A2(n16780), .ZN(n16794) );
  NAND4_X1 U19628 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16794), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16775) );
  NOR2_X1 U19629 ( .A1(n18740), .A2(n16775), .ZN(n16765) );
  NAND2_X1 U19630 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16765), .ZN(n16706) );
  NOR2_X1 U19631 ( .A1(n18745), .A2(n16706), .ZN(n16683) );
  NAND4_X1 U19632 ( .A1(n16683), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16672) );
  NAND2_X1 U19633 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16688) );
  NOR3_X1 U19634 ( .A1(n18757), .A2(n16672), .A3(n16688), .ZN(n16653) );
  NAND4_X1 U19635 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16653), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n16635) );
  NOR2_X1 U19636 ( .A1(n18763), .A2(n16635), .ZN(n16628) );
  NAND2_X1 U19637 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16628), .ZN(n16613) );
  NOR2_X1 U19638 ( .A1(n18767), .A2(n16613), .ZN(n16559) );
  NAND2_X1 U19639 ( .A1(n16900), .A2(n16559), .ZN(n16594) );
  NOR2_X1 U19640 ( .A1(n18769), .A2(n16594), .ZN(n16593) );
  NAND3_X1 U19641 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16593), .ZN(n16561) );
  NOR3_X1 U19642 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18779), .A3(n16561), 
        .ZN(n16545) );
  AOI21_X1 U19643 ( .B1(n16886), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16545), .ZN(
        n16566) );
  NAND2_X1 U19644 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18203), .ZN(n16546) );
  AOI211_X4 U19645 ( .C1(n18840), .C2(n18842), .A(n16547), .B(n16546), .ZN(
        n16897) );
  NOR3_X1 U19646 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16895) );
  NAND2_X1 U19647 ( .A1(n16895), .A2(n16882), .ZN(n16881) );
  NOR2_X1 U19648 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16881), .ZN(n16866) );
  INV_X1 U19649 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17204) );
  NAND2_X1 U19650 ( .A1(n16866), .A2(n17204), .ZN(n16855) );
  INV_X1 U19651 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16833) );
  NAND2_X1 U19652 ( .A1(n16838), .A2(n16833), .ZN(n16832) );
  INV_X1 U19653 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16804) );
  NAND2_X1 U19654 ( .A1(n16812), .A2(n16804), .ZN(n16792) );
  INV_X1 U19655 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16788) );
  NAND2_X1 U19656 ( .A1(n16791), .A2(n16788), .ZN(n16787) );
  NAND2_X1 U19657 ( .A1(n16770), .A2(n16758), .ZN(n16756) );
  NAND2_X1 U19658 ( .A1(n16749), .A2(n16743), .ZN(n16740) );
  INV_X1 U19659 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16716) );
  NAND2_X1 U19660 ( .A1(n16720), .A2(n16716), .ZN(n16715) );
  INV_X1 U19661 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16693) );
  NAND2_X1 U19662 ( .A1(n16699), .A2(n16693), .ZN(n16692) );
  INV_X1 U19663 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17019) );
  NAND2_X1 U19664 ( .A1(n16673), .A2(n17019), .ZN(n16662) );
  NAND2_X1 U19665 ( .A1(n16654), .A2(n16647), .ZN(n16646) );
  NAND2_X1 U19666 ( .A1(n16633), .A2(n16624), .ZN(n16611) );
  NOR2_X1 U19667 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16611), .ZN(n16610) );
  NAND2_X1 U19668 ( .A1(n16610), .A2(n16969), .ZN(n16603) );
  NOR2_X1 U19669 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16603), .ZN(n16588) );
  INV_X1 U19670 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16957) );
  NAND2_X1 U19671 ( .A1(n16588), .A2(n16957), .ZN(n16568) );
  NOR2_X1 U19672 ( .A1(n16919), .A2(n16568), .ZN(n16574) );
  INV_X1 U19673 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16931) );
  INV_X1 U19674 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16590) );
  INV_X1 U19675 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16614) );
  INV_X1 U19676 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17556) );
  INV_X1 U19677 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17613) );
  NAND2_X1 U19678 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17610), .ZN(
        n16558) );
  NOR2_X1 U19679 ( .A1(n17613), .A2(n16558), .ZN(n16556) );
  INV_X1 U19680 ( .A(n16556), .ZN(n16557) );
  NOR2_X1 U19681 ( .A1(n17586), .A2(n16557), .ZN(n16554) );
  NAND2_X1 U19682 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16554), .ZN(
        n16553) );
  NOR2_X1 U19683 ( .A1(n17556), .A2(n16553), .ZN(n16551) );
  NAND2_X1 U19684 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16551), .ZN(
        n17496) );
  NOR2_X1 U19685 ( .A1(n16614), .A2(n17496), .ZN(n16550) );
  NAND2_X1 U19686 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16550), .ZN(
        n16549) );
  AOI21_X1 U19687 ( .B1(n16590), .B2(n16549), .A(n16548), .ZN(n17498) );
  INV_X1 U19688 ( .A(n17498), .ZN(n16597) );
  OAI21_X1 U19689 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16550), .A(
        n16549), .ZN(n17518) );
  AOI21_X1 U19690 ( .B1(n16614), .B2(n17496), .A(n16550), .ZN(n17531) );
  INV_X1 U19691 ( .A(n17531), .ZN(n16619) );
  OAI21_X1 U19692 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16551), .A(
        n17496), .ZN(n17543) );
  AOI21_X1 U19693 ( .B1(n17556), .B2(n16553), .A(n16551), .ZN(n16552) );
  INV_X1 U19694 ( .A(n16552), .ZN(n17559) );
  OAI21_X1 U19695 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n16554), .A(
        n16553), .ZN(n17581) );
  INV_X1 U19696 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17601) );
  NOR2_X1 U19697 ( .A1(n17601), .A2(n16557), .ZN(n16555) );
  INV_X1 U19698 ( .A(n16554), .ZN(n17564) );
  OAI21_X1 U19699 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16555), .A(
        n17564), .ZN(n17588) );
  AOI22_X1 U19700 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16557), .B1(
        n16556), .B2(n17601), .ZN(n17598) );
  INV_X1 U19701 ( .A(n16558), .ZN(n17582) );
  OAI21_X1 U19702 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17582), .A(
        n16557), .ZN(n17616) );
  INV_X1 U19703 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17675) );
  NOR2_X1 U19704 ( .A1(n17864), .A2(n17662), .ZN(n17661) );
  INV_X1 U19705 ( .A(n17661), .ZN(n16747) );
  NOR2_X1 U19706 ( .A1(n17675), .A2(n16747), .ZN(n16732) );
  INV_X1 U19707 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16912) );
  NAND2_X1 U19708 ( .A1(n16732), .A2(n16912), .ZN(n16724) );
  OAI21_X1 U19709 ( .B1(n16558), .B2(n16724), .A(n16352), .ZN(n16675) );
  NAND2_X1 U19710 ( .A1(n17616), .A2(n16675), .ZN(n16674) );
  NAND2_X1 U19711 ( .A1(n17588), .A2(n16659), .ZN(n16658) );
  NAND2_X1 U19712 ( .A1(n16909), .A2(n16658), .ZN(n16649) );
  NAND2_X1 U19713 ( .A1(n17581), .A2(n16649), .ZN(n16648) );
  NAND2_X1 U19714 ( .A1(n16909), .A2(n16648), .ZN(n16639) );
  NAND2_X1 U19715 ( .A1(n17559), .A2(n16639), .ZN(n16638) );
  NAND2_X1 U19716 ( .A1(n16909), .A2(n16638), .ZN(n16627) );
  NAND2_X1 U19717 ( .A1(n17543), .A2(n16627), .ZN(n16626) );
  NAND2_X1 U19718 ( .A1(n16909), .A2(n16626), .ZN(n16618) );
  NAND2_X1 U19719 ( .A1(n16619), .A2(n16618), .ZN(n16617) );
  NAND2_X1 U19720 ( .A1(n16909), .A2(n16617), .ZN(n16605) );
  NAND2_X1 U19721 ( .A1(n17518), .A2(n16605), .ZN(n16604) );
  NAND2_X1 U19722 ( .A1(n16909), .A2(n16604), .ZN(n16596) );
  NAND2_X1 U19723 ( .A1(n16597), .A2(n16596), .ZN(n16595) );
  NAND2_X1 U19724 ( .A1(n16909), .A2(n16595), .ZN(n16583) );
  NAND2_X1 U19725 ( .A1(n16584), .A2(n16583), .ZN(n16582) );
  NOR4_X1 U19726 ( .A1(n16570), .A2(n16861), .A3(n18696), .A4(n16582), .ZN(
        n16564) );
  NAND2_X1 U19727 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n16560) );
  OR2_X1 U19728 ( .A1(n16913), .A2(n16559), .ZN(n16612) );
  NAND2_X1 U19729 ( .A1(n16923), .A2(n16612), .ZN(n16609) );
  AOI221_X1 U19730 ( .B1(n18769), .B2(n16900), .C1(n16560), .C2(n16900), .A(
        n16609), .ZN(n16587) );
  NOR2_X1 U19731 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16561), .ZN(n16572) );
  INV_X1 U19732 ( .A(n16572), .ZN(n16562) );
  AOI21_X1 U19733 ( .B1(n16587), .B2(n16562), .A(n18776), .ZN(n16563) );
  AOI211_X1 U19734 ( .C1(n16574), .C2(n16931), .A(n16564), .B(n16563), .ZN(
        n16565) );
  OAI211_X1 U19735 ( .C1(n16567), .C2(n16910), .A(n16566), .B(n16565), .ZN(
        P3_U2640) );
  NAND2_X1 U19736 ( .A1(n16897), .A2(n16568), .ZN(n16577) );
  NAND2_X1 U19737 ( .A1(n16909), .A2(n16582), .ZN(n16569) );
  XNOR2_X1 U19738 ( .A(n16570), .B(n16569), .ZN(n16573) );
  OAI22_X1 U19739 ( .A1(n16587), .A2(n18779), .B1(n9886), .B2(n16910), .ZN(
        n16571) );
  AOI211_X1 U19740 ( .C1(n16573), .C2(n16908), .A(n16572), .B(n16571), .ZN(
        n16576) );
  OAI21_X1 U19741 ( .B1(n16886), .B2(n16574), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16575) );
  INV_X1 U19742 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18773) );
  INV_X1 U19743 ( .A(n16588), .ZN(n16578) );
  AOI21_X1 U19744 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16578), .A(n16577), .ZN(
        n16581) );
  NAND2_X1 U19745 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16593), .ZN(n16579) );
  OAI22_X1 U19746 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16579), .B1(n16957), 
        .B2(n16920), .ZN(n16580) );
  AOI211_X1 U19747 ( .C1(n16887), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16581), .B(n16580), .ZN(n16586) );
  OAI211_X1 U19748 ( .C1(n16584), .C2(n16583), .A(n16908), .B(n16582), .ZN(
        n16585) );
  OAI211_X1 U19749 ( .C1(n16587), .C2(n18773), .A(n16586), .B(n16585), .ZN(
        P3_U2642) );
  INV_X1 U19750 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18772) );
  AOI211_X1 U19751 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16603), .A(n16588), .B(
        n16919), .ZN(n16592) );
  OAI22_X1 U19752 ( .A1(n16590), .A2(n16910), .B1(n16920), .B2(n16589), .ZN(
        n16591) );
  AOI211_X1 U19753 ( .C1(n16593), .C2(n18772), .A(n16592), .B(n16591), .ZN(
        n16600) );
  NOR2_X1 U19754 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16594), .ZN(n16602) );
  OAI21_X1 U19755 ( .B1(n16602), .B2(n16609), .A(P3_REIP_REG_28__SCAN_IN), 
        .ZN(n16599) );
  OAI211_X1 U19756 ( .C1(n16597), .C2(n16596), .A(n16908), .B(n16595), .ZN(
        n16598) );
  NAND3_X1 U19757 ( .A1(n16600), .A2(n16599), .A3(n16598), .ZN(P3_U2643) );
  INV_X1 U19758 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17521) );
  OAI22_X1 U19759 ( .A1(n17521), .A2(n16910), .B1(n16920), .B2(n16969), .ZN(
        n16601) );
  AOI211_X1 U19760 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16609), .A(n16602), 
        .B(n16601), .ZN(n16608) );
  OAI211_X1 U19761 ( .C1(n16610), .C2(n16969), .A(n16897), .B(n16603), .ZN(
        n16607) );
  OAI211_X1 U19762 ( .C1(n17518), .C2(n16605), .A(n16908), .B(n16604), .ZN(
        n16606) );
  NAND3_X1 U19763 ( .A1(n16608), .A2(n16607), .A3(n16606), .ZN(P3_U2644) );
  INV_X1 U19764 ( .A(n16609), .ZN(n16622) );
  AOI211_X1 U19765 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16611), .A(n16610), .B(
        n16919), .ZN(n16616) );
  OAI22_X1 U19766 ( .A1(n16614), .A2(n16910), .B1(n16613), .B2(n16612), .ZN(
        n16615) );
  AOI211_X1 U19767 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16886), .A(n16616), .B(
        n16615), .ZN(n16621) );
  OAI211_X1 U19768 ( .C1(n16619), .C2(n16618), .A(n16908), .B(n16617), .ZN(
        n16620) );
  OAI211_X1 U19769 ( .C1(n16622), .C2(n18767), .A(n16621), .B(n16620), .ZN(
        P3_U2645) );
  AOI21_X1 U19770 ( .B1(n16900), .B2(n16635), .A(n16907), .ZN(n16642) );
  OAI21_X1 U19771 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16913), .A(n16642), 
        .ZN(n16623) );
  AOI22_X1 U19772 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16887), .B1(
        P3_REIP_REG_25__SCAN_IN), .B2(n16623), .ZN(n16632) );
  XOR2_X1 U19773 ( .A(n16624), .B(n16633), .Z(n16625) );
  AOI22_X1 U19774 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16886), .B1(n16897), 
        .B2(n16625), .ZN(n16631) );
  OAI211_X1 U19775 ( .C1(n17543), .C2(n16627), .A(n16908), .B(n16626), .ZN(
        n16630) );
  INV_X1 U19776 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18765) );
  NAND3_X1 U19777 ( .A1(n16900), .A2(n16628), .A3(n18765), .ZN(n16629) );
  NAND4_X1 U19778 ( .A1(n16632), .A2(n16631), .A3(n16630), .A4(n16629), .ZN(
        P3_U2646) );
  AOI211_X1 U19779 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16646), .A(n16633), .B(
        n16919), .ZN(n16637) );
  NAND2_X1 U19780 ( .A1(n16900), .A2(n18763), .ZN(n16634) );
  OAI22_X1 U19781 ( .A1(n17556), .A2(n16910), .B1(n16635), .B2(n16634), .ZN(
        n16636) );
  AOI211_X1 U19782 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16886), .A(n16637), .B(
        n16636), .ZN(n16641) );
  OAI211_X1 U19783 ( .C1(n17559), .C2(n16639), .A(n16908), .B(n16638), .ZN(
        n16640) );
  OAI211_X1 U19784 ( .C1(n16642), .C2(n18763), .A(n16641), .B(n16640), .ZN(
        P3_U2647) );
  INV_X1 U19785 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18759) );
  INV_X1 U19786 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18758) );
  NAND2_X1 U19787 ( .A1(n16900), .A2(n16653), .ZN(n16664) );
  NOR3_X1 U19788 ( .A1(n18759), .A2(n18758), .A3(n16664), .ZN(n16645) );
  INV_X1 U19789 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18761) );
  INV_X1 U19790 ( .A(n16642), .ZN(n16644) );
  INV_X1 U19791 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17565) );
  OAI22_X1 U19792 ( .A1(n17565), .A2(n16910), .B1(n16920), .B2(n16647), .ZN(
        n16643) );
  AOI221_X1 U19793 ( .B1(n16645), .B2(n18761), .C1(n16644), .C2(
        P3_REIP_REG_23__SCAN_IN), .A(n16643), .ZN(n16652) );
  OAI211_X1 U19794 ( .C1(n16654), .C2(n16647), .A(n16897), .B(n16646), .ZN(
        n16651) );
  OAI211_X1 U19795 ( .C1(n17581), .C2(n16649), .A(n16908), .B(n16648), .ZN(
        n16650) );
  NAND3_X1 U19796 ( .A1(n16652), .A2(n16651), .A3(n16650), .ZN(P3_U2648) );
  NAND2_X1 U19797 ( .A1(n16653), .A2(n16923), .ZN(n16676) );
  NOR2_X1 U19798 ( .A1(n16900), .A2(n16907), .ZN(n16722) );
  INV_X1 U19799 ( .A(n16722), .ZN(n16921) );
  OAI21_X1 U19800 ( .B1(n18758), .B2(n16676), .A(n16921), .ZN(n16663) );
  AOI211_X1 U19801 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16662), .A(n16654), .B(
        n16919), .ZN(n16657) );
  INV_X1 U19802 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16976) );
  NAND2_X1 U19803 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n18759), .ZN(n16655) );
  OAI22_X1 U19804 ( .A1(n16920), .A2(n16976), .B1(n16664), .B2(n16655), .ZN(
        n16656) );
  AOI211_X1 U19805 ( .C1(n16887), .C2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16657), .B(n16656), .ZN(n16661) );
  OAI211_X1 U19806 ( .C1(n17588), .C2(n16659), .A(n16908), .B(n16658), .ZN(
        n16660) );
  OAI211_X1 U19807 ( .C1(n16663), .C2(n18759), .A(n16661), .B(n16660), .ZN(
        P3_U2649) );
  AOI22_X1 U19808 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16887), .B1(
        n16886), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16671) );
  OAI211_X1 U19809 ( .C1(n16673), .C2(n17019), .A(n16897), .B(n16662), .ZN(
        n16670) );
  AOI21_X1 U19810 ( .B1(n18758), .B2(n16664), .A(n16663), .ZN(n16665) );
  INV_X1 U19811 ( .A(n16665), .ZN(n16669) );
  OAI211_X1 U19812 ( .C1(n17598), .C2(n16667), .A(n16908), .B(n16666), .ZN(
        n16668) );
  NAND4_X1 U19813 ( .A1(n16671), .A2(n16670), .A3(n16669), .A4(n16668), .ZN(
        P3_U2650) );
  NOR2_X1 U19814 ( .A1(n16913), .A2(n16672), .ZN(n16702) );
  NAND2_X1 U19815 ( .A1(n16702), .A2(n18757), .ZN(n16682) );
  AOI211_X1 U19816 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16692), .A(n16673), .B(
        n16919), .ZN(n16680) );
  INV_X1 U19817 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17017) );
  OAI211_X1 U19818 ( .C1(n17616), .C2(n16675), .A(n16908), .B(n16674), .ZN(
        n16678) );
  NAND3_X1 U19819 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16921), .A3(n16676), 
        .ZN(n16677) );
  OAI211_X1 U19820 ( .C1(n17017), .C2(n16920), .A(n16678), .B(n16677), .ZN(
        n16679) );
  AOI211_X1 U19821 ( .C1(n16887), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16680), .B(n16679), .ZN(n16681) );
  OAI21_X1 U19822 ( .B1(n16688), .B2(n16682), .A(n16681), .ZN(P3_U2651) );
  INV_X1 U19823 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16696) );
  INV_X1 U19824 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18751) );
  NAND2_X1 U19825 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16707) );
  NOR2_X1 U19826 ( .A1(n18751), .A2(n16707), .ZN(n16684) );
  AND2_X1 U19827 ( .A1(n16683), .A2(n16923), .ZN(n16755) );
  AOI21_X1 U19828 ( .B1(n16684), .B2(n16755), .A(n16722), .ZN(n16714) );
  NAND2_X1 U19829 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17648), .ZN(
        n16723) );
  INV_X1 U19830 ( .A(n16723), .ZN(n16709) );
  NAND2_X1 U19831 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16709), .ZN(
        n16708) );
  INV_X1 U19832 ( .A(n16708), .ZN(n17627) );
  NAND2_X1 U19833 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17627), .ZN(
        n16697) );
  OAI21_X1 U19834 ( .B1(n16724), .B2(n16697), .A(n16352), .ZN(n16687) );
  AOI21_X1 U19835 ( .B1(n16696), .B2(n16697), .A(n17582), .ZN(n16685) );
  INV_X1 U19836 ( .A(n16685), .ZN(n17631) );
  OAI21_X1 U19837 ( .B1(n16687), .B2(n17631), .A(n16908), .ZN(n16686) );
  AOI21_X1 U19838 ( .B1(n16687), .B2(n17631), .A(n16686), .ZN(n16691) );
  OAI211_X1 U19839 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16702), .B(n16688), .ZN(n16689) );
  OAI211_X1 U19840 ( .C1(n16920), .C2(n16693), .A(n18132), .B(n16689), .ZN(
        n16690) );
  AOI211_X1 U19841 ( .C1(n16714), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16691), 
        .B(n16690), .ZN(n16695) );
  OAI211_X1 U19842 ( .C1(n16699), .C2(n16693), .A(n16897), .B(n16692), .ZN(
        n16694) );
  OAI211_X1 U19843 ( .C1(n16910), .C2(n16696), .A(n16695), .B(n16694), .ZN(
        P3_U2652) );
  OAI21_X1 U19844 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17627), .A(
        n16697), .ZN(n17638) );
  NAND2_X1 U19845 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16912), .ZN(
        n16890) );
  OAI21_X1 U19846 ( .B1(n17628), .B2(n16890), .A(n16909), .ZN(n16698) );
  XNOR2_X1 U19847 ( .A(n17638), .B(n16698), .ZN(n16705) );
  AOI211_X1 U19848 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16715), .A(n16699), .B(
        n16919), .ZN(n16700) );
  AOI21_X1 U19849 ( .B1(n16887), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16700), .ZN(n16704) );
  INV_X1 U19850 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18752) );
  OAI21_X1 U19851 ( .B1(n16920), .B2(n17060), .A(n18132), .ZN(n16701) );
  AOI221_X1 U19852 ( .B1(n16714), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16702), 
        .C2(n18752), .A(n16701), .ZN(n16703) );
  OAI211_X1 U19853 ( .C1(n18696), .C2(n16705), .A(n16704), .B(n16703), .ZN(
        P3_U2653) );
  AOI22_X1 U19854 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16887), .B1(
        n16886), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16719) );
  NOR2_X1 U19855 ( .A1(n16913), .A2(n16706), .ZN(n16744) );
  NAND2_X1 U19856 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16744), .ZN(n16731) );
  NOR2_X1 U19857 ( .A1(n16707), .A2(n16731), .ZN(n16713) );
  OAI21_X1 U19858 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16709), .A(
        n16708), .ZN(n17649) );
  OAI21_X1 U19859 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16723), .A(
        n16352), .ZN(n16711) );
  OAI21_X1 U19860 ( .B1(n17649), .B2(n16711), .A(n16908), .ZN(n16710) );
  AOI21_X1 U19861 ( .B1(n17649), .B2(n16711), .A(n16710), .ZN(n16712) );
  AOI221_X1 U19862 ( .B1(n16714), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16713), 
        .C2(n18751), .A(n16712), .ZN(n16718) );
  OAI211_X1 U19863 ( .C1(n16720), .C2(n16716), .A(n16897), .B(n16715), .ZN(
        n16717) );
  NAND4_X1 U19864 ( .A1(n16719), .A2(n16718), .A3(n18132), .A4(n16717), .ZN(
        P3_U2654) );
  INV_X1 U19865 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17089) );
  AOI211_X1 U19866 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16740), .A(n16720), .B(
        n16919), .ZN(n16721) );
  AOI211_X1 U19867 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16887), .A(
        n18174), .B(n16721), .ZN(n16730) );
  AOI21_X1 U19868 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16755), .A(n16722), 
        .ZN(n16739) );
  INV_X1 U19869 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18746) );
  NOR3_X1 U19870 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18746), .A3(n16731), 
        .ZN(n16728) );
  OAI21_X1 U19871 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16732), .A(
        n16723), .ZN(n17666) );
  INV_X1 U19872 ( .A(n17666), .ZN(n16726) );
  NAND2_X1 U19873 ( .A1(n16352), .A2(n16724), .ZN(n16725) );
  INV_X1 U19874 ( .A(n16725), .ZN(n16734) );
  AOI221_X1 U19875 ( .B1(n16726), .B2(n16734), .C1(n17666), .C2(n16725), .A(
        n18696), .ZN(n16727) );
  AOI211_X1 U19876 ( .C1(n16739), .C2(P3_REIP_REG_16__SCAN_IN), .A(n16728), 
        .B(n16727), .ZN(n16729) );
  OAI211_X1 U19877 ( .C1(n16920), .C2(n17089), .A(n16730), .B(n16729), .ZN(
        P3_U2655) );
  NAND2_X1 U19878 ( .A1(n18746), .A2(n16731), .ZN(n16738) );
  INV_X1 U19879 ( .A(n16732), .ZN(n16733) );
  OAI21_X1 U19880 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17661), .A(
        n16733), .ZN(n17671) );
  OAI21_X1 U19881 ( .B1(n16861), .B2(n16912), .A(n16908), .ZN(n16762) );
  AOI211_X1 U19882 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16909), .A(
        n17671), .B(n16762), .ZN(n16737) );
  NAND3_X1 U19883 ( .A1(n16908), .A2(n16734), .A3(n17671), .ZN(n16735) );
  OAI211_X1 U19884 ( .C1(n17675), .C2(n16910), .A(n18132), .B(n16735), .ZN(
        n16736) );
  AOI211_X1 U19885 ( .C1(n16739), .C2(n16738), .A(n16737), .B(n16736), .ZN(
        n16742) );
  OAI211_X1 U19886 ( .C1(n16749), .C2(n16743), .A(n16897), .B(n16740), .ZN(
        n16741) );
  OAI211_X1 U19887 ( .C1(n16743), .C2(n16920), .A(n16742), .B(n16741), .ZN(
        P3_U2656) );
  AOI21_X1 U19888 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16921), .A(n16744), 
        .ZN(n16754) );
  AOI22_X1 U19889 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16887), .B1(
        n16886), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16753) );
  NAND2_X1 U19890 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16745), .ZN(
        n16839) );
  NOR2_X1 U19891 ( .A1(n16746), .A2(n16839), .ZN(n17698) );
  NAND2_X1 U19892 ( .A1(n17702), .A2(n17698), .ZN(n16761) );
  INV_X1 U19893 ( .A(n16761), .ZN(n16748) );
  AOI21_X1 U19894 ( .B1(n16748), .B2(n16912), .A(n16861), .ZN(n16764) );
  OAI21_X1 U19895 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16748), .A(
        n16747), .ZN(n17689) );
  XNOR2_X1 U19896 ( .A(n16764), .B(n17689), .ZN(n16751) );
  AOI211_X1 U19897 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16756), .A(n16749), .B(
        n16919), .ZN(n16750) );
  AOI211_X1 U19898 ( .C1(n16908), .C2(n16751), .A(n18174), .B(n16750), .ZN(
        n16752) );
  OAI211_X1 U19899 ( .C1(n16755), .C2(n16754), .A(n16753), .B(n16752), .ZN(
        P3_U2657) );
  AOI21_X1 U19900 ( .B1(n16900), .B2(n16775), .A(n16907), .ZN(n16784) );
  NAND2_X1 U19901 ( .A1(n16900), .A2(n18740), .ZN(n16774) );
  INV_X1 U19902 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18742) );
  AOI21_X1 U19903 ( .B1(n16784), .B2(n16774), .A(n18742), .ZN(n16760) );
  OAI211_X1 U19904 ( .C1(n16770), .C2(n16758), .A(n16897), .B(n16756), .ZN(
        n16757) );
  OAI211_X1 U19905 ( .C1(n16920), .C2(n16758), .A(n18132), .B(n16757), .ZN(
        n16759) );
  AOI211_X1 U19906 ( .C1(n16887), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16760), .B(n16759), .ZN(n16769) );
  INV_X1 U19907 ( .A(n17698), .ZN(n16781) );
  NOR2_X1 U19908 ( .A1(n17721), .A2(n16781), .ZN(n16772) );
  OAI21_X1 U19909 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16772), .A(
        n16761), .ZN(n16763) );
  INV_X1 U19910 ( .A(n16763), .ZN(n17705) );
  INV_X1 U19911 ( .A(n16762), .ZN(n16916) );
  OAI211_X1 U19912 ( .C1(n16772), .C2(n16861), .A(n17705), .B(n16916), .ZN(
        n16768) );
  NAND3_X1 U19913 ( .A1(n16908), .A2(n16764), .A3(n16763), .ZN(n16767) );
  NAND3_X1 U19914 ( .A1(n16900), .A2(n16765), .A3(n18742), .ZN(n16766) );
  NAND4_X1 U19915 ( .A1(n16769), .A2(n16768), .A3(n16767), .A4(n16766), .ZN(
        P3_U2658) );
  AOI211_X1 U19916 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16787), .A(n16770), .B(
        n16919), .ZN(n16771) );
  AOI21_X1 U19917 ( .B1(n16887), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16771), .ZN(n16779) );
  AOI21_X1 U19918 ( .B1(n17721), .B2(n16781), .A(n16772), .ZN(n17729) );
  OAI21_X1 U19919 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16781), .A(
        n16352), .ZN(n16773) );
  XNOR2_X1 U19920 ( .A(n17729), .B(n16773), .ZN(n16777) );
  OAI22_X1 U19921 ( .A1(n16920), .A2(n17124), .B1(n16775), .B2(n16774), .ZN(
        n16776) );
  AOI211_X1 U19922 ( .C1(n16908), .C2(n16777), .A(n18174), .B(n16776), .ZN(
        n16778) );
  OAI211_X1 U19923 ( .C1(n16784), .C2(n18740), .A(n16779), .B(n16778), .ZN(
        P3_U2659) );
  INV_X1 U19924 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17737) );
  INV_X1 U19925 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18736) );
  INV_X1 U19926 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18734) );
  NOR2_X1 U19927 ( .A1(n18736), .A2(n18734), .ZN(n16799) );
  NOR2_X1 U19928 ( .A1(n16913), .A2(n16828), .ZN(n16834) );
  INV_X1 U19929 ( .A(n16834), .ZN(n16816) );
  NOR2_X1 U19930 ( .A1(n16780), .A2(n16816), .ZN(n16811) );
  AOI21_X1 U19931 ( .B1(n16799), .B2(n16811), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16785) );
  INV_X1 U19932 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17746) );
  NOR2_X1 U19933 ( .A1(n17772), .A2(n16839), .ZN(n16806) );
  NAND2_X1 U19934 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16806), .ZN(
        n16805) );
  NOR2_X1 U19935 ( .A1(n17746), .A2(n16805), .ZN(n16795) );
  AOI21_X1 U19936 ( .B1(n16795), .B2(n16912), .A(n16861), .ZN(n16782) );
  OAI21_X1 U19937 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16795), .A(
        n16781), .ZN(n17735) );
  XOR2_X1 U19938 ( .A(n16782), .B(n17735), .Z(n16783) );
  OAI22_X1 U19939 ( .A1(n16785), .A2(n16784), .B1(n18696), .B2(n16783), .ZN(
        n16786) );
  AOI211_X1 U19940 ( .C1(n16886), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18174), .B(
        n16786), .ZN(n16790) );
  OAI211_X1 U19941 ( .C1(n16791), .C2(n16788), .A(n16897), .B(n16787), .ZN(
        n16789) );
  OAI211_X1 U19942 ( .C1(n16910), .C2(n17737), .A(n16790), .B(n16789), .ZN(
        P3_U2660) );
  AOI211_X1 U19943 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16792), .A(n16791), .B(
        n16919), .ZN(n16793) );
  AOI211_X1 U19944 ( .C1(n16886), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18174), .B(
        n16793), .ZN(n16803) );
  OAI21_X1 U19945 ( .B1(n16794), .B2(n16913), .A(n16923), .ZN(n16822) );
  AOI21_X1 U19946 ( .B1(n17746), .B2(n16805), .A(n16795), .ZN(n17751) );
  INV_X1 U19947 ( .A(n16806), .ZN(n16820) );
  NOR2_X1 U19948 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16820), .ZN(
        n16808) );
  AOI21_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16808), .A(
        n16861), .ZN(n16807) );
  INV_X1 U19950 ( .A(n17751), .ZN(n16797) );
  INV_X1 U19951 ( .A(n16807), .ZN(n16796) );
  AOI221_X1 U19952 ( .B1(n17751), .B2(n16807), .C1(n16797), .C2(n16796), .A(
        n18696), .ZN(n16801) );
  INV_X1 U19953 ( .A(n16811), .ZN(n16798) );
  AOI211_X1 U19954 ( .C1(n18736), .C2(n18734), .A(n16799), .B(n16798), .ZN(
        n16800) );
  AOI211_X1 U19955 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16822), .A(n16801), 
        .B(n16800), .ZN(n16802) );
  OAI211_X1 U19956 ( .C1(n17746), .C2(n16910), .A(n16803), .B(n16802), .ZN(
        P3_U2661) );
  NOR2_X1 U19957 ( .A1(n16812), .A2(n16919), .ZN(n16819) );
  AOI22_X1 U19958 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16887), .B1(
        n16819), .B2(n16804), .ZN(n16815) );
  OAI21_X1 U19959 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16806), .A(
        n16805), .ZN(n17764) );
  OAI21_X1 U19960 ( .B1(n16808), .B2(n17764), .A(n16807), .ZN(n16809) );
  AOI221_X1 U19961 ( .B1(n16352), .B2(n16809), .C1(n17764), .C2(n16809), .A(
        n18696), .ZN(n16810) );
  AOI221_X1 U19962 ( .B1(n16811), .B2(n18734), .C1(n16822), .C2(
        P3_REIP_REG_9__SCAN_IN), .A(n16810), .ZN(n16814) );
  OAI221_X1 U19963 ( .B1(n16886), .B2(n16897), .C1(n16886), .C2(n16812), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16813) );
  NAND4_X1 U19964 ( .A1(n16815), .A2(n16814), .A3(n18132), .A4(n16813), .ZN(
        P3_U2662) );
  INV_X1 U19965 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18730) );
  INV_X1 U19966 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18728) );
  NOR4_X1 U19967 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18730), .A3(n18728), .A4(
        n16816), .ZN(n16817) );
  AOI21_X1 U19968 ( .B1(n16887), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16817), .ZN(n16826) );
  NAND2_X1 U19969 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16832), .ZN(n16818) );
  AOI22_X1 U19970 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16886), .B1(n16819), .B2(
        n16818), .ZN(n16825) );
  INV_X1 U19971 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17789) );
  NOR3_X1 U19972 ( .A1(n17864), .A2(n17787), .A3(n17789), .ZN(n16827) );
  AOI21_X1 U19973 ( .B1(n16827), .B2(n16912), .A(n16861), .ZN(n16821) );
  OAI21_X1 U19974 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16827), .A(
        n16820), .ZN(n17776) );
  XNOR2_X1 U19975 ( .A(n16821), .B(n17776), .ZN(n16823) );
  AOI22_X1 U19976 ( .A1(n16908), .A2(n16823), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n16822), .ZN(n16824) );
  NAND4_X1 U19977 ( .A1(n16826), .A2(n16825), .A3(n16824), .A4(n18132), .ZN(
        P3_U2663) );
  AOI21_X1 U19978 ( .B1(n17789), .B2(n16839), .A(n16827), .ZN(n17793) );
  OAI21_X1 U19979 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16839), .A(
        n16352), .ZN(n16840) );
  XNOR2_X1 U19980 ( .A(n17793), .B(n16840), .ZN(n16831) );
  AOI21_X1 U19981 ( .B1(n16900), .B2(n16828), .A(n16907), .ZN(n16853) );
  NAND2_X1 U19982 ( .A1(n16834), .A2(n18728), .ZN(n16843) );
  AOI21_X1 U19983 ( .B1(n16853), .B2(n16843), .A(n18730), .ZN(n16830) );
  OAI22_X1 U19984 ( .A1(n17789), .A2(n16910), .B1(n16920), .B2(n16833), .ZN(
        n16829) );
  AOI211_X1 U19985 ( .C1(n16831), .C2(n16908), .A(n16830), .B(n16829), .ZN(
        n16837) );
  OAI211_X1 U19986 ( .C1(n16838), .C2(n16833), .A(n16897), .B(n16832), .ZN(
        n16836) );
  NAND3_X1 U19987 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16834), .A3(n18730), 
        .ZN(n16835) );
  NAND4_X1 U19988 ( .A1(n16837), .A2(n18132), .A3(n16836), .A4(n16835), .ZN(
        P3_U2664) );
  AOI211_X1 U19989 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16855), .A(n16838), .B(
        n16919), .ZN(n16846) );
  NOR2_X1 U19990 ( .A1(n17864), .A2(n17799), .ZN(n16850) );
  OAI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16850), .A(
        n16839), .ZN(n16847) );
  INV_X1 U19992 ( .A(n16840), .ZN(n16841) );
  NAND3_X1 U19993 ( .A1(n16908), .A2(n16847), .A3(n16841), .ZN(n16842) );
  NAND2_X1 U19994 ( .A1(n16843), .A2(n16842), .ZN(n16845) );
  INV_X1 U19995 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17199) );
  OAI22_X1 U19996 ( .A1(n17806), .A2(n16910), .B1(n16920), .B2(n17199), .ZN(
        n16844) );
  NOR4_X1 U19997 ( .A1(n18174), .A2(n16846), .A3(n16845), .A4(n16844), .ZN(
        n16849) );
  INV_X1 U19998 ( .A(n16847), .ZN(n17803) );
  OAI211_X1 U19999 ( .C1(n16850), .C2(n16861), .A(n17803), .B(n16916), .ZN(
        n16848) );
  OAI211_X1 U20000 ( .C1(n16853), .C2(n18728), .A(n16849), .B(n16848), .ZN(
        P3_U2665) );
  NOR2_X1 U20001 ( .A1(n16913), .A2(n16874), .ZN(n16862) );
  AOI21_X1 U20002 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16862), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16852) );
  INV_X1 U20003 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20912) );
  NAND3_X1 U20004 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16859), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16858) );
  AOI21_X1 U20005 ( .B1(n20912), .B2(n16858), .A(n16850), .ZN(n17815) );
  OAI21_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16858), .A(
        n16352), .ZN(n16860) );
  XOR2_X1 U20007 ( .A(n17815), .B(n16860), .Z(n16851) );
  OAI22_X1 U20008 ( .A1(n16853), .A2(n16852), .B1(n18696), .B2(n16851), .ZN(
        n16854) );
  AOI211_X1 U20009 ( .C1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n16887), .A(
        n18174), .B(n16854), .ZN(n16857) );
  OAI211_X1 U20010 ( .C1(n16866), .C2(n17204), .A(n16897), .B(n16855), .ZN(
        n16856) );
  OAI211_X1 U20011 ( .C1(n17204), .C2(n16920), .A(n16857), .B(n16856), .ZN(
        P3_U2666) );
  AOI21_X1 U20012 ( .B1(n16900), .B2(n16874), .A(n16907), .ZN(n16878) );
  NOR2_X1 U20013 ( .A1(n17864), .A2(n17830), .ZN(n16876) );
  OAI21_X1 U20014 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16876), .A(
        n16858), .ZN(n17833) );
  INV_X1 U20015 ( .A(n17833), .ZN(n16863) );
  INV_X1 U20016 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17832) );
  NAND2_X1 U20017 ( .A1(n16859), .A2(n17832), .ZN(n17828) );
  OAI22_X1 U20018 ( .A1(n16863), .A2(n16860), .B1(n16890), .B2(n17828), .ZN(
        n16872) );
  NAND2_X1 U20019 ( .A1(n16861), .A2(n16908), .ZN(n16892) );
  INV_X1 U20020 ( .A(n16892), .ZN(n16864) );
  AOI22_X1 U20021 ( .A1(n16864), .A2(n16863), .B1(n16862), .B2(n18725), .ZN(
        n16870) );
  NOR2_X1 U20022 ( .A1(n18195), .A2(n18853), .ZN(n16906) );
  INV_X1 U20023 ( .A(n16906), .ZN(n18855) );
  AOI21_X1 U20024 ( .B1(n9694), .B2(n16865), .A(n18855), .ZN(n16868) );
  AOI211_X1 U20025 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16881), .A(n16866), .B(
        n16919), .ZN(n16867) );
  AOI211_X1 U20026 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16886), .A(n16868), .B(
        n16867), .ZN(n16869) );
  OAI211_X1 U20027 ( .C1(n17832), .C2(n16910), .A(n16870), .B(n16869), .ZN(
        n16871) );
  AOI211_X1 U20028 ( .C1(n16908), .C2(n16872), .A(n18174), .B(n16871), .ZN(
        n16873) );
  OAI21_X1 U20029 ( .B1(n16878), .B2(n18725), .A(n16873), .ZN(P3_U2667) );
  INV_X1 U20030 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16885) );
  NAND2_X1 U20031 ( .A1(n18649), .A2(n18638), .ZN(n18636) );
  AOI21_X1 U20032 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18636), .A(
        n17188), .ZN(n18793) );
  NAND2_X1 U20033 ( .A1(n16900), .A2(n16874), .ZN(n16875) );
  OAI22_X1 U20034 ( .A1(n18793), .A2(n18855), .B1(n16899), .B2(n16875), .ZN(
        n16880) );
  NAND2_X1 U20035 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16888) );
  AOI21_X1 U20036 ( .B1(n16885), .B2(n16888), .A(n16876), .ZN(n17841) );
  INV_X1 U20037 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17855) );
  OAI21_X1 U20038 ( .B1(n17855), .B2(n16890), .A(n16352), .ZN(n16889) );
  XOR2_X1 U20039 ( .A(n17841), .B(n16889), .Z(n16877) );
  OAI22_X1 U20040 ( .A1(n16878), .A2(n18722), .B1(n18696), .B2(n16877), .ZN(
        n16879) );
  AOI211_X1 U20041 ( .C1(n16886), .C2(P3_EBX_REG_3__SCAN_IN), .A(n16880), .B(
        n16879), .ZN(n16884) );
  OAI211_X1 U20042 ( .C1(n16895), .C2(n16882), .A(n16897), .B(n16881), .ZN(
        n16883) );
  OAI211_X1 U20043 ( .C1(n16910), .C2(n16885), .A(n16884), .B(n16883), .ZN(
        P3_U2668) );
  AOI22_X1 U20044 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16887), .B1(
        n16886), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20045 ( .A1(n18638), .A2(n18649), .B1(n18808), .B2(n18661), .ZN(
        n18804) );
  OAI21_X1 U20046 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16888), .ZN(n17851) );
  INV_X1 U20047 ( .A(n17851), .ZN(n16891) );
  AOI211_X1 U20048 ( .C1(n16891), .C2(n16890), .A(n18696), .B(n16889), .ZN(
        n16894) );
  INV_X1 U20049 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18720) );
  OAI22_X1 U20050 ( .A1(n18720), .A2(n16923), .B1(n17851), .B2(n16892), .ZN(
        n16893) );
  AOI211_X1 U20051 ( .C1(n16906), .C2(n18804), .A(n16894), .B(n16893), .ZN(
        n16903) );
  NOR2_X1 U20052 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16898) );
  INV_X1 U20053 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17221) );
  INV_X1 U20054 ( .A(n16895), .ZN(n16896) );
  OAI211_X1 U20055 ( .C1(n16898), .C2(n17221), .A(n16897), .B(n16896), .ZN(
        n16902) );
  OAI211_X1 U20056 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16900), .B(n16899), .ZN(n16901) );
  NAND4_X1 U20057 ( .A1(n16904), .A2(n16903), .A3(n16902), .A4(n16901), .ZN(
        P3_U2669) );
  NAND2_X1 U20058 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17222) );
  OAI21_X1 U20059 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17222), .ZN(n17231) );
  AND2_X1 U20060 ( .A1(n18661), .A2(n16905), .ZN(n18812) );
  AOI22_X1 U20061 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16907), .B1(n18812), 
        .B2(n16906), .ZN(n16918) );
  NAND2_X1 U20062 ( .A1(n16909), .A2(n16908), .ZN(n16911) );
  OAI21_X1 U20063 ( .B1(n16912), .B2(n16911), .A(n16910), .ZN(n16915) );
  INV_X1 U20064 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17230) );
  OAI22_X1 U20065 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16913), .B1(n16920), 
        .B2(n17230), .ZN(n16914) );
  AOI221_X1 U20066 ( .B1(n16916), .B2(n17864), .C1(n16915), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16914), .ZN(n16917) );
  OAI211_X1 U20067 ( .C1(n16919), .C2(n17231), .A(n16918), .B(n16917), .ZN(
        P3_U2670) );
  NAND2_X1 U20068 ( .A1(n16920), .A2(n16919), .ZN(n16922) );
  AOI22_X1 U20069 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16922), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16921), .ZN(n16925) );
  NAND3_X1 U20070 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18851), .A3(
        n16923), .ZN(n16924) );
  OAI211_X1 U20071 ( .C1(n18649), .C2(n18855), .A(n16925), .B(n16924), .ZN(
        P3_U2671) );
  NOR3_X1 U20072 ( .A1(n17017), .A2(n17045), .A3(n16926), .ZN(n16927) );
  NAND4_X1 U20073 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(n16958), .A4(n16927), .ZN(n16930) );
  NOR2_X1 U20074 ( .A1(n16931), .A2(n16930), .ZN(n16956) );
  NAND2_X1 U20075 ( .A1(n17219), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16929) );
  NAND2_X1 U20076 ( .A1(n16956), .A2(n17342), .ZN(n16928) );
  OAI22_X1 U20077 ( .A1(n16956), .A2(n16929), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16928), .ZN(P3_U2672) );
  NAND2_X1 U20078 ( .A1(n16931), .A2(n16930), .ZN(n16932) );
  NAND2_X1 U20079 ( .A1(n16932), .A2(n17219), .ZN(n16955) );
  AOI22_X1 U20080 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20081 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20082 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20083 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16933) );
  NAND4_X1 U20084 ( .A1(n16936), .A2(n16935), .A3(n16934), .A4(n16933), .ZN(
        n16943) );
  AOI22_X1 U20085 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20086 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20087 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20088 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16937), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16938) );
  NAND4_X1 U20089 ( .A1(n16941), .A2(n16940), .A3(n16939), .A4(n16938), .ZN(
        n16942) );
  NOR2_X1 U20090 ( .A1(n16943), .A2(n16942), .ZN(n16961) );
  NOR2_X1 U20091 ( .A1(n16961), .A2(n16960), .ZN(n16959) );
  AOI22_X1 U20092 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20093 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n9647), .ZN(n16946) );
  AOI22_X1 U20094 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17138), .B1(
        n17099), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20095 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17181), .ZN(n16944) );
  NAND4_X1 U20096 ( .A1(n16947), .A2(n16946), .A3(n16945), .A4(n16944), .ZN(
        n16953) );
  AOI22_X1 U20097 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U20098 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16950) );
  AOI22_X1 U20099 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17188), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20100 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9654), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17186), .ZN(n16948) );
  NAND4_X1 U20101 ( .A1(n16951), .A2(n16950), .A3(n16949), .A4(n16948), .ZN(
        n16952) );
  NOR2_X1 U20102 ( .A1(n16953), .A2(n16952), .ZN(n16954) );
  XOR2_X1 U20103 ( .A(n16959), .B(n16954), .Z(n17243) );
  OAI22_X1 U20104 ( .A1(n16956), .A2(n16955), .B1(n17243), .B2(n17219), .ZN(
        P3_U2673) );
  NAND2_X1 U20105 ( .A1(n16958), .A2(n16957), .ZN(n16964) );
  AOI21_X1 U20106 ( .B1(n16961), .B2(n16960), .A(n16959), .ZN(n17247) );
  AOI22_X1 U20107 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16962), .B1(n17247), 
        .B2(n17233), .ZN(n16963) );
  OAI21_X1 U20108 ( .B1(n16970), .B2(n16964), .A(n16963), .ZN(P3_U2674) );
  AOI21_X1 U20109 ( .B1(n16966), .B2(n16971), .A(n16965), .ZN(n17256) );
  NAND2_X1 U20110 ( .A1(n17256), .A2(n17233), .ZN(n16967) );
  OAI221_X1 U20111 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16970), .C1(n16969), 
        .C2(n16968), .A(n16967), .ZN(P3_U2676) );
  INV_X1 U20112 ( .A(n16970), .ZN(n16974) );
  AOI21_X1 U20113 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17219), .A(n16981), .ZN(
        n16973) );
  OAI21_X1 U20114 ( .B1(n16977), .B2(n16972), .A(n16971), .ZN(n17264) );
  OAI22_X1 U20115 ( .A1(n16974), .A2(n16973), .B1(n17264), .B2(n17219), .ZN(
        P3_U2677) );
  INV_X1 U20116 ( .A(n16975), .ZN(n17020) );
  NAND2_X1 U20117 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17020), .ZN(n17006) );
  NOR2_X1 U20118 ( .A1(n16976), .A2(n17006), .ZN(n16986) );
  AND2_X1 U20119 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16986), .ZN(n16992) );
  AND2_X1 U20120 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16992), .ZN(n16985) );
  AOI21_X1 U20121 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17219), .A(n16985), .ZN(
        n16980) );
  AOI21_X1 U20122 ( .B1(n16978), .B2(n16982), .A(n16977), .ZN(n17266) );
  INV_X1 U20123 ( .A(n17266), .ZN(n16979) );
  OAI22_X1 U20124 ( .A1(n16981), .A2(n16980), .B1(n16979), .B2(n17219), .ZN(
        P3_U2678) );
  AOI21_X1 U20125 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17219), .A(n16992), .ZN(
        n16984) );
  OAI21_X1 U20126 ( .B1(n16987), .B2(n16983), .A(n16982), .ZN(n17275) );
  OAI22_X1 U20127 ( .A1(n16985), .A2(n16984), .B1(n17219), .B2(n17275), .ZN(
        P3_U2679) );
  AOI21_X1 U20128 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17219), .A(n16986), .ZN(
        n16991) );
  AOI21_X1 U20129 ( .B1(n16989), .B2(n16988), .A(n16987), .ZN(n17276) );
  INV_X1 U20130 ( .A(n17276), .ZN(n16990) );
  OAI22_X1 U20131 ( .A1(n16992), .A2(n16991), .B1(n17219), .B2(n16990), .ZN(
        P3_U2680) );
  AOI22_X1 U20132 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20133 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17002) );
  INV_X1 U20134 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20135 ( .A1(n15482), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16993) );
  OAI21_X1 U20136 ( .B1(n9699), .B2(n16994), .A(n16993), .ZN(n17000) );
  AOI22_X1 U20137 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20138 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20139 ( .A1(n14111), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20140 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16995) );
  NAND4_X1 U20141 ( .A1(n16998), .A2(n16997), .A3(n16996), .A4(n16995), .ZN(
        n16999) );
  AOI211_X1 U20142 ( .C1(n16937), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17000), .B(n16999), .ZN(n17001) );
  NAND3_X1 U20143 ( .A1(n17003), .A2(n17002), .A3(n17001), .ZN(n17282) );
  INV_X1 U20144 ( .A(n17282), .ZN(n17005) );
  NAND3_X1 U20145 ( .A1(n17006), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17219), 
        .ZN(n17004) );
  OAI221_X1 U20146 ( .B1(n17006), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17219), 
        .C2(n17005), .A(n17004), .ZN(P3_U2681) );
  AOI22_X1 U20147 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20148 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20149 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20150 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17007) );
  NAND4_X1 U20151 ( .A1(n17010), .A2(n17009), .A3(n17008), .A4(n17007), .ZN(
        n17016) );
  AOI22_X1 U20152 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20153 ( .A1(n15518), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20154 ( .A1(n14111), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20155 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20156 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  NOR2_X1 U20157 ( .A1(n17016), .A2(n17015), .ZN(n17288) );
  NOR2_X1 U20158 ( .A1(n17017), .A2(n17045), .ZN(n17018) );
  NOR2_X1 U20159 ( .A1(n17233), .A2(n17018), .ZN(n17032) );
  AOI22_X1 U20160 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17032), .B1(n17020), 
        .B2(n17019), .ZN(n17021) );
  OAI21_X1 U20161 ( .B1(n17288), .B2(n17219), .A(n17021), .ZN(P3_U2682) );
  AOI22_X1 U20162 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20163 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20164 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15355), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20165 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17022) );
  NAND4_X1 U20166 ( .A1(n17025), .A2(n17024), .A3(n17023), .A4(n17022), .ZN(
        n17031) );
  AOI22_X1 U20167 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20168 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20169 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17099), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20170 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17026) );
  NAND4_X1 U20171 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17030) );
  NOR2_X1 U20172 ( .A1(n17031), .A2(n17030), .ZN(n17295) );
  OAI21_X1 U20173 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17033), .A(n17032), .ZN(
        n17034) );
  OAI21_X1 U20174 ( .B1(n17295), .B2(n17219), .A(n17034), .ZN(P3_U2683) );
  AOI22_X1 U20175 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20176 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20177 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17036) );
  AOI22_X1 U20178 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17035) );
  NAND4_X1 U20179 ( .A1(n17038), .A2(n17037), .A3(n17036), .A4(n17035), .ZN(
        n17044) );
  AOI22_X1 U20180 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20181 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17099), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20182 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20183 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17039) );
  NAND4_X1 U20184 ( .A1(n17042), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17043) );
  NOR2_X1 U20185 ( .A1(n17044), .A2(n17043), .ZN(n17301) );
  OAI21_X1 U20186 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17046), .A(n17045), .ZN(
        n17047) );
  AOI22_X1 U20187 ( .A1(n17233), .A2(n17301), .B1(n17047), .B2(n17219), .ZN(
        P3_U2684) );
  NAND2_X1 U20188 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17048), .ZN(n17062) );
  AOI22_X1 U20189 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20190 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20191 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20192 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17049) );
  NAND4_X1 U20193 ( .A1(n17052), .A2(n17051), .A3(n17050), .A4(n17049), .ZN(
        n17059) );
  AOI22_X1 U20194 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15355), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20195 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20196 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20197 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17054) );
  NAND4_X1 U20198 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17058) );
  NOR2_X1 U20199 ( .A1(n17059), .A2(n17058), .ZN(n17306) );
  NAND4_X1 U20200 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17073), .A3(n17223), 
        .A4(n17060), .ZN(n17061) );
  OAI221_X1 U20201 ( .B1(n17233), .B2(n17062), .C1(n17219), .C2(n17306), .A(
        n17061), .ZN(P3_U2685) );
  AOI22_X1 U20202 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15355), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20203 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20204 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20205 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17063) );
  NAND4_X1 U20206 ( .A1(n17066), .A2(n17065), .A3(n17064), .A4(n17063), .ZN(
        n17072) );
  AOI22_X1 U20207 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20208 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20209 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20210 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17067) );
  NAND4_X1 U20211 ( .A1(n17070), .A2(n17069), .A3(n17068), .A4(n17067), .ZN(
        n17071) );
  NOR2_X1 U20212 ( .A1(n17072), .A2(n17071), .ZN(n17311) );
  AND2_X1 U20213 ( .A1(n17073), .A2(n17223), .ZN(n17075) );
  NOR2_X1 U20214 ( .A1(n18234), .A2(n17073), .ZN(n17077) );
  NAND2_X1 U20215 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17229), .ZN(n17074) );
  OAI22_X1 U20216 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17075), .B1(n17077), 
        .B2(n17074), .ZN(n17076) );
  OAI21_X1 U20217 ( .B1(n17311), .B2(n17219), .A(n17076), .ZN(P3_U2686) );
  INV_X1 U20218 ( .A(n17077), .ZN(n17091) );
  INV_X1 U20219 ( .A(n17078), .ZN(n17108) );
  NAND2_X1 U20220 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17123), .ZN(n17090) );
  AOI22_X1 U20221 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20222 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20223 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20224 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17079) );
  NAND4_X1 U20225 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        n17088) );
  AOI22_X1 U20226 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20227 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20228 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20229 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17099), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17083) );
  NAND4_X1 U20230 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17087) );
  NOR2_X1 U20231 ( .A1(n17088), .A2(n17087), .ZN(n17317) );
  NAND2_X1 U20232 ( .A1(n17219), .A2(n17090), .ZN(n17106) );
  OAI222_X1 U20233 ( .A1(n17091), .A2(n17090), .B1(n17219), .B2(n17317), .C1(
        n17089), .C2(n17106), .ZN(P3_U2687) );
  NOR2_X1 U20234 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17123), .ZN(n17107) );
  AOI22_X1 U20235 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15517), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20236 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17092), .ZN(n17095) );
  AOI22_X1 U20237 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n9653), .ZN(n17094) );
  AOI22_X1 U20238 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17186), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17181), .ZN(n17093) );
  NAND4_X1 U20239 ( .A1(n17096), .A2(n17095), .A3(n17094), .A4(n17093), .ZN(
        n17105) );
  AOI22_X1 U20240 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20241 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9654), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n15518), .ZN(n17102) );
  AOI22_X1 U20242 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17098), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17097), .ZN(n17101) );
  AOI22_X1 U20243 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17099), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17188), .ZN(n17100) );
  NAND4_X1 U20244 ( .A1(n17103), .A2(n17102), .A3(n17101), .A4(n17100), .ZN(
        n17104) );
  NOR2_X1 U20245 ( .A1(n17105), .A2(n17104), .ZN(n17321) );
  OAI22_X1 U20246 ( .A1(n17107), .A2(n17106), .B1(n17321), .B2(n17219), .ZN(
        P3_U2688) );
  OAI21_X1 U20247 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17108), .A(n17219), .ZN(
        n17122) );
  AOI22_X1 U20248 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20249 ( .A1(n9654), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20250 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20251 ( .A1(n17110), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17111) );
  NAND4_X1 U20252 ( .A1(n17114), .A2(n17113), .A3(n17112), .A4(n17111), .ZN(
        n17121) );
  AOI22_X1 U20253 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20254 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20255 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20256 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17116) );
  NAND4_X1 U20257 ( .A1(n17119), .A2(n17118), .A3(n17117), .A4(n17116), .ZN(
        n17120) );
  NOR2_X1 U20258 ( .A1(n17121), .A2(n17120), .ZN(n17325) );
  OAI22_X1 U20259 ( .A1(n17123), .A2(n17122), .B1(n17325), .B2(n17219), .ZN(
        P3_U2689) );
  AOI21_X1 U20260 ( .B1(n17124), .B2(n17150), .A(n17233), .ZN(n17125) );
  INV_X1 U20261 ( .A(n17125), .ZN(n17136) );
  AOI22_X1 U20262 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17129) );
  AOI22_X1 U20263 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20264 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20265 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17126) );
  NAND4_X1 U20266 ( .A1(n17129), .A2(n17128), .A3(n17127), .A4(n17126), .ZN(
        n17135) );
  AOI22_X1 U20267 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20268 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20269 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20270 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17130) );
  NAND4_X1 U20271 ( .A1(n17133), .A2(n17132), .A3(n17131), .A4(n17130), .ZN(
        n17134) );
  NOR2_X1 U20272 ( .A1(n17135), .A2(n17134), .ZN(n17331) );
  OAI22_X1 U20273 ( .A1(n17137), .A2(n17136), .B1(n17331), .B2(n17219), .ZN(
        P3_U2691) );
  AOI22_X1 U20274 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20275 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20276 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17139) );
  OAI21_X1 U20277 ( .B1(n17140), .B2(n17218), .A(n17139), .ZN(n17146) );
  AOI22_X1 U20278 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17187), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20279 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20280 ( .A1(n17099), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20281 ( .A1(n9654), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17141) );
  NAND4_X1 U20282 ( .A1(n17144), .A2(n17143), .A3(n17142), .A4(n17141), .ZN(
        n17145) );
  AOI211_X1 U20283 ( .C1(n17053), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17146), .B(n17145), .ZN(n17147) );
  NAND3_X1 U20284 ( .A1(n17149), .A2(n17148), .A3(n17147), .ZN(n17335) );
  INV_X1 U20285 ( .A(n17335), .ZN(n17152) );
  OAI21_X1 U20286 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17168), .A(n17150), .ZN(
        n17151) );
  AOI22_X1 U20287 ( .A1(n17233), .A2(n17152), .B1(n17151), .B2(n17219), .ZN(
        P3_U2692) );
  OAI21_X1 U20288 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17153), .A(n17219), .ZN(
        n17167) );
  AOI22_X1 U20289 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20290 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20291 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U20292 ( .B1(n17156), .B2(n17155), .A(n17154), .ZN(n17162) );
  AOI22_X1 U20293 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9647), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20294 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15482), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20295 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20296 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17157) );
  NAND4_X1 U20297 ( .A1(n17160), .A2(n17159), .A3(n17158), .A4(n17157), .ZN(
        n17161) );
  AOI211_X1 U20298 ( .C1(n15517), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17162), .B(n17161), .ZN(n17163) );
  NAND3_X1 U20299 ( .A1(n17165), .A2(n17164), .A3(n17163), .ZN(n17338) );
  INV_X1 U20300 ( .A(n17338), .ZN(n17166) );
  OAI22_X1 U20301 ( .A1(n17168), .A2(n17167), .B1(n17166), .B2(n17219), .ZN(
        P3_U2693) );
  AOI22_X1 U20302 ( .A1(n15482), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17098), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U20303 ( .A1(n17092), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20304 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20305 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17169) );
  NAND4_X1 U20306 ( .A1(n17172), .A2(n17171), .A3(n17170), .A4(n17169), .ZN(
        n17178) );
  AOI22_X1 U20307 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20308 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9654), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20309 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20310 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17173) );
  NAND4_X1 U20311 ( .A1(n17176), .A2(n17175), .A3(n17174), .A4(n17173), .ZN(
        n17177) );
  NOR2_X1 U20312 ( .A1(n17178), .A2(n17177), .ZN(n17343) );
  OAI221_X1 U20313 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(P3_EBX_REG_8__SCAN_IN), 
        .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17195), .A(n17179), .ZN(n17180) );
  AOI22_X1 U20314 ( .A1(n17233), .A2(n17343), .B1(n17180), .B2(n17219), .ZN(
        P3_U2694) );
  AOI22_X1 U20315 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20316 ( .A1(n15482), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20317 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15355), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20318 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17182) );
  NAND4_X1 U20319 ( .A1(n17185), .A2(n17184), .A3(n17183), .A4(n17182), .ZN(
        n17194) );
  AOI22_X1 U20320 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15518), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20321 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20322 ( .A1(n15517), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9654), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20323 ( .A1(n15423), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17189) );
  NAND4_X1 U20324 ( .A1(n17192), .A2(n17191), .A3(n17190), .A4(n17189), .ZN(
        n17193) );
  NOR2_X1 U20325 ( .A1(n17194), .A2(n17193), .ZN(n17351) );
  NOR2_X1 U20326 ( .A1(n17233), .A2(n17195), .ZN(n17200) );
  NOR2_X1 U20327 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17235), .ZN(n17196) );
  AOI22_X1 U20328 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17200), .B1(n17197), .B2(
        n17196), .ZN(n17198) );
  OAI21_X1 U20329 ( .B1(n17351), .B2(n17219), .A(n17198), .ZN(P3_U2695) );
  INV_X1 U20330 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17202) );
  NOR3_X1 U20331 ( .A1(n17199), .A2(n17204), .A3(n17203), .ZN(n17207) );
  OAI21_X1 U20332 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17207), .A(n17200), .ZN(
        n17201) );
  OAI21_X1 U20333 ( .B1(n17219), .B2(n17202), .A(n17201), .ZN(P3_U2696) );
  NOR2_X1 U20334 ( .A1(n17204), .A2(n17203), .ZN(n17211) );
  OAI21_X1 U20335 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17211), .A(n17219), .ZN(
        n17206) );
  INV_X1 U20336 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17205) );
  OAI22_X1 U20337 ( .A1(n17207), .A2(n17206), .B1(n17205), .B2(n17219), .ZN(
        P3_U2697) );
  OAI21_X1 U20338 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17208), .A(n17219), .ZN(
        n17210) );
  INV_X1 U20339 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17209) );
  OAI22_X1 U20340 ( .A1(n17211), .A2(n17210), .B1(n17209), .B2(n17219), .ZN(
        P3_U2698) );
  AOI22_X1 U20341 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n17233), .B1(
        P3_EBX_REG_4__SCAN_IN), .B2(n17232), .ZN(n17215) );
  OAI211_X1 U20342 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17213), .A(n17223), .B(
        n17212), .ZN(n17214) );
  NAND2_X1 U20343 ( .A1(n17215), .A2(n17214), .ZN(P3_U2699) );
  INV_X1 U20344 ( .A(n17216), .ZN(n17224) );
  NAND2_X1 U20345 ( .A1(n17224), .A2(n17223), .ZN(n17220) );
  NAND3_X1 U20346 ( .A1(n17220), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17219), .ZN(
        n17217) );
  OAI221_X1 U20347 ( .B1(n17220), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17219), 
        .C2(n17218), .A(n17217), .ZN(P3_U2700) );
  OAI21_X1 U20348 ( .B1(n17232), .B2(n17222), .A(n17221), .ZN(n17226) );
  AOI21_X1 U20349 ( .B1(n17224), .B2(n17223), .A(n17233), .ZN(n17225) );
  AOI22_X1 U20350 ( .A1(n17226), .A2(n17225), .B1(
        P3_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n17233), .ZN(n17227) );
  INV_X1 U20351 ( .A(n17227), .ZN(P3_U2701) );
  INV_X1 U20352 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17228) );
  OAI222_X1 U20353 ( .A1(n17231), .A2(n17235), .B1(n17230), .B2(n17229), .C1(
        n17228), .C2(n17219), .ZN(P3_U2702) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17233), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17232), .ZN(n17234) );
  OAI21_X1 U20355 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17235), .A(n17234), .ZN(
        P3_U2703) );
  INV_X1 U20356 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17457) );
  INV_X1 U20357 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17450) );
  INV_X1 U20358 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17495) );
  INV_X1 U20359 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17479) );
  NAND4_X1 U20360 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_1__SCAN_IN), .ZN(n17353) );
  NAND4_X1 U20361 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_7__SCAN_IN), .A4(P3_EAX_REG_6__SCAN_IN), .ZN(n17236) );
  NOR2_X1 U20362 ( .A1(n17353), .A2(n17236), .ZN(n17357) );
  NAND2_X1 U20363 ( .A1(n17357), .A2(n17384), .ZN(n17348) );
  INV_X1 U20364 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17492) );
  INV_X1 U20365 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17490) );
  INV_X1 U20366 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17483) );
  INV_X1 U20367 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17481) );
  NOR4_X1 U20368 ( .A1(n17492), .A2(n17490), .A3(n17483), .A4(n17481), .ZN(
        n17237) );
  NAND4_X1 U20369 ( .A1(n17347), .A2(P3_EAX_REG_12__SCAN_IN), .A3(
        P3_EAX_REG_11__SCAN_IN), .A4(n17237), .ZN(n17322) );
  NOR2_X2 U20370 ( .A1(n17495), .A2(n17322), .ZN(n17318) );
  NAND2_X1 U20371 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n17281) );
  NAND4_X1 U20372 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_22__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17238)
         );
  NAND2_X1 U20373 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17278), .ZN(n17277) );
  NAND2_X1 U20374 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17272), .ZN(n17271) );
  NAND2_X1 U20375 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17270), .ZN(n17261) );
  NOR2_X2 U20376 ( .A1(n17457), .A2(n17257), .ZN(n17251) );
  NAND2_X1 U20377 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17251), .ZN(n17248) );
  INV_X1 U20378 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17460) );
  OR2_X1 U20379 ( .A1(n17248), .A2(n17460), .ZN(n17242) );
  NAND2_X2 U20380 ( .A1(n18234), .A2(n17384), .ZN(n17370) );
  NAND2_X1 U20381 ( .A1(n17370), .A2(n17248), .ZN(n17246) );
  OAI21_X1 U20382 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17352), .A(n17246), .ZN(
        n17240) );
  AOI22_X1 U20383 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17312), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17240), .ZN(n17241) );
  OAI21_X1 U20384 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17242), .A(n17241), .ZN(
        P3_U2704) );
  NOR2_X2 U20385 ( .A1(n18224), .A2(n17370), .ZN(n17313) );
  INV_X1 U20386 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18230) );
  INV_X1 U20387 ( .A(n17312), .ZN(n17287) );
  OAI22_X1 U20388 ( .A1(n17243), .A2(n17376), .B1(n18230), .B2(n17287), .ZN(
        n17244) );
  AOI21_X1 U20389 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17313), .A(n17244), .ZN(
        n17245) );
  OAI221_X1 U20390 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17248), .C1(n17460), 
        .C2(n17246), .A(n17245), .ZN(P3_U2705) );
  INV_X1 U20391 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U20392 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17313), .B1(n17381), .B2(
        n17247), .ZN(n17250) );
  OAI211_X1 U20393 ( .C1(n17251), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17370), .B(
        n17248), .ZN(n17249) );
  OAI211_X1 U20394 ( .C1(n17287), .C2(n18225), .A(n17250), .B(n17249), .ZN(
        P3_U2706) );
  AOI22_X1 U20395 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17312), .ZN(n17254) );
  AOI211_X1 U20396 ( .C1(n17457), .C2(n17257), .A(n17251), .B(n17296), .ZN(
        n17252) );
  INV_X1 U20397 ( .A(n17252), .ZN(n17253) );
  OAI211_X1 U20398 ( .C1(n17255), .C2(n17376), .A(n17254), .B(n17253), .ZN(
        P3_U2707) );
  INV_X1 U20399 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U20400 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17313), .B1(n17381), .B2(
        n17256), .ZN(n17260) );
  OAI211_X1 U20401 ( .C1(n17258), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17370), .B(
        n17257), .ZN(n17259) );
  OAI211_X1 U20402 ( .C1(n17287), .C2(n18216), .A(n17260), .B(n17259), .ZN(
        P3_U2708) );
  AOI22_X1 U20403 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17312), .ZN(n17263) );
  OAI211_X1 U20404 ( .C1(n17270), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17370), .B(
        n17261), .ZN(n17262) );
  OAI211_X1 U20405 ( .C1(n17264), .C2(n17376), .A(n17263), .B(n17262), .ZN(
        P3_U2709) );
  OAI21_X1 U20406 ( .B1(n17450), .B2(n17296), .A(n17271), .ZN(n17265) );
  INV_X1 U20407 ( .A(n17265), .ZN(n17269) );
  AOI22_X1 U20408 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17312), .ZN(n17268) );
  NAND2_X1 U20409 ( .A1(n17381), .A2(n17266), .ZN(n17267) );
  OAI211_X1 U20410 ( .C1(n17270), .C2(n17269), .A(n17268), .B(n17267), .ZN(
        P3_U2710) );
  AOI22_X1 U20411 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17312), .ZN(n17274) );
  OAI211_X1 U20412 ( .C1(n17272), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17370), .B(
        n17271), .ZN(n17273) );
  OAI211_X1 U20413 ( .C1(n17275), .C2(n17376), .A(n17274), .B(n17273), .ZN(
        P3_U2711) );
  INV_X1 U20414 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18239) );
  AOI22_X1 U20415 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17313), .B1(n17381), .B2(
        n17276), .ZN(n17280) );
  OAI211_X1 U20416 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17278), .A(n17370), .B(
        n17277), .ZN(n17279) );
  OAI211_X1 U20417 ( .C1(n17287), .C2(n18239), .A(n17280), .B(n17279), .ZN(
        P3_U2712) );
  NOR2_X1 U20418 ( .A1(n18234), .A2(n17314), .ZN(n17308) );
  NAND2_X1 U20419 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17308), .ZN(n17307) );
  NAND3_X1 U20420 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(n17297), .ZN(n17286) );
  AOI22_X1 U20421 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17312), .B1(n17381), .B2(
        n17282), .ZN(n17285) );
  NAND2_X1 U20422 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17297), .ZN(n17292) );
  NAND2_X1 U20423 ( .A1(n17370), .A2(n17292), .ZN(n17291) );
  OAI21_X1 U20424 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17352), .A(n17291), .ZN(
        n17283) );
  AOI22_X1 U20425 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17313), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17283), .ZN(n17284) );
  OAI211_X1 U20426 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17286), .A(n17285), .B(
        n17284), .ZN(P3_U2713) );
  INV_X1 U20427 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17442) );
  INV_X1 U20428 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19252) );
  OAI22_X1 U20429 ( .A1(n17288), .A2(n17376), .B1(n19252), .B2(n17287), .ZN(
        n17289) );
  AOI21_X1 U20430 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17313), .A(n17289), .ZN(
        n17290) );
  OAI221_X1 U20431 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17292), .C1(n17442), 
        .C2(n17291), .A(n17290), .ZN(P3_U2714) );
  AOI22_X1 U20432 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17312), .ZN(n17294) );
  OAI211_X1 U20433 ( .C1(n17297), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17370), .B(
        n17292), .ZN(n17293) );
  OAI211_X1 U20434 ( .C1(n17295), .C2(n17376), .A(n17294), .B(n17293), .ZN(
        P3_U2715) );
  AOI22_X1 U20435 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17312), .ZN(n17300) );
  INV_X1 U20436 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17438) );
  INV_X1 U20437 ( .A(n17307), .ZN(n17303) );
  NAND2_X1 U20438 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17303), .ZN(n17302) );
  AOI211_X1 U20439 ( .C1(n17438), .C2(n17302), .A(n17297), .B(n17296), .ZN(
        n17298) );
  INV_X1 U20440 ( .A(n17298), .ZN(n17299) );
  OAI211_X1 U20441 ( .C1(n17301), .C2(n17376), .A(n17300), .B(n17299), .ZN(
        P3_U2716) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17312), .ZN(n17305) );
  OAI211_X1 U20443 ( .C1(n17303), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17370), .B(
        n17302), .ZN(n17304) );
  OAI211_X1 U20444 ( .C1(n17306), .C2(n17376), .A(n17305), .B(n17304), .ZN(
        P3_U2717) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17312), .ZN(n17310) );
  OAI211_X1 U20446 ( .C1(n17308), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17370), .B(
        n17307), .ZN(n17309) );
  OAI211_X1 U20447 ( .C1(n17311), .C2(n17376), .A(n17310), .B(n17309), .ZN(
        P3_U2718) );
  AOI22_X1 U20448 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17313), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17312), .ZN(n17316) );
  OAI211_X1 U20449 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17318), .A(n17370), .B(
        n17314), .ZN(n17315) );
  OAI211_X1 U20450 ( .C1(n17317), .C2(n17376), .A(n17316), .B(n17315), .ZN(
        P3_U2719) );
  AOI21_X1 U20451 ( .B1(n17495), .B2(n17322), .A(n17318), .ZN(n17319) );
  AOI22_X1 U20452 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17382), .B1(n17319), .B2(
        n17370), .ZN(n17320) );
  OAI21_X1 U20453 ( .B1(n17321), .B2(n17376), .A(n17320), .ZN(P3_U2720) );
  INV_X1 U20454 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17488) );
  INV_X1 U20455 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17485) );
  NAND3_X1 U20456 ( .A1(n17342), .A2(n17347), .A3(P3_EAX_REG_9__SCAN_IN), .ZN(
        n17340) );
  INV_X1 U20457 ( .A(n17340), .ZN(n17345) );
  NAND2_X1 U20458 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17345), .ZN(n17337) );
  NOR3_X1 U20459 ( .A1(n17488), .A2(n17485), .A3(n17337), .ZN(n17333) );
  AND2_X1 U20460 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17333), .ZN(n17328) );
  AOI22_X1 U20461 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17382), .B1(n17328), .B2(
        n17492), .ZN(n17324) );
  NAND3_X1 U20462 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17370), .A3(n17322), 
        .ZN(n17323) );
  OAI211_X1 U20463 ( .C1(n17325), .C2(n17376), .A(n17324), .B(n17323), .ZN(
        P3_U2721) );
  INV_X1 U20464 ( .A(n17382), .ZN(n17379) );
  AOI21_X1 U20465 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17370), .A(n17333), .ZN(
        n17327) );
  OAI222_X1 U20466 ( .A1(n17379), .A2(n17329), .B1(n17328), .B2(n17327), .C1(
        n17376), .C2(n17326), .ZN(P3_U2722) );
  INV_X1 U20467 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17334) );
  INV_X1 U20468 ( .A(n17337), .ZN(n17330) );
  AOI22_X1 U20469 ( .A1(n17330), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17370), .ZN(n17332) );
  OAI222_X1 U20470 ( .A1(n17379), .A2(n17334), .B1(n17333), .B2(n17332), .C1(
        n17376), .C2(n17331), .ZN(P3_U2723) );
  NAND2_X1 U20471 ( .A1(n17370), .A2(n17337), .ZN(n17341) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17382), .B1(n17381), .B2(
        n17335), .ZN(n17336) );
  OAI221_X1 U20473 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17337), .C1(n17485), 
        .C2(n17341), .A(n17336), .ZN(P3_U2724) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17382), .B1(n17381), .B2(
        n17338), .ZN(n17339) );
  OAI221_X1 U20475 ( .B1(n17341), .B2(n17483), .C1(n17341), .C2(n17340), .A(
        n17339), .ZN(P3_U2725) );
  AOI22_X1 U20476 ( .A1(n17342), .A2(n17347), .B1(P3_EAX_REG_9__SCAN_IN), .B2(
        n17370), .ZN(n17344) );
  OAI222_X1 U20477 ( .A1(n17379), .A2(n17346), .B1(n17345), .B2(n17344), .C1(
        n17376), .C2(n17343), .ZN(P3_U2726) );
  AOI21_X1 U20478 ( .B1(n17479), .B2(n17348), .A(n17347), .ZN(n17349) );
  AOI22_X1 U20479 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17382), .B1(n17349), .B2(
        n17370), .ZN(n17350) );
  OAI21_X1 U20480 ( .B1(n17351), .B2(n17376), .A(n17350), .ZN(P3_U2727) );
  INV_X1 U20481 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17474) );
  NOR2_X1 U20482 ( .A1(n17353), .A2(n17388), .ZN(n17369) );
  NAND2_X1 U20483 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17369), .ZN(n17359) );
  NOR2_X1 U20484 ( .A1(n17474), .A2(n17359), .ZN(n17361) );
  AOI21_X1 U20485 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17370), .A(n17361), .ZN(
        n17358) );
  AOI22_X1 U20486 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17382), .B1(n17381), .B2(
        n17354), .ZN(n17355) );
  OAI221_X1 U20487 ( .B1(n17358), .B2(n17357), .C1(n17358), .C2(n17356), .A(
        n17355), .ZN(P3_U2728) );
  INV_X1 U20488 ( .A(n17359), .ZN(n17365) );
  AOI21_X1 U20489 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17370), .A(n17365), .ZN(
        n17362) );
  OAI222_X1 U20490 ( .A1(n17379), .A2(n18231), .B1(n17362), .B2(n17361), .C1(
        n17376), .C2(n17360), .ZN(P3_U2729) );
  AOI21_X1 U20491 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17370), .A(n17369), .ZN(
        n17364) );
  OAI222_X1 U20492 ( .A1(n18226), .A2(n17379), .B1(n17365), .B2(n17364), .C1(
        n17376), .C2(n17363), .ZN(P3_U2730) );
  INV_X1 U20493 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17466) );
  INV_X1 U20494 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17464) );
  NOR3_X1 U20495 ( .A1(n17466), .A2(n17464), .A3(n17388), .ZN(n17378) );
  AND2_X1 U20496 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17378), .ZN(n17373) );
  AOI21_X1 U20497 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17370), .A(n17373), .ZN(
        n17368) );
  INV_X1 U20498 ( .A(n17366), .ZN(n17367) );
  OAI222_X1 U20499 ( .A1(n18221), .A2(n17379), .B1(n17369), .B2(n17368), .C1(
        n17376), .C2(n17367), .ZN(P3_U2731) );
  AOI21_X1 U20500 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17370), .A(n17378), .ZN(
        n17372) );
  OAI222_X1 U20501 ( .A1(n18215), .A2(n17379), .B1(n17373), .B2(n17372), .C1(
        n17376), .C2(n17371), .ZN(P3_U2732) );
  AOI22_X1 U20502 ( .A1(n17374), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n17370), .ZN(n17377) );
  OAI222_X1 U20503 ( .A1(n18210), .A2(n17379), .B1(n17378), .B2(n17377), .C1(
        n17376), .C2(n17375), .ZN(P3_U2733) );
  AOI22_X1 U20504 ( .A1(n17382), .A2(BUF2_REG_1__SCAN_IN), .B1(n17381), .B2(
        n17380), .ZN(n17387) );
  AOI21_X1 U20505 ( .B1(n17384), .B2(n17383), .A(n17464), .ZN(n17385) );
  INV_X1 U20506 ( .A(n17385), .ZN(n17386) );
  OAI211_X1 U20507 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17388), .A(n17387), .B(
        n17386), .ZN(P3_U2734) );
  AND2_X1 U20508 ( .A1(n17416), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20509 ( .A1(n17406), .A2(n18195), .ZN(n17405) );
  AOI22_X1 U20510 ( .A1(n18838), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20511 ( .B1(n17460), .B2(n17405), .A(n17390), .ZN(P3_U2737) );
  INV_X1 U20512 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U20513 ( .A1(n18838), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20514 ( .B1(n20905), .B2(n17405), .A(n17391), .ZN(P3_U2738) );
  AOI22_X1 U20515 ( .A1(n18838), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20516 ( .B1(n17457), .B2(n17405), .A(n17392), .ZN(P3_U2739) );
  INV_X1 U20517 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20518 ( .A1(n18838), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20519 ( .B1(n17454), .B2(n17405), .A(n17393), .ZN(P3_U2740) );
  INV_X1 U20520 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20521 ( .A1(n18838), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17394) );
  OAI21_X1 U20522 ( .B1(n17452), .B2(n17405), .A(n17394), .ZN(P3_U2741) );
  AOI22_X1 U20523 ( .A1(n18838), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20524 ( .B1(n17450), .B2(n17405), .A(n17395), .ZN(P3_U2742) );
  INV_X1 U20525 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20526 ( .A1(n18838), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20527 ( .B1(n17448), .B2(n17405), .A(n17396), .ZN(P3_U2743) );
  INV_X1 U20528 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17446) );
  CLKBUF_X1 U20529 ( .A(n18838), .Z(n17424) );
  AOI22_X1 U20530 ( .A1(n17424), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17397) );
  OAI21_X1 U20531 ( .B1(n17446), .B2(n17405), .A(n17397), .ZN(P3_U2744) );
  INV_X1 U20532 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20533 ( .A1(n17424), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20534 ( .B1(n17444), .B2(n17405), .A(n17398), .ZN(P3_U2745) );
  AOI22_X1 U20535 ( .A1(n17424), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20536 ( .B1(n17442), .B2(n17405), .A(n17399), .ZN(P3_U2746) );
  INV_X1 U20537 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20538 ( .A1(n17424), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20539 ( .B1(n17440), .B2(n17405), .A(n17400), .ZN(P3_U2747) );
  AOI22_X1 U20540 ( .A1(n17424), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U20541 ( .B1(n17438), .B2(n17405), .A(n17401), .ZN(P3_U2748) );
  INV_X1 U20542 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20543 ( .A1(n17424), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20544 ( .B1(n17436), .B2(n17405), .A(n17402), .ZN(P3_U2749) );
  INV_X1 U20545 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20546 ( .A1(n17424), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20547 ( .B1(n17434), .B2(n17405), .A(n17403), .ZN(P3_U2750) );
  INV_X1 U20548 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20549 ( .A1(n17424), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20550 ( .B1(n17432), .B2(n17405), .A(n17404), .ZN(P3_U2751) );
  AOI22_X1 U20551 ( .A1(n17424), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20552 ( .B1(n17495), .B2(n17426), .A(n17407), .ZN(P3_U2752) );
  AOI22_X1 U20553 ( .A1(n17424), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20554 ( .B1(n17492), .B2(n17426), .A(n17408), .ZN(P3_U2753) );
  AOI22_X1 U20555 ( .A1(n17424), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20556 ( .B1(n17490), .B2(n17426), .A(n17409), .ZN(P3_U2754) );
  AOI22_X1 U20557 ( .A1(n17424), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20558 ( .B1(n17488), .B2(n17426), .A(n17410), .ZN(P3_U2755) );
  AOI22_X1 U20559 ( .A1(n17424), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20560 ( .B1(n17485), .B2(n17426), .A(n17411), .ZN(P3_U2756) );
  AOI22_X1 U20561 ( .A1(n17424), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20562 ( .B1(n17483), .B2(n17426), .A(n17412), .ZN(P3_U2757) );
  AOI22_X1 U20563 ( .A1(n17424), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17413) );
  OAI21_X1 U20564 ( .B1(n17481), .B2(n17426), .A(n17413), .ZN(P3_U2758) );
  AOI22_X1 U20565 ( .A1(n17424), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20566 ( .B1(n17479), .B2(n17426), .A(n17414), .ZN(P3_U2759) );
  INV_X1 U20567 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20568 ( .A1(n17424), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20569 ( .B1(n17476), .B2(n17426), .A(n17415), .ZN(P3_U2760) );
  AOI22_X1 U20570 ( .A1(n17424), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17416), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17417) );
  OAI21_X1 U20571 ( .B1(n17474), .B2(n17426), .A(n17417), .ZN(P3_U2761) );
  INV_X1 U20572 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20573 ( .A1(n17424), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20574 ( .B1(n17472), .B2(n17426), .A(n17418), .ZN(P3_U2762) );
  INV_X1 U20575 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20576 ( .A1(n17424), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17419) );
  OAI21_X1 U20577 ( .B1(n17470), .B2(n17426), .A(n17419), .ZN(P3_U2763) );
  INV_X1 U20578 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20579 ( .A1(n17424), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20580 ( .B1(n17468), .B2(n17426), .A(n17420), .ZN(P3_U2764) );
  AOI22_X1 U20581 ( .A1(n17424), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20582 ( .B1(n17466), .B2(n17426), .A(n17421), .ZN(P3_U2765) );
  AOI22_X1 U20583 ( .A1(n17424), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17422) );
  OAI21_X1 U20584 ( .B1(n17464), .B2(n17426), .A(n17422), .ZN(P3_U2766) );
  AOI22_X1 U20585 ( .A1(n17424), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17423), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20586 ( .B1(n17462), .B2(n17426), .A(n17425), .ZN(P3_U2767) );
  NOR3_X1 U20587 ( .A1(n18841), .A2(n17429), .A3(n17428), .ZN(n17455) );
  OAI21_X1 U20588 ( .B1(n18841), .B2(n18842), .A(n17430), .ZN(n17486) );
  AOI22_X1 U20589 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17493), .ZN(n17431) );
  OAI21_X1 U20590 ( .B1(n17432), .B2(n17478), .A(n17431), .ZN(P3_U2768) );
  AOI22_X1 U20591 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17493), .ZN(n17433) );
  OAI21_X1 U20592 ( .B1(n17434), .B2(n17478), .A(n17433), .ZN(P3_U2769) );
  AOI22_X1 U20593 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17493), .ZN(n17435) );
  OAI21_X1 U20594 ( .B1(n17436), .B2(n17478), .A(n17435), .ZN(P3_U2770) );
  AOI22_X1 U20595 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17493), .ZN(n17437) );
  OAI21_X1 U20596 ( .B1(n17438), .B2(n17478), .A(n17437), .ZN(P3_U2771) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17493), .ZN(n17439) );
  OAI21_X1 U20598 ( .B1(n17440), .B2(n17478), .A(n17439), .ZN(P3_U2772) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17493), .ZN(n17441) );
  OAI21_X1 U20600 ( .B1(n17442), .B2(n17478), .A(n17441), .ZN(P3_U2773) );
  AOI22_X1 U20601 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17486), .ZN(n17443) );
  OAI21_X1 U20602 ( .B1(n17444), .B2(n17478), .A(n17443), .ZN(P3_U2774) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17486), .ZN(n17445) );
  OAI21_X1 U20604 ( .B1(n17446), .B2(n17478), .A(n17445), .ZN(P3_U2775) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17486), .ZN(n17447) );
  OAI21_X1 U20606 ( .B1(n17448), .B2(n17478), .A(n17447), .ZN(P3_U2776) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17486), .ZN(n17449) );
  OAI21_X1 U20608 ( .B1(n17450), .B2(n17478), .A(n17449), .ZN(P3_U2777) );
  AOI22_X1 U20609 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17486), .ZN(n17451) );
  OAI21_X1 U20610 ( .B1(n17452), .B2(n17478), .A(n17451), .ZN(P3_U2778) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17486), .ZN(n17453) );
  OAI21_X1 U20612 ( .B1(n17454), .B2(n17478), .A(n17453), .ZN(P3_U2779) );
  AOI22_X1 U20613 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17493), .ZN(n17456) );
  OAI21_X1 U20614 ( .B1(n17457), .B2(n17478), .A(n17456), .ZN(P3_U2780) );
  AOI22_X1 U20615 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17493), .ZN(n17458) );
  OAI21_X1 U20616 ( .B1(n20905), .B2(n17478), .A(n17458), .ZN(P3_U2781) );
  AOI22_X1 U20617 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n9649), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17493), .ZN(n17459) );
  OAI21_X1 U20618 ( .B1(n17460), .B2(n17478), .A(n17459), .ZN(P3_U2782) );
  AOI22_X1 U20619 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17493), .ZN(n17461) );
  OAI21_X1 U20620 ( .B1(n17462), .B2(n17478), .A(n17461), .ZN(P3_U2783) );
  AOI22_X1 U20621 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17493), .ZN(n17463) );
  OAI21_X1 U20622 ( .B1(n17464), .B2(n17478), .A(n17463), .ZN(P3_U2784) );
  AOI22_X1 U20623 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17493), .ZN(n17465) );
  OAI21_X1 U20624 ( .B1(n17466), .B2(n17478), .A(n17465), .ZN(P3_U2785) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17493), .ZN(n17467) );
  OAI21_X1 U20626 ( .B1(n17468), .B2(n17478), .A(n17467), .ZN(P3_U2786) );
  AOI22_X1 U20627 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17493), .ZN(n17469) );
  OAI21_X1 U20628 ( .B1(n17470), .B2(n17478), .A(n17469), .ZN(P3_U2787) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17493), .ZN(n17471) );
  OAI21_X1 U20630 ( .B1(n17472), .B2(n17478), .A(n17471), .ZN(P3_U2788) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17493), .ZN(n17473) );
  OAI21_X1 U20632 ( .B1(n17474), .B2(n17478), .A(n17473), .ZN(P3_U2789) );
  AOI22_X1 U20633 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17493), .ZN(n17475) );
  OAI21_X1 U20634 ( .B1(n17476), .B2(n17478), .A(n17475), .ZN(P3_U2790) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17493), .ZN(n17477) );
  OAI21_X1 U20636 ( .B1(n17479), .B2(n17478), .A(n17477), .ZN(P3_U2791) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17486), .ZN(n17480) );
  OAI21_X1 U20638 ( .B1(n17481), .B2(n17478), .A(n17480), .ZN(P3_U2792) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17486), .ZN(n17482) );
  OAI21_X1 U20640 ( .B1(n17483), .B2(n17478), .A(n17482), .ZN(P3_U2793) );
  AOI22_X1 U20641 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17486), .ZN(n17484) );
  OAI21_X1 U20642 ( .B1(n17485), .B2(n17478), .A(n17484), .ZN(P3_U2794) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17486), .ZN(n17487) );
  OAI21_X1 U20644 ( .B1(n17488), .B2(n17478), .A(n17487), .ZN(P3_U2795) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17493), .ZN(n17489) );
  OAI21_X1 U20646 ( .B1(n17490), .B2(n17478), .A(n17489), .ZN(P3_U2796) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17493), .ZN(n17491) );
  OAI21_X1 U20648 ( .B1(n17492), .B2(n17478), .A(n17491), .ZN(P3_U2797) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n9649), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17493), .ZN(n17494) );
  OAI21_X1 U20650 ( .B1(n17495), .B2(n17478), .A(n17494), .ZN(P3_U2798) );
  INV_X1 U20651 ( .A(n18700), .ZN(n17539) );
  AND2_X1 U20652 ( .A1(n17496), .A2(n17539), .ZN(n17497) );
  AOI211_X1 U20653 ( .C1(n17831), .C2(n17508), .A(n17829), .B(n17497), .ZN(
        n17534) );
  OAI21_X1 U20654 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17617), .A(
        n17534), .ZN(n17520) );
  AOI22_X1 U20655 ( .A1(n17730), .A2(n17498), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17520), .ZN(n17513) );
  NOR2_X1 U20656 ( .A1(n17780), .A2(n17842), .ZN(n17620) );
  AOI22_X1 U20657 ( .A1(n17883), .A2(n17780), .B1(n17875), .B2(n17842), .ZN(
        n17499) );
  INV_X1 U20658 ( .A(n17499), .ZN(n17536) );
  NOR2_X1 U20659 ( .A1(n17524), .A2(n17536), .ZN(n17501) );
  NOR3_X1 U20660 ( .A1(n17620), .A2(n17501), .A3(n17500), .ZN(n17507) );
  NOR3_X1 U20661 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17524), .A3(
        n17523), .ZN(n17506) );
  AOI211_X1 U20662 ( .C1(n17504), .C2(n17503), .A(n17502), .B(n17783), .ZN(
        n17505) );
  NOR3_X1 U20663 ( .A1(n17507), .A2(n17506), .A3(n17505), .ZN(n17512) );
  NAND2_X1 U20664 ( .A1(n18174), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17511) );
  NOR2_X1 U20665 ( .A1(n17700), .A2(n17508), .ZN(n17522) );
  OAI211_X1 U20666 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17522), .B(n17509), .ZN(n17510) );
  NAND4_X1 U20667 ( .A1(n17513), .A2(n17512), .A3(n17511), .A4(n17510), .ZN(
        P3_U2802) );
  INV_X1 U20668 ( .A(n17514), .ZN(n17515) );
  NAND2_X1 U20669 ( .A1(n17516), .A2(n17515), .ZN(n17517) );
  XOR2_X1 U20670 ( .A(n17770), .B(n17517), .Z(n17889) );
  OAI22_X1 U20671 ( .A1(n18132), .A2(n18769), .B1(n17672), .B2(n17518), .ZN(
        n17519) );
  AOI221_X1 U20672 ( .B1(n17522), .B2(n17521), .C1(n17520), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17519), .ZN(n17527) );
  INV_X1 U20673 ( .A(n17523), .ZN(n17525) );
  AOI22_X1 U20674 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17536), .B1(
        n17525), .B2(n17524), .ZN(n17526) );
  OAI211_X1 U20675 ( .C1(n17889), .C2(n17783), .A(n17527), .B(n17526), .ZN(
        P3_U2803) );
  AOI21_X1 U20676 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17529), .A(
        n17528), .ZN(n17896) );
  INV_X1 U20677 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17892) );
  AOI21_X1 U20678 ( .B1(n17530), .B2(n18570), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20679 ( .B1(n17730), .B2(n17615), .A(n17531), .ZN(n17532) );
  NAND2_X1 U20680 ( .A1(n18174), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17894) );
  OAI211_X1 U20681 ( .C1(n17534), .C2(n17533), .A(n17532), .B(n17894), .ZN(
        n17535) );
  AOI221_X1 U20682 ( .B1(n9707), .B2(n17892), .C1(n17536), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17535), .ZN(n17537) );
  OAI21_X1 U20683 ( .B1(n17896), .B2(n17783), .A(n17537), .ZN(P3_U2804) );
  XOR2_X1 U20684 ( .A(n17898), .B(n17538), .Z(n17905) );
  AND2_X1 U20685 ( .A1(n17540), .A2(n18570), .ZN(n17569) );
  AOI211_X1 U20686 ( .C1(n17539), .C2(n17564), .A(n17829), .B(n17569), .ZN(
        n17566) );
  OAI21_X1 U20687 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17617), .A(
        n17566), .ZN(n17555) );
  NOR2_X1 U20688 ( .A1(n17700), .A2(n17540), .ZN(n17557) );
  OAI211_X1 U20689 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17557), .B(n17541), .ZN(n17542) );
  NAND2_X1 U20690 ( .A1(n18174), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17902) );
  OAI211_X1 U20691 ( .C1(n17672), .C2(n17543), .A(n17542), .B(n17902), .ZN(
        n17549) );
  XOR2_X1 U20692 ( .A(n17544), .B(n17898), .Z(n17909) );
  OAI21_X1 U20693 ( .B1(n17770), .B2(n17546), .A(n17545), .ZN(n17547) );
  XOR2_X1 U20694 ( .A(n17547), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17904) );
  OAI22_X1 U20695 ( .A1(n17733), .A2(n17909), .B1(n17783), .B2(n17904), .ZN(
        n17548) );
  AOI211_X1 U20696 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17555), .A(
        n17549), .B(n17548), .ZN(n17550) );
  OAI21_X1 U20697 ( .B1(n17872), .B2(n17905), .A(n17550), .ZN(P3_U2805) );
  AOI22_X1 U20698 ( .A1(n17780), .A2(n17912), .B1(n17842), .B2(n17910), .ZN(
        n17575) );
  AOI21_X1 U20699 ( .B1(n17552), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n17551), .ZN(n17553) );
  INV_X1 U20700 ( .A(n17553), .ZN(n17918) );
  NOR2_X1 U20701 ( .A1(n18132), .A2(n18763), .ZN(n17554) );
  AOI221_X1 U20702 ( .B1(n17557), .B2(n17556), .C1(n17555), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17554), .ZN(n17558) );
  OAI21_X1 U20703 ( .B1(n17672), .B2(n17559), .A(n17558), .ZN(n17560) );
  AOI21_X1 U20704 ( .B1(n17752), .B2(n17918), .A(n17560), .ZN(n17561) );
  OAI221_X1 U20705 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17562), 
        .C1(n17919), .C2(n17575), .A(n17561), .ZN(P3_U2806) );
  NOR2_X1 U20706 ( .A1(n18132), .A2(n18761), .ZN(n17927) );
  NAND2_X1 U20707 ( .A1(n17615), .A2(n17565), .ZN(n17563) );
  OAI22_X1 U20708 ( .A1(n17566), .A2(n17565), .B1(n17564), .B2(n17563), .ZN(
        n17567) );
  AOI211_X1 U20709 ( .C1(n17569), .C2(n17568), .A(n17927), .B(n17567), .ZN(
        n17580) );
  AOI22_X1 U20710 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17770), .B1(
        n17571), .B2(n17592), .ZN(n17572) );
  NAND2_X1 U20711 ( .A1(n17570), .A2(n17572), .ZN(n17573) );
  XOR2_X1 U20712 ( .A(n17573), .B(n17924), .Z(n17928) );
  NOR2_X1 U20713 ( .A1(n17574), .A2(n17670), .ZN(n17577) );
  INV_X1 U20714 ( .A(n17575), .ZN(n17576) );
  MUX2_X1 U20715 ( .A(n17577), .B(n17576), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17578) );
  AOI21_X1 U20716 ( .B1(n17752), .B2(n17928), .A(n17578), .ZN(n17579) );
  OAI211_X1 U20717 ( .C1(n17672), .C2(n17581), .A(n17580), .B(n17579), .ZN(
        P3_U2807) );
  OAI21_X1 U20718 ( .B1(n17582), .B2(n18700), .A(n17868), .ZN(n17583) );
  AOI21_X1 U20719 ( .B1(n17831), .B2(n17585), .A(n17583), .ZN(n17612) );
  OAI21_X1 U20720 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17617), .A(
        n17612), .ZN(n17600) );
  NAND2_X1 U20721 ( .A1(n17979), .A2(n17584), .ZN(n17941) );
  NOR3_X1 U20722 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17670), .A3(
        n17941), .ZN(n17590) );
  NAND2_X1 U20723 ( .A1(n18174), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17945) );
  NOR2_X1 U20724 ( .A1(n17700), .A2(n17585), .ZN(n17602) );
  OAI211_X1 U20725 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17602), .B(n17586), .ZN(n17587) );
  OAI211_X1 U20726 ( .C1(n17588), .C2(n17672), .A(n17945), .B(n17587), .ZN(
        n17589) );
  AOI211_X1 U20727 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17600), .A(
        n17590), .B(n17589), .ZN(n17597) );
  INV_X1 U20728 ( .A(n17941), .ZN(n17943) );
  NOR2_X1 U20729 ( .A1(n17591), .A2(n17733), .ZN(n17682) );
  AOI21_X1 U20730 ( .B1(n17842), .B2(n17932), .A(n17682), .ZN(n17669) );
  OAI21_X1 U20731 ( .B1(n17620), .B2(n17943), .A(n17669), .ZN(n17607) );
  INV_X1 U20732 ( .A(n17592), .ZN(n17594) );
  OAI221_X1 U20733 ( .B1(n17594), .B2(n17593), .C1(n17594), .C2(n17943), .A(
        n17570), .ZN(n17595) );
  XNOR2_X1 U20734 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17595), .ZN(
        n17944) );
  AOI22_X1 U20735 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17607), .B1(
        n17752), .B2(n17944), .ZN(n17596) );
  NAND2_X1 U20736 ( .A1(n17597), .A2(n17596), .ZN(P3_U2808) );
  INV_X1 U20737 ( .A(n17938), .ZN(n17953) );
  NAND4_X1 U20738 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17979), .A3(
        n17953), .A4(n17937), .ZN(n17957) );
  OAI22_X1 U20739 ( .A1(n18132), .A2(n18758), .B1(n17672), .B2(n17598), .ZN(
        n17599) );
  AOI221_X1 U20740 ( .B1(n17602), .B2(n17601), .C1(n17600), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17599), .ZN(n17609) );
  NOR3_X1 U20741 ( .A1(n17770), .A2(n17637), .A3(n17603), .ZN(n17625) );
  INV_X1 U20742 ( .A(n17604), .ZN(n17644) );
  AOI22_X1 U20743 ( .A1(n17953), .A2(n17625), .B1(n17644), .B2(n17605), .ZN(
        n17606) );
  XOR2_X1 U20744 ( .A(n17937), .B(n17606), .Z(n17949) );
  AOI22_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17607), .B1(
        n17752), .B2(n17949), .ZN(n17608) );
  OAI211_X1 U20746 ( .C1(n17670), .C2(n17957), .A(n17609), .B(n17608), .ZN(
        P3_U2809) );
  NAND2_X1 U20747 ( .A1(n17979), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17951) );
  NOR2_X1 U20748 ( .A1(n17621), .A2(n17951), .ZN(n17935) );
  INV_X1 U20749 ( .A(n17935), .ZN(n17960) );
  OR2_X1 U20750 ( .A1(n17960), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17967) );
  INV_X1 U20751 ( .A(n17610), .ZN(n17614) );
  AOI221_X1 U20752 ( .B1(n17614), .B2(n17613), .C1(n18266), .C2(n17613), .A(
        n17612), .ZN(n17619) );
  INV_X1 U20753 ( .A(n17615), .ZN(n17617) );
  AOI21_X1 U20754 ( .B1(n17672), .B2(n17617), .A(n17616), .ZN(n17618) );
  AOI211_X1 U20755 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n18174), .A(n17619), 
        .B(n17618), .ZN(n17624) );
  OAI21_X1 U20756 ( .B1(n17620), .B2(n17935), .A(n17669), .ZN(n17634) );
  OAI221_X1 U20757 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17643), 
        .C1(n17621), .C2(n17625), .A(n17570), .ZN(n17622) );
  XNOR2_X1 U20758 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17622), .ZN(
        n17958) );
  AOI22_X1 U20759 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17634), .B1(
        n17752), .B2(n17958), .ZN(n17623) );
  OAI211_X1 U20760 ( .C1(n17670), .C2(n17967), .A(n17624), .B(n17623), .ZN(
        P3_U2810) );
  AOI21_X1 U20761 ( .B1(n17644), .B2(n17643), .A(n17625), .ZN(n17626) );
  XOR2_X1 U20762 ( .A(n17626), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17973) );
  AOI21_X1 U20763 ( .B1(n17831), .B2(n17628), .A(n17829), .ZN(n17650) );
  OAI21_X1 U20764 ( .B1(n17627), .B2(n18700), .A(n17650), .ZN(n17640) );
  NOR2_X1 U20765 ( .A1(n17700), .A2(n17628), .ZN(n17642) );
  OAI211_X1 U20766 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17642), .B(n17629), .ZN(n17630) );
  NAND2_X1 U20767 ( .A1(n18174), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17971) );
  OAI211_X1 U20768 ( .C1(n17672), .C2(n17631), .A(n17630), .B(n17971), .ZN(
        n17632) );
  AOI21_X1 U20769 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17640), .A(
        n17632), .ZN(n17636) );
  NOR2_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17951), .ZN(
        n17969) );
  AOI22_X1 U20771 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17634), .B1(
        n17633), .B2(n17969), .ZN(n17635) );
  OAI211_X1 U20772 ( .C1(n17973), .C2(n17783), .A(n17636), .B(n17635), .ZN(
        P3_U2811) );
  NAND2_X1 U20773 ( .A1(n17979), .A2(n17637), .ZN(n17986) );
  INV_X1 U20774 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17641) );
  NAND2_X1 U20775 ( .A1(n18174), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17984) );
  OAI21_X1 U20776 ( .B1(n17672), .B2(n17638), .A(n17984), .ZN(n17639) );
  AOI221_X1 U20777 ( .B1(n17642), .B2(n17641), .C1(n17640), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17639), .ZN(n17647) );
  OAI21_X1 U20778 ( .B1(n17979), .B2(n17670), .A(n17669), .ZN(n17655) );
  AOI21_X1 U20779 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17758), .A(
        n17643), .ZN(n17645) );
  XOR2_X1 U20780 ( .A(n17645), .B(n17644), .Z(n17982) );
  AOI22_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17655), .B1(
        n17752), .B2(n17982), .ZN(n17646) );
  OAI211_X1 U20782 ( .C1(n17670), .C2(n17986), .A(n17647), .B(n17646), .ZN(
        P3_U2812) );
  NAND2_X1 U20783 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17987), .ZN(
        n17993) );
  AOI21_X1 U20784 ( .B1(n17648), .B2(n18570), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17651) );
  OAI22_X1 U20785 ( .A1(n17651), .A2(n17650), .B1(n17852), .B2(n17649), .ZN(
        n17652) );
  AOI21_X1 U20786 ( .B1(n18174), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17652), 
        .ZN(n17657) );
  OAI21_X1 U20787 ( .B1(n17654), .B2(n17987), .A(n17653), .ZN(n17990) );
  AOI22_X1 U20788 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17655), .B1(
        n17752), .B2(n17990), .ZN(n17656) );
  OAI211_X1 U20789 ( .C1(n17670), .C2(n17993), .A(n17657), .B(n17656), .ZN(
        P3_U2813) );
  AOI21_X1 U20790 ( .B1(n17758), .B2(n17659), .A(n17658), .ZN(n17660) );
  XOR2_X1 U20791 ( .A(n17660), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n18001) );
  AOI21_X1 U20792 ( .B1(n17831), .B2(n17662), .A(n17829), .ZN(n17691) );
  OAI21_X1 U20793 ( .B1(n17661), .B2(n18700), .A(n17691), .ZN(n17674) );
  AOI22_X1 U20794 ( .A1(n18174), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17674), .ZN(n17665) );
  NOR2_X1 U20795 ( .A1(n17700), .A2(n17662), .ZN(n17676) );
  OAI211_X1 U20796 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17676), .B(n17663), .ZN(n17664) );
  OAI211_X1 U20797 ( .C1(n17666), .C2(n17672), .A(n17665), .B(n17664), .ZN(
        n17667) );
  AOI21_X1 U20798 ( .B1(n17752), .B2(n18001), .A(n17667), .ZN(n17668) );
  OAI221_X1 U20799 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17670), 
        .C1(n18004), .C2(n17669), .A(n17668), .ZN(P3_U2814) );
  NOR3_X1 U20800 ( .A1(n18053), .A2(n17677), .A3(n17708), .ZN(n17694) );
  NOR2_X1 U20801 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17694), .ZN(
        n18013) );
  NAND2_X1 U20802 ( .A1(n17842), .A2(n17932), .ZN(n17685) );
  NAND2_X1 U20803 ( .A1(n18174), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18018) );
  OAI21_X1 U20804 ( .B1(n17672), .B2(n17671), .A(n18018), .ZN(n17673) );
  AOI221_X1 U20805 ( .B1(n17676), .B2(n17675), .C1(n17674), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17673), .ZN(n17684) );
  INV_X1 U20806 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18020) );
  INV_X1 U20807 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18024) );
  NAND2_X1 U20808 ( .A1(n17710), .A2(n17770), .ZN(n17717) );
  NAND2_X1 U20809 ( .A1(n17706), .A2(n18060), .ZN(n17678) );
  OAI22_X1 U20810 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17717), .B1(
        n17678), .B2(n17677), .ZN(n17679) );
  OAI221_X1 U20811 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18024), 
        .C1(n17718), .C2(n17758), .A(n17679), .ZN(n17680) );
  XOR2_X1 U20812 ( .A(n18020), .B(n17680), .Z(n18017) );
  AOI21_X1 U20813 ( .B1(n17999), .B2(n17734), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18012) );
  INV_X1 U20814 ( .A(n18012), .ZN(n17681) );
  AOI22_X1 U20815 ( .A1(n17752), .A2(n18017), .B1(n17682), .B2(n17681), .ZN(
        n17683) );
  OAI211_X1 U20816 ( .C1(n18013), .C2(n17685), .A(n17684), .B(n17683), .ZN(
        P3_U2815) );
  INV_X1 U20817 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17712) );
  NAND2_X1 U20818 ( .A1(n17718), .A2(n17712), .ZN(n17686) );
  NAND2_X1 U20819 ( .A1(n18021), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18022) );
  NAND2_X1 U20820 ( .A1(n17758), .A2(n17706), .ZN(n17757) );
  OAI22_X1 U20821 ( .A1(n17686), .A2(n17717), .B1(n18022), .B2(n17757), .ZN(
        n17687) );
  XOR2_X1 U20822 ( .A(n18024), .B(n17687), .Z(n18033) );
  AOI21_X1 U20823 ( .B1(n17688), .B2(n18570), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17690) );
  OAI22_X1 U20824 ( .A1(n17691), .A2(n17690), .B1(n17852), .B2(n17689), .ZN(
        n17692) );
  AOI21_X1 U20825 ( .B1(n18174), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17692), 
        .ZN(n17696) );
  AND2_X1 U20826 ( .A1(n17734), .A2(n17999), .ZN(n17693) );
  AOI221_X1 U20827 ( .B1(n18051), .B2(n18024), .C1(n18022), .C2(n18024), .A(
        n17693), .ZN(n18030) );
  AOI221_X1 U20828 ( .B1(n18053), .B2(n18024), .C1(n18022), .C2(n18024), .A(
        n17694), .ZN(n18029) );
  AOI22_X1 U20829 ( .A1(n17780), .A2(n18030), .B1(n17842), .B2(n18029), .ZN(
        n17695) );
  OAI211_X1 U20830 ( .C1(n18033), .C2(n17783), .A(n17696), .B(n17695), .ZN(
        P3_U2816) );
  INV_X1 U20831 ( .A(n17697), .ZN(n17701) );
  NOR2_X1 U20832 ( .A1(n17698), .A2(n18700), .ZN(n17699) );
  AOI211_X1 U20833 ( .C1(n17831), .C2(n17701), .A(n17829), .B(n17699), .ZN(
        n17720) );
  OR2_X1 U20834 ( .A1(n17701), .A2(n17700), .ZN(n17722) );
  AOI211_X1 U20835 ( .C1(n17716), .C2(n17721), .A(n17702), .B(n17722), .ZN(
        n17704) );
  NOR2_X1 U20836 ( .A1(n18132), .A2(n18742), .ZN(n17703) );
  AOI211_X1 U20837 ( .C1(n17730), .C2(n17705), .A(n17704), .B(n17703), .ZN(
        n17715) );
  NOR2_X1 U20838 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17708), .ZN(
        n18034) );
  NAND2_X1 U20839 ( .A1(n17734), .A2(n18021), .ZN(n18040) );
  NAND2_X1 U20840 ( .A1(n17732), .A2(n18021), .ZN(n18035) );
  AOI22_X1 U20841 ( .A1(n17780), .A2(n18040), .B1(n17842), .B2(n18035), .ZN(
        n17724) );
  INV_X1 U20842 ( .A(n17706), .ZN(n17707) );
  OAI22_X1 U20843 ( .A1(n17758), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17708), .B2(n17707), .ZN(n17709) );
  OAI21_X1 U20844 ( .B1(n17758), .B2(n17710), .A(n17709), .ZN(n17711) );
  XOR2_X1 U20845 ( .A(n17711), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18044) );
  OAI22_X1 U20846 ( .A1(n17724), .A2(n17712), .B1(n17783), .B2(n18044), .ZN(
        n17713) );
  AOI21_X1 U20847 ( .B1(n18034), .B2(n17766), .A(n17713), .ZN(n17714) );
  OAI211_X1 U20848 ( .C1(n17720), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        P3_U2817) );
  OR3_X1 U20849 ( .A1(n10139), .A2(n10140), .A3(n17757), .ZN(n17740) );
  OAI21_X1 U20850 ( .B1(n17744), .B2(n17740), .A(n17717), .ZN(n17719) );
  XOR2_X1 U20851 ( .A(n17719), .B(n17718), .Z(n18050) );
  NAND2_X1 U20852 ( .A1(n18174), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18048) );
  OAI221_X1 U20853 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17722), .C1(
        n17721), .C2(n17720), .A(n18048), .ZN(n17728) );
  INV_X1 U20854 ( .A(n17766), .ZN(n17723) );
  NOR2_X1 U20855 ( .A1(n17723), .A2(n18036), .ZN(n17726) );
  INV_X1 U20856 ( .A(n17724), .ZN(n17725) );
  MUX2_X1 U20857 ( .A(n17726), .B(n17725), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17727) );
  AOI211_X1 U20858 ( .C1(n17730), .C2(n17729), .A(n17728), .B(n17727), .ZN(
        n17731) );
  OAI21_X1 U20859 ( .B1(n18050), .B2(n17783), .A(n17731), .ZN(P3_U2818) );
  OAI22_X1 U20860 ( .A1(n17734), .A2(n17733), .B1(n17872), .B2(n17732), .ZN(
        n17767) );
  AOI21_X1 U20861 ( .B1(n18058), .B2(n17766), .A(n17767), .ZN(n17756) );
  INV_X1 U20862 ( .A(n17865), .ZN(n17796) );
  NOR3_X1 U20863 ( .A1(n17787), .A2(n17772), .A3(n18266), .ZN(n17762) );
  NAND2_X1 U20864 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17762), .ZN(
        n17761) );
  NOR2_X1 U20865 ( .A1(n17746), .A2(n17761), .ZN(n17745) );
  NOR2_X1 U20866 ( .A1(n17737), .A2(n17745), .ZN(n17738) );
  INV_X1 U20867 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18738) );
  OAI22_X1 U20868 ( .A1(n17852), .A2(n17735), .B1(n18132), .B2(n18738), .ZN(
        n17736) );
  AOI221_X1 U20869 ( .B1(n17796), .B2(n17738), .C1(n17737), .C2(n17745), .A(
        n17736), .ZN(n17743) );
  NAND3_X1 U20870 ( .A1(n17739), .A2(n17770), .A3(n10139), .ZN(n17749) );
  OAI21_X1 U20871 ( .B1(n17749), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17740), .ZN(n17741) );
  XOR2_X1 U20872 ( .A(n17741), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18064) );
  NOR2_X1 U20873 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18058), .ZN(
        n18063) );
  AOI22_X1 U20874 ( .A1(n17752), .A2(n18064), .B1(n18063), .B2(n17766), .ZN(
        n17742) );
  OAI211_X1 U20875 ( .C1(n17756), .C2(n17744), .A(n17743), .B(n17742), .ZN(
        P3_U2819) );
  AOI21_X1 U20876 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17766), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17755) );
  INV_X1 U20877 ( .A(n17745), .ZN(n17748) );
  OAI21_X1 U20878 ( .B1(n17865), .B2(n17746), .A(n17761), .ZN(n17747) );
  AOI22_X1 U20879 ( .A1(n18174), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17748), 
        .B2(n17747), .ZN(n17754) );
  OAI21_X1 U20880 ( .B1(n17757), .B2(n10139), .A(n17749), .ZN(n17750) );
  XNOR2_X1 U20881 ( .A(n10140), .B(n17750), .ZN(n18069) );
  AOI22_X1 U20882 ( .A1(n17752), .A2(n18069), .B1(n17751), .B2(n17860), .ZN(
        n17753) );
  OAI211_X1 U20883 ( .C1(n17756), .C2(n17755), .A(n17754), .B(n17753), .ZN(
        P3_U2820) );
  OAI21_X1 U20884 ( .B1(n17759), .B2(n17758), .A(n17757), .ZN(n17760) );
  XOR2_X1 U20885 ( .A(n17760), .B(n10139), .Z(n18073) );
  OAI211_X1 U20886 ( .C1(n17762), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17796), .B(n17761), .ZN(n17763) );
  NAND2_X1 U20887 ( .A1(n18174), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18082) );
  OAI211_X1 U20888 ( .C1(n17852), .C2(n17764), .A(n17763), .B(n18082), .ZN(
        n17765) );
  AOI221_X1 U20889 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17767), .C1(
        n10139), .C2(n17766), .A(n17765), .ZN(n17768) );
  OAI21_X1 U20890 ( .B1(n18073), .B2(n17783), .A(n17768), .ZN(P3_U2821) );
  OAI21_X1 U20891 ( .B1(n18094), .B2(n17770), .A(n17769), .ZN(n18097) );
  AOI21_X1 U20892 ( .B1(n17787), .B2(n17831), .A(n17829), .ZN(n17771) );
  INV_X1 U20893 ( .A(n17771), .ZN(n17788) );
  NOR2_X1 U20894 ( .A1(n17787), .A2(n17789), .ZN(n17773) );
  OAI211_X1 U20895 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17773), .A(
        n18570), .B(n17772), .ZN(n17775) );
  INV_X1 U20896 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18733) );
  NOR2_X1 U20897 ( .A1(n18132), .A2(n18733), .ZN(n18088) );
  INV_X1 U20898 ( .A(n18088), .ZN(n17774) );
  OAI211_X1 U20899 ( .C1(n17852), .C2(n17776), .A(n17775), .B(n17774), .ZN(
        n17777) );
  AOI21_X1 U20900 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17788), .A(
        n17777), .ZN(n17782) );
  AOI21_X1 U20901 ( .B1(n17779), .B2(n18090), .A(n17778), .ZN(n18092) );
  AOI22_X1 U20902 ( .A1(n17780), .A2(n18094), .B1(n17842), .B2(n18092), .ZN(
        n17781) );
  OAI211_X1 U20903 ( .C1(n17783), .C2(n18097), .A(n17782), .B(n17781), .ZN(
        P3_U2822) );
  NAND2_X1 U20904 ( .A1(n17785), .A2(n17784), .ZN(n17786) );
  XOR2_X1 U20905 ( .A(n17786), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18110) );
  NOR2_X1 U20906 ( .A1(n17787), .A2(n18266), .ZN(n17790) );
  NOR2_X1 U20907 ( .A1(n18132), .A2(n18730), .ZN(n18099) );
  AOI221_X1 U20908 ( .B1(n17790), .B2(n17789), .C1(n17788), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18099), .ZN(n17795) );
  AOI21_X1 U20909 ( .B1(n18104), .B2(n17792), .A(n17791), .ZN(n18106) );
  AOI22_X1 U20910 ( .A1(n17861), .A2(n18106), .B1(n17793), .B2(n17860), .ZN(
        n17794) );
  OAI211_X1 U20911 ( .C1(n17872), .C2(n18110), .A(n17795), .B(n17794), .ZN(
        P3_U2823) );
  OAI21_X1 U20912 ( .B1(n17799), .B2(n18266), .A(n17796), .ZN(n17818) );
  AOI21_X1 U20913 ( .B1(n18105), .B2(n17798), .A(n17797), .ZN(n18114) );
  NOR2_X1 U20914 ( .A1(n18132), .A2(n18728), .ZN(n18113) );
  NOR3_X1 U20915 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17799), .A3(
        n18266), .ZN(n17800) );
  AOI211_X1 U20916 ( .C1(n17842), .C2(n18114), .A(n18113), .B(n17800), .ZN(
        n17805) );
  AOI21_X1 U20917 ( .B1(n9767), .B2(n17802), .A(n17801), .ZN(n18115) );
  AOI22_X1 U20918 ( .A1(n17861), .A2(n18115), .B1(n17803), .B2(n17860), .ZN(
        n17804) );
  OAI211_X1 U20919 ( .C1(n17806), .C2(n17818), .A(n17805), .B(n17804), .ZN(
        P3_U2824) );
  NOR2_X1 U20920 ( .A1(n17830), .A2(n17832), .ZN(n17807) );
  AOI21_X1 U20921 ( .B1(n17807), .B2(n17868), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17819) );
  AOI21_X1 U20922 ( .B1(n17810), .B2(n17809), .A(n17808), .ZN(n18119) );
  AOI22_X1 U20923 ( .A1(n17842), .A2(n18119), .B1(n18174), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17817) );
  AOI21_X1 U20924 ( .B1(n17813), .B2(n17812), .A(n17811), .ZN(n17814) );
  XOR2_X1 U20925 ( .A(n17814), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18120) );
  AOI22_X1 U20926 ( .A1(n17861), .A2(n18120), .B1(n17815), .B2(n17860), .ZN(
        n17816) );
  OAI211_X1 U20927 ( .C1(n17819), .C2(n17818), .A(n17817), .B(n17816), .ZN(
        P3_U2825) );
  OAI21_X1 U20928 ( .B1(n17822), .B2(n17821), .A(n17820), .ZN(n17823) );
  XOR2_X1 U20929 ( .A(n17823), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18137) );
  OAI21_X1 U20930 ( .B1(n17826), .B2(n17825), .A(n17824), .ZN(n17827) );
  XOR2_X1 U20931 ( .A(n17827), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18131) );
  OAI22_X1 U20932 ( .A1(n17872), .A2(n18131), .B1(n18266), .B2(n17828), .ZN(
        n17835) );
  AOI21_X1 U20933 ( .B1(n17831), .B2(n17830), .A(n17829), .ZN(n17845) );
  OAI22_X1 U20934 ( .A1(n17852), .A2(n17833), .B1(n17832), .B2(n17845), .ZN(
        n17834) );
  AOI211_X1 U20935 ( .C1(n18174), .C2(P3_REIP_REG_4__SCAN_IN), .A(n17835), .B(
        n17834), .ZN(n17836) );
  OAI21_X1 U20936 ( .B1(n17871), .B2(n18137), .A(n17836), .ZN(P3_U2826) );
  AOI21_X1 U20937 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17868), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17846) );
  AOI22_X1 U20938 ( .A1(n17861), .A2(n18140), .B1(n18174), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17844) );
  AOI21_X1 U20939 ( .B1(n17840), .B2(n17839), .A(n17838), .ZN(n18139) );
  AOI22_X1 U20940 ( .A1(n17842), .A2(n18139), .B1(n17841), .B2(n17860), .ZN(
        n17843) );
  OAI211_X1 U20941 ( .C1(n17846), .C2(n17845), .A(n17844), .B(n17843), .ZN(
        P3_U2827) );
  AOI21_X1 U20942 ( .B1(n9778), .B2(n17848), .A(n17847), .ZN(n18153) );
  NOR2_X1 U20943 ( .A1(n18132), .A2(n18720), .ZN(n18159) );
  XNOR2_X1 U20944 ( .A(n17850), .B(n17849), .ZN(n18161) );
  OAI22_X1 U20945 ( .A1(n17852), .A2(n17851), .B1(n17872), .B2(n18161), .ZN(
        n17853) );
  AOI211_X1 U20946 ( .C1(n17861), .C2(n18153), .A(n18159), .B(n17853), .ZN(
        n17854) );
  OAI221_X1 U20947 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18266), .C1(
        n17855), .C2(n17868), .A(n17854), .ZN(P3_U2828) );
  NOR2_X1 U20948 ( .A1(n17867), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17856) );
  XOR2_X1 U20949 ( .A(n17856), .B(n17859), .Z(n18173) );
  OAI22_X1 U20950 ( .A1(n17872), .A2(n18173), .B1(n18132), .B2(n18823), .ZN(
        n17857) );
  INV_X1 U20951 ( .A(n17857), .ZN(n17863) );
  AOI21_X1 U20952 ( .B1(n17866), .B2(n17859), .A(n17858), .ZN(n18166) );
  AOI22_X1 U20953 ( .A1(n17861), .A2(n18166), .B1(n17864), .B2(n17860), .ZN(
        n17862) );
  OAI211_X1 U20954 ( .C1(n17865), .C2(n17864), .A(n17863), .B(n17862), .ZN(
        P3_U2829) );
  OAI21_X1 U20955 ( .B1(n17867), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17866), .ZN(n18181) );
  INV_X1 U20956 ( .A(n18181), .ZN(n17873) );
  OAI21_X1 U20957 ( .B1(n18692), .B2(n18844), .A(n17868), .ZN(n17869) );
  AOI22_X1 U20958 ( .A1(n18174), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17869), .ZN(n17870) );
  OAI221_X1 U20959 ( .B1(n17873), .B2(n17872), .C1(n18181), .C2(n17871), .A(
        n17870), .ZN(P3_U2830) );
  NAND2_X1 U20960 ( .A1(n18132), .A2(n18167), .ZN(n18130) );
  NOR2_X1 U20961 ( .A1(n17874), .A2(n17925), .ZN(n17885) );
  INV_X1 U20962 ( .A(n17875), .ZN(n17881) );
  NOR2_X1 U20963 ( .A1(n18648), .A2(n17997), .ZN(n18126) );
  INV_X1 U20964 ( .A(n18126), .ZN(n18146) );
  INV_X1 U20965 ( .A(n17900), .ZN(n17877) );
  NOR2_X1 U20966 ( .A1(n18657), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18129) );
  INV_X1 U20967 ( .A(n18129), .ZN(n18149) );
  AOI21_X1 U20968 ( .B1(n17876), .B2(n18149), .A(n18126), .ZN(n17911) );
  AOI21_X1 U20969 ( .B1(n18146), .B2(n17877), .A(n17911), .ZN(n17897) );
  AOI21_X1 U20970 ( .B1(n17879), .B2(n18146), .A(n17878), .ZN(n17880) );
  OAI211_X1 U20971 ( .C1(n17881), .C2(n18629), .A(n17897), .B(n17880), .ZN(
        n17882) );
  AOI21_X1 U20972 ( .B1(n18052), .B2(n17883), .A(n17882), .ZN(n17890) );
  INV_X1 U20973 ( .A(n17890), .ZN(n17884) );
  MUX2_X1 U20974 ( .A(n17885), .B(n17884), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17886) );
  AOI22_X1 U20975 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18169), .B1(
        n18175), .B2(n17886), .ZN(n17888) );
  NAND2_X1 U20976 ( .A1(n18174), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17887) );
  OAI211_X1 U20977 ( .C1(n17889), .C2(n18098), .A(n17888), .B(n17887), .ZN(
        P3_U2835) );
  NAND4_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17920), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A4(n17942), .ZN(n17891) );
  AOI211_X1 U20979 ( .C1(n17892), .C2(n17891), .A(n17890), .B(n18167), .ZN(
        n17893) );
  AOI21_X1 U20980 ( .B1(n18169), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17893), .ZN(n17895) );
  OAI211_X1 U20981 ( .C1(n17896), .C2(n18098), .A(n17895), .B(n17894), .ZN(
        P3_U2836) );
  OAI221_X1 U20982 ( .B1(n18665), .B2(n17900), .C1(n18665), .C2(n17915), .A(
        n17897), .ZN(n17899) );
  OAI222_X1 U20983 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17901), 
        .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17900), .C1(n17899), 
        .C2(n17898), .ZN(n17903) );
  OAI21_X1 U20984 ( .B1(n18167), .B2(n17903), .A(n17902), .ZN(n17907) );
  OAI22_X1 U20985 ( .A1(n18172), .A2(n17905), .B1(n18098), .B2(n17904), .ZN(
        n17906) );
  AOI211_X1 U20986 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18169), .A(
        n17907), .B(n17906), .ZN(n17908) );
  OAI21_X1 U20987 ( .B1(n17974), .B2(n17909), .A(n17908), .ZN(P3_U2837) );
  INV_X1 U20988 ( .A(n17910), .ZN(n17914) );
  AOI211_X1 U20989 ( .C1(n18052), .C2(n17912), .A(n17911), .B(n18169), .ZN(
        n17913) );
  OAI21_X1 U20990 ( .B1(n17914), .B2(n18629), .A(n17913), .ZN(n17917) );
  OAI21_X1 U20991 ( .B1(n18087), .B2(n17917), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17923) );
  OAI21_X1 U20992 ( .B1(n17915), .B2(n18665), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17916) );
  OAI21_X1 U20993 ( .B1(n17917), .B2(n17916), .A(n18132), .ZN(n17930) );
  AOI22_X1 U20994 ( .A1(n18174), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18076), 
        .B2(n17918), .ZN(n17922) );
  NAND2_X1 U20995 ( .A1(n18175), .A2(n17942), .ZN(n17966) );
  INV_X1 U20996 ( .A(n17966), .ZN(n17968) );
  NAND3_X1 U20997 ( .A1(n17920), .A2(n17968), .A3(n17919), .ZN(n17921) );
  OAI211_X1 U20998 ( .C1(n17923), .C2(n17930), .A(n17922), .B(n17921), .ZN(
        P3_U2838) );
  OAI21_X1 U20999 ( .B1(n17925), .B2(n18169), .A(n17924), .ZN(n17926) );
  INV_X1 U21000 ( .A(n17926), .ZN(n17931) );
  AOI21_X1 U21001 ( .B1(n17928), .B2(n18076), .A(n17927), .ZN(n17929) );
  OAI21_X1 U21002 ( .B1(n17931), .B2(n17930), .A(n17929), .ZN(P3_U2839) );
  AND2_X1 U21003 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17994), .ZN(
        n18077) );
  NAND2_X1 U21004 ( .A1(n17975), .A2(n18077), .ZN(n17996) );
  AOI22_X1 U21005 ( .A1(n18054), .A2(n17932), .B1(n18052), .B2(n18009), .ZN(
        n17950) );
  OAI21_X1 U21006 ( .B1(n17933), .B2(n17951), .A(n18148), .ZN(n17934) );
  OAI221_X1 U21007 ( .B1(n18639), .B2(n17976), .C1(n18639), .C2(n17935), .A(
        n17934), .ZN(n17959) );
  NOR2_X1 U21008 ( .A1(n18054), .A2(n18052), .ZN(n17977) );
  OAI22_X1 U21009 ( .A1(n18639), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17943), .B2(n17977), .ZN(n17936) );
  NOR2_X1 U21010 ( .A1(n17959), .A2(n17936), .ZN(n17952) );
  AOI22_X1 U21011 ( .A1(n18148), .A2(n17938), .B1(n18067), .B2(n17937), .ZN(
        n17939) );
  NAND4_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17950), .A3(
        n17952), .A4(n17939), .ZN(n17940) );
  AOI221_X1 U21013 ( .B1(n17941), .B2(n17997), .C1(n17996), .C2(n17997), .A(
        n17940), .ZN(n17948) );
  OAI221_X1 U21014 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17943), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17942), .A(n18175), .ZN(
        n17947) );
  AOI22_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18169), .B1(
        n18076), .B2(n17944), .ZN(n17946) );
  OAI211_X1 U21016 ( .C1(n17948), .C2(n17947), .A(n17946), .B(n17945), .ZN(
        P3_U2840) );
  AOI22_X1 U21017 ( .A1(n18174), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18076), 
        .B2(n17949), .ZN(n17956) );
  NAND2_X1 U21018 ( .A1(n18175), .A2(n17950), .ZN(n18000) );
  NOR2_X1 U21019 ( .A1(n18148), .A2(n17997), .ZN(n18168) );
  OAI21_X1 U21020 ( .B1(n17951), .B2(n17996), .A(n17997), .ZN(n17961) );
  OAI211_X1 U21021 ( .C1(n18168), .C2(n17953), .A(n17961), .B(n17952), .ZN(
        n17954) );
  OAI211_X1 U21022 ( .C1(n18000), .C2(n17954), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18132), .ZN(n17955) );
  OAI211_X1 U21023 ( .C1(n17966), .C2(n17957), .A(n17956), .B(n17955), .ZN(
        P3_U2841) );
  AOI22_X1 U21024 ( .A1(n18174), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18076), 
        .B2(n17958), .ZN(n17965) );
  INV_X1 U21025 ( .A(n17977), .ZN(n18057) );
  AOI211_X1 U21026 ( .C1(n17960), .C2(n18057), .A(n18000), .B(n17959), .ZN(
        n17962) );
  AOI21_X1 U21027 ( .B1(n17962), .B2(n17961), .A(n18174), .ZN(n17970) );
  NOR3_X1 U21028 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18168), .A3(
        n18682), .ZN(n17963) );
  OAI21_X1 U21029 ( .B1(n17970), .B2(n17963), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17964) );
  OAI211_X1 U21030 ( .C1(n17967), .C2(n17966), .A(n17965), .B(n17964), .ZN(
        P3_U2842) );
  AOI22_X1 U21031 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17970), .B1(
        n17969), .B2(n17968), .ZN(n17972) );
  OAI211_X1 U21032 ( .C1(n17973), .C2(n18098), .A(n17972), .B(n17971), .ZN(
        P3_U2843) );
  AOI22_X1 U21033 ( .A1(n18148), .A2(n18145), .B1(n18155), .B2(n18125), .ZN(
        n18100) );
  NOR3_X1 U21034 ( .A1(n18100), .A2(n18167), .A3(n18128), .ZN(n18135) );
  NAND3_X1 U21035 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n18135), .ZN(n18118) );
  OAI222_X1 U21036 ( .A1(n18118), .A2(n18007), .B1(n18172), .B2(n18053), .C1(
        n18051), .C2(n17974), .ZN(n18074) );
  NAND2_X1 U21037 ( .A1(n17975), .A2(n18074), .ZN(n18005) );
  NAND3_X1 U21038 ( .A1(n17976), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18149), .ZN(n17981) );
  AOI222_X1 U21039 ( .A1(n17979), .A2(n18665), .B1(n17979), .B2(n17978), .C1(
        n18665), .C2(n17977), .ZN(n17980) );
  AOI211_X1 U21040 ( .C1(n18146), .C2(n17981), .A(n17980), .B(n18000), .ZN(
        n17988) );
  AOI221_X1 U21041 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17988), 
        .C1(n18126), .C2(n17988), .A(n18174), .ZN(n17983) );
  AOI22_X1 U21042 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17983), .B1(
        n18076), .B2(n17982), .ZN(n17985) );
  OAI211_X1 U21043 ( .C1(n18005), .C2(n17986), .A(n17985), .B(n17984), .ZN(
        P3_U2844) );
  NOR3_X1 U21044 ( .A1(n18174), .A2(n17988), .A3(n17987), .ZN(n17989) );
  AOI21_X1 U21045 ( .B1(n18076), .B2(n17990), .A(n17989), .ZN(n17992) );
  NAND2_X1 U21046 ( .A1(n18174), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17991) );
  OAI211_X1 U21047 ( .C1(n17993), .C2(n18005), .A(n17992), .B(n17991), .ZN(
        P3_U2845) );
  OAI22_X1 U21048 ( .A1(n18665), .A2(n17995), .B1(n18639), .B2(n17994), .ZN(
        n18056) );
  INV_X1 U21049 ( .A(n18056), .ZN(n18078) );
  OAI21_X1 U21050 ( .B1(n18020), .B2(n17997), .A(n17996), .ZN(n17998) );
  OAI211_X1 U21051 ( .C1(n18061), .C2(n17999), .A(n18078), .B(n17998), .ZN(
        n18008) );
  OAI221_X1 U21052 ( .B1(n18000), .B2(n18087), .C1(n18000), .C2(n18008), .A(
        n18132), .ZN(n18003) );
  AOI22_X1 U21053 ( .A1(n18174), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18076), 
        .B2(n18001), .ZN(n18002) );
  OAI221_X1 U21054 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18005), 
        .C1(n18004), .C2(n18003), .A(n18002), .ZN(P3_U2846) );
  NOR4_X1 U21055 ( .A1(n18100), .A2(n18007), .A3(n18006), .A4(n18022), .ZN(
        n18023) );
  OAI221_X1 U21056 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18023), .A(n18008), .ZN(
        n18011) );
  NAND2_X1 U21057 ( .A1(n18052), .A2(n18009), .ZN(n18010) );
  AOI221_X1 U21058 ( .B1(n18012), .B2(n18011), .C1(n18010), .C2(n18011), .A(
        n18167), .ZN(n18016) );
  NOR3_X1 U21059 ( .A1(n18014), .A2(n18013), .A3(n18172), .ZN(n18015) );
  AOI211_X1 U21060 ( .C1(n18076), .C2(n18017), .A(n18016), .B(n18015), .ZN(
        n18019) );
  OAI211_X1 U21061 ( .C1(n18130), .C2(n18020), .A(n18019), .B(n18018), .ZN(
        P3_U2847) );
  NOR2_X1 U21062 ( .A1(n18132), .A2(n18745), .ZN(n18028) );
  OAI221_X1 U21063 ( .B1(n18657), .B2(n18021), .C1(n18657), .C2(n18077), .A(
        n18078), .ZN(n18039) );
  AOI21_X1 U21064 ( .B1(n18087), .B2(n18022), .A(n18039), .ZN(n18026) );
  INV_X1 U21065 ( .A(n18023), .ZN(n18025) );
  AOI221_X1 U21066 ( .B1(n18026), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n18025), .C2(n18024), .A(n18167), .ZN(n18027) );
  AOI211_X1 U21067 ( .C1(n18169), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18028), .B(n18027), .ZN(n18032) );
  AOI22_X1 U21068 ( .A1(n18093), .A2(n18030), .B1(n18178), .B2(n18029), .ZN(
        n18031) );
  OAI211_X1 U21069 ( .C1(n18033), .C2(n18098), .A(n18032), .B(n18031), .ZN(
        P3_U2848) );
  AOI22_X1 U21070 ( .A1(n18174), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18034), 
        .B2(n18074), .ZN(n18043) );
  AOI22_X1 U21071 ( .A1(n18067), .A2(n18036), .B1(n18035), .B2(n18054), .ZN(
        n18037) );
  INV_X1 U21072 ( .A(n18037), .ZN(n18038) );
  AOI211_X1 U21073 ( .C1(n18052), .C2(n18040), .A(n18039), .B(n18038), .ZN(
        n18046) );
  OAI211_X1 U21074 ( .C1(n18061), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18175), .B(n18046), .ZN(n18041) );
  NAND3_X1 U21075 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18132), .A3(
        n18041), .ZN(n18042) );
  OAI211_X1 U21076 ( .C1(n18044), .C2(n18098), .A(n18043), .B(n18042), .ZN(
        P3_U2849) );
  AOI22_X1 U21077 ( .A1(n18060), .A2(n18074), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18175), .ZN(n18045) );
  AOI21_X1 U21078 ( .B1(n18046), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18045), .ZN(n18047) );
  AOI21_X1 U21079 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18169), .A(
        n18047), .ZN(n18049) );
  OAI211_X1 U21080 ( .C1(n18050), .C2(n18098), .A(n18049), .B(n18048), .ZN(
        P3_U2850) );
  AOI22_X1 U21081 ( .A1(n18054), .A2(n18053), .B1(n18052), .B2(n18051), .ZN(
        n18055) );
  NAND2_X1 U21082 ( .A1(n18175), .A2(n18055), .ZN(n18079) );
  AOI211_X1 U21083 ( .C1(n18058), .C2(n18057), .A(n18056), .B(n18079), .ZN(
        n18059) );
  OAI221_X1 U21084 ( .B1(n18657), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18657), .C2(n18077), .A(n18059), .ZN(n18068) );
  OAI22_X1 U21085 ( .A1(n18061), .A2(n18060), .B1(n18657), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18062) );
  OAI21_X1 U21086 ( .B1(n18068), .B2(n18062), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U21087 ( .A1(n18076), .A2(n18064), .B1(n18063), .B2(n18074), .ZN(
        n18065) );
  OAI221_X1 U21088 ( .B1(n18174), .B2(n18066), .C1(n18132), .C2(n18738), .A(
        n18065), .ZN(P3_U2851) );
  NAND2_X1 U21089 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18074), .ZN(
        n18072) );
  OAI221_X1 U21090 ( .B1(n18068), .B2(n18067), .C1(n18068), .C2(n10139), .A(
        n18132), .ZN(n18071) );
  AOI22_X1 U21091 ( .A1(n18174), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18076), 
        .B2(n18069), .ZN(n18070) );
  OAI221_X1 U21092 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18072), 
        .C1(n10140), .C2(n18071), .A(n18070), .ZN(P3_U2852) );
  INV_X1 U21093 ( .A(n18073), .ZN(n18075) );
  AOI22_X1 U21094 ( .A1(n18076), .A2(n18075), .B1(n10139), .B2(n18074), .ZN(
        n18083) );
  AOI21_X1 U21095 ( .B1(n18657), .B2(n18078), .A(n18077), .ZN(n18080) );
  OAI211_X1 U21096 ( .C1(n18080), .C2(n18079), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18132), .ZN(n18081) );
  NAND3_X1 U21097 ( .A1(n18083), .A2(n18082), .A3(n18081), .ZN(P3_U2853) );
  NOR3_X1 U21098 ( .A1(n18105), .A2(n18104), .A3(n18118), .ZN(n18091) );
  AOI22_X1 U21099 ( .A1(n18148), .A2(n18085), .B1(n18146), .B2(n18084), .ZN(
        n18086) );
  NAND2_X1 U21100 ( .A1(n18086), .A2(n18149), .ZN(n18111) );
  AOI211_X1 U21101 ( .C1(n18087), .C2(n18105), .A(n18104), .B(n18111), .ZN(
        n18102) );
  OAI21_X1 U21102 ( .B1(n18102), .B2(n18162), .A(n18130), .ZN(n18089) );
  AOI221_X1 U21103 ( .B1(n18091), .B2(n18090), .C1(n18089), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18088), .ZN(n18096) );
  AOI22_X1 U21104 ( .A1(n18094), .A2(n18093), .B1(n18178), .B2(n18092), .ZN(
        n18095) );
  OAI211_X1 U21105 ( .C1(n18098), .C2(n18097), .A(n18096), .B(n18095), .ZN(
        P3_U2854) );
  AOI21_X1 U21106 ( .B1(n18169), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18099), .ZN(n18109) );
  INV_X1 U21107 ( .A(n18100), .ZN(n18138) );
  NAND2_X1 U21108 ( .A1(n18101), .A2(n18138), .ZN(n18103) );
  AOI221_X1 U21109 ( .B1(n18105), .B2(n18104), .C1(n18103), .C2(n18104), .A(
        n18102), .ZN(n18107) );
  AOI22_X1 U21110 ( .A1(n18175), .A2(n18107), .B1(n18165), .B2(n18106), .ZN(
        n18108) );
  OAI211_X1 U21111 ( .C1(n18172), .C2(n18110), .A(n18109), .B(n18108), .ZN(
        P3_U2855) );
  OAI21_X1 U21112 ( .B1(n18167), .B2(n18111), .A(n18132), .ZN(n18112) );
  INV_X1 U21113 ( .A(n18112), .ZN(n18121) );
  AOI21_X1 U21114 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18121), .A(
        n18113), .ZN(n18117) );
  AOI22_X1 U21115 ( .A1(n18165), .A2(n18115), .B1(n18178), .B2(n18114), .ZN(
        n18116) );
  OAI211_X1 U21116 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18118), .A(
        n18117), .B(n18116), .ZN(P3_U2856) );
  AOI22_X1 U21117 ( .A1(n18174), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18178), 
        .B2(n18119), .ZN(n18124) );
  AOI22_X1 U21118 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18121), .B1(
        n18165), .B2(n18120), .ZN(n18123) );
  NAND3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18135), .A3(
        n10148), .ZN(n18122) );
  NAND3_X1 U21120 ( .A1(n18124), .A2(n18123), .A3(n18122), .ZN(P3_U2857) );
  OAI22_X1 U21121 ( .A1(n18126), .A2(n18125), .B1(n18665), .B2(n18145), .ZN(
        n18127) );
  NOR3_X1 U21122 ( .A1(n18129), .A2(n18128), .A3(n18127), .ZN(n18144) );
  OAI21_X1 U21123 ( .B1(n18144), .B2(n18162), .A(n18130), .ZN(n18134) );
  OAI22_X1 U21124 ( .A1(n18132), .A2(n18725), .B1(n18172), .B2(n18131), .ZN(
        n18133) );
  AOI221_X1 U21125 ( .B1(n18135), .B2(n15535), .C1(n18134), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18133), .ZN(n18136) );
  OAI21_X1 U21126 ( .B1(n18182), .B2(n18137), .A(n18136), .ZN(P3_U2858) );
  OAI21_X1 U21127 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18138), .A(
        n18175), .ZN(n18143) );
  AOI22_X1 U21128 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18169), .B1(
        n18174), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U21129 ( .A1(n18165), .A2(n18140), .B1(n18178), .B2(n18139), .ZN(
        n18141) );
  OAI211_X1 U21130 ( .C1(n18144), .C2(n18143), .A(n18142), .B(n18141), .ZN(
        P3_U2859) );
  NOR2_X1 U21131 ( .A1(n18665), .A2(n18145), .ZN(n18152) );
  NOR2_X1 U21132 ( .A1(n18802), .A2(n18819), .ZN(n18147) );
  AOI22_X1 U21133 ( .A1(n18148), .A2(n18147), .B1(n18802), .B2(n18146), .ZN(
        n18150) );
  AOI21_X1 U21134 ( .B1(n18150), .B2(n18149), .A(n18154), .ZN(n18151) );
  AOI211_X1 U21135 ( .C1(n18153), .C2(n18627), .A(n18152), .B(n18151), .ZN(
        n18157) );
  NAND3_X1 U21136 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18155), .A3(
        n18154), .ZN(n18156) );
  AOI21_X1 U21137 ( .B1(n18157), .B2(n18156), .A(n18167), .ZN(n18158) );
  AOI211_X1 U21138 ( .C1(n18169), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18159), .B(n18158), .ZN(n18160) );
  OAI21_X1 U21139 ( .B1(n18172), .B2(n18161), .A(n18160), .ZN(P3_U2860) );
  NOR2_X1 U21140 ( .A1(n18132), .A2(n18823), .ZN(n18164) );
  AOI211_X1 U21141 ( .C1(n18639), .C2(n18819), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18162), .ZN(n18163) );
  AOI211_X1 U21142 ( .C1(n18166), .C2(n18165), .A(n18164), .B(n18163), .ZN(
        n18171) );
  NOR3_X1 U21143 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18168), .A3(
        n18167), .ZN(n18177) );
  OAI21_X1 U21144 ( .B1(n18169), .B2(n18177), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18170) );
  OAI211_X1 U21145 ( .C1(n18173), .C2(n18172), .A(n18171), .B(n18170), .ZN(
        P3_U2861) );
  AOI211_X1 U21146 ( .C1(n18639), .C2(n18175), .A(n18174), .B(n18819), .ZN(
        n18176) );
  AOI211_X1 U21147 ( .C1(n18178), .C2(n18181), .A(n18177), .B(n18176), .ZN(
        n18180) );
  NAND2_X1 U21148 ( .A1(n18174), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18179) );
  OAI211_X1 U21149 ( .C1(n18182), .C2(n18181), .A(n18180), .B(n18179), .ZN(
        P3_U2862) );
  OAI211_X1 U21150 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18183), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18683)
         );
  OAI21_X1 U21151 ( .B1(n18186), .B2(n18184), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18185) );
  OAI221_X1 U21152 ( .B1(n18186), .B2(n18683), .C1(n18186), .C2(n18243), .A(
        n18185), .ZN(P3_U2863) );
  INV_X1 U21153 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18670) );
  NAND2_X1 U21154 ( .A1(n18670), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18352) );
  NAND2_X1 U21155 ( .A1(n18192), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18469) );
  INV_X1 U21156 ( .A(n18469), .ZN(n18420) );
  NAND2_X1 U21157 ( .A1(n18447), .A2(n18420), .ZN(n18492) );
  AND2_X1 U21158 ( .A1(n18352), .A2(n18492), .ZN(n18188) );
  OAI22_X1 U21159 ( .A1(n18189), .A2(n18670), .B1(n18188), .B2(n18187), .ZN(
        P3_U2866) );
  NOR2_X1 U21160 ( .A1(n18191), .A2(n18190), .ZN(P3_U2867) );
  NOR2_X1 U21161 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18654) );
  NAND2_X1 U21162 ( .A1(n18192), .A2(n18670), .ZN(n18289) );
  INV_X1 U21163 ( .A(n18289), .ZN(n18244) );
  NAND2_X1 U21164 ( .A1(n18654), .A2(n18244), .ZN(n18263) );
  NOR2_X1 U21165 ( .A1(n18194), .A2(n18193), .ZN(n18235) );
  NAND2_X1 U21166 ( .A1(n18235), .A2(n18195), .ZN(n18574) );
  NAND2_X1 U21167 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18200) );
  NOR2_X1 U21168 ( .A1(n18200), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18569) );
  NAND2_X1 U21169 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18569), .ZN(
        n18536) );
  INV_X1 U21170 ( .A(n18536), .ZN(n18614) );
  AND2_X1 U21171 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18570), .ZN(n18571) );
  NOR2_X2 U21172 ( .A1(n18265), .A2(n18196), .ZN(n18565) );
  NOR2_X1 U21173 ( .A1(n18670), .A2(n18378), .ZN(n18568) );
  NAND2_X1 U21174 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18568), .ZN(
        n18621) );
  NAND2_X1 U21175 ( .A1(n18621), .A2(n18263), .ZN(n18198) );
  INV_X1 U21176 ( .A(n18198), .ZN(n18267) );
  NOR2_X1 U21177 ( .A1(n18538), .A2(n18267), .ZN(n18238) );
  AOI22_X1 U21178 ( .A1(n18614), .A2(n18571), .B1(n18565), .B2(n18238), .ZN(
        n18202) );
  NAND2_X1 U21179 ( .A1(n18650), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18443) );
  INV_X1 U21180 ( .A(n18443), .ZN(n18197) );
  NOR2_X1 U21181 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18650), .ZN(
        n18421) );
  NOR2_X1 U21182 ( .A1(n18197), .A2(n18421), .ZN(n18493) );
  NOR2_X1 U21183 ( .A1(n18493), .A2(n18200), .ZN(n18537) );
  AOI21_X1 U21184 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18265), .ZN(n18445) );
  AOI22_X1 U21185 ( .A1(n18570), .A2(n18537), .B1(n18445), .B2(n18198), .ZN(
        n18240) );
  INV_X1 U21186 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18199) );
  NOR2_X2 U21187 ( .A1(n18266), .A2(n18199), .ZN(n18566) );
  NOR2_X2 U21188 ( .A1(n18200), .A2(n18443), .ZN(n18544) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18240), .B1(
        n18566), .B2(n18544), .ZN(n18201) );
  OAI211_X1 U21190 ( .C1(n18263), .C2(n18574), .A(n18202), .B(n18201), .ZN(
        P3_U2868) );
  NAND2_X1 U21191 ( .A1(n18235), .A2(n18203), .ZN(n18580) );
  INV_X1 U21192 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18204) );
  NOR2_X2 U21193 ( .A1(n18266), .A2(n18204), .ZN(n18577) );
  INV_X1 U21194 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18205) );
  NOR2_X2 U21195 ( .A1(n18265), .A2(n18205), .ZN(n18575) );
  AOI22_X1 U21196 ( .A1(n18544), .A2(n18577), .B1(n18238), .B2(n18575), .ZN(
        n18207) );
  AND2_X1 U21197 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18570), .ZN(n18576) );
  AOI22_X1 U21198 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18240), .B1(
        n18614), .B2(n18576), .ZN(n18206) );
  OAI211_X1 U21199 ( .C1(n18263), .C2(n18580), .A(n18207), .B(n18206), .ZN(
        P3_U2869) );
  NAND2_X1 U21200 ( .A1(n18235), .A2(n18208), .ZN(n18586) );
  INV_X1 U21201 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18209) );
  NOR2_X2 U21202 ( .A1(n18266), .A2(n18209), .ZN(n18582) );
  NOR2_X2 U21203 ( .A1(n18265), .A2(n18210), .ZN(n18581) );
  AOI22_X1 U21204 ( .A1(n18544), .A2(n18582), .B1(n18238), .B2(n18581), .ZN(
        n18212) );
  AND2_X1 U21205 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18570), .ZN(n18583) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18240), .B1(
        n18614), .B2(n18583), .ZN(n18211) );
  OAI211_X1 U21207 ( .C1(n18263), .C2(n18586), .A(n18212), .B(n18211), .ZN(
        P3_U2870) );
  INV_X1 U21208 ( .A(n18213), .ZN(n18214) );
  NAND2_X1 U21209 ( .A1(n18235), .A2(n18214), .ZN(n18592) );
  AND2_X1 U21210 ( .A1(n18570), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18588) );
  NOR2_X2 U21211 ( .A1(n18265), .A2(n18215), .ZN(n18587) );
  AOI22_X1 U21212 ( .A1(n18544), .A2(n18588), .B1(n18238), .B2(n18587), .ZN(
        n18218) );
  NOR2_X2 U21213 ( .A1(n18216), .A2(n18266), .ZN(n18589) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18240), .B1(
        n18614), .B2(n18589), .ZN(n18217) );
  OAI211_X1 U21215 ( .C1(n18263), .C2(n18592), .A(n18218), .B(n18217), .ZN(
        P3_U2871) );
  NAND2_X1 U21216 ( .A1(n18235), .A2(n18219), .ZN(n18598) );
  INV_X1 U21217 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18220) );
  NOR2_X2 U21218 ( .A1(n18266), .A2(n18220), .ZN(n18594) );
  NOR2_X2 U21219 ( .A1(n18265), .A2(n18221), .ZN(n18593) );
  AOI22_X1 U21220 ( .A1(n18544), .A2(n18594), .B1(n18238), .B2(n18593), .ZN(
        n18223) );
  AND2_X1 U21221 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18570), .ZN(n18595) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18240), .B1(
        n18614), .B2(n18595), .ZN(n18222) );
  OAI211_X1 U21223 ( .C1(n18263), .C2(n18598), .A(n18223), .B(n18222), .ZN(
        P3_U2872) );
  NAND2_X1 U21224 ( .A1(n18235), .A2(n18224), .ZN(n18604) );
  NOR2_X2 U21225 ( .A1(n18225), .A2(n18266), .ZN(n18600) );
  NOR2_X2 U21226 ( .A1(n18265), .A2(n18226), .ZN(n18599) );
  AOI22_X1 U21227 ( .A1(n18614), .A2(n18600), .B1(n18238), .B2(n18599), .ZN(
        n18228) );
  NOR2_X2 U21228 ( .A1(n18266), .A2(n19252), .ZN(n18601) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18240), .B1(
        n18544), .B2(n18601), .ZN(n18227) );
  OAI211_X1 U21230 ( .C1(n18263), .C2(n18604), .A(n18228), .B(n18227), .ZN(
        P3_U2873) );
  NAND2_X1 U21231 ( .A1(n18235), .A2(n18229), .ZN(n18610) );
  NOR2_X2 U21232 ( .A1(n18230), .A2(n18266), .ZN(n18606) );
  NOR2_X2 U21233 ( .A1(n18231), .A2(n18265), .ZN(n18605) );
  AOI22_X1 U21234 ( .A1(n18614), .A2(n18606), .B1(n18238), .B2(n18605), .ZN(
        n18233) );
  AND2_X1 U21235 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18570), .ZN(n18607) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18240), .B1(
        n18544), .B2(n18607), .ZN(n18232) );
  OAI211_X1 U21237 ( .C1(n18263), .C2(n18610), .A(n18233), .B(n18232), .ZN(
        P3_U2874) );
  NAND2_X1 U21238 ( .A1(n18235), .A2(n18234), .ZN(n18620) );
  NOR2_X2 U21239 ( .A1(n18266), .A2(n18236), .ZN(n18616) );
  NOR2_X2 U21240 ( .A1(n18237), .A2(n18265), .ZN(n18612) );
  AOI22_X1 U21241 ( .A1(n18614), .A2(n18616), .B1(n18238), .B2(n18612), .ZN(
        n18242) );
  NOR2_X2 U21242 ( .A1(n18239), .A2(n18266), .ZN(n18613) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18240), .B1(
        n18544), .B2(n18613), .ZN(n18241) );
  OAI211_X1 U21244 ( .C1(n18263), .C2(n18620), .A(n18242), .B(n18241), .ZN(
        P3_U2875) );
  NAND2_X1 U21245 ( .A1(n18244), .A2(n18421), .ZN(n18264) );
  INV_X1 U21246 ( .A(n18621), .ZN(n18284) );
  NAND2_X1 U21247 ( .A1(n18651), .A2(n18690), .ZN(n18422) );
  NOR2_X1 U21248 ( .A1(n18289), .A2(n18422), .ZN(n18259) );
  AOI22_X1 U21249 ( .A1(n18284), .A2(n18566), .B1(n18565), .B2(n18259), .ZN(
        n18246) );
  NAND2_X1 U21250 ( .A1(n18543), .A2(n18243), .ZN(n18376) );
  NOR2_X1 U21251 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18376), .ZN(
        n18331) );
  AOI22_X1 U21252 ( .A1(n18570), .A2(n18568), .B1(n18244), .B2(n18331), .ZN(
        n18260) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18260), .B1(
        n18544), .B2(n18571), .ZN(n18245) );
  OAI211_X1 U21254 ( .C1(n18574), .C2(n18264), .A(n18246), .B(n18245), .ZN(
        P3_U2876) );
  AOI22_X1 U21255 ( .A1(n18544), .A2(n18576), .B1(n18575), .B2(n18259), .ZN(
        n18248) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18260), .B1(
        n18284), .B2(n18577), .ZN(n18247) );
  OAI211_X1 U21257 ( .C1(n18580), .C2(n18264), .A(n18248), .B(n18247), .ZN(
        P3_U2877) );
  AOI22_X1 U21258 ( .A1(n18284), .A2(n18582), .B1(n18581), .B2(n18259), .ZN(
        n18250) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18260), .B1(
        n18544), .B2(n18583), .ZN(n18249) );
  OAI211_X1 U21260 ( .C1(n18586), .C2(n18264), .A(n18250), .B(n18249), .ZN(
        P3_U2878) );
  AOI22_X1 U21261 ( .A1(n18284), .A2(n18588), .B1(n18587), .B2(n18259), .ZN(
        n18252) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18260), .B1(
        n18544), .B2(n18589), .ZN(n18251) );
  OAI211_X1 U21263 ( .C1(n18592), .C2(n18264), .A(n18252), .B(n18251), .ZN(
        P3_U2879) );
  AOI22_X1 U21264 ( .A1(n18544), .A2(n18595), .B1(n18593), .B2(n18259), .ZN(
        n18254) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18260), .B1(
        n18284), .B2(n18594), .ZN(n18253) );
  OAI211_X1 U21266 ( .C1(n18598), .C2(n18264), .A(n18254), .B(n18253), .ZN(
        P3_U2880) );
  AOI22_X1 U21267 ( .A1(n18284), .A2(n18601), .B1(n18599), .B2(n18259), .ZN(
        n18256) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18260), .B1(
        n18544), .B2(n18600), .ZN(n18255) );
  OAI211_X1 U21269 ( .C1(n18604), .C2(n18264), .A(n18256), .B(n18255), .ZN(
        P3_U2881) );
  AOI22_X1 U21270 ( .A1(n18544), .A2(n18606), .B1(n18605), .B2(n18259), .ZN(
        n18258) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18260), .B1(
        n18284), .B2(n18607), .ZN(n18257) );
  OAI211_X1 U21272 ( .C1(n18610), .C2(n18264), .A(n18258), .B(n18257), .ZN(
        P3_U2882) );
  AOI22_X1 U21273 ( .A1(n18284), .A2(n18613), .B1(n18612), .B2(n18259), .ZN(
        n18262) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18260), .B1(
        n18544), .B2(n18616), .ZN(n18261) );
  OAI211_X1 U21275 ( .C1(n18620), .C2(n18264), .A(n18262), .B(n18261), .ZN(
        P3_U2883) );
  NOR2_X2 U21276 ( .A1(n18289), .A2(n18443), .ZN(n18348) );
  INV_X1 U21277 ( .A(n18348), .ZN(n18288) );
  INV_X1 U21278 ( .A(n18263), .ZN(n18306) );
  NOR2_X1 U21279 ( .A1(n18327), .A2(n18348), .ZN(n18310) );
  NOR2_X1 U21280 ( .A1(n18538), .A2(n18310), .ZN(n18283) );
  AOI22_X1 U21281 ( .A1(n18306), .A2(n18566), .B1(n18565), .B2(n18283), .ZN(
        n18270) );
  OAI22_X1 U21282 ( .A1(n18267), .A2(n18266), .B1(n18310), .B2(n18265), .ZN(
        n18268) );
  OAI21_X1 U21283 ( .B1(n18348), .B2(n18791), .A(n18268), .ZN(n18285) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18285), .B1(
        n18284), .B2(n18571), .ZN(n18269) );
  OAI211_X1 U21285 ( .C1(n18574), .C2(n18288), .A(n18270), .B(n18269), .ZN(
        P3_U2884) );
  AOI22_X1 U21286 ( .A1(n18284), .A2(n18576), .B1(n18575), .B2(n18283), .ZN(
        n18272) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18285), .B1(
        n18306), .B2(n18577), .ZN(n18271) );
  OAI211_X1 U21288 ( .C1(n18580), .C2(n18288), .A(n18272), .B(n18271), .ZN(
        P3_U2885) );
  AOI22_X1 U21289 ( .A1(n18306), .A2(n18582), .B1(n18581), .B2(n18283), .ZN(
        n18274) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18285), .B1(
        n18284), .B2(n18583), .ZN(n18273) );
  OAI211_X1 U21291 ( .C1(n18586), .C2(n18288), .A(n18274), .B(n18273), .ZN(
        P3_U2886) );
  AOI22_X1 U21292 ( .A1(n18306), .A2(n18588), .B1(n18587), .B2(n18283), .ZN(
        n18276) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18285), .B1(
        n18284), .B2(n18589), .ZN(n18275) );
  OAI211_X1 U21294 ( .C1(n18592), .C2(n18288), .A(n18276), .B(n18275), .ZN(
        P3_U2887) );
  AOI22_X1 U21295 ( .A1(n18284), .A2(n18595), .B1(n18593), .B2(n18283), .ZN(
        n18278) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18285), .B1(
        n18306), .B2(n18594), .ZN(n18277) );
  OAI211_X1 U21297 ( .C1(n18598), .C2(n18288), .A(n18278), .B(n18277), .ZN(
        P3_U2888) );
  AOI22_X1 U21298 ( .A1(n18284), .A2(n18600), .B1(n18599), .B2(n18283), .ZN(
        n18280) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18285), .B1(
        n18306), .B2(n18601), .ZN(n18279) );
  OAI211_X1 U21300 ( .C1(n18604), .C2(n18288), .A(n18280), .B(n18279), .ZN(
        P3_U2889) );
  AOI22_X1 U21301 ( .A1(n18306), .A2(n18607), .B1(n18605), .B2(n18283), .ZN(
        n18282) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18285), .B1(
        n18284), .B2(n18606), .ZN(n18281) );
  OAI211_X1 U21303 ( .C1(n18610), .C2(n18288), .A(n18282), .B(n18281), .ZN(
        P3_U2890) );
  AOI22_X1 U21304 ( .A1(n18306), .A2(n18613), .B1(n18612), .B2(n18283), .ZN(
        n18287) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18285), .B1(
        n18284), .B2(n18616), .ZN(n18286) );
  OAI211_X1 U21306 ( .C1(n18620), .C2(n18288), .A(n18287), .B(n18286), .ZN(
        P3_U2891) );
  NOR2_X1 U21307 ( .A1(n18651), .A2(n18289), .ZN(n18332) );
  NAND2_X1 U21308 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18332), .ZN(
        n18354) );
  AND2_X1 U21309 ( .A1(n18690), .A2(n18332), .ZN(n18305) );
  AOI22_X1 U21310 ( .A1(n18306), .A2(n18571), .B1(n18565), .B2(n18305), .ZN(
        n18292) );
  OAI21_X1 U21311 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18289), .A(n18354), 
        .ZN(n18290) );
  OAI211_X1 U21312 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18447), .A(
        n18543), .B(n18290), .ZN(n18307) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18307), .B1(
        n18566), .B2(n18327), .ZN(n18291) );
  OAI211_X1 U21314 ( .C1(n18574), .C2(n18354), .A(n18292), .B(n18291), .ZN(
        P3_U2892) );
  AOI22_X1 U21315 ( .A1(n18577), .A2(n18327), .B1(n18575), .B2(n18305), .ZN(
        n18294) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18576), .ZN(n18293) );
  OAI211_X1 U21317 ( .C1(n18580), .C2(n18354), .A(n18294), .B(n18293), .ZN(
        P3_U2893) );
  AOI22_X1 U21318 ( .A1(n18581), .A2(n18305), .B1(n18582), .B2(n18327), .ZN(
        n18296) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18583), .ZN(n18295) );
  OAI211_X1 U21320 ( .C1(n18586), .C2(n18354), .A(n18296), .B(n18295), .ZN(
        P3_U2894) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18307), .B1(
        n18587), .B2(n18305), .ZN(n18298) );
  AOI22_X1 U21322 ( .A1(n18306), .A2(n18589), .B1(n18588), .B2(n18327), .ZN(
        n18297) );
  OAI211_X1 U21323 ( .C1(n18592), .C2(n18354), .A(n18298), .B(n18297), .ZN(
        P3_U2895) );
  AOI22_X1 U21324 ( .A1(n18593), .A2(n18305), .B1(n18594), .B2(n18327), .ZN(
        n18300) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18595), .ZN(n18299) );
  OAI211_X1 U21326 ( .C1(n18598), .C2(n18354), .A(n18300), .B(n18299), .ZN(
        P3_U2896) );
  AOI22_X1 U21327 ( .A1(n18601), .A2(n18327), .B1(n18599), .B2(n18305), .ZN(
        n18302) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18600), .ZN(n18301) );
  OAI211_X1 U21329 ( .C1(n18604), .C2(n18354), .A(n18302), .B(n18301), .ZN(
        P3_U2897) );
  AOI22_X1 U21330 ( .A1(n18607), .A2(n18327), .B1(n18605), .B2(n18305), .ZN(
        n18304) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18606), .ZN(n18303) );
  OAI211_X1 U21332 ( .C1(n18610), .C2(n18354), .A(n18304), .B(n18303), .ZN(
        P3_U2898) );
  AOI22_X1 U21333 ( .A1(n18613), .A2(n18327), .B1(n18612), .B2(n18305), .ZN(
        n18309) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18616), .ZN(n18308) );
  OAI211_X1 U21335 ( .C1(n18620), .C2(n18354), .A(n18309), .B(n18308), .ZN(
        P3_U2899) );
  INV_X1 U21336 ( .A(n18352), .ZN(n18377) );
  NAND2_X1 U21337 ( .A1(n18654), .A2(n18377), .ZN(n18353) );
  AOI21_X1 U21338 ( .B1(n18354), .B2(n18353), .A(n18538), .ZN(n18326) );
  AOI22_X1 U21339 ( .A1(n18566), .A2(n18348), .B1(n18565), .B2(n18326), .ZN(
        n18313) );
  INV_X1 U21340 ( .A(n18353), .ZN(n18396) );
  AOI221_X1 U21341 ( .B1(n18310), .B2(n18354), .C1(n18540), .C2(n18354), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18311) );
  OAI21_X1 U21342 ( .B1(n18396), .B2(n18311), .A(n18543), .ZN(n18328) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18328), .B1(
        n18571), .B2(n18327), .ZN(n18312) );
  OAI211_X1 U21344 ( .C1(n18574), .C2(n18353), .A(n18313), .B(n18312), .ZN(
        P3_U2900) );
  AOI22_X1 U21345 ( .A1(n18577), .A2(n18348), .B1(n18575), .B2(n18326), .ZN(
        n18315) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18328), .B1(
        n18576), .B2(n18327), .ZN(n18314) );
  OAI211_X1 U21347 ( .C1(n18580), .C2(n18353), .A(n18315), .B(n18314), .ZN(
        P3_U2901) );
  AOI22_X1 U21348 ( .A1(n18583), .A2(n18327), .B1(n18581), .B2(n18326), .ZN(
        n18317) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18328), .B1(
        n18582), .B2(n18348), .ZN(n18316) );
  OAI211_X1 U21350 ( .C1(n18586), .C2(n18353), .A(n18317), .B(n18316), .ZN(
        P3_U2902) );
  AOI22_X1 U21351 ( .A1(n18589), .A2(n18327), .B1(n18587), .B2(n18326), .ZN(
        n18319) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18328), .B1(
        n18588), .B2(n18348), .ZN(n18318) );
  OAI211_X1 U21353 ( .C1(n18592), .C2(n18353), .A(n18319), .B(n18318), .ZN(
        P3_U2903) );
  AOI22_X1 U21354 ( .A1(n18593), .A2(n18326), .B1(n18594), .B2(n18348), .ZN(
        n18321) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18328), .B1(
        n18595), .B2(n18327), .ZN(n18320) );
  OAI211_X1 U21356 ( .C1(n18598), .C2(n18353), .A(n18321), .B(n18320), .ZN(
        P3_U2904) );
  AOI22_X1 U21357 ( .A1(n18600), .A2(n18327), .B1(n18599), .B2(n18326), .ZN(
        n18323) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18328), .B1(
        n18601), .B2(n18348), .ZN(n18322) );
  OAI211_X1 U21359 ( .C1(n18604), .C2(n18353), .A(n18323), .B(n18322), .ZN(
        P3_U2905) );
  AOI22_X1 U21360 ( .A1(n18607), .A2(n18348), .B1(n18605), .B2(n18326), .ZN(
        n18325) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18328), .B1(
        n18606), .B2(n18327), .ZN(n18324) );
  OAI211_X1 U21362 ( .C1(n18610), .C2(n18353), .A(n18325), .B(n18324), .ZN(
        P3_U2906) );
  AOI22_X1 U21363 ( .A1(n18613), .A2(n18348), .B1(n18612), .B2(n18326), .ZN(
        n18330) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18328), .B1(
        n18616), .B2(n18327), .ZN(n18329) );
  OAI211_X1 U21365 ( .C1(n18620), .C2(n18353), .A(n18330), .B(n18329), .ZN(
        P3_U2907) );
  NAND2_X1 U21366 ( .A1(n18421), .A2(n18377), .ZN(n18379) );
  NOR2_X1 U21367 ( .A1(n18422), .A2(n18352), .ZN(n18347) );
  AOI22_X1 U21368 ( .A1(n18571), .A2(n18348), .B1(n18565), .B2(n18347), .ZN(
        n18334) );
  AOI22_X1 U21369 ( .A1(n18570), .A2(n18332), .B1(n18331), .B2(n18377), .ZN(
        n18349) );
  INV_X1 U21370 ( .A(n18354), .ZN(n18371) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18349), .B1(
        n18566), .B2(n18371), .ZN(n18333) );
  OAI211_X1 U21372 ( .C1(n18574), .C2(n18379), .A(n18334), .B(n18333), .ZN(
        P3_U2908) );
  AOI22_X1 U21373 ( .A1(n18576), .A2(n18348), .B1(n18575), .B2(n18347), .ZN(
        n18336) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18349), .B1(
        n18577), .B2(n18371), .ZN(n18335) );
  OAI211_X1 U21375 ( .C1(n18580), .C2(n18379), .A(n18336), .B(n18335), .ZN(
        P3_U2909) );
  AOI22_X1 U21376 ( .A1(n18581), .A2(n18347), .B1(n18582), .B2(n18371), .ZN(
        n18338) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18349), .B1(
        n18583), .B2(n18348), .ZN(n18337) );
  OAI211_X1 U21378 ( .C1(n18586), .C2(n18379), .A(n18338), .B(n18337), .ZN(
        P3_U2910) );
  AOI22_X1 U21379 ( .A1(n18589), .A2(n18348), .B1(n18587), .B2(n18347), .ZN(
        n18340) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18349), .B1(
        n18588), .B2(n18371), .ZN(n18339) );
  OAI211_X1 U21381 ( .C1(n18592), .C2(n18379), .A(n18340), .B(n18339), .ZN(
        P3_U2911) );
  AOI22_X1 U21382 ( .A1(n18593), .A2(n18347), .B1(n18594), .B2(n18371), .ZN(
        n18342) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18349), .B1(
        n18595), .B2(n18348), .ZN(n18341) );
  OAI211_X1 U21384 ( .C1(n18598), .C2(n18379), .A(n18342), .B(n18341), .ZN(
        P3_U2912) );
  AOI22_X1 U21385 ( .A1(n18601), .A2(n18371), .B1(n18599), .B2(n18347), .ZN(
        n18344) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18349), .B1(
        n18600), .B2(n18348), .ZN(n18343) );
  OAI211_X1 U21387 ( .C1(n18604), .C2(n18379), .A(n18344), .B(n18343), .ZN(
        P3_U2913) );
  AOI22_X1 U21388 ( .A1(n18607), .A2(n18371), .B1(n18605), .B2(n18347), .ZN(
        n18346) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18349), .B1(
        n18606), .B2(n18348), .ZN(n18345) );
  OAI211_X1 U21390 ( .C1(n18610), .C2(n18379), .A(n18346), .B(n18345), .ZN(
        P3_U2914) );
  AOI22_X1 U21391 ( .A1(n18613), .A2(n18371), .B1(n18612), .B2(n18347), .ZN(
        n18351) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18349), .B1(
        n18616), .B2(n18348), .ZN(n18350) );
  OAI211_X1 U21393 ( .C1(n18620), .C2(n18379), .A(n18351), .B(n18350), .ZN(
        P3_U2915) );
  NOR2_X2 U21394 ( .A1(n18443), .A2(n18352), .ZN(n18439) );
  INV_X1 U21395 ( .A(n18439), .ZN(n18375) );
  NAND2_X1 U21396 ( .A1(n18379), .A2(n18375), .ZN(n18400) );
  AND2_X1 U21397 ( .A1(n18690), .A2(n18400), .ZN(n18370) );
  AOI22_X1 U21398 ( .A1(n18571), .A2(n18371), .B1(n18565), .B2(n18370), .ZN(
        n18357) );
  NAND2_X1 U21399 ( .A1(n18354), .A2(n18353), .ZN(n18355) );
  OAI221_X1 U21400 ( .B1(n18400), .B2(n18447), .C1(n18400), .C2(n18355), .A(
        n18445), .ZN(n18372) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18372), .B1(
        n18566), .B2(n18396), .ZN(n18356) );
  OAI211_X1 U21402 ( .C1(n18574), .C2(n18375), .A(n18357), .B(n18356), .ZN(
        P3_U2916) );
  AOI22_X1 U21403 ( .A1(n18576), .A2(n18371), .B1(n18575), .B2(n18370), .ZN(
        n18359) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18372), .B1(
        n18577), .B2(n18396), .ZN(n18358) );
  OAI211_X1 U21405 ( .C1(n18580), .C2(n18375), .A(n18359), .B(n18358), .ZN(
        P3_U2917) );
  AOI22_X1 U21406 ( .A1(n18581), .A2(n18370), .B1(n18582), .B2(n18396), .ZN(
        n18361) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18372), .B1(
        n18583), .B2(n18371), .ZN(n18360) );
  OAI211_X1 U21408 ( .C1(n18586), .C2(n18375), .A(n18361), .B(n18360), .ZN(
        P3_U2918) );
  AOI22_X1 U21409 ( .A1(n18588), .A2(n18396), .B1(n18587), .B2(n18370), .ZN(
        n18363) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18372), .B1(
        n18589), .B2(n18371), .ZN(n18362) );
  OAI211_X1 U21411 ( .C1(n18592), .C2(n18375), .A(n18363), .B(n18362), .ZN(
        P3_U2919) );
  AOI22_X1 U21412 ( .A1(n18595), .A2(n18371), .B1(n18593), .B2(n18370), .ZN(
        n18365) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18372), .B1(
        n18594), .B2(n18396), .ZN(n18364) );
  OAI211_X1 U21414 ( .C1(n18598), .C2(n18375), .A(n18365), .B(n18364), .ZN(
        P3_U2920) );
  AOI22_X1 U21415 ( .A1(n18600), .A2(n18371), .B1(n18599), .B2(n18370), .ZN(
        n18367) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18372), .B1(
        n18601), .B2(n18396), .ZN(n18366) );
  OAI211_X1 U21417 ( .C1(n18604), .C2(n18375), .A(n18367), .B(n18366), .ZN(
        P3_U2921) );
  AOI22_X1 U21418 ( .A1(n18607), .A2(n18396), .B1(n18605), .B2(n18370), .ZN(
        n18369) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18372), .B1(
        n18606), .B2(n18371), .ZN(n18368) );
  OAI211_X1 U21420 ( .C1(n18610), .C2(n18375), .A(n18369), .B(n18368), .ZN(
        P3_U2922) );
  AOI22_X1 U21421 ( .A1(n18613), .A2(n18396), .B1(n18612), .B2(n18370), .ZN(
        n18374) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18372), .B1(
        n18616), .B2(n18371), .ZN(n18373) );
  OAI211_X1 U21423 ( .C1(n18620), .C2(n18375), .A(n18374), .B(n18373), .ZN(
        P3_U2923) );
  INV_X1 U21424 ( .A(n18464), .ZN(n18399) );
  INV_X1 U21425 ( .A(n18376), .ZN(n18567) );
  OAI211_X1 U21426 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18447), .A(
        n18567), .B(n18377), .ZN(n18395) );
  NOR2_X1 U21427 ( .A1(n18378), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18423) );
  AND2_X1 U21428 ( .A1(n18690), .A2(n18423), .ZN(n18394) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18395), .B1(
        n18565), .B2(n18394), .ZN(n18381) );
  INV_X1 U21430 ( .A(n18379), .ZN(n18416) );
  AOI22_X1 U21431 ( .A1(n18566), .A2(n18416), .B1(n18571), .B2(n18396), .ZN(
        n18380) );
  OAI211_X1 U21432 ( .C1(n18574), .C2(n18399), .A(n18381), .B(n18380), .ZN(
        P3_U2924) );
  AOI22_X1 U21433 ( .A1(n18576), .A2(n18396), .B1(n18575), .B2(n18394), .ZN(
        n18383) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18395), .B1(
        n18577), .B2(n18416), .ZN(n18382) );
  OAI211_X1 U21435 ( .C1(n18580), .C2(n18399), .A(n18383), .B(n18382), .ZN(
        P3_U2925) );
  AOI22_X1 U21436 ( .A1(n18583), .A2(n18396), .B1(n18581), .B2(n18394), .ZN(
        n18385) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18395), .B1(
        n18582), .B2(n18416), .ZN(n18384) );
  OAI211_X1 U21438 ( .C1(n18586), .C2(n18399), .A(n18385), .B(n18384), .ZN(
        P3_U2926) );
  AOI22_X1 U21439 ( .A1(n18588), .A2(n18416), .B1(n18587), .B2(n18394), .ZN(
        n18387) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18395), .B1(
        n18589), .B2(n18396), .ZN(n18386) );
  OAI211_X1 U21441 ( .C1(n18592), .C2(n18399), .A(n18387), .B(n18386), .ZN(
        P3_U2927) );
  AOI22_X1 U21442 ( .A1(n18593), .A2(n18394), .B1(n18594), .B2(n18416), .ZN(
        n18389) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18395), .B1(
        n18595), .B2(n18396), .ZN(n18388) );
  OAI211_X1 U21444 ( .C1(n18598), .C2(n18399), .A(n18389), .B(n18388), .ZN(
        P3_U2928) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18395), .B1(
        n18599), .B2(n18394), .ZN(n18391) );
  AOI22_X1 U21446 ( .A1(n18601), .A2(n18416), .B1(n18600), .B2(n18396), .ZN(
        n18390) );
  OAI211_X1 U21447 ( .C1(n18604), .C2(n18399), .A(n18391), .B(n18390), .ZN(
        P3_U2929) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18395), .B1(
        n18605), .B2(n18394), .ZN(n18393) );
  AOI22_X1 U21449 ( .A1(n18607), .A2(n18416), .B1(n18606), .B2(n18396), .ZN(
        n18392) );
  OAI211_X1 U21450 ( .C1(n18610), .C2(n18399), .A(n18393), .B(n18392), .ZN(
        P3_U2930) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18395), .B1(
        n18612), .B2(n18394), .ZN(n18398) );
  AOI22_X1 U21452 ( .A1(n18613), .A2(n18416), .B1(n18616), .B2(n18396), .ZN(
        n18397) );
  OAI211_X1 U21453 ( .C1(n18620), .C2(n18399), .A(n18398), .B(n18397), .ZN(
        P3_U2931) );
  NAND2_X1 U21454 ( .A1(n18654), .A2(n18420), .ZN(n18444) );
  NAND2_X1 U21455 ( .A1(n18399), .A2(n18444), .ZN(n18446) );
  AND2_X1 U21456 ( .A1(n18690), .A2(n18446), .ZN(n18415) );
  AOI22_X1 U21457 ( .A1(n18571), .A2(n18416), .B1(n18565), .B2(n18415), .ZN(
        n18402) );
  OAI221_X1 U21458 ( .B1(n18446), .B2(n18447), .C1(n18446), .C2(n18400), .A(
        n18445), .ZN(n18417) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18417), .B1(
        n18566), .B2(n18439), .ZN(n18401) );
  OAI211_X1 U21460 ( .C1(n18574), .C2(n18444), .A(n18402), .B(n18401), .ZN(
        P3_U2932) );
  AOI22_X1 U21461 ( .A1(n18576), .A2(n18416), .B1(n18575), .B2(n18415), .ZN(
        n18404) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18417), .B1(
        n18577), .B2(n18439), .ZN(n18403) );
  OAI211_X1 U21463 ( .C1(n18580), .C2(n18444), .A(n18404), .B(n18403), .ZN(
        P3_U2933) );
  AOI22_X1 U21464 ( .A1(n18583), .A2(n18416), .B1(n18581), .B2(n18415), .ZN(
        n18406) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18417), .B1(
        n18582), .B2(n18439), .ZN(n18405) );
  OAI211_X1 U21466 ( .C1(n18586), .C2(n18444), .A(n18406), .B(n18405), .ZN(
        P3_U2934) );
  AOI22_X1 U21467 ( .A1(n18588), .A2(n18439), .B1(n18587), .B2(n18415), .ZN(
        n18408) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18417), .B1(
        n18589), .B2(n18416), .ZN(n18407) );
  OAI211_X1 U21469 ( .C1(n18592), .C2(n18444), .A(n18408), .B(n18407), .ZN(
        P3_U2935) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18417), .B1(
        n18593), .B2(n18415), .ZN(n18410) );
  AOI22_X1 U21471 ( .A1(n18595), .A2(n18416), .B1(n18594), .B2(n18439), .ZN(
        n18409) );
  OAI211_X1 U21472 ( .C1(n18598), .C2(n18444), .A(n18410), .B(n18409), .ZN(
        P3_U2936) );
  AOI22_X1 U21473 ( .A1(n18600), .A2(n18416), .B1(n18599), .B2(n18415), .ZN(
        n18412) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18417), .B1(
        n18601), .B2(n18439), .ZN(n18411) );
  OAI211_X1 U21475 ( .C1(n18604), .C2(n18444), .A(n18412), .B(n18411), .ZN(
        P3_U2937) );
  AOI22_X1 U21476 ( .A1(n18606), .A2(n18416), .B1(n18605), .B2(n18415), .ZN(
        n18414) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18417), .B1(
        n18607), .B2(n18439), .ZN(n18413) );
  OAI211_X1 U21478 ( .C1(n18610), .C2(n18444), .A(n18414), .B(n18413), .ZN(
        P3_U2938) );
  AOI22_X1 U21479 ( .A1(n18616), .A2(n18416), .B1(n18612), .B2(n18415), .ZN(
        n18419) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18417), .B1(
        n18613), .B2(n18439), .ZN(n18418) );
  OAI211_X1 U21481 ( .C1(n18620), .C2(n18444), .A(n18419), .B(n18418), .ZN(
        P3_U2939) );
  NAND2_X1 U21482 ( .A1(n18421), .A2(n18420), .ZN(n18470) );
  NOR2_X1 U21483 ( .A1(n18422), .A2(n18469), .ZN(n18438) );
  AOI22_X1 U21484 ( .A1(n18566), .A2(n18464), .B1(n18565), .B2(n18438), .ZN(
        n18425) );
  NOR2_X1 U21485 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18469), .ZN(
        n18471) );
  AOI22_X1 U21486 ( .A1(n18570), .A2(n18423), .B1(n18567), .B2(n18471), .ZN(
        n18440) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18440), .B1(
        n18571), .B2(n18439), .ZN(n18424) );
  OAI211_X1 U21488 ( .C1(n18574), .C2(n18470), .A(n18425), .B(n18424), .ZN(
        P3_U2940) );
  AOI22_X1 U21489 ( .A1(n18576), .A2(n18439), .B1(n18575), .B2(n18438), .ZN(
        n18427) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18440), .B1(
        n18577), .B2(n18464), .ZN(n18426) );
  OAI211_X1 U21491 ( .C1(n18580), .C2(n18470), .A(n18427), .B(n18426), .ZN(
        P3_U2941) );
  AOI22_X1 U21492 ( .A1(n18581), .A2(n18438), .B1(n18582), .B2(n18464), .ZN(
        n18429) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18440), .B1(
        n18583), .B2(n18439), .ZN(n18428) );
  OAI211_X1 U21494 ( .C1(n18586), .C2(n18470), .A(n18429), .B(n18428), .ZN(
        P3_U2942) );
  AOI22_X1 U21495 ( .A1(n18588), .A2(n18464), .B1(n18587), .B2(n18438), .ZN(
        n18431) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18440), .B1(
        n18589), .B2(n18439), .ZN(n18430) );
  OAI211_X1 U21497 ( .C1(n18592), .C2(n18470), .A(n18431), .B(n18430), .ZN(
        P3_U2943) );
  AOI22_X1 U21498 ( .A1(n18593), .A2(n18438), .B1(n18594), .B2(n18464), .ZN(
        n18433) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18440), .B1(
        n18595), .B2(n18439), .ZN(n18432) );
  OAI211_X1 U21500 ( .C1(n18598), .C2(n18470), .A(n18433), .B(n18432), .ZN(
        P3_U2944) );
  AOI22_X1 U21501 ( .A1(n18600), .A2(n18439), .B1(n18599), .B2(n18438), .ZN(
        n18435) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18440), .B1(
        n18601), .B2(n18464), .ZN(n18434) );
  OAI211_X1 U21503 ( .C1(n18604), .C2(n18470), .A(n18435), .B(n18434), .ZN(
        P3_U2945) );
  AOI22_X1 U21504 ( .A1(n18607), .A2(n18464), .B1(n18605), .B2(n18438), .ZN(
        n18437) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18440), .B1(
        n18606), .B2(n18439), .ZN(n18436) );
  OAI211_X1 U21506 ( .C1(n18610), .C2(n18470), .A(n18437), .B(n18436), .ZN(
        P3_U2946) );
  AOI22_X1 U21507 ( .A1(n18613), .A2(n18464), .B1(n18612), .B2(n18438), .ZN(
        n18442) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18440), .B1(
        n18616), .B2(n18439), .ZN(n18441) );
  OAI211_X1 U21509 ( .C1(n18620), .C2(n18470), .A(n18442), .B(n18441), .ZN(
        P3_U2947) );
  NOR2_X2 U21510 ( .A1(n18443), .A2(n18469), .ZN(n18532) );
  INV_X1 U21511 ( .A(n18532), .ZN(n18468) );
  INV_X1 U21512 ( .A(n18444), .ZN(n18487) );
  AOI21_X1 U21513 ( .B1(n18470), .B2(n18468), .A(n18538), .ZN(n18463) );
  AOI22_X1 U21514 ( .A1(n18566), .A2(n18487), .B1(n18565), .B2(n18463), .ZN(
        n18450) );
  NAND2_X1 U21515 ( .A1(n18470), .A2(n18468), .ZN(n18448) );
  OAI221_X1 U21516 ( .B1(n18448), .B2(n18447), .C1(n18448), .C2(n18446), .A(
        n18445), .ZN(n18465) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18465), .B1(
        n18571), .B2(n18464), .ZN(n18449) );
  OAI211_X1 U21518 ( .C1(n18574), .C2(n18468), .A(n18450), .B(n18449), .ZN(
        P3_U2948) );
  AOI22_X1 U21519 ( .A1(n18576), .A2(n18464), .B1(n18575), .B2(n18463), .ZN(
        n18452) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18465), .B1(
        n18577), .B2(n18487), .ZN(n18451) );
  OAI211_X1 U21521 ( .C1(n18580), .C2(n18468), .A(n18452), .B(n18451), .ZN(
        P3_U2949) );
  AOI22_X1 U21522 ( .A1(n18583), .A2(n18464), .B1(n18581), .B2(n18463), .ZN(
        n18454) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18465), .B1(
        n18582), .B2(n18487), .ZN(n18453) );
  OAI211_X1 U21524 ( .C1(n18586), .C2(n18468), .A(n18454), .B(n18453), .ZN(
        P3_U2950) );
  AOI22_X1 U21525 ( .A1(n18589), .A2(n18464), .B1(n18587), .B2(n18463), .ZN(
        n18456) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18465), .B1(
        n18588), .B2(n18487), .ZN(n18455) );
  OAI211_X1 U21527 ( .C1(n18592), .C2(n18468), .A(n18456), .B(n18455), .ZN(
        P3_U2951) );
  AOI22_X1 U21528 ( .A1(n18595), .A2(n18464), .B1(n18593), .B2(n18463), .ZN(
        n18458) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18465), .B1(
        n18594), .B2(n18487), .ZN(n18457) );
  OAI211_X1 U21530 ( .C1(n18598), .C2(n18468), .A(n18458), .B(n18457), .ZN(
        P3_U2952) );
  AOI22_X1 U21531 ( .A1(n18600), .A2(n18464), .B1(n18599), .B2(n18463), .ZN(
        n18460) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18465), .B1(
        n18601), .B2(n18487), .ZN(n18459) );
  OAI211_X1 U21533 ( .C1(n18604), .C2(n18468), .A(n18460), .B(n18459), .ZN(
        P3_U2953) );
  AOI22_X1 U21534 ( .A1(n18607), .A2(n18487), .B1(n18605), .B2(n18463), .ZN(
        n18462) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18465), .B1(
        n18606), .B2(n18464), .ZN(n18461) );
  OAI211_X1 U21536 ( .C1(n18610), .C2(n18468), .A(n18462), .B(n18461), .ZN(
        P3_U2954) );
  AOI22_X1 U21537 ( .A1(n18613), .A2(n18487), .B1(n18612), .B2(n18463), .ZN(
        n18467) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18465), .B1(
        n18616), .B2(n18464), .ZN(n18466) );
  OAI211_X1 U21539 ( .C1(n18620), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2955) );
  NOR2_X1 U21540 ( .A1(n18651), .A2(n18469), .ZN(n18516) );
  NAND2_X1 U21541 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18516), .ZN(
        n18491) );
  INV_X1 U21542 ( .A(n18470), .ZN(n18511) );
  AND2_X1 U21543 ( .A1(n18690), .A2(n18516), .ZN(n18486) );
  AOI22_X1 U21544 ( .A1(n18566), .A2(n18511), .B1(n18565), .B2(n18486), .ZN(
        n18473) );
  AOI22_X1 U21545 ( .A1(n18570), .A2(n18471), .B1(n18567), .B2(n18516), .ZN(
        n18488) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18488), .B1(
        n18571), .B2(n18487), .ZN(n18472) );
  OAI211_X1 U21547 ( .C1(n18574), .C2(n18491), .A(n18473), .B(n18472), .ZN(
        P3_U2956) );
  AOI22_X1 U21548 ( .A1(n18576), .A2(n18487), .B1(n18575), .B2(n18486), .ZN(
        n18475) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18488), .B1(
        n18577), .B2(n18511), .ZN(n18474) );
  OAI211_X1 U21550 ( .C1(n18580), .C2(n18491), .A(n18475), .B(n18474), .ZN(
        P3_U2957) );
  AOI22_X1 U21551 ( .A1(n18583), .A2(n18487), .B1(n18581), .B2(n18486), .ZN(
        n18477) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18488), .B1(
        n18582), .B2(n18511), .ZN(n18476) );
  OAI211_X1 U21553 ( .C1(n18586), .C2(n18491), .A(n18477), .B(n18476), .ZN(
        P3_U2958) );
  AOI22_X1 U21554 ( .A1(n18589), .A2(n18487), .B1(n18587), .B2(n18486), .ZN(
        n18479) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18488), .B1(
        n18588), .B2(n18511), .ZN(n18478) );
  OAI211_X1 U21556 ( .C1(n18592), .C2(n18491), .A(n18479), .B(n18478), .ZN(
        P3_U2959) );
  AOI22_X1 U21557 ( .A1(n18595), .A2(n18487), .B1(n18593), .B2(n18486), .ZN(
        n18481) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18488), .B1(
        n18594), .B2(n18511), .ZN(n18480) );
  OAI211_X1 U21559 ( .C1(n18598), .C2(n18491), .A(n18481), .B(n18480), .ZN(
        P3_U2960) );
  AOI22_X1 U21560 ( .A1(n18600), .A2(n18487), .B1(n18599), .B2(n18486), .ZN(
        n18483) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18488), .B1(
        n18601), .B2(n18511), .ZN(n18482) );
  OAI211_X1 U21562 ( .C1(n18604), .C2(n18491), .A(n18483), .B(n18482), .ZN(
        P3_U2961) );
  AOI22_X1 U21563 ( .A1(n18606), .A2(n18487), .B1(n18605), .B2(n18486), .ZN(
        n18485) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18488), .B1(
        n18607), .B2(n18511), .ZN(n18484) );
  OAI211_X1 U21565 ( .C1(n18610), .C2(n18491), .A(n18485), .B(n18484), .ZN(
        P3_U2962) );
  AOI22_X1 U21566 ( .A1(n18613), .A2(n18511), .B1(n18612), .B2(n18486), .ZN(
        n18490) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18488), .B1(
        n18616), .B2(n18487), .ZN(n18489) );
  OAI211_X1 U21568 ( .C1(n18620), .C2(n18491), .A(n18490), .B(n18489), .ZN(
        P3_U2963) );
  INV_X1 U21569 ( .A(n18569), .ZN(n18515) );
  NOR2_X2 U21570 ( .A1(n18515), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18615) );
  INV_X1 U21571 ( .A(n18615), .ZN(n18514) );
  NOR2_X1 U21572 ( .A1(n18560), .A2(n18615), .ZN(n18541) );
  NOR2_X1 U21573 ( .A1(n18538), .A2(n18541), .ZN(n18509) );
  AOI22_X1 U21574 ( .A1(n18566), .A2(n18532), .B1(n18565), .B2(n18509), .ZN(
        n18496) );
  OAI21_X1 U21575 ( .B1(n18493), .B2(n18492), .A(n18541), .ZN(n18494) );
  OAI211_X1 U21576 ( .C1(n18615), .C2(n18791), .A(n18543), .B(n18494), .ZN(
        n18510) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18510), .B1(
        n18571), .B2(n18511), .ZN(n18495) );
  OAI211_X1 U21578 ( .C1(n18574), .C2(n18514), .A(n18496), .B(n18495), .ZN(
        P3_U2964) );
  AOI22_X1 U21579 ( .A1(n18576), .A2(n18511), .B1(n18575), .B2(n18509), .ZN(
        n18498) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18510), .B1(
        n18577), .B2(n18532), .ZN(n18497) );
  OAI211_X1 U21581 ( .C1(n18580), .C2(n18514), .A(n18498), .B(n18497), .ZN(
        P3_U2965) );
  AOI22_X1 U21582 ( .A1(n18581), .A2(n18509), .B1(n18582), .B2(n18532), .ZN(
        n18500) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18510), .B1(
        n18583), .B2(n18511), .ZN(n18499) );
  OAI211_X1 U21584 ( .C1(n18586), .C2(n18514), .A(n18500), .B(n18499), .ZN(
        P3_U2966) );
  AOI22_X1 U21585 ( .A1(n18588), .A2(n18532), .B1(n18587), .B2(n18509), .ZN(
        n18502) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18510), .B1(
        n18589), .B2(n18511), .ZN(n18501) );
  OAI211_X1 U21587 ( .C1(n18592), .C2(n18514), .A(n18502), .B(n18501), .ZN(
        P3_U2967) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18510), .B1(
        n18593), .B2(n18509), .ZN(n18504) );
  AOI22_X1 U21589 ( .A1(n18595), .A2(n18511), .B1(n18594), .B2(n18532), .ZN(
        n18503) );
  OAI211_X1 U21590 ( .C1(n18598), .C2(n18514), .A(n18504), .B(n18503), .ZN(
        P3_U2968) );
  AOI22_X1 U21591 ( .A1(n18600), .A2(n18511), .B1(n18599), .B2(n18509), .ZN(
        n18506) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18510), .B1(
        n18601), .B2(n18532), .ZN(n18505) );
  OAI211_X1 U21593 ( .C1(n18604), .C2(n18514), .A(n18506), .B(n18505), .ZN(
        P3_U2969) );
  AOI22_X1 U21594 ( .A1(n18606), .A2(n18511), .B1(n18605), .B2(n18509), .ZN(
        n18508) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18510), .B1(
        n18607), .B2(n18532), .ZN(n18507) );
  OAI211_X1 U21596 ( .C1(n18610), .C2(n18514), .A(n18508), .B(n18507), .ZN(
        P3_U2970) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18510), .B1(
        n18612), .B2(n18509), .ZN(n18513) );
  AOI22_X1 U21598 ( .A1(n18613), .A2(n18532), .B1(n18616), .B2(n18511), .ZN(
        n18512) );
  OAI211_X1 U21599 ( .C1(n18620), .C2(n18514), .A(n18513), .B(n18512), .ZN(
        P3_U2971) );
  NOR2_X1 U21600 ( .A1(n18538), .A2(n18515), .ZN(n18531) );
  AOI22_X1 U21601 ( .A1(n18566), .A2(n18560), .B1(n18565), .B2(n18531), .ZN(
        n18518) );
  AOI22_X1 U21602 ( .A1(n18570), .A2(n18516), .B1(n18569), .B2(n18567), .ZN(
        n18533) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18533), .B1(
        n18571), .B2(n18532), .ZN(n18517) );
  OAI211_X1 U21604 ( .C1(n18574), .C2(n18536), .A(n18518), .B(n18517), .ZN(
        P3_U2972) );
  AOI22_X1 U21605 ( .A1(n18577), .A2(n18560), .B1(n18575), .B2(n18531), .ZN(
        n18520) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18533), .B1(
        n18576), .B2(n18532), .ZN(n18519) );
  OAI211_X1 U21607 ( .C1(n18536), .C2(n18580), .A(n18520), .B(n18519), .ZN(
        P3_U2973) );
  AOI22_X1 U21608 ( .A1(n18583), .A2(n18532), .B1(n18581), .B2(n18531), .ZN(
        n18522) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18533), .B1(
        n18582), .B2(n18560), .ZN(n18521) );
  OAI211_X1 U21610 ( .C1(n18536), .C2(n18586), .A(n18522), .B(n18521), .ZN(
        P3_U2974) );
  AOI22_X1 U21611 ( .A1(n18589), .A2(n18532), .B1(n18587), .B2(n18531), .ZN(
        n18524) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18533), .B1(
        n18588), .B2(n18560), .ZN(n18523) );
  OAI211_X1 U21613 ( .C1(n18536), .C2(n18592), .A(n18524), .B(n18523), .ZN(
        P3_U2975) );
  AOI22_X1 U21614 ( .A1(n18595), .A2(n18532), .B1(n18593), .B2(n18531), .ZN(
        n18526) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18533), .B1(
        n18594), .B2(n18560), .ZN(n18525) );
  OAI211_X1 U21616 ( .C1(n18536), .C2(n18598), .A(n18526), .B(n18525), .ZN(
        P3_U2976) );
  AOI22_X1 U21617 ( .A1(n18600), .A2(n18532), .B1(n18599), .B2(n18531), .ZN(
        n18528) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18533), .B1(
        n18601), .B2(n18560), .ZN(n18527) );
  OAI211_X1 U21619 ( .C1(n18536), .C2(n18604), .A(n18528), .B(n18527), .ZN(
        P3_U2977) );
  AOI22_X1 U21620 ( .A1(n18606), .A2(n18532), .B1(n18605), .B2(n18531), .ZN(
        n18530) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18533), .B1(
        n18607), .B2(n18560), .ZN(n18529) );
  OAI211_X1 U21622 ( .C1(n18536), .C2(n18610), .A(n18530), .B(n18529), .ZN(
        P3_U2978) );
  AOI22_X1 U21623 ( .A1(n18613), .A2(n18560), .B1(n18612), .B2(n18531), .ZN(
        n18535) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18533), .B1(
        n18616), .B2(n18532), .ZN(n18534) );
  OAI211_X1 U21625 ( .C1(n18536), .C2(n18620), .A(n18535), .B(n18534), .ZN(
        P3_U2979) );
  INV_X1 U21626 ( .A(n18544), .ZN(n18564) );
  INV_X1 U21627 ( .A(n18537), .ZN(n18539) );
  NOR2_X1 U21628 ( .A1(n18538), .A2(n18539), .ZN(n18559) );
  AOI22_X1 U21629 ( .A1(n18571), .A2(n18560), .B1(n18565), .B2(n18559), .ZN(
        n18546) );
  OAI21_X1 U21630 ( .B1(n18541), .B2(n18540), .A(n18539), .ZN(n18542) );
  OAI211_X1 U21631 ( .C1(n18544), .C2(n18791), .A(n18543), .B(n18542), .ZN(
        n18561) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18561), .B1(
        n18566), .B2(n18615), .ZN(n18545) );
  OAI211_X1 U21633 ( .C1(n18564), .C2(n18574), .A(n18546), .B(n18545), .ZN(
        P3_U2980) );
  AOI22_X1 U21634 ( .A1(n18576), .A2(n18560), .B1(n18575), .B2(n18559), .ZN(
        n18548) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18561), .B1(
        n18577), .B2(n18615), .ZN(n18547) );
  OAI211_X1 U21636 ( .C1(n18564), .C2(n18580), .A(n18548), .B(n18547), .ZN(
        P3_U2981) );
  AOI22_X1 U21637 ( .A1(n18581), .A2(n18559), .B1(n18582), .B2(n18615), .ZN(
        n18550) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18561), .B1(
        n18583), .B2(n18560), .ZN(n18549) );
  OAI211_X1 U21639 ( .C1(n18564), .C2(n18586), .A(n18550), .B(n18549), .ZN(
        P3_U2982) );
  AOI22_X1 U21640 ( .A1(n18589), .A2(n18560), .B1(n18587), .B2(n18559), .ZN(
        n18552) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18561), .B1(
        n18588), .B2(n18615), .ZN(n18551) );
  OAI211_X1 U21642 ( .C1(n18564), .C2(n18592), .A(n18552), .B(n18551), .ZN(
        P3_U2983) );
  AOI22_X1 U21643 ( .A1(n18593), .A2(n18559), .B1(n18594), .B2(n18615), .ZN(
        n18554) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18561), .B1(
        n18595), .B2(n18560), .ZN(n18553) );
  OAI211_X1 U21645 ( .C1(n18564), .C2(n18598), .A(n18554), .B(n18553), .ZN(
        P3_U2984) );
  AOI22_X1 U21646 ( .A1(n18601), .A2(n18615), .B1(n18599), .B2(n18559), .ZN(
        n18556) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18561), .B1(
        n18600), .B2(n18560), .ZN(n18555) );
  OAI211_X1 U21648 ( .C1(n18564), .C2(n18604), .A(n18556), .B(n18555), .ZN(
        P3_U2985) );
  AOI22_X1 U21649 ( .A1(n18607), .A2(n18615), .B1(n18605), .B2(n18559), .ZN(
        n18558) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18561), .B1(
        n18606), .B2(n18560), .ZN(n18557) );
  OAI211_X1 U21651 ( .C1(n18564), .C2(n18610), .A(n18558), .B(n18557), .ZN(
        P3_U2986) );
  AOI22_X1 U21652 ( .A1(n18613), .A2(n18615), .B1(n18612), .B2(n18559), .ZN(
        n18563) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18561), .B1(
        n18616), .B2(n18560), .ZN(n18562) );
  OAI211_X1 U21654 ( .C1(n18564), .C2(n18620), .A(n18563), .B(n18562), .ZN(
        P3_U2987) );
  AND2_X1 U21655 ( .A1(n18690), .A2(n18568), .ZN(n18611) );
  AOI22_X1 U21656 ( .A1(n18566), .A2(n18614), .B1(n18565), .B2(n18611), .ZN(
        n18573) );
  AOI22_X1 U21657 ( .A1(n18570), .A2(n18569), .B1(n18568), .B2(n18567), .ZN(
        n18617) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18617), .B1(
        n18571), .B2(n18615), .ZN(n18572) );
  OAI211_X1 U21659 ( .C1(n18621), .C2(n18574), .A(n18573), .B(n18572), .ZN(
        P3_U2988) );
  AOI22_X1 U21660 ( .A1(n18576), .A2(n18615), .B1(n18575), .B2(n18611), .ZN(
        n18579) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18617), .B1(
        n18614), .B2(n18577), .ZN(n18578) );
  OAI211_X1 U21662 ( .C1(n18621), .C2(n18580), .A(n18579), .B(n18578), .ZN(
        P3_U2989) );
  AOI22_X1 U21663 ( .A1(n18614), .A2(n18582), .B1(n18581), .B2(n18611), .ZN(
        n18585) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18617), .B1(
        n18583), .B2(n18615), .ZN(n18584) );
  OAI211_X1 U21665 ( .C1(n18621), .C2(n18586), .A(n18585), .B(n18584), .ZN(
        P3_U2990) );
  AOI22_X1 U21666 ( .A1(n18614), .A2(n18588), .B1(n18587), .B2(n18611), .ZN(
        n18591) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18617), .B1(
        n18589), .B2(n18615), .ZN(n18590) );
  OAI211_X1 U21668 ( .C1(n18621), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U2991) );
  AOI22_X1 U21669 ( .A1(n18614), .A2(n18594), .B1(n18593), .B2(n18611), .ZN(
        n18597) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18617), .B1(
        n18595), .B2(n18615), .ZN(n18596) );
  OAI211_X1 U21671 ( .C1(n18621), .C2(n18598), .A(n18597), .B(n18596), .ZN(
        P3_U2992) );
  AOI22_X1 U21672 ( .A1(n18600), .A2(n18615), .B1(n18599), .B2(n18611), .ZN(
        n18603) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18617), .B1(
        n18614), .B2(n18601), .ZN(n18602) );
  OAI211_X1 U21674 ( .C1(n18621), .C2(n18604), .A(n18603), .B(n18602), .ZN(
        P3_U2993) );
  AOI22_X1 U21675 ( .A1(n18606), .A2(n18615), .B1(n18605), .B2(n18611), .ZN(
        n18609) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18617), .B1(
        n18614), .B2(n18607), .ZN(n18608) );
  OAI211_X1 U21677 ( .C1(n18621), .C2(n18610), .A(n18609), .B(n18608), .ZN(
        P3_U2994) );
  AOI22_X1 U21678 ( .A1(n18614), .A2(n18613), .B1(n18612), .B2(n18611), .ZN(
        n18619) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18617), .B1(
        n18616), .B2(n18615), .ZN(n18618) );
  OAI211_X1 U21680 ( .C1(n18621), .C2(n18620), .A(n18619), .B(n18618), .ZN(
        P3_U2995) );
  AOI21_X1 U21681 ( .B1(n18624), .B2(n18623), .A(n18622), .ZN(n18626) );
  OAI21_X1 U21682 ( .B1(n18627), .B2(n18626), .A(n18625), .ZN(n18628) );
  OAI221_X1 U21683 ( .B1(n18630), .B2(n18665), .C1(n18630), .C2(n18629), .A(
        n18628), .ZN(n18834) );
  AOI221_X1 U21684 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18632), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18632), .A(n18631), .ZN(n18676) );
  INV_X1 U21685 ( .A(n18678), .ZN(n18666) );
  OAI21_X1 U21686 ( .B1(n18635), .B2(n18634), .A(n18633), .ZN(n18662) );
  AOI22_X1 U21687 ( .A1(n18808), .A2(n18661), .B1(n18636), .B2(n18662), .ZN(
        n18637) );
  OAI21_X1 U21688 ( .B1(n18638), .B2(n18639), .A(n18637), .ZN(n18797) );
  NOR2_X1 U21689 ( .A1(n18798), .A2(n18797), .ZN(n18644) );
  AND2_X1 U21690 ( .A1(n18808), .A2(n18661), .ZN(n18642) );
  NAND2_X1 U21691 ( .A1(n18639), .A2(n20913), .ZN(n18646) );
  INV_X1 U21692 ( .A(n18646), .ZN(n18641) );
  OAI22_X1 U21693 ( .A1(n18642), .A2(n18665), .B1(n18641), .B2(n18640), .ZN(
        n18794) );
  AOI21_X1 U21694 ( .B1(n18794), .B2(n18666), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18643) );
  AOI21_X1 U21695 ( .B1(n18666), .B2(n18644), .A(n18643), .ZN(n18673) );
  NAND2_X1 U21696 ( .A1(n18657), .A2(n18645), .ZN(n18647) );
  AOI22_X1 U21697 ( .A1(n18812), .A2(n18647), .B1(n18815), .B2(n18646), .ZN(
        n18809) );
  AOI22_X1 U21698 ( .A1(n18649), .A2(n18648), .B1(n18647), .B2(n20913), .ZN(
        n18652) );
  INV_X1 U21699 ( .A(n18652), .ZN(n18817) );
  NOR3_X1 U21700 ( .A1(n18651), .A2(n18650), .A3(n18817), .ZN(n18653) );
  OAI22_X1 U21701 ( .A1(n18809), .A2(n18653), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18652), .ZN(n18655) );
  AOI21_X1 U21702 ( .B1(n18655), .B2(n18666), .A(n18654), .ZN(n18668) );
  OAI21_X1 U21703 ( .B1(n18657), .B2(n20913), .A(n18656), .ZN(n18659) );
  NAND2_X1 U21704 ( .A1(n18815), .A2(n18808), .ZN(n18658) );
  OAI221_X1 U21705 ( .B1(n18815), .B2(n18808), .C1(n18660), .C2(n18659), .A(
        n18658), .ZN(n18664) );
  NAND3_X1 U21706 ( .A1(n18662), .A2(n18661), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18663) );
  OAI211_X1 U21707 ( .C1(n18804), .C2(n18665), .A(n18664), .B(n18663), .ZN(
        n18806) );
  AOI22_X1 U21708 ( .A1(n18678), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18806), .B2(n18666), .ZN(n18669) );
  OR2_X1 U21709 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18669), .ZN(
        n18667) );
  AOI221_X1 U21710 ( .B1(n18668), .B2(n18667), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18669), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18672) );
  OAI21_X1 U21711 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18669), .ZN(n18671) );
  AOI222_X1 U21712 ( .A1(n18673), .A2(n18672), .B1(n18673), .B2(n18671), .C1(
        n18672), .C2(n18670), .ZN(n18675) );
  NAND3_X1 U21713 ( .A1(n18676), .A2(n18675), .A3(n18674), .ZN(n18677) );
  AOI211_X1 U21714 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18678), .A(
        n18834), .B(n18677), .ZN(n18689) );
  INV_X1 U21715 ( .A(n18689), .ZN(n18679) );
  AOI211_X1 U21716 ( .C1(n18681), .C2(n18680), .A(n18688), .B(n18679), .ZN(
        n18789) );
  AOI21_X1 U21717 ( .B1(n18708), .B2(n18682), .A(n18789), .ZN(n18691) );
  NAND3_X1 U21718 ( .A1(n18691), .A2(n18684), .A3(n18683), .ZN(n18686) );
  AOI22_X1 U21719 ( .A1(n18816), .A2(n18844), .B1(n18708), .B2(n18838), .ZN(
        n18685) );
  AOI22_X1 U21720 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18686), .B1(n18685), 
        .B2(n18788), .ZN(n18687) );
  OAI21_X1 U21721 ( .B1(n18689), .B2(n18688), .A(n18687), .ZN(P3_U2996) );
  NAND2_X1 U21722 ( .A1(n18708), .A2(n18838), .ZN(n18695) );
  NOR4_X1 U21723 ( .A1(n18788), .A2(n18801), .A3(n18842), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18698) );
  INV_X1 U21724 ( .A(n18698), .ZN(n18694) );
  NAND3_X1 U21725 ( .A1(n18692), .A2(n18691), .A3(n18690), .ZN(n18693) );
  NAND4_X1 U21726 ( .A1(n18696), .A2(n18695), .A3(n18694), .A4(n18693), .ZN(
        P3_U2997) );
  OAI21_X1 U21727 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18697), .ZN(n18699) );
  AOI21_X1 U21728 ( .B1(n18700), .B2(n18699), .A(n18698), .ZN(P3_U2998) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18701), .ZN(
        P3_U2999) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18701), .ZN(
        P3_U3000) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18701), .ZN(
        P3_U3001) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18701), .ZN(
        P3_U3002) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18701), .ZN(
        P3_U3003) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18701), .ZN(
        P3_U3004) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18701), .ZN(
        P3_U3005) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18701), .ZN(
        P3_U3006) );
  AND2_X1 U21737 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18701), .ZN(
        P3_U3007) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18701), .ZN(
        P3_U3008) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18701), .ZN(
        P3_U3009) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18701), .ZN(
        P3_U3010) );
  AND2_X1 U21741 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18701), .ZN(
        P3_U3011) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18701), .ZN(
        P3_U3012) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18701), .ZN(
        P3_U3013) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18701), .ZN(
        P3_U3014) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18701), .ZN(
        P3_U3015) );
  AND2_X1 U21746 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18701), .ZN(
        P3_U3016) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18701), .ZN(
        P3_U3017) );
  AND2_X1 U21748 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18701), .ZN(
        P3_U3018) );
  AND2_X1 U21749 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18701), .ZN(
        P3_U3019) );
  AND2_X1 U21750 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18701), .ZN(
        P3_U3020) );
  AND2_X1 U21751 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18701), .ZN(P3_U3021) );
  AND2_X1 U21752 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18701), .ZN(P3_U3022) );
  AND2_X1 U21753 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18701), .ZN(P3_U3023) );
  AND2_X1 U21754 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18701), .ZN(P3_U3024) );
  AND2_X1 U21755 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18701), .ZN(P3_U3025) );
  AND2_X1 U21756 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18701), .ZN(P3_U3026) );
  AND2_X1 U21757 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18701), .ZN(P3_U3027) );
  AND2_X1 U21758 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18701), .ZN(P3_U3028) );
  OAI21_X1 U21759 ( .B1(n18702), .B2(n20648), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18703) );
  AOI22_X1 U21760 ( .A1(n18716), .A2(n18718), .B1(n18849), .B2(n18703), .ZN(
        n18704) );
  NAND3_X1 U21761 ( .A1(NA), .A2(n18716), .A3(n20897), .ZN(n18711) );
  OAI211_X1 U21762 ( .C1(n18842), .C2(n18705), .A(n18704), .B(n18711), .ZN(
        P3_U3029) );
  INV_X1 U21763 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18706) );
  NOR2_X1 U21764 ( .A1(n18718), .A2(n20648), .ZN(n18714) );
  OAI22_X1 U21765 ( .A1(n18706), .A2(n18714), .B1(n20648), .B2(n18705), .ZN(
        n18707) );
  INV_X1 U21766 ( .A(n18707), .ZN(n18709) );
  NAND2_X1 U21767 ( .A1(n18708), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18712) );
  OAI211_X1 U21768 ( .C1(n18709), .C2(n18716), .A(n18712), .B(n18839), .ZN(
        P3_U3030) );
  INV_X1 U21769 ( .A(n18712), .ZN(n18710) );
  AOI21_X1 U21770 ( .B1(n18716), .B2(n18711), .A(n18710), .ZN(n18717) );
  OAI22_X1 U21771 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18712), .ZN(n18713) );
  OAI22_X1 U21772 ( .A1(n18714), .A2(n18713), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18715) );
  OAI22_X1 U21773 ( .A1(n18717), .A2(n18718), .B1(n18716), .B2(n18715), .ZN(
        P3_U3031) );
  OAI222_X1 U21774 ( .A1(n18823), .A2(n9650), .B1(n18719), .B2(n18777), .C1(
        n18720), .C2(n18775), .ZN(P3_U3032) );
  OAI222_X1 U21775 ( .A1(n18775), .A2(n18722), .B1(n18721), .B2(n18777), .C1(
        n18720), .C2(n9650), .ZN(P3_U3033) );
  OAI222_X1 U21776 ( .A1(n18775), .A2(n18725), .B1(n18723), .B2(n18777), .C1(
        n18722), .C2(n9650), .ZN(P3_U3034) );
  OAI222_X1 U21777 ( .A1(n18775), .A2(n18727), .B1(n20898), .B2(n18777), .C1(
        n18725), .C2(n9650), .ZN(P3_U3035) );
  OAI222_X1 U21778 ( .A1(n18727), .A2(n9650), .B1(n18726), .B2(n18777), .C1(
        n18728), .C2(n18775), .ZN(P3_U3036) );
  OAI222_X1 U21779 ( .A1(n18775), .A2(n18730), .B1(n18729), .B2(n18777), .C1(
        n18728), .C2(n9650), .ZN(P3_U3037) );
  OAI222_X1 U21780 ( .A1(n18775), .A2(n18733), .B1(n18731), .B2(n18777), .C1(
        n18730), .C2(n9650), .ZN(P3_U3038) );
  OAI222_X1 U21781 ( .A1(n18733), .A2(n9650), .B1(n18732), .B2(n18777), .C1(
        n18734), .C2(n18775), .ZN(P3_U3039) );
  OAI222_X1 U21782 ( .A1(n18775), .A2(n18736), .B1(n18735), .B2(n18777), .C1(
        n18734), .C2(n9650), .ZN(P3_U3040) );
  OAI222_X1 U21783 ( .A1(n18775), .A2(n18738), .B1(n18737), .B2(n18777), .C1(
        n18736), .C2(n9650), .ZN(P3_U3041) );
  OAI222_X1 U21784 ( .A1(n18775), .A2(n18740), .B1(n18739), .B2(n18777), .C1(
        n18738), .C2(n9650), .ZN(P3_U3042) );
  OAI222_X1 U21785 ( .A1(n18775), .A2(n18742), .B1(n18741), .B2(n18832), .C1(
        n18740), .C2(n9650), .ZN(P3_U3043) );
  OAI222_X1 U21786 ( .A1(n18775), .A2(n18745), .B1(n18743), .B2(n18832), .C1(
        n18742), .C2(n9650), .ZN(P3_U3044) );
  OAI222_X1 U21787 ( .A1(n18745), .A2(n9650), .B1(n18744), .B2(n18832), .C1(
        n18746), .C2(n18775), .ZN(P3_U3045) );
  INV_X1 U21788 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18748) );
  OAI222_X1 U21789 ( .A1(n18775), .A2(n18748), .B1(n18747), .B2(n18832), .C1(
        n18746), .C2(n9650), .ZN(P3_U3046) );
  OAI222_X1 U21790 ( .A1(n18775), .A2(n18751), .B1(n18749), .B2(n18832), .C1(
        n18748), .C2(n9650), .ZN(P3_U3047) );
  OAI222_X1 U21791 ( .A1(n18751), .A2(n9650), .B1(n18750), .B2(n18832), .C1(
        n18752), .C2(n18775), .ZN(P3_U3048) );
  INV_X1 U21792 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18754) );
  OAI222_X1 U21793 ( .A1(n18775), .A2(n18754), .B1(n18753), .B2(n18832), .C1(
        n18752), .C2(n9650), .ZN(P3_U3049) );
  OAI222_X1 U21794 ( .A1(n18775), .A2(n18757), .B1(n18755), .B2(n18832), .C1(
        n18754), .C2(n9650), .ZN(P3_U3050) );
  OAI222_X1 U21795 ( .A1(n18757), .A2(n9650), .B1(n18756), .B2(n18832), .C1(
        n18758), .C2(n18775), .ZN(P3_U3051) );
  OAI222_X1 U21796 ( .A1(n18775), .A2(n18759), .B1(n20900), .B2(n18832), .C1(
        n18758), .C2(n9650), .ZN(P3_U3052) );
  OAI222_X1 U21797 ( .A1(n18775), .A2(n18761), .B1(n18760), .B2(n18832), .C1(
        n18759), .C2(n9650), .ZN(P3_U3053) );
  OAI222_X1 U21798 ( .A1(n18775), .A2(n18763), .B1(n18762), .B2(n18832), .C1(
        n18761), .C2(n9650), .ZN(P3_U3054) );
  OAI222_X1 U21799 ( .A1(n18775), .A2(n18765), .B1(n18764), .B2(n18777), .C1(
        n18763), .C2(n9650), .ZN(P3_U3055) );
  OAI222_X1 U21800 ( .A1(n18775), .A2(n18767), .B1(n18766), .B2(n18777), .C1(
        n18765), .C2(n9650), .ZN(P3_U3056) );
  OAI222_X1 U21801 ( .A1(n18775), .A2(n18769), .B1(n18768), .B2(n18777), .C1(
        n18767), .C2(n9650), .ZN(P3_U3057) );
  OAI222_X1 U21802 ( .A1(n18775), .A2(n18772), .B1(n18770), .B2(n18777), .C1(
        n18769), .C2(n9650), .ZN(P3_U3058) );
  OAI222_X1 U21803 ( .A1(n18772), .A2(n9650), .B1(n18771), .B2(n18777), .C1(
        n18773), .C2(n18775), .ZN(P3_U3059) );
  OAI222_X1 U21804 ( .A1(n18775), .A2(n18779), .B1(n18774), .B2(n18777), .C1(
        n18773), .C2(n9650), .ZN(P3_U3060) );
  OAI222_X1 U21805 ( .A1(n9650), .A2(n18779), .B1(n18778), .B2(n18777), .C1(
        n18776), .C2(n18775), .ZN(P3_U3061) );
  INV_X1 U21806 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n20920) );
  AOI22_X1 U21807 ( .A1(n18832), .A2(n18780), .B1(n20920), .B2(n18849), .ZN(
        P3_U3274) );
  OAI22_X1 U21808 ( .A1(n18849), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18777), .ZN(n18781) );
  INV_X1 U21809 ( .A(n18781), .ZN(P3_U3275) );
  OAI22_X1 U21810 ( .A1(n18849), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18832), .ZN(n18782) );
  INV_X1 U21811 ( .A(n18782), .ZN(P3_U3276) );
  OAI22_X1 U21812 ( .A1(n18849), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18832), .ZN(n18783) );
  INV_X1 U21813 ( .A(n18783), .ZN(P3_U3277) );
  OAI21_X1 U21814 ( .B1(n18787), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18785), 
        .ZN(n18784) );
  INV_X1 U21815 ( .A(n18784), .ZN(P3_U3280) );
  OAI21_X1 U21816 ( .B1(n18787), .B2(n18786), .A(n18785), .ZN(P3_U3281) );
  NOR2_X1 U21817 ( .A1(n18789), .A2(n18788), .ZN(n18792) );
  OAI21_X1 U21818 ( .B1(n18792), .B2(n18791), .A(n18790), .ZN(P3_U3282) );
  INV_X1 U21819 ( .A(n18793), .ZN(n18796) );
  NOR2_X1 U21820 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18851), .ZN(
        n18795) );
  AOI22_X1 U21821 ( .A1(n18816), .A2(n18796), .B1(n18795), .B2(n18794), .ZN(
        n18800) );
  INV_X1 U21822 ( .A(n18851), .ZN(n18818) );
  AOI21_X1 U21823 ( .B1(n18818), .B2(n18797), .A(n18822), .ZN(n18799) );
  OAI22_X1 U21824 ( .A1(n18822), .A2(n18800), .B1(n18799), .B2(n18798), .ZN(
        P3_U3285) );
  NOR2_X1 U21825 ( .A1(n18801), .A2(n18819), .ZN(n18810) );
  OAI22_X1 U21826 ( .A1(n18803), .A2(n18802), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18811) );
  INV_X1 U21827 ( .A(n18811), .ZN(n18805) );
  AOI222_X1 U21828 ( .A1(n18806), .A2(n18818), .B1(n18810), .B2(n18805), .C1(
        n18816), .C2(n18804), .ZN(n18807) );
  AOI22_X1 U21829 ( .A1(n18822), .A2(n18808), .B1(n18807), .B2(n18820), .ZN(
        P3_U3288) );
  INV_X1 U21830 ( .A(n18809), .ZN(n18813) );
  AOI222_X1 U21831 ( .A1(n18813), .A2(n18818), .B1(n18816), .B2(n18812), .C1(
        n18811), .C2(n18810), .ZN(n18814) );
  AOI22_X1 U21832 ( .A1(n18822), .A2(n18815), .B1(n18814), .B2(n18820), .ZN(
        P3_U3289) );
  AOI222_X1 U21833 ( .A1(n18819), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18818), 
        .B2(n18817), .C1(n20913), .C2(n18816), .ZN(n18821) );
  AOI22_X1 U21834 ( .A1(n18822), .A2(n20913), .B1(n18821), .B2(n18820), .ZN(
        P3_U3290) );
  AOI21_X1 U21835 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18824) );
  AOI22_X1 U21836 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18824), .B2(n18823), .ZN(n18827) );
  INV_X1 U21837 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18826) );
  AOI22_X1 U21838 ( .A1(n18830), .A2(n18827), .B1(n18826), .B2(n18825), .ZN(
        P3_U3292) );
  INV_X1 U21839 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18829) );
  OAI21_X1 U21840 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18830), .ZN(n18828) );
  OAI21_X1 U21841 ( .B1(n18830), .B2(n18829), .A(n18828), .ZN(P3_U3293) );
  INV_X1 U21842 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18831) );
  AOI22_X1 U21843 ( .A1(n18832), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18831), 
        .B2(n18849), .ZN(P3_U3294) );
  MUX2_X1 U21844 ( .A(P3_MORE_REG_SCAN_IN), .B(n18834), .S(n18833), .Z(
        P3_U3295) );
  OAI21_X1 U21845 ( .B1(n18836), .B2(n18835), .A(n18853), .ZN(n18837) );
  AOI21_X1 U21846 ( .B1(n18838), .B2(n18842), .A(n18837), .ZN(n18848) );
  AOI21_X1 U21847 ( .B1(n18841), .B2(n18840), .A(n18839), .ZN(n18843) );
  OAI211_X1 U21848 ( .C1(n18852), .C2(n18843), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18842), .ZN(n18845) );
  AOI21_X1 U21849 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18845), .A(n18844), 
        .ZN(n18847) );
  NAND2_X1 U21850 ( .A1(n18848), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18846) );
  OAI21_X1 U21851 ( .B1(n18848), .B2(n18847), .A(n18846), .ZN(P3_U3296) );
  OAI22_X1 U21852 ( .A1(n18849), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18777), .ZN(n18850) );
  INV_X1 U21853 ( .A(n18850), .ZN(P3_U3297) );
  OAI21_X1 U21854 ( .B1(n18851), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18853), 
        .ZN(n18856) );
  OAI22_X1 U21855 ( .A1(n18856), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18853), 
        .B2(n18852), .ZN(n18854) );
  INV_X1 U21856 ( .A(n18854), .ZN(P3_U3298) );
  OAI21_X1 U21857 ( .B1(n18856), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18855), 
        .ZN(n18857) );
  INV_X1 U21858 ( .A(n18857), .ZN(P3_U3299) );
  INV_X1 U21859 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19784) );
  NAND2_X1 U21860 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19784), .ZN(n19772) );
  AOI22_X1 U21861 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19772), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19765), .ZN(n19845) );
  AOI21_X1 U21862 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19845), .ZN(n18858) );
  INV_X1 U21863 ( .A(n18858), .ZN(P2_U2815) );
  INV_X1 U21864 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18861) );
  INV_X1 U21865 ( .A(n18859), .ZN(n18860) );
  OAI22_X1 U21866 ( .A1(n18862), .A2(n18861), .B1(n12960), .B2(n18860), .ZN(
        P2_U2816) );
  NAND2_X1 U21867 ( .A1(n19765), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19910) );
  INV_X2 U21868 ( .A(n19910), .ZN(n19835) );
  OR2_X1 U21869 ( .A1(n19775), .A2(n19835), .ZN(n19768) );
  AOI21_X1 U21870 ( .B1(n19765), .B2(n19768), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18863) );
  AOI21_X1 U21871 ( .B1(n19835), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n18863), 
        .ZN(P2_U2817) );
  OAI21_X1 U21872 ( .B1(n19775), .B2(BS16), .A(n19845), .ZN(n19843) );
  OAI21_X1 U21873 ( .B1(n19845), .B2(n19470), .A(n19843), .ZN(P2_U2818) );
  NOR4_X1 U21874 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18867) );
  NOR4_X1 U21875 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18866) );
  NOR4_X1 U21876 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18865) );
  NOR4_X1 U21877 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18864) );
  NAND4_X1 U21878 ( .A1(n18867), .A2(n18866), .A3(n18865), .A4(n18864), .ZN(
        n18873) );
  NOR4_X1 U21879 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18871) );
  AOI211_X1 U21880 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_19__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18870) );
  NOR4_X1 U21881 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18869) );
  NOR4_X1 U21882 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18868) );
  NAND4_X1 U21883 ( .A1(n18871), .A2(n18870), .A3(n18869), .A4(n18868), .ZN(
        n18872) );
  NOR2_X1 U21884 ( .A1(n18873), .A2(n18872), .ZN(n18884) );
  INV_X1 U21885 ( .A(n18884), .ZN(n18882) );
  NOR2_X1 U21886 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18882), .ZN(n18876) );
  INV_X1 U21887 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18874) );
  AOI22_X1 U21888 ( .A1(n18876), .A2(n18877), .B1(n18882), .B2(n18874), .ZN(
        P2_U2820) );
  OR3_X1 U21889 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18881) );
  INV_X1 U21890 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18875) );
  AOI22_X1 U21891 ( .A1(n18876), .A2(n18881), .B1(n18882), .B2(n18875), .ZN(
        P2_U2821) );
  INV_X1 U21892 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19844) );
  NAND2_X1 U21893 ( .A1(n18876), .A2(n19844), .ZN(n18880) );
  OAI21_X1 U21894 ( .B1(n18877), .B2(n10419), .A(n18884), .ZN(n18878) );
  OAI21_X1 U21895 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18884), .A(n18878), 
        .ZN(n18879) );
  OAI221_X1 U21896 ( .B1(n18880), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18880), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18879), .ZN(P2_U2822) );
  INV_X1 U21897 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18883) );
  OAI221_X1 U21898 ( .B1(n18884), .B2(n18883), .C1(n18882), .C2(n18881), .A(
        n18880), .ZN(P2_U2823) );
  AOI22_X1 U21899 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19038), .ZN(n18896) );
  AOI22_X1 U21900 ( .A1(n18885), .A2(n19062), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19055), .ZN(n18895) );
  INV_X1 U21901 ( .A(n18886), .ZN(n18887) );
  AOI22_X1 U21902 ( .A1(n18888), .A2(n19067), .B1(n18887), .B2(n18972), .ZN(
        n18894) );
  AOI21_X1 U21903 ( .B1(n18891), .B2(n18890), .A(n18889), .ZN(n18892) );
  NAND2_X1 U21904 ( .A1(n12968), .A2(n18892), .ZN(n18893) );
  NAND4_X1 U21905 ( .A1(n18896), .A2(n18895), .A3(n18894), .A4(n18893), .ZN(
        P2_U2835) );
  INV_X1 U21906 ( .A(n18897), .ZN(n18899) );
  OAI22_X1 U21907 ( .A1(n18899), .A2(n19024), .B1(n19042), .B2(n18898), .ZN(
        n18900) );
  AOI211_X1 U21908 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19045), .A(n19044), 
        .B(n18900), .ZN(n18901) );
  OAI21_X1 U21909 ( .B1(n18902), .B2(n19057), .A(n18901), .ZN(n18903) );
  INV_X1 U21910 ( .A(n18903), .ZN(n18910) );
  NAND2_X1 U21911 ( .A1(n18905), .A2(n18904), .ZN(n18908) );
  NOR2_X1 U21912 ( .A1(n19759), .A2(n18906), .ZN(n18907) );
  NAND2_X1 U21913 ( .A1(n18908), .A2(n18907), .ZN(n18909) );
  OAI211_X1 U21914 ( .C1(n18958), .C2(n18911), .A(n18910), .B(n18909), .ZN(
        n18912) );
  INV_X1 U21915 ( .A(n18912), .ZN(n18913) );
  OAI21_X1 U21916 ( .B1(n18914), .B2(n19065), .A(n18913), .ZN(P2_U2836) );
  XNOR2_X1 U21917 ( .A(n18916), .B(n18915), .ZN(n18926) );
  INV_X1 U21918 ( .A(n18917), .ZN(n18919) );
  AOI22_X1 U21919 ( .A1(n19055), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19038), .ZN(n18918) );
  OAI21_X1 U21920 ( .B1(n18919), .B2(n19024), .A(n18918), .ZN(n18920) );
  AOI211_X1 U21921 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19045), .A(n19044), 
        .B(n18920), .ZN(n18925) );
  OAI22_X1 U21922 ( .A1(n18922), .A2(n18958), .B1(n18921), .B2(n19065), .ZN(
        n18923) );
  INV_X1 U21923 ( .A(n18923), .ZN(n18924) );
  OAI211_X1 U21924 ( .C1(n19759), .C2(n18926), .A(n18925), .B(n18924), .ZN(
        P2_U2837) );
  AOI22_X1 U21925 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19055), .ZN(n18937) );
  INV_X1 U21926 ( .A(n18956), .ZN(n19075) );
  OAI22_X1 U21927 ( .A1(n18927), .A2(n19024), .B1(n19075), .B2(n18932), .ZN(
        n18928) );
  AOI211_X1 U21928 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19045), .A(n19044), 
        .B(n18928), .ZN(n18936) );
  AOI22_X1 U21929 ( .A1(n18930), .A2(n19067), .B1(n18972), .B2(n18929), .ZN(
        n18935) );
  OAI211_X1 U21930 ( .C1(n18933), .C2(n18932), .A(n18942), .B(n18931), .ZN(
        n18934) );
  NAND4_X1 U21931 ( .A1(n18937), .A2(n18936), .A3(n18935), .A4(n18934), .ZN(
        P2_U2838) );
  NOR2_X1 U21932 ( .A1(n19059), .A2(n15090), .ZN(n18938) );
  AOI211_X1 U21933 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19038), .A(
        n19044), .B(n18938), .ZN(n18939) );
  OAI21_X1 U21934 ( .B1(n19042), .B2(n18940), .A(n18939), .ZN(n18946) );
  OAI211_X1 U21935 ( .C1(n18943), .C2(n18952), .A(n18942), .B(n18941), .ZN(
        n18944) );
  INV_X1 U21936 ( .A(n18944), .ZN(n18945) );
  AOI211_X1 U21937 ( .C1(n19062), .C2(n18947), .A(n18946), .B(n18945), .ZN(
        n18951) );
  INV_X1 U21938 ( .A(n19089), .ZN(n18948) );
  AOI22_X1 U21939 ( .A1(n18949), .A2(n19067), .B1(n18972), .B2(n18948), .ZN(
        n18950) );
  OAI211_X1 U21940 ( .C1(n18952), .C2(n19075), .A(n18951), .B(n18950), .ZN(
        P2_U2840) );
  AOI22_X1 U21941 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19055), .ZN(n18953) );
  OAI211_X1 U21942 ( .C1(n19059), .C2(n11342), .A(n18953), .B(n19023), .ZN(
        n18954) );
  AOI21_X1 U21943 ( .B1(n18956), .B2(n18955), .A(n18954), .ZN(n18957) );
  OAI21_X1 U21944 ( .B1(n19082), .B2(n18958), .A(n18957), .ZN(n18959) );
  AOI21_X1 U21945 ( .B1(n18960), .B2(n19062), .A(n18959), .ZN(n18966) );
  INV_X1 U21946 ( .A(n18961), .ZN(n18962) );
  OAI211_X1 U21947 ( .C1(n18964), .C2(n18963), .A(n12968), .B(n18962), .ZN(
        n18965) );
  OAI211_X1 U21948 ( .C1(n19065), .C2(n19094), .A(n18966), .B(n18965), .ZN(
        P2_U2842) );
  NAND2_X1 U21949 ( .A1(n19029), .A2(n18967), .ZN(n18986) );
  XOR2_X1 U21950 ( .A(n18968), .B(n18986), .Z(n18976) );
  AOI22_X1 U21951 ( .A1(n19055), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19038), .ZN(n18969) );
  OAI21_X1 U21952 ( .B1(n18970), .B2(n19024), .A(n18969), .ZN(n18971) );
  AOI211_X1 U21953 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19045), .A(n19044), 
        .B(n18971), .ZN(n18975) );
  AOI22_X1 U21954 ( .A1(n18973), .A2(n19067), .B1(n18972), .B2(n19095), .ZN(
        n18974) );
  OAI211_X1 U21955 ( .C1(n19759), .C2(n18976), .A(n18975), .B(n18974), .ZN(
        P2_U2843) );
  AOI22_X1 U21956 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19055), .ZN(n18977) );
  OAI211_X1 U21957 ( .C1(n19065), .C2(n19101), .A(n18977), .B(n19023), .ZN(
        n18978) );
  INV_X1 U21958 ( .A(n18978), .ZN(n18979) );
  OAI21_X1 U21959 ( .B1(n11310), .B2(n19059), .A(n18979), .ZN(n18984) );
  INV_X1 U21960 ( .A(n18980), .ZN(n18981) );
  NOR3_X1 U21961 ( .A1(n18982), .A2(n18981), .A3(n19024), .ZN(n18983) );
  AOI211_X1 U21962 ( .C1(n18985), .C2(n19067), .A(n18984), .B(n18983), .ZN(
        n18990) );
  INV_X1 U21963 ( .A(n18986), .ZN(n18987) );
  OAI211_X1 U21964 ( .C1(n18988), .C2(n18991), .A(n12968), .B(n18987), .ZN(
        n18989) );
  OAI211_X1 U21965 ( .C1(n19075), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P2_U2844) );
  OAI21_X1 U21966 ( .B1(n19799), .B2(n19059), .A(n19023), .ZN(n18994) );
  OAI22_X1 U21967 ( .A1(n18992), .A2(n19024), .B1(n19042), .B2(n10040), .ZN(
        n18993) );
  AOI211_X1 U21968 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19038), .A(
        n18994), .B(n18993), .ZN(n19001) );
  NAND2_X1 U21969 ( .A1(n19029), .A2(n18995), .ZN(n18996) );
  XOR2_X1 U21970 ( .A(n18997), .B(n18996), .Z(n18999) );
  AOI22_X1 U21971 ( .A1(n18999), .A2(n12968), .B1(n19067), .B2(n18998), .ZN(
        n19000) );
  OAI211_X1 U21972 ( .C1(n19103), .C2(n19065), .A(n19001), .B(n19000), .ZN(
        P2_U2845) );
  AOI22_X1 U21973 ( .A1(n19002), .A2(n19062), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19055), .ZN(n19003) );
  OAI21_X1 U21974 ( .B1(n19004), .B2(n19057), .A(n19003), .ZN(n19005) );
  AOI211_X1 U21975 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19045), .A(n19044), .B(
        n19005), .ZN(n19012) );
  NOR2_X1 U21976 ( .A1(n19047), .A2(n19006), .ZN(n19008) );
  XNOR2_X1 U21977 ( .A(n19008), .B(n19007), .ZN(n19010) );
  AOI22_X1 U21978 ( .A1(n19010), .A2(n12968), .B1(n19067), .B2(n19009), .ZN(
        n19011) );
  OAI211_X1 U21979 ( .C1(n19065), .C2(n19105), .A(n19012), .B(n19011), .ZN(
        P2_U2846) );
  AOI22_X1 U21980 ( .A1(n19013), .A2(n19062), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19055), .ZN(n19014) );
  OAI211_X1 U21981 ( .C1(n19794), .C2(n19059), .A(n19014), .B(n19023), .ZN(
        n19015) );
  AOI21_X1 U21982 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19038), .A(
        n19015), .ZN(n19022) );
  NOR2_X1 U21983 ( .A1(n19047), .A2(n19016), .ZN(n19018) );
  XNOR2_X1 U21984 ( .A(n19018), .B(n19017), .ZN(n19020) );
  AOI22_X1 U21985 ( .A1(n19020), .A2(n12968), .B1(n19067), .B2(n19019), .ZN(
        n19021) );
  OAI211_X1 U21986 ( .C1(n19065), .C2(n19109), .A(n19022), .B(n19021), .ZN(
        P2_U2848) );
  OAI21_X1 U21987 ( .B1(n19792), .B2(n19059), .A(n19023), .ZN(n19027) );
  OAI22_X1 U21988 ( .A1(n19042), .A2(n13370), .B1(n19025), .B2(n19024), .ZN(
        n19026) );
  AOI211_X1 U21989 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19038), .A(
        n19027), .B(n19026), .ZN(n19036) );
  NAND2_X1 U21990 ( .A1(n19029), .A2(n19028), .ZN(n19030) );
  XNOR2_X1 U21991 ( .A(n19031), .B(n19030), .ZN(n19034) );
  INV_X1 U21992 ( .A(n19032), .ZN(n19033) );
  AOI22_X1 U21993 ( .A1(n19034), .A2(n12968), .B1(n19067), .B2(n19033), .ZN(
        n19035) );
  OAI211_X1 U21994 ( .C1(n19065), .C2(n19110), .A(n19036), .B(n19035), .ZN(
        P2_U2849) );
  INV_X1 U21995 ( .A(n19037), .ZN(n19039) );
  AOI22_X1 U21996 ( .A1(n19039), .A2(n19062), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19038), .ZN(n19040) );
  OAI21_X1 U21997 ( .B1(n19042), .B2(n19041), .A(n19040), .ZN(n19043) );
  AOI211_X1 U21998 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19045), .A(n19044), .B(
        n19043), .ZN(n19053) );
  NOR2_X1 U21999 ( .A1(n19047), .A2(n19046), .ZN(n19049) );
  XNOR2_X1 U22000 ( .A(n19049), .B(n19048), .ZN(n19051) );
  AOI22_X1 U22001 ( .A1(n19051), .A2(n12968), .B1(n19067), .B2(n19050), .ZN(
        n19052) );
  OAI211_X1 U22002 ( .C1(n19065), .C2(n19122), .A(n19053), .B(n19052), .ZN(
        P2_U2850) );
  NAND2_X1 U22003 ( .A1(n19055), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19064) );
  INV_X1 U22004 ( .A(n19056), .ZN(n19061) );
  OAI22_X1 U22005 ( .A1(n10419), .A2(n19059), .B1(n19058), .B2(n19057), .ZN(
        n19060) );
  AOI21_X1 U22006 ( .B1(n19062), .B2(n19061), .A(n19060), .ZN(n19063) );
  OAI211_X1 U22007 ( .C1(n19879), .C2(n19065), .A(n19064), .B(n19063), .ZN(
        n19066) );
  AOI21_X1 U22008 ( .B1(n19068), .B2(n19067), .A(n19066), .ZN(n19071) );
  NAND2_X1 U22009 ( .A1(n19883), .A2(n19069), .ZN(n19070) );
  OAI211_X1 U22010 ( .C1(n19072), .C2(n19759), .A(n19071), .B(n19070), .ZN(
        n19073) );
  INV_X1 U22011 ( .A(n19073), .ZN(n19074) );
  OAI21_X1 U22012 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19075), .A(
        n19074), .ZN(P2_U2854) );
  XOR2_X1 U22013 ( .A(n19077), .B(n19076), .Z(n19080) );
  AOI22_X1 U22014 ( .A1(n19080), .A2(n19079), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n19078), .ZN(n19081) );
  OAI21_X1 U22015 ( .B1(n19082), .B2(n19078), .A(n19081), .ZN(P2_U2874) );
  AOI22_X1 U22016 ( .A1(n19084), .A2(BUF2_REG_31__SCAN_IN), .B1(n19138), .B2(
        n19083), .ZN(n19087) );
  AOI22_X1 U22017 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19137), .B1(n19085), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19086) );
  NAND2_X1 U22018 ( .A1(n19087), .A2(n19086), .ZN(P2_U2888) );
  OAI222_X1 U22019 ( .A1(n19089), .A2(n19123), .B1(n13055), .B2(n19111), .C1(
        n19088), .C2(n19145), .ZN(P2_U2904) );
  AOI22_X1 U22020 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19137), .B1(n19090), 
        .B2(n19096), .ZN(n19091) );
  OAI21_X1 U22021 ( .B1(n19123), .B2(n19092), .A(n19091), .ZN(P2_U2905) );
  INV_X1 U22022 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19189) );
  OAI222_X1 U22023 ( .A1(n19094), .A2(n19123), .B1(n19189), .B2(n19111), .C1(
        n19145), .C2(n19093), .ZN(P2_U2906) );
  INV_X1 U22024 ( .A(n19095), .ZN(n19099) );
  AOI22_X1 U22025 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19137), .B1(n19097), 
        .B2(n19096), .ZN(n19098) );
  OAI21_X1 U22026 ( .B1(n19123), .B2(n19099), .A(n19098), .ZN(P2_U2907) );
  INV_X1 U22027 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19193) );
  OAI222_X1 U22028 ( .A1(n19101), .A2(n19123), .B1(n19193), .B2(n19111), .C1(
        n19145), .C2(n19100), .ZN(P2_U2908) );
  INV_X1 U22029 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19195) );
  OAI222_X1 U22030 ( .A1(n19103), .A2(n19123), .B1(n19195), .B2(n19111), .C1(
        n19145), .C2(n19102), .ZN(P2_U2909) );
  INV_X1 U22031 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19197) );
  OAI222_X1 U22032 ( .A1(n19105), .A2(n19123), .B1(n19197), .B2(n19111), .C1(
        n19145), .C2(n19104), .ZN(P2_U2910) );
  INV_X1 U22033 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19199) );
  OAI222_X1 U22034 ( .A1(n19107), .A2(n19123), .B1(n19199), .B2(n19111), .C1(
        n19145), .C2(n19106), .ZN(P2_U2911) );
  INV_X1 U22035 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19203) );
  OAI222_X1 U22036 ( .A1(n19109), .A2(n19123), .B1(n19203), .B2(n19111), .C1(
        n19145), .C2(n19108), .ZN(P2_U2912) );
  INV_X1 U22037 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19205) );
  OAI222_X1 U22038 ( .A1(n19110), .A2(n19123), .B1(n19205), .B2(n19111), .C1(
        n19145), .C2(n19260), .ZN(P2_U2913) );
  INV_X1 U22039 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20871) );
  OAI22_X1 U22040 ( .A1(n20871), .A2(n19111), .B1(n19250), .B2(n19145), .ZN(
        n19112) );
  INV_X1 U22041 ( .A(n19112), .ZN(n19121) );
  XNOR2_X1 U22042 ( .A(n19113), .B(n19865), .ZN(n19132) );
  NAND2_X1 U22043 ( .A1(n19872), .A2(n19114), .ZN(n19116) );
  NAND2_X1 U22044 ( .A1(n19116), .A2(n19115), .ZN(n19131) );
  NAND2_X1 U22045 ( .A1(n19132), .A2(n19131), .ZN(n19130) );
  OAI21_X1 U22046 ( .B1(n19866), .B2(n19865), .A(n19130), .ZN(n19118) );
  NAND2_X1 U22047 ( .A1(n19118), .A2(n19117), .ZN(n19126) );
  INV_X1 U22048 ( .A(n19125), .ZN(n19119) );
  NAND3_X1 U22049 ( .A1(n19126), .A2(n19119), .A3(n19139), .ZN(n19120) );
  OAI211_X1 U22050 ( .C1(n19123), .C2(n19122), .A(n19121), .B(n19120), .ZN(
        P2_U2914) );
  AOI22_X1 U22051 ( .A1(n19138), .A2(n19124), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19137), .ZN(n19129) );
  XNOR2_X1 U22052 ( .A(n19126), .B(n19125), .ZN(n19127) );
  NAND2_X1 U22053 ( .A1(n19127), .A2(n19139), .ZN(n19128) );
  OAI211_X1 U22054 ( .C1(n19246), .C2(n19145), .A(n19129), .B(n19128), .ZN(
        P2_U2915) );
  OAI21_X1 U22055 ( .B1(n19132), .B2(n19131), .A(n19130), .ZN(n19133) );
  NAND2_X1 U22056 ( .A1(n19133), .A2(n19139), .ZN(n19135) );
  AOI22_X1 U22057 ( .A1(n19865), .A2(n19138), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19137), .ZN(n19134) );
  OAI211_X1 U22058 ( .C1(n19136), .C2(n19145), .A(n19135), .B(n19134), .ZN(
        P2_U2916) );
  AOI22_X1 U22059 ( .A1(n19138), .A2(n19141), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19137), .ZN(n19144) );
  OAI211_X1 U22060 ( .C1(n19142), .C2(n19141), .A(n19140), .B(n19139), .ZN(
        n19143) );
  OAI211_X1 U22061 ( .C1(n19146), .C2(n19145), .A(n19144), .B(n19143), .ZN(
        P2_U2919) );
  OAI21_X1 U22062 ( .B1(n19149), .B2(n19148), .A(n19147), .ZN(n19151) );
  NOR2_X4 U22063 ( .A1(n19184), .A2(n19201), .ZN(n19200) );
  AND2_X1 U22064 ( .A1(n19200), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22065 ( .A1(n19201), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19153) );
  OAI21_X1 U22066 ( .B1(n19154), .B2(n19182), .A(n19153), .ZN(P2_U2921) );
  AOI22_X1 U22067 ( .A1(n19201), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19155) );
  OAI21_X1 U22068 ( .B1(n19156), .B2(n19182), .A(n19155), .ZN(P2_U2922) );
  AOI22_X1 U22069 ( .A1(n19201), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19157) );
  OAI21_X1 U22070 ( .B1(n19158), .B2(n19182), .A(n19157), .ZN(P2_U2923) );
  AOI22_X1 U22071 ( .A1(n19201), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19159) );
  OAI21_X1 U22072 ( .B1(n19160), .B2(n19182), .A(n19159), .ZN(P2_U2924) );
  AOI22_X1 U22073 ( .A1(n19201), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19161) );
  OAI21_X1 U22074 ( .B1(n19162), .B2(n19182), .A(n19161), .ZN(P2_U2925) );
  INV_X1 U22075 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U22076 ( .A1(n19201), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19163) );
  OAI21_X1 U22077 ( .B1(n19164), .B2(n19182), .A(n19163), .ZN(P2_U2926) );
  AOI22_X1 U22078 ( .A1(n19201), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19165) );
  OAI21_X1 U22079 ( .B1(n19166), .B2(n19182), .A(n19165), .ZN(P2_U2927) );
  INV_X1 U22080 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19168) );
  AOI22_X1 U22081 ( .A1(n19201), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19167) );
  OAI21_X1 U22082 ( .B1(n19168), .B2(n19182), .A(n19167), .ZN(P2_U2928) );
  INV_X1 U22083 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19170) );
  AOI22_X1 U22084 ( .A1(n19201), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19169) );
  OAI21_X1 U22085 ( .B1(n19170), .B2(n19182), .A(n19169), .ZN(P2_U2929) );
  AOI22_X1 U22086 ( .A1(n19201), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19171) );
  OAI21_X1 U22087 ( .B1(n19172), .B2(n19182), .A(n19171), .ZN(P2_U2930) );
  INV_X1 U22088 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19174) );
  AOI22_X1 U22089 ( .A1(n19201), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19173) );
  OAI21_X1 U22090 ( .B1(n19174), .B2(n19182), .A(n19173), .ZN(P2_U2931) );
  INV_X1 U22091 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19176) );
  AOI22_X1 U22092 ( .A1(n19215), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19175) );
  OAI21_X1 U22093 ( .B1(n19176), .B2(n19182), .A(n19175), .ZN(P2_U2932) );
  INV_X1 U22094 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19178) );
  AOI22_X1 U22095 ( .A1(n19215), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19177) );
  OAI21_X1 U22096 ( .B1(n19178), .B2(n19182), .A(n19177), .ZN(P2_U2933) );
  INV_X1 U22097 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19180) );
  AOI22_X1 U22098 ( .A1(n19215), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U22099 ( .B1(n19180), .B2(n19182), .A(n19179), .ZN(P2_U2934) );
  INV_X1 U22100 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19183) );
  AOI22_X1 U22101 ( .A1(n19201), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22102 ( .B1(n19183), .B2(n19182), .A(n19181), .ZN(P2_U2935) );
  AOI22_X1 U22103 ( .A1(n19201), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U22104 ( .B1(n13055), .B2(n19217), .A(n19185), .ZN(P2_U2936) );
  AOI22_X1 U22105 ( .A1(n19201), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U22106 ( .B1(n19187), .B2(n19217), .A(n19186), .ZN(P2_U2937) );
  AOI22_X1 U22107 ( .A1(n19201), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U22108 ( .B1(n19189), .B2(n19217), .A(n19188), .ZN(P2_U2938) );
  AOI22_X1 U22109 ( .A1(n19201), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U22110 ( .B1(n19191), .B2(n19217), .A(n19190), .ZN(P2_U2939) );
  AOI22_X1 U22111 ( .A1(n19201), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U22112 ( .B1(n19193), .B2(n19217), .A(n19192), .ZN(P2_U2940) );
  AOI22_X1 U22113 ( .A1(n19201), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22114 ( .B1(n19195), .B2(n19217), .A(n19194), .ZN(P2_U2941) );
  AOI22_X1 U22115 ( .A1(n19201), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22116 ( .B1(n19197), .B2(n19217), .A(n19196), .ZN(P2_U2942) );
  AOI22_X1 U22117 ( .A1(n19201), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22118 ( .B1(n19199), .B2(n19217), .A(n19198), .ZN(P2_U2943) );
  AOI22_X1 U22119 ( .A1(n19201), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22120 ( .B1(n19203), .B2(n19217), .A(n19202), .ZN(P2_U2944) );
  AOI22_X1 U22121 ( .A1(n19215), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22122 ( .B1(n19205), .B2(n19217), .A(n19204), .ZN(P2_U2945) );
  AOI22_X1 U22123 ( .A1(n19215), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19206) );
  OAI21_X1 U22124 ( .B1(n20871), .B2(n19217), .A(n19206), .ZN(P2_U2946) );
  INV_X1 U22125 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19208) );
  AOI22_X1 U22126 ( .A1(n19215), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22127 ( .B1(n19208), .B2(n19217), .A(n19207), .ZN(P2_U2947) );
  INV_X1 U22128 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19210) );
  AOI22_X1 U22129 ( .A1(n19215), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22130 ( .B1(n19210), .B2(n19217), .A(n19209), .ZN(P2_U2948) );
  INV_X1 U22131 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19212) );
  AOI22_X1 U22132 ( .A1(n19215), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22133 ( .B1(n19212), .B2(n19217), .A(n19211), .ZN(P2_U2949) );
  AOI22_X1 U22134 ( .A1(n19215), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22135 ( .B1(n19214), .B2(n19217), .A(n19213), .ZN(P2_U2950) );
  INV_X1 U22136 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19218) );
  AOI22_X1 U22137 ( .A1(n19215), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19200), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19216) );
  OAI21_X1 U22138 ( .B1(n19218), .B2(n19217), .A(n19216), .ZN(P2_U2951) );
  AOI22_X1 U22139 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19044), .B1(n19220), 
        .B2(n19219), .ZN(n19227) );
  AOI222_X1 U22140 ( .A1(n19225), .A2(n19224), .B1(n19239), .B2(n19223), .C1(
        n19222), .C2(n19221), .ZN(n19226) );
  OAI211_X1 U22141 ( .C1(n19229), .C2(n19228), .A(n19227), .B(n19226), .ZN(
        P2_U3010) );
  OAI21_X1 U22142 ( .B1(n19231), .B2(n19230), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19241) );
  OAI21_X1 U22143 ( .B1(n19234), .B2(n19233), .A(n19232), .ZN(n19238) );
  NOR2_X1 U22144 ( .A1(n19236), .A2(n19235), .ZN(n19237) );
  AOI211_X1 U22145 ( .C1(n19239), .C2(n10461), .A(n19238), .B(n19237), .ZN(
        n19240) );
  NAND2_X1 U22146 ( .A1(n19241), .A2(n19240), .ZN(P2_U3014) );
  AOI22_X1 U22147 ( .A1(n19649), .A2(n19749), .B1(n19695), .B2(n19259), .ZN(
        n19244) );
  INV_X1 U22148 ( .A(n19663), .ZN(n19704) );
  AOI22_X1 U22149 ( .A1(n19696), .A2(n19263), .B1(n19292), .B2(n19704), .ZN(
        n19243) );
  OAI211_X1 U22150 ( .C1(n19266), .C2(n12737), .A(n19244), .B(n19243), .ZN(
        P2_U3048) );
  AOI22_X1 U22151 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19261), .ZN(n19731) );
  INV_X1 U22152 ( .A(n19731), .ZN(n19602) );
  AOI22_X1 U22153 ( .A1(n19602), .A2(n19749), .B1(n19259), .B2(n19726), .ZN(
        n19248) );
  NOR2_X2 U22154 ( .A1(n19246), .A2(n19447), .ZN(n19727) );
  AOI22_X1 U22155 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19261), .ZN(n19605) );
  AOI22_X1 U22156 ( .A1(n19727), .A2(n19263), .B1(n19292), .B2(n19728), .ZN(
        n19247) );
  OAI211_X1 U22157 ( .C1(n19266), .C2(n19249), .A(n19248), .B(n19247), .ZN(
        P2_U3052) );
  AOI22_X1 U22158 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19261), .ZN(n19737) );
  AOI22_X1 U22159 ( .A1(n19606), .A2(n19749), .B1(n19259), .B2(n19732), .ZN(
        n19256) );
  NOR2_X2 U22160 ( .A1(n19250), .A2(n19447), .ZN(n19733) );
  AOI22_X1 U22161 ( .A1(n19733), .A2(n19263), .B1(n19292), .B2(n19734), .ZN(
        n19255) );
  OAI211_X1 U22162 ( .C1(n19266), .C2(n19257), .A(n19256), .B(n19255), .ZN(
        P2_U3053) );
  AOI22_X1 U22163 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19261), .ZN(n19743) );
  AOI22_X1 U22164 ( .A1(n19639), .A2(n19749), .B1(n19259), .B2(n19738), .ZN(
        n19265) );
  NOR2_X2 U22165 ( .A1(n19260), .A2(n19447), .ZN(n19739) );
  AOI22_X1 U22166 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19262), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19261), .ZN(n19642) );
  INV_X1 U22167 ( .A(n19642), .ZN(n19740) );
  AOI22_X1 U22168 ( .A1(n19739), .A2(n19263), .B1(n19292), .B2(n19740), .ZN(
        n19264) );
  OAI211_X1 U22169 ( .C1(n19266), .C2(n13474), .A(n19265), .B(n19264), .ZN(
        P2_U3054) );
  INV_X1 U22170 ( .A(n10711), .ZN(n19267) );
  NAND2_X1 U22171 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19886), .ZN(
        n19501) );
  NOR2_X1 U22172 ( .A1(n19501), .A2(n19328), .ZN(n19290) );
  OAI21_X1 U22173 ( .B1(n19267), .B2(n19290), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19268) );
  OAI21_X1 U22174 ( .B1(n19269), .B2(n19652), .A(n19268), .ZN(n19291) );
  AOI22_X1 U22175 ( .A1(n19291), .A2(n19696), .B1(n19695), .B2(n19290), .ZN(
        n19273) );
  AOI21_X1 U22176 ( .B1(n10711), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19271) );
  OAI21_X1 U22177 ( .B1(n19445), .B2(n19502), .A(n19269), .ZN(n19270) );
  OAI211_X1 U22178 ( .C1(n19290), .C2(n19271), .A(n19270), .B(n19702), .ZN(
        n19293) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19649), .ZN(n19272) );
  OAI211_X1 U22180 ( .C1(n19663), .C2(n19327), .A(n19273), .B(n19272), .ZN(
        P2_U3056) );
  AOI22_X1 U22181 ( .A1(n19291), .A2(n19709), .B1(n19708), .B2(n19290), .ZN(
        n19276) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19594), .ZN(n19275) );
  OAI211_X1 U22183 ( .C1(n19597), .C2(n19327), .A(n19276), .B(n19275), .ZN(
        P2_U3057) );
  AOI22_X1 U22184 ( .A1(n19291), .A2(n19715), .B1(n19714), .B2(n19290), .ZN(
        n19279) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19666), .ZN(n19278) );
  OAI211_X1 U22186 ( .C1(n19669), .C2(n19327), .A(n19279), .B(n19278), .ZN(
        P2_U3058) );
  AOI22_X1 U22187 ( .A1(n19291), .A2(n19721), .B1(n19720), .B2(n19290), .ZN(
        n19282) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19670), .ZN(n19281) );
  OAI211_X1 U22189 ( .C1(n19673), .C2(n19327), .A(n19282), .B(n19281), .ZN(
        P2_U3059) );
  AOI22_X1 U22190 ( .A1(n19291), .A2(n19727), .B1(n19726), .B2(n19290), .ZN(
        n19284) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19602), .ZN(n19283) );
  OAI211_X1 U22192 ( .C1(n19605), .C2(n19327), .A(n19284), .B(n19283), .ZN(
        P2_U3060) );
  AOI22_X1 U22193 ( .A1(n19291), .A2(n19733), .B1(n19732), .B2(n19290), .ZN(
        n19286) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19606), .ZN(n19285) );
  OAI211_X1 U22195 ( .C1(n19609), .C2(n19327), .A(n19286), .B(n19285), .ZN(
        P2_U3061) );
  AOI22_X1 U22196 ( .A1(n19291), .A2(n19739), .B1(n19738), .B2(n19290), .ZN(
        n19288) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19639), .ZN(n19287) );
  OAI211_X1 U22198 ( .C1(n19642), .C2(n19327), .A(n19288), .B(n19287), .ZN(
        P2_U3062) );
  AOI22_X1 U22199 ( .A1(n19291), .A2(n19746), .B1(n19744), .B2(n19290), .ZN(
        n19295) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19293), .B1(
        n19292), .B2(n19684), .ZN(n19294) );
  OAI211_X1 U22201 ( .C1(n19689), .C2(n19327), .A(n19295), .B(n19294), .ZN(
        P2_U3063) );
  INV_X1 U22202 ( .A(n19301), .ZN(n19297) );
  NOR2_X1 U22203 ( .A1(n19296), .A2(n19328), .ZN(n19322) );
  OAI21_X1 U22204 ( .B1(n19297), .B2(n19322), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19299) );
  OR2_X1 U22205 ( .A1(n19298), .A2(n19328), .ZN(n19302) );
  NAND2_X1 U22206 ( .A1(n19299), .A2(n19302), .ZN(n19323) );
  AOI22_X1 U22207 ( .A1(n19323), .A2(n19696), .B1(n19695), .B2(n19322), .ZN(
        n19308) );
  INV_X1 U22208 ( .A(n19322), .ZN(n19300) );
  OAI21_X1 U22209 ( .B1(n19301), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19300), 
        .ZN(n19305) );
  OAI21_X1 U22210 ( .B1(n19353), .B2(n19319), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19303) );
  NAND2_X1 U22211 ( .A1(n19303), .A2(n19302), .ZN(n19304) );
  MUX2_X1 U22212 ( .A(n19305), .B(n19304), .S(n19864), .Z(n19306) );
  NAND2_X1 U22213 ( .A1(n19306), .A2(n19702), .ZN(n19324) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19324), .B1(
        n19353), .B2(n19704), .ZN(n19307) );
  OAI211_X1 U22215 ( .C1(n19707), .C2(n19327), .A(n19308), .B(n19307), .ZN(
        P2_U3064) );
  AOI22_X1 U22216 ( .A1(n19323), .A2(n19709), .B1(n19708), .B2(n19322), .ZN(
        n19310) );
  AOI22_X1 U22217 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19324), .B1(
        n19353), .B2(n19710), .ZN(n19309) );
  OAI211_X1 U22218 ( .C1(n19713), .C2(n19327), .A(n19310), .B(n19309), .ZN(
        P2_U3065) );
  AOI22_X1 U22219 ( .A1(n19323), .A2(n19715), .B1(n19714), .B2(n19322), .ZN(
        n19312) );
  AOI22_X1 U22220 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19324), .B1(
        n19353), .B2(n19716), .ZN(n19311) );
  OAI211_X1 U22221 ( .C1(n19719), .C2(n19327), .A(n19312), .B(n19311), .ZN(
        P2_U3066) );
  AOI22_X1 U22222 ( .A1(n19323), .A2(n19721), .B1(n19720), .B2(n19322), .ZN(
        n19314) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19324), .B1(
        n19319), .B2(n19670), .ZN(n19313) );
  OAI211_X1 U22224 ( .C1(n19673), .C2(n19351), .A(n19314), .B(n19313), .ZN(
        P2_U3067) );
  AOI22_X1 U22225 ( .A1(n19323), .A2(n19727), .B1(n19726), .B2(n19322), .ZN(
        n19316) );
  AOI22_X1 U22226 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19324), .B1(
        n19353), .B2(n19728), .ZN(n19315) );
  OAI211_X1 U22227 ( .C1(n19731), .C2(n19327), .A(n19316), .B(n19315), .ZN(
        P2_U3068) );
  AOI22_X1 U22228 ( .A1(n19323), .A2(n19733), .B1(n19732), .B2(n19322), .ZN(
        n19318) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19324), .B1(
        n19353), .B2(n19734), .ZN(n19317) );
  OAI211_X1 U22230 ( .C1(n19737), .C2(n19327), .A(n19318), .B(n19317), .ZN(
        P2_U3069) );
  AOI22_X1 U22231 ( .A1(n19323), .A2(n19739), .B1(n19738), .B2(n19322), .ZN(
        n19321) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19324), .B1(
        n19319), .B2(n19639), .ZN(n19320) );
  OAI211_X1 U22233 ( .C1(n19642), .C2(n19351), .A(n19321), .B(n19320), .ZN(
        P2_U3070) );
  INV_X1 U22234 ( .A(n19684), .ZN(n19754) );
  AOI22_X1 U22235 ( .A1(n19323), .A2(n19746), .B1(n19744), .B2(n19322), .ZN(
        n19326) );
  INV_X1 U22236 ( .A(n19689), .ZN(n19748) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19324), .B1(
        n19353), .B2(n19748), .ZN(n19325) );
  OAI211_X1 U22238 ( .C1(n19754), .C2(n19327), .A(n19326), .B(n19325), .ZN(
        P2_U3071) );
  NOR2_X1 U22239 ( .A1(n19554), .A2(n19328), .ZN(n19352) );
  AOI22_X1 U22240 ( .A1(n19649), .A2(n19353), .B1(n19695), .B2(n19352), .ZN(
        n19338) );
  OAI21_X1 U22241 ( .B1(n19445), .B2(n19859), .A(n19864), .ZN(n19336) );
  NOR2_X1 U22242 ( .A1(n19886), .A2(n19328), .ZN(n19332) );
  INV_X1 U22243 ( .A(n19352), .ZN(n19329) );
  OAI211_X1 U22244 ( .C1(n19330), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19329), 
        .B(n19652), .ZN(n19331) );
  OAI211_X1 U22245 ( .C1(n19336), .C2(n19332), .A(n19702), .B(n19331), .ZN(
        n19355) );
  INV_X1 U22246 ( .A(n19332), .ZN(n19335) );
  OAI21_X1 U22247 ( .B1(n19333), .B2(n19352), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19334) );
  OAI21_X1 U22248 ( .B1(n19336), .B2(n19335), .A(n19334), .ZN(n19354) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19355), .B1(
        n19696), .B2(n19354), .ZN(n19337) );
  OAI211_X1 U22250 ( .C1(n19663), .C2(n19388), .A(n19338), .B(n19337), .ZN(
        P2_U3072) );
  AOI22_X1 U22251 ( .A1(n19594), .A2(n19353), .B1(n19708), .B2(n19352), .ZN(
        n19340) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19355), .B1(
        n19709), .B2(n19354), .ZN(n19339) );
  OAI211_X1 U22253 ( .C1(n19597), .C2(n19388), .A(n19340), .B(n19339), .ZN(
        P2_U3073) );
  AOI22_X1 U22254 ( .A1(n19716), .A2(n19364), .B1(n19714), .B2(n19352), .ZN(
        n19342) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19355), .B1(
        n19715), .B2(n19354), .ZN(n19341) );
  OAI211_X1 U22256 ( .C1(n19719), .C2(n19351), .A(n19342), .B(n19341), .ZN(
        P2_U3074) );
  INV_X1 U22257 ( .A(n19673), .ZN(n19722) );
  AOI22_X1 U22258 ( .A1(n19722), .A2(n19364), .B1(n19720), .B2(n19352), .ZN(
        n19344) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19355), .B1(
        n19721), .B2(n19354), .ZN(n19343) );
  OAI211_X1 U22260 ( .C1(n19725), .C2(n19351), .A(n19344), .B(n19343), .ZN(
        P2_U3075) );
  AOI22_X1 U22261 ( .A1(n19602), .A2(n19353), .B1(n19352), .B2(n19726), .ZN(
        n19346) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19355), .B1(
        n19727), .B2(n19354), .ZN(n19345) );
  OAI211_X1 U22263 ( .C1(n19605), .C2(n19388), .A(n19346), .B(n19345), .ZN(
        P2_U3076) );
  AOI22_X1 U22264 ( .A1(n19606), .A2(n19353), .B1(n19352), .B2(n19732), .ZN(
        n19348) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19355), .B1(
        n19733), .B2(n19354), .ZN(n19347) );
  OAI211_X1 U22266 ( .C1(n19609), .C2(n19388), .A(n19348), .B(n19347), .ZN(
        P2_U3077) );
  AOI22_X1 U22267 ( .A1(n19740), .A2(n19364), .B1(n19352), .B2(n19738), .ZN(
        n19350) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19355), .B1(
        n19739), .B2(n19354), .ZN(n19349) );
  OAI211_X1 U22269 ( .C1(n19743), .C2(n19351), .A(n19350), .B(n19349), .ZN(
        P2_U3078) );
  AOI22_X1 U22270 ( .A1(n19684), .A2(n19353), .B1(n19744), .B2(n19352), .ZN(
        n19357) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19355), .B1(
        n19746), .B2(n19354), .ZN(n19356) );
  OAI211_X1 U22272 ( .C1(n19689), .C2(n19388), .A(n19357), .B(n19356), .ZN(
        P2_U3079) );
  OR2_X1 U22273 ( .A1(n19359), .A2(n19358), .ZN(n19588) );
  INV_X1 U22274 ( .A(n19588), .ZN(n19360) );
  NAND2_X1 U22275 ( .A1(n19360), .A2(n19869), .ZN(n19367) );
  INV_X1 U22276 ( .A(n19361), .ZN(n19363) );
  NOR2_X1 U22277 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19362), .ZN(
        n19383) );
  NOR3_X1 U22278 ( .A1(n19363), .A2(n19383), .A3(n19693), .ZN(n19365) );
  AOI211_X2 U22279 ( .C1(n19367), .C2(n19693), .A(n19443), .B(n19365), .ZN(
        n19384) );
  AOI22_X1 U22280 ( .A1(n19384), .A2(n19696), .B1(n19695), .B2(n19383), .ZN(
        n19370) );
  OAI21_X1 U22281 ( .B1(n19364), .B2(n19405), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19366) );
  AOI211_X1 U22282 ( .C1(n19367), .C2(n19366), .A(n19447), .B(n19365), .ZN(
        n19368) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19704), .ZN(n19369) );
  OAI211_X1 U22284 ( .C1(n19707), .C2(n19388), .A(n19370), .B(n19369), .ZN(
        P2_U3080) );
  AOI22_X1 U22285 ( .A1(n19384), .A2(n19709), .B1(n19708), .B2(n19383), .ZN(
        n19372) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19710), .ZN(n19371) );
  OAI211_X1 U22287 ( .C1(n19713), .C2(n19388), .A(n19372), .B(n19371), .ZN(
        P2_U3081) );
  AOI22_X1 U22288 ( .A1(n19384), .A2(n19715), .B1(n19714), .B2(n19383), .ZN(
        n19374) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19716), .ZN(n19373) );
  OAI211_X1 U22290 ( .C1(n19719), .C2(n19388), .A(n19374), .B(n19373), .ZN(
        P2_U3082) );
  AOI22_X1 U22291 ( .A1(n19384), .A2(n19721), .B1(n19720), .B2(n19383), .ZN(
        n19376) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19722), .ZN(n19375) );
  OAI211_X1 U22293 ( .C1(n19725), .C2(n19388), .A(n19376), .B(n19375), .ZN(
        P2_U3083) );
  AOI22_X1 U22294 ( .A1(n19384), .A2(n19727), .B1(n19726), .B2(n19383), .ZN(
        n19378) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19728), .ZN(n19377) );
  OAI211_X1 U22296 ( .C1(n19731), .C2(n19388), .A(n19378), .B(n19377), .ZN(
        P2_U3084) );
  AOI22_X1 U22297 ( .A1(n19384), .A2(n19733), .B1(n19732), .B2(n19383), .ZN(
        n19380) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19734), .ZN(n19379) );
  OAI211_X1 U22299 ( .C1(n19737), .C2(n19388), .A(n19380), .B(n19379), .ZN(
        P2_U3085) );
  AOI22_X1 U22300 ( .A1(n19384), .A2(n19739), .B1(n19738), .B2(n19383), .ZN(
        n19382) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19740), .ZN(n19381) );
  OAI211_X1 U22302 ( .C1(n19743), .C2(n19388), .A(n19382), .B(n19381), .ZN(
        P2_U3086) );
  AOI22_X1 U22303 ( .A1(n19384), .A2(n19746), .B1(n19744), .B2(n19383), .ZN(
        n19387) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19385), .B1(
        n19405), .B2(n19748), .ZN(n19386) );
  OAI211_X1 U22305 ( .C1(n19754), .C2(n19388), .A(n19387), .B(n19386), .ZN(
        P2_U3087) );
  INV_X1 U22306 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19392) );
  AOI22_X1 U22307 ( .A1(n19710), .A2(n19437), .B1(n19708), .B2(n19412), .ZN(
        n19391) );
  AOI22_X1 U22308 ( .A1(n19709), .A2(n19406), .B1(n19405), .B2(n19594), .ZN(
        n19390) );
  OAI211_X1 U22309 ( .C1(n19410), .C2(n19392), .A(n19391), .B(n19390), .ZN(
        P2_U3089) );
  INV_X1 U22310 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19395) );
  AOI22_X1 U22311 ( .A1(n19716), .A2(n19437), .B1(n19714), .B2(n19412), .ZN(
        n19394) );
  AOI22_X1 U22312 ( .A1(n19715), .A2(n19406), .B1(n19405), .B2(n19666), .ZN(
        n19393) );
  OAI211_X1 U22313 ( .C1(n19410), .C2(n19395), .A(n19394), .B(n19393), .ZN(
        P2_U3090) );
  AOI22_X1 U22314 ( .A1(n19722), .A2(n19437), .B1(n19720), .B2(n19412), .ZN(
        n19397) );
  AOI22_X1 U22315 ( .A1(n19721), .A2(n19406), .B1(n19405), .B2(n19670), .ZN(
        n19396) );
  OAI211_X1 U22316 ( .C1(n19410), .C2(n10496), .A(n19397), .B(n19396), .ZN(
        P2_U3091) );
  INV_X1 U22317 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19400) );
  AOI22_X1 U22318 ( .A1(n19728), .A2(n19437), .B1(n19412), .B2(n19726), .ZN(
        n19399) );
  AOI22_X1 U22319 ( .A1(n19727), .A2(n19406), .B1(n19405), .B2(n19602), .ZN(
        n19398) );
  OAI211_X1 U22320 ( .C1(n19410), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        P2_U3092) );
  AOI22_X1 U22321 ( .A1(n19606), .A2(n19405), .B1(n19412), .B2(n19732), .ZN(
        n19402) );
  AOI22_X1 U22322 ( .A1(n19733), .A2(n19406), .B1(n19437), .B2(n19734), .ZN(
        n19401) );
  OAI211_X1 U22323 ( .C1(n19410), .C2(n12862), .A(n19402), .B(n19401), .ZN(
        P2_U3093) );
  AOI22_X1 U22324 ( .A1(n19639), .A2(n19405), .B1(n19412), .B2(n19738), .ZN(
        n19404) );
  AOI22_X1 U22325 ( .A1(n19739), .A2(n19406), .B1(n19437), .B2(n19740), .ZN(
        n19403) );
  OAI211_X1 U22326 ( .C1(n19410), .C2(n12880), .A(n19404), .B(n19403), .ZN(
        P2_U3094) );
  INV_X1 U22327 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19409) );
  AOI22_X1 U22328 ( .A1(n19748), .A2(n19437), .B1(n19744), .B2(n19412), .ZN(
        n19408) );
  AOI22_X1 U22329 ( .A1(n19746), .A2(n19406), .B1(n19405), .B2(n19684), .ZN(
        n19407) );
  OAI211_X1 U22330 ( .C1(n19410), .C2(n19409), .A(n19408), .B(n19407), .ZN(
        P2_U3095) );
  NAND2_X1 U22331 ( .A1(n19869), .A2(n19692), .ZN(n19444) );
  NOR2_X1 U22332 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19444), .ZN(
        n19435) );
  NOR2_X1 U22333 ( .A1(n19412), .A2(n19435), .ZN(n19418) );
  INV_X1 U22334 ( .A(n19413), .ZN(n19416) );
  OAI21_X1 U22335 ( .B1(n19416), .B2(n19435), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19414) );
  OAI21_X1 U22336 ( .B1(n19418), .B2(n19652), .A(n19414), .ZN(n19436) );
  AOI22_X1 U22337 ( .A1(n19436), .A2(n19696), .B1(n19695), .B2(n19435), .ZN(
        n19422) );
  OAI21_X1 U22338 ( .B1(n19437), .B2(n19415), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19419) );
  AOI211_X1 U22339 ( .C1(n19416), .C2(n19888), .A(n19435), .B(n19864), .ZN(
        n19417) );
  AOI211_X1 U22340 ( .C1(n19419), .C2(n19418), .A(n19447), .B(n19417), .ZN(
        n19420) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19649), .ZN(n19421) );
  OAI211_X1 U22342 ( .C1(n19663), .C2(n19469), .A(n19422), .B(n19421), .ZN(
        P2_U3096) );
  AOI22_X1 U22343 ( .A1(n19436), .A2(n19709), .B1(n19708), .B2(n19435), .ZN(
        n19424) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19594), .ZN(n19423) );
  OAI211_X1 U22345 ( .C1(n19597), .C2(n19469), .A(n19424), .B(n19423), .ZN(
        P2_U3097) );
  AOI22_X1 U22346 ( .A1(n19436), .A2(n19715), .B1(n19714), .B2(n19435), .ZN(
        n19426) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19666), .ZN(n19425) );
  OAI211_X1 U22348 ( .C1(n19669), .C2(n19469), .A(n19426), .B(n19425), .ZN(
        P2_U3098) );
  AOI22_X1 U22349 ( .A1(n19436), .A2(n19721), .B1(n19720), .B2(n19435), .ZN(
        n19428) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19670), .ZN(n19427) );
  OAI211_X1 U22351 ( .C1(n19673), .C2(n19469), .A(n19428), .B(n19427), .ZN(
        P2_U3099) );
  AOI22_X1 U22352 ( .A1(n19436), .A2(n19727), .B1(n19726), .B2(n19435), .ZN(
        n19430) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19602), .ZN(n19429) );
  OAI211_X1 U22354 ( .C1(n19605), .C2(n19469), .A(n19430), .B(n19429), .ZN(
        P2_U3100) );
  AOI22_X1 U22355 ( .A1(n19436), .A2(n19733), .B1(n19732), .B2(n19435), .ZN(
        n19432) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19606), .ZN(n19431) );
  OAI211_X1 U22357 ( .C1(n19609), .C2(n19469), .A(n19432), .B(n19431), .ZN(
        P2_U3101) );
  AOI22_X1 U22358 ( .A1(n19436), .A2(n19739), .B1(n19738), .B2(n19435), .ZN(
        n19434) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19639), .ZN(n19433) );
  OAI211_X1 U22360 ( .C1(n19642), .C2(n19469), .A(n19434), .B(n19433), .ZN(
        P2_U3102) );
  AOI22_X1 U22361 ( .A1(n19436), .A2(n19746), .B1(n19744), .B2(n19435), .ZN(
        n19440) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19684), .ZN(n19439) );
  OAI211_X1 U22363 ( .C1(n19689), .C2(n19469), .A(n19440), .B(n19439), .ZN(
        P2_U3103) );
  NOR2_X1 U22364 ( .A1(n19896), .A2(n19444), .ZN(n19476) );
  INV_X1 U22365 ( .A(n19476), .ZN(n19473) );
  AND2_X1 U22366 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19473), .ZN(n19441) );
  AOI211_X2 U22367 ( .C1(n19444), .C2(n19693), .A(n19443), .B(n19446), .ZN(
        n19465) );
  AOI22_X1 U22368 ( .A1(n19465), .A2(n19696), .B1(n19695), .B2(n19476), .ZN(
        n19452) );
  INV_X1 U22369 ( .A(n19444), .ZN(n19449) );
  NOR2_X1 U22370 ( .A1(n19445), .A2(n19698), .ZN(n19863) );
  AOI211_X1 U22371 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19473), .A(n19447), 
        .B(n19446), .ZN(n19448) );
  OAI21_X1 U22372 ( .B1(n19449), .B2(n19863), .A(n19448), .ZN(n19466) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19704), .ZN(n19451) );
  OAI211_X1 U22374 ( .C1(n19707), .C2(n19469), .A(n19452), .B(n19451), .ZN(
        P2_U3104) );
  AOI22_X1 U22375 ( .A1(n19465), .A2(n19709), .B1(n19708), .B2(n19476), .ZN(
        n19454) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19710), .ZN(n19453) );
  OAI211_X1 U22377 ( .C1(n19713), .C2(n19469), .A(n19454), .B(n19453), .ZN(
        P2_U3105) );
  AOI22_X1 U22378 ( .A1(n19465), .A2(n19715), .B1(n19714), .B2(n19476), .ZN(
        n19456) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19716), .ZN(n19455) );
  OAI211_X1 U22380 ( .C1(n19719), .C2(n19469), .A(n19456), .B(n19455), .ZN(
        P2_U3106) );
  AOI22_X1 U22381 ( .A1(n19465), .A2(n19721), .B1(n19720), .B2(n19476), .ZN(
        n19458) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19722), .ZN(n19457) );
  OAI211_X1 U22383 ( .C1(n19725), .C2(n19469), .A(n19458), .B(n19457), .ZN(
        P2_U3107) );
  AOI22_X1 U22384 ( .A1(n19465), .A2(n19727), .B1(n19726), .B2(n19476), .ZN(
        n19460) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19728), .ZN(n19459) );
  OAI211_X1 U22386 ( .C1(n19731), .C2(n19469), .A(n19460), .B(n19459), .ZN(
        P2_U3108) );
  AOI22_X1 U22387 ( .A1(n19465), .A2(n19733), .B1(n19732), .B2(n19476), .ZN(
        n19462) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19734), .ZN(n19461) );
  OAI211_X1 U22389 ( .C1(n19737), .C2(n19469), .A(n19462), .B(n19461), .ZN(
        P2_U3109) );
  AOI22_X1 U22390 ( .A1(n19465), .A2(n19739), .B1(n19738), .B2(n19476), .ZN(
        n19464) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19740), .ZN(n19463) );
  OAI211_X1 U22392 ( .C1(n19743), .C2(n19469), .A(n19464), .B(n19463), .ZN(
        P2_U3110) );
  AOI22_X1 U22393 ( .A1(n19465), .A2(n19746), .B1(n19744), .B2(n19476), .ZN(
        n19468) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19466), .B1(
        n19492), .B2(n19748), .ZN(n19467) );
  OAI211_X1 U22395 ( .C1(n19754), .C2(n19469), .A(n19468), .B(n19467), .ZN(
        P2_U3111) );
  NOR2_X1 U22396 ( .A1(n19553), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19503) );
  INV_X1 U22397 ( .A(n19503), .ZN(n19508) );
  NOR2_X1 U22398 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19508), .ZN(
        n19495) );
  AOI22_X1 U22399 ( .A1(n19704), .A2(n19520), .B1(n19695), .B2(n19495), .ZN(
        n19481) );
  AOI21_X1 U22400 ( .B1(n19531), .B2(n19500), .A(n19470), .ZN(n19471) );
  NOR2_X1 U22401 ( .A1(n19471), .A2(n19652), .ZN(n19475) );
  INV_X1 U22402 ( .A(n10699), .ZN(n19477) );
  OAI21_X1 U22403 ( .B1(n19477), .B2(n19693), .A(n19888), .ZN(n19472) );
  AOI21_X1 U22404 ( .B1(n19475), .B2(n19473), .A(n19472), .ZN(n19474) );
  OAI21_X1 U22405 ( .B1(n19495), .B2(n19474), .A(n19702), .ZN(n19497) );
  OAI21_X1 U22406 ( .B1(n19495), .B2(n19476), .A(n19475), .ZN(n19479) );
  OAI21_X1 U22407 ( .B1(n19477), .B2(n19495), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19478) );
  NAND2_X1 U22408 ( .A1(n19479), .A2(n19478), .ZN(n19496) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19497), .B1(
        n19696), .B2(n19496), .ZN(n19480) );
  OAI211_X1 U22410 ( .C1(n19707), .C2(n19500), .A(n19481), .B(n19480), .ZN(
        P2_U3112) );
  AOI22_X1 U22411 ( .A1(n19710), .A2(n19520), .B1(n19708), .B2(n19495), .ZN(
        n19483) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19709), .ZN(n19482) );
  OAI211_X1 U22413 ( .C1(n19713), .C2(n19500), .A(n19483), .B(n19482), .ZN(
        P2_U3113) );
  AOI22_X1 U22414 ( .A1(n19716), .A2(n19520), .B1(n19714), .B2(n19495), .ZN(
        n19485) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19715), .ZN(n19484) );
  OAI211_X1 U22416 ( .C1(n19719), .C2(n19500), .A(n19485), .B(n19484), .ZN(
        P2_U3114) );
  AOI22_X1 U22417 ( .A1(n19670), .A2(n19492), .B1(n19720), .B2(n19495), .ZN(
        n19487) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19721), .ZN(n19486) );
  OAI211_X1 U22419 ( .C1(n19673), .C2(n19531), .A(n19487), .B(n19486), .ZN(
        P2_U3115) );
  AOI22_X1 U22420 ( .A1(n19728), .A2(n19520), .B1(n19495), .B2(n19726), .ZN(
        n19489) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19727), .ZN(n19488) );
  OAI211_X1 U22422 ( .C1(n19731), .C2(n19500), .A(n19489), .B(n19488), .ZN(
        P2_U3116) );
  AOI22_X1 U22423 ( .A1(n19606), .A2(n19492), .B1(n19495), .B2(n19732), .ZN(
        n19491) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19733), .ZN(n19490) );
  OAI211_X1 U22425 ( .C1(n19609), .C2(n19531), .A(n19491), .B(n19490), .ZN(
        P2_U3117) );
  AOI22_X1 U22426 ( .A1(n19639), .A2(n19492), .B1(n19495), .B2(n19738), .ZN(
        n19494) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19739), .ZN(n19493) );
  OAI211_X1 U22428 ( .C1(n19642), .C2(n19531), .A(n19494), .B(n19493), .ZN(
        P2_U3118) );
  AOI22_X1 U22429 ( .A1(n19748), .A2(n19520), .B1(n19744), .B2(n19495), .ZN(
        n19499) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19746), .ZN(n19498) );
  OAI211_X1 U22431 ( .C1(n19754), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P2_U3119) );
  NOR2_X1 U22432 ( .A1(n19501), .A2(n19553), .ZN(n19526) );
  AOI22_X1 U22433 ( .A1(n19704), .A2(n19547), .B1(n19695), .B2(n19526), .ZN(
        n19511) );
  AOI21_X1 U22434 ( .B1(n10707), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19505) );
  NAND2_X1 U22435 ( .A1(n19866), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19699) );
  OAI21_X1 U22436 ( .B1(n19699), .B2(n19502), .A(n19864), .ZN(n19509) );
  OR2_X1 U22437 ( .A1(n19509), .A2(n19503), .ZN(n19504) );
  OAI211_X1 U22438 ( .C1(n19526), .C2(n19505), .A(n19504), .B(n19702), .ZN(
        n19528) );
  INV_X1 U22439 ( .A(n10707), .ZN(n19506) );
  OAI21_X1 U22440 ( .B1(n19506), .B2(n19526), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19507) );
  OAI21_X1 U22441 ( .B1(n19509), .B2(n19508), .A(n19507), .ZN(n19527) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19528), .B1(
        n19696), .B2(n19527), .ZN(n19510) );
  OAI211_X1 U22443 ( .C1(n19707), .C2(n19531), .A(n19511), .B(n19510), .ZN(
        P2_U3120) );
  AOI22_X1 U22444 ( .A1(n19594), .A2(n19520), .B1(n19708), .B2(n19526), .ZN(
        n19513) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19528), .B1(
        n19709), .B2(n19527), .ZN(n19512) );
  OAI211_X1 U22446 ( .C1(n19597), .C2(n19523), .A(n19513), .B(n19512), .ZN(
        P2_U3121) );
  AOI22_X1 U22447 ( .A1(n19716), .A2(n19547), .B1(n19714), .B2(n19526), .ZN(
        n19515) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19528), .B1(
        n19715), .B2(n19527), .ZN(n19514) );
  OAI211_X1 U22449 ( .C1(n19719), .C2(n19531), .A(n19515), .B(n19514), .ZN(
        P2_U3122) );
  AOI22_X1 U22450 ( .A1(n19722), .A2(n19547), .B1(n19720), .B2(n19526), .ZN(
        n19517) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19528), .B1(
        n19721), .B2(n19527), .ZN(n19516) );
  OAI211_X1 U22452 ( .C1(n19725), .C2(n19531), .A(n19517), .B(n19516), .ZN(
        P2_U3123) );
  AOI22_X1 U22453 ( .A1(n19728), .A2(n19547), .B1(n19726), .B2(n19526), .ZN(
        n19519) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19528), .B1(
        n19727), .B2(n19527), .ZN(n19518) );
  OAI211_X1 U22455 ( .C1(n19731), .C2(n19531), .A(n19519), .B(n19518), .ZN(
        P2_U3124) );
  AOI22_X1 U22456 ( .A1(n19606), .A2(n19520), .B1(n19526), .B2(n19732), .ZN(
        n19522) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19528), .B1(
        n19733), .B2(n19527), .ZN(n19521) );
  OAI211_X1 U22458 ( .C1(n19609), .C2(n19523), .A(n19522), .B(n19521), .ZN(
        P2_U3125) );
  AOI22_X1 U22459 ( .A1(n19740), .A2(n19547), .B1(n19526), .B2(n19738), .ZN(
        n19525) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19528), .B1(
        n19739), .B2(n19527), .ZN(n19524) );
  OAI211_X1 U22461 ( .C1(n19743), .C2(n19531), .A(n19525), .B(n19524), .ZN(
        P2_U3126) );
  AOI22_X1 U22462 ( .A1(n19748), .A2(n19547), .B1(n19744), .B2(n19526), .ZN(
        n19530) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19528), .B1(
        n19746), .B2(n19527), .ZN(n19529) );
  OAI211_X1 U22464 ( .C1(n19754), .C2(n19531), .A(n19530), .B(n19529), .ZN(
        P2_U3127) );
  AOI22_X1 U22465 ( .A1(n19594), .A2(n19547), .B1(n19546), .B2(n19708), .ZN(
        n19533) );
  AOI22_X1 U22466 ( .A1(n19709), .A2(n19548), .B1(n19579), .B2(n19710), .ZN(
        n19532) );
  OAI211_X1 U22467 ( .C1(n19552), .C2(n12630), .A(n19533), .B(n19532), .ZN(
        P2_U3129) );
  INV_X1 U22468 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n19536) );
  AOI22_X1 U22469 ( .A1(n19716), .A2(n19579), .B1(n19546), .B2(n19714), .ZN(
        n19535) );
  AOI22_X1 U22470 ( .A1(n19715), .A2(n19548), .B1(n19547), .B2(n19666), .ZN(
        n19534) );
  OAI211_X1 U22471 ( .C1(n19552), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P2_U3130) );
  AOI22_X1 U22472 ( .A1(n19722), .A2(n19579), .B1(n19546), .B2(n19720), .ZN(
        n19538) );
  AOI22_X1 U22473 ( .A1(n19721), .A2(n19548), .B1(n19547), .B2(n19670), .ZN(
        n19537) );
  OAI211_X1 U22474 ( .C1(n19552), .C2(n10478), .A(n19538), .B(n19537), .ZN(
        P2_U3131) );
  INV_X1 U22475 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n19541) );
  AOI22_X1 U22476 ( .A1(n19728), .A2(n19579), .B1(n19546), .B2(n19726), .ZN(
        n19540) );
  AOI22_X1 U22477 ( .A1(n19727), .A2(n19548), .B1(n19547), .B2(n19602), .ZN(
        n19539) );
  OAI211_X1 U22478 ( .C1(n19552), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3132) );
  AOI22_X1 U22479 ( .A1(n19734), .A2(n19579), .B1(n19546), .B2(n19732), .ZN(
        n19543) );
  AOI22_X1 U22480 ( .A1(n19733), .A2(n19548), .B1(n19547), .B2(n19606), .ZN(
        n19542) );
  OAI211_X1 U22481 ( .C1(n19552), .C2(n10700), .A(n19543), .B(n19542), .ZN(
        P2_U3133) );
  AOI22_X1 U22482 ( .A1(n19740), .A2(n19579), .B1(n19546), .B2(n19738), .ZN(
        n19545) );
  AOI22_X1 U22483 ( .A1(n19739), .A2(n19548), .B1(n19547), .B2(n19639), .ZN(
        n19544) );
  OAI211_X1 U22484 ( .C1(n19552), .C2(n12896), .A(n19545), .B(n19544), .ZN(
        P2_U3134) );
  INV_X1 U22485 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19551) );
  AOI22_X1 U22486 ( .A1(n19684), .A2(n19547), .B1(n19546), .B2(n19744), .ZN(
        n19550) );
  AOI22_X1 U22487 ( .A1(n19746), .A2(n19548), .B1(n19579), .B2(n19748), .ZN(
        n19549) );
  OAI211_X1 U22488 ( .C1(n19552), .C2(n19551), .A(n19550), .B(n19549), .ZN(
        P2_U3135) );
  NOR2_X1 U22489 ( .A1(n19554), .A2(n19553), .ZN(n19577) );
  NOR2_X1 U22490 ( .A1(n19577), .A2(n19693), .ZN(n19555) );
  NAND2_X1 U22491 ( .A1(n19556), .A2(n19555), .ZN(n19560) );
  NAND2_X1 U22492 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19557), .ZN(
        n19559) );
  OAI21_X1 U22493 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19559), .A(n19693), 
        .ZN(n19558) );
  AND2_X1 U22494 ( .A1(n19560), .A2(n19558), .ZN(n19578) );
  AOI22_X1 U22495 ( .A1(n19578), .A2(n19696), .B1(n19695), .B2(n19577), .ZN(
        n19564) );
  OAI21_X1 U22496 ( .B1(n19699), .B2(n19859), .A(n19559), .ZN(n19561) );
  AND2_X1 U22497 ( .A1(n19561), .A2(n19560), .ZN(n19562) );
  OAI211_X1 U22498 ( .C1(n19577), .C2(n19888), .A(n19562), .B(n19702), .ZN(
        n19580) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19649), .ZN(n19563) );
  OAI211_X1 U22500 ( .C1(n19663), .C2(n19583), .A(n19564), .B(n19563), .ZN(
        P2_U3136) );
  AOI22_X1 U22501 ( .A1(n19578), .A2(n19709), .B1(n19708), .B2(n19577), .ZN(
        n19566) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19594), .ZN(n19565) );
  OAI211_X1 U22503 ( .C1(n19597), .C2(n19583), .A(n19566), .B(n19565), .ZN(
        P2_U3137) );
  AOI22_X1 U22504 ( .A1(n19578), .A2(n19715), .B1(n19714), .B2(n19577), .ZN(
        n19568) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19666), .ZN(n19567) );
  OAI211_X1 U22506 ( .C1(n19669), .C2(n19583), .A(n19568), .B(n19567), .ZN(
        P2_U3138) );
  AOI22_X1 U22507 ( .A1(n19578), .A2(n19721), .B1(n19720), .B2(n19577), .ZN(
        n19570) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19670), .ZN(n19569) );
  OAI211_X1 U22509 ( .C1(n19673), .C2(n19583), .A(n19570), .B(n19569), .ZN(
        P2_U3139) );
  AOI22_X1 U22510 ( .A1(n19578), .A2(n19727), .B1(n19726), .B2(n19577), .ZN(
        n19572) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19602), .ZN(n19571) );
  OAI211_X1 U22512 ( .C1(n19605), .C2(n19583), .A(n19572), .B(n19571), .ZN(
        P2_U3140) );
  AOI22_X1 U22513 ( .A1(n19578), .A2(n19733), .B1(n19732), .B2(n19577), .ZN(
        n19574) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19606), .ZN(n19573) );
  OAI211_X1 U22515 ( .C1(n19609), .C2(n19583), .A(n19574), .B(n19573), .ZN(
        P2_U3141) );
  AOI22_X1 U22516 ( .A1(n19578), .A2(n19739), .B1(n19738), .B2(n19577), .ZN(
        n19576) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19639), .ZN(n19575) );
  OAI211_X1 U22518 ( .C1(n19642), .C2(n19583), .A(n19576), .B(n19575), .ZN(
        P2_U3142) );
  AOI22_X1 U22519 ( .A1(n19578), .A2(n19746), .B1(n19744), .B2(n19577), .ZN(
        n19582) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19580), .B1(
        n19579), .B2(n19684), .ZN(n19581) );
  OAI211_X1 U22521 ( .C1(n19689), .C2(n19583), .A(n19582), .B(n19581), .ZN(
        P2_U3143) );
  INV_X1 U22522 ( .A(n19584), .ZN(n19586) );
  NAND3_X1 U22523 ( .A1(n19886), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19619) );
  NOR2_X1 U22524 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19619), .ZN(
        n19612) );
  OAI21_X1 U22525 ( .B1(n10557), .B2(n19612), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19585) );
  OAI21_X1 U22526 ( .B1(n19586), .B2(n19588), .A(n19585), .ZN(n19613) );
  AOI22_X1 U22527 ( .A1(n19613), .A2(n19696), .B1(n19695), .B2(n19612), .ZN(
        n19593) );
  OAI21_X1 U22528 ( .B1(n19644), .B2(n19614), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19587) );
  OAI21_X1 U22529 ( .B1(n19588), .B2(n19869), .A(n19587), .ZN(n19591) );
  INV_X1 U22530 ( .A(n19612), .ZN(n19589) );
  OAI211_X1 U22531 ( .C1(n10696), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19589), 
        .B(n19652), .ZN(n19590) );
  NAND3_X1 U22532 ( .A1(n19591), .A2(n19702), .A3(n19590), .ZN(n19615) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19649), .ZN(n19592) );
  OAI211_X1 U22534 ( .C1(n19663), .C2(n19638), .A(n19593), .B(n19592), .ZN(
        P2_U3144) );
  AOI22_X1 U22535 ( .A1(n19613), .A2(n19709), .B1(n19708), .B2(n19612), .ZN(
        n19596) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19594), .ZN(n19595) );
  OAI211_X1 U22537 ( .C1(n19597), .C2(n19638), .A(n19596), .B(n19595), .ZN(
        P2_U3145) );
  AOI22_X1 U22538 ( .A1(n19613), .A2(n19715), .B1(n19714), .B2(n19612), .ZN(
        n19599) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19666), .ZN(n19598) );
  OAI211_X1 U22540 ( .C1(n19669), .C2(n19638), .A(n19599), .B(n19598), .ZN(
        P2_U3146) );
  AOI22_X1 U22541 ( .A1(n19613), .A2(n19721), .B1(n19720), .B2(n19612), .ZN(
        n19601) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19670), .ZN(n19600) );
  OAI211_X1 U22543 ( .C1(n19673), .C2(n19638), .A(n19601), .B(n19600), .ZN(
        P2_U3147) );
  AOI22_X1 U22544 ( .A1(n19613), .A2(n19727), .B1(n19726), .B2(n19612), .ZN(
        n19604) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19602), .ZN(n19603) );
  OAI211_X1 U22546 ( .C1(n19605), .C2(n19638), .A(n19604), .B(n19603), .ZN(
        P2_U3148) );
  AOI22_X1 U22547 ( .A1(n19613), .A2(n19733), .B1(n19732), .B2(n19612), .ZN(
        n19608) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19606), .ZN(n19607) );
  OAI211_X1 U22549 ( .C1(n19609), .C2(n19638), .A(n19608), .B(n19607), .ZN(
        P2_U3149) );
  AOI22_X1 U22550 ( .A1(n19613), .A2(n19739), .B1(n19738), .B2(n19612), .ZN(
        n19611) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19639), .ZN(n19610) );
  OAI211_X1 U22552 ( .C1(n19642), .C2(n19638), .A(n19611), .B(n19610), .ZN(
        P2_U3150) );
  AOI22_X1 U22553 ( .A1(n19613), .A2(n19746), .B1(n19744), .B2(n19612), .ZN(
        n19617) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19684), .ZN(n19616) );
  OAI211_X1 U22555 ( .C1(n19689), .C2(n19638), .A(n19617), .B(n19616), .ZN(
        P2_U3151) );
  INV_X1 U22556 ( .A(n10708), .ZN(n19620) );
  NOR2_X1 U22557 ( .A1(n19896), .A2(n19619), .ZN(n19651) );
  OAI21_X1 U22558 ( .B1(n19620), .B2(n19651), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19618) );
  OAI21_X1 U22559 ( .B1(n19619), .B2(n19652), .A(n19618), .ZN(n19643) );
  AOI22_X1 U22560 ( .A1(n19643), .A2(n19696), .B1(n19695), .B2(n19651), .ZN(
        n19627) );
  OAI21_X1 U22561 ( .B1(n19699), .B2(n19624), .A(n19619), .ZN(n19623) );
  INV_X1 U22562 ( .A(n19651), .ZN(n19621) );
  OAI211_X1 U22563 ( .C1(n10708), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19621), 
        .B(n19652), .ZN(n19622) );
  NAND3_X1 U22564 ( .A1(n19623), .A2(n19702), .A3(n19622), .ZN(n19645) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19645), .B1(
        n19683), .B2(n19704), .ZN(n19626) );
  OAI211_X1 U22566 ( .C1(n19707), .C2(n19638), .A(n19627), .B(n19626), .ZN(
        P2_U3152) );
  AOI22_X1 U22567 ( .A1(n19643), .A2(n19709), .B1(n19708), .B2(n19651), .ZN(
        n19629) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19645), .B1(
        n19683), .B2(n19710), .ZN(n19628) );
  OAI211_X1 U22569 ( .C1(n19713), .C2(n19638), .A(n19629), .B(n19628), .ZN(
        P2_U3153) );
  AOI22_X1 U22570 ( .A1(n19643), .A2(n19715), .B1(n19714), .B2(n19651), .ZN(
        n19631) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19645), .B1(
        n19683), .B2(n19716), .ZN(n19630) );
  OAI211_X1 U22572 ( .C1(n19719), .C2(n19638), .A(n19631), .B(n19630), .ZN(
        P2_U3154) );
  AOI22_X1 U22573 ( .A1(n19643), .A2(n19721), .B1(n19720), .B2(n19651), .ZN(
        n19633) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19645), .B1(
        n19644), .B2(n19670), .ZN(n19632) );
  OAI211_X1 U22575 ( .C1(n19673), .C2(n19681), .A(n19633), .B(n19632), .ZN(
        P2_U3155) );
  AOI22_X1 U22576 ( .A1(n19643), .A2(n19727), .B1(n19726), .B2(n19651), .ZN(
        n19635) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19645), .B1(
        n19683), .B2(n19728), .ZN(n19634) );
  OAI211_X1 U22578 ( .C1(n19731), .C2(n19638), .A(n19635), .B(n19634), .ZN(
        P2_U3156) );
  AOI22_X1 U22579 ( .A1(n19643), .A2(n19733), .B1(n19732), .B2(n19651), .ZN(
        n19637) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19645), .B1(
        n19683), .B2(n19734), .ZN(n19636) );
  OAI211_X1 U22581 ( .C1(n19737), .C2(n19638), .A(n19637), .B(n19636), .ZN(
        P2_U3157) );
  AOI22_X1 U22582 ( .A1(n19643), .A2(n19739), .B1(n19738), .B2(n19651), .ZN(
        n19641) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19645), .B1(
        n19644), .B2(n19639), .ZN(n19640) );
  OAI211_X1 U22584 ( .C1(n19642), .C2(n19681), .A(n19641), .B(n19640), .ZN(
        P2_U3158) );
  AOI22_X1 U22585 ( .A1(n19643), .A2(n19746), .B1(n19744), .B2(n19651), .ZN(
        n19647) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19645), .B1(
        n19644), .B2(n19684), .ZN(n19646) );
  OAI211_X1 U22587 ( .C1(n19689), .C2(n19681), .A(n19647), .B(n19646), .ZN(
        P2_U3159) );
  AND3_X1 U22588 ( .A1(n19896), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19692), .ZN(n19682) );
  AOI22_X1 U22589 ( .A1(n19649), .A2(n19683), .B1(n19695), .B2(n19682), .ZN(
        n19662) );
  OAI21_X1 U22590 ( .B1(n19683), .B2(n19678), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19650) );
  NAND2_X1 U22591 ( .A1(n19650), .A2(n19864), .ZN(n19660) );
  NOR2_X1 U22592 ( .A1(n19682), .A2(n19651), .ZN(n19659) );
  INV_X1 U22593 ( .A(n19659), .ZN(n19655) );
  INV_X1 U22594 ( .A(n19682), .ZN(n19653) );
  OAI211_X1 U22595 ( .C1(n19656), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19653), 
        .B(n19652), .ZN(n19654) );
  OAI211_X1 U22596 ( .C1(n19660), .C2(n19655), .A(n19702), .B(n19654), .ZN(
        n19686) );
  INV_X1 U22597 ( .A(n19656), .ZN(n19657) );
  OAI21_X1 U22598 ( .B1(n19657), .B2(n19682), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19658) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19686), .B1(
        n19696), .B2(n19685), .ZN(n19661) );
  OAI211_X1 U22600 ( .C1(n19663), .C2(n19753), .A(n19662), .B(n19661), .ZN(
        P2_U3160) );
  AOI22_X1 U22601 ( .A1(n19710), .A2(n19678), .B1(n19708), .B2(n19682), .ZN(
        n19665) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19686), .B1(
        n19709), .B2(n19685), .ZN(n19664) );
  OAI211_X1 U22603 ( .C1(n19713), .C2(n19681), .A(n19665), .B(n19664), .ZN(
        P2_U3161) );
  AOI22_X1 U22604 ( .A1(n19666), .A2(n19683), .B1(n19714), .B2(n19682), .ZN(
        n19668) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19686), .B1(
        n19715), .B2(n19685), .ZN(n19667) );
  OAI211_X1 U22606 ( .C1(n19669), .C2(n19753), .A(n19668), .B(n19667), .ZN(
        P2_U3162) );
  AOI22_X1 U22607 ( .A1(n19670), .A2(n19683), .B1(n19720), .B2(n19682), .ZN(
        n19672) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19686), .B1(
        n19721), .B2(n19685), .ZN(n19671) );
  OAI211_X1 U22609 ( .C1(n19673), .C2(n19753), .A(n19672), .B(n19671), .ZN(
        P2_U3163) );
  AOI22_X1 U22610 ( .A1(n19728), .A2(n19678), .B1(n19726), .B2(n19682), .ZN(
        n19675) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19686), .B1(
        n19727), .B2(n19685), .ZN(n19674) );
  OAI211_X1 U22612 ( .C1(n19731), .C2(n19681), .A(n19675), .B(n19674), .ZN(
        P2_U3164) );
  AOI22_X1 U22613 ( .A1(n19734), .A2(n19678), .B1(n19732), .B2(n19682), .ZN(
        n19677) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19686), .B1(
        n19733), .B2(n19685), .ZN(n19676) );
  OAI211_X1 U22615 ( .C1(n19737), .C2(n19681), .A(n19677), .B(n19676), .ZN(
        P2_U3165) );
  AOI22_X1 U22616 ( .A1(n19740), .A2(n19678), .B1(n19682), .B2(n19738), .ZN(
        n19680) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19686), .B1(
        n19739), .B2(n19685), .ZN(n19679) );
  OAI211_X1 U22618 ( .C1(n19743), .C2(n19681), .A(n19680), .B(n19679), .ZN(
        P2_U3166) );
  AOI22_X1 U22619 ( .A1(n19684), .A2(n19683), .B1(n19744), .B2(n19682), .ZN(
        n19688) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19686), .B1(
        n19746), .B2(n19685), .ZN(n19687) );
  OAI211_X1 U22621 ( .C1(n19689), .C2(n19753), .A(n19688), .B(n19687), .ZN(
        P2_U3167) );
  NOR2_X1 U22622 ( .A1(n19745), .A2(n19693), .ZN(n19690) );
  NAND2_X1 U22623 ( .A1(n19691), .A2(n19690), .ZN(n19700) );
  NAND2_X1 U22624 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19692), .ZN(
        n19697) );
  OAI21_X1 U22625 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19697), .A(n19693), 
        .ZN(n19694) );
  AND2_X1 U22626 ( .A1(n19700), .A2(n19694), .ZN(n19747) );
  AOI22_X1 U22627 ( .A1(n19747), .A2(n19696), .B1(n19745), .B2(n19695), .ZN(
        n19706) );
  OAI21_X1 U22628 ( .B1(n19699), .B2(n19698), .A(n19697), .ZN(n19701) );
  AND2_X1 U22629 ( .A1(n19701), .A2(n19700), .ZN(n19703) );
  OAI211_X1 U22630 ( .C1(n19745), .C2(n19888), .A(n19703), .B(n19702), .ZN(
        n19750) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19704), .ZN(n19705) );
  OAI211_X1 U22632 ( .C1(n19707), .C2(n19753), .A(n19706), .B(n19705), .ZN(
        P2_U3168) );
  AOI22_X1 U22633 ( .A1(n19747), .A2(n19709), .B1(n19745), .B2(n19708), .ZN(
        n19712) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19710), .ZN(n19711) );
  OAI211_X1 U22635 ( .C1(n19713), .C2(n19753), .A(n19712), .B(n19711), .ZN(
        P2_U3169) );
  AOI22_X1 U22636 ( .A1(n19747), .A2(n19715), .B1(n19745), .B2(n19714), .ZN(
        n19718) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19716), .ZN(n19717) );
  OAI211_X1 U22638 ( .C1(n19719), .C2(n19753), .A(n19718), .B(n19717), .ZN(
        P2_U3170) );
  AOI22_X1 U22639 ( .A1(n19747), .A2(n19721), .B1(n19745), .B2(n19720), .ZN(
        n19724) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19722), .ZN(n19723) );
  OAI211_X1 U22641 ( .C1(n19725), .C2(n19753), .A(n19724), .B(n19723), .ZN(
        P2_U3171) );
  AOI22_X1 U22642 ( .A1(n19747), .A2(n19727), .B1(n19745), .B2(n19726), .ZN(
        n19730) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19728), .ZN(n19729) );
  OAI211_X1 U22644 ( .C1(n19731), .C2(n19753), .A(n19730), .B(n19729), .ZN(
        P2_U3172) );
  AOI22_X1 U22645 ( .A1(n19747), .A2(n19733), .B1(n19745), .B2(n19732), .ZN(
        n19736) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19734), .ZN(n19735) );
  OAI211_X1 U22647 ( .C1(n19737), .C2(n19753), .A(n19736), .B(n19735), .ZN(
        P2_U3173) );
  AOI22_X1 U22648 ( .A1(n19747), .A2(n19739), .B1(n19745), .B2(n19738), .ZN(
        n19742) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19740), .ZN(n19741) );
  OAI211_X1 U22650 ( .C1(n19743), .C2(n19753), .A(n19742), .B(n19741), .ZN(
        P2_U3174) );
  AOI22_X1 U22651 ( .A1(n19747), .A2(n19746), .B1(n19745), .B2(n19744), .ZN(
        n19752) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n19748), .ZN(n19751) );
  OAI211_X1 U22653 ( .C1(n19754), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        P2_U3175) );
  OAI211_X1 U22654 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19764), .A(n19756), 
        .B(n19755), .ZN(n19761) );
  OAI21_X1 U22655 ( .B1(n19758), .B2(n19757), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19760) );
  OAI211_X1 U22656 ( .C1(n19762), .C2(n19761), .A(n19760), .B(n19759), .ZN(
        P2_U3177) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19763), .ZN(
        P2_U3179) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19763), .ZN(
        P2_U3180) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19763), .ZN(
        P2_U3181) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19763), .ZN(
        P2_U3182) );
  AND2_X1 U22661 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19763), .ZN(
        P2_U3183) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19763), .ZN(
        P2_U3184) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19763), .ZN(
        P2_U3185) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19763), .ZN(
        P2_U3186) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19763), .ZN(
        P2_U3187) );
  AND2_X1 U22666 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19763), .ZN(
        P2_U3188) );
  AND2_X1 U22667 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19763), .ZN(
        P2_U3189) );
  AND2_X1 U22668 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19763), .ZN(
        P2_U3190) );
  INV_X1 U22669 ( .A(P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20782) );
  NOR2_X1 U22670 ( .A1(n20782), .A2(n19845), .ZN(P2_U3191) );
  AND2_X1 U22671 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19763), .ZN(
        P2_U3192) );
  AND2_X1 U22672 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19763), .ZN(
        P2_U3193) );
  AND2_X1 U22673 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19763), .ZN(
        P2_U3194) );
  AND2_X1 U22674 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19763), .ZN(
        P2_U3195) );
  AND2_X1 U22675 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19763), .ZN(
        P2_U3196) );
  AND2_X1 U22676 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19763), .ZN(
        P2_U3197) );
  AND2_X1 U22677 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19763), .ZN(
        P2_U3198) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19763), .ZN(
        P2_U3199) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19763), .ZN(
        P2_U3200) );
  AND2_X1 U22680 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19763), .ZN(P2_U3201) );
  AND2_X1 U22681 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19763), .ZN(P2_U3202) );
  AND2_X1 U22682 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19763), .ZN(P2_U3203) );
  AND2_X1 U22683 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19763), .ZN(P2_U3204) );
  AND2_X1 U22684 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19763), .ZN(P2_U3205) );
  AND2_X1 U22685 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19763), .ZN(P2_U3206) );
  AND2_X1 U22686 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19763), .ZN(P2_U3207) );
  AND2_X1 U22687 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19763), .ZN(P2_U3208) );
  INV_X1 U22688 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19776) );
  NOR2_X1 U22689 ( .A1(n19764), .A2(n19776), .ZN(n19773) );
  OR3_X1 U22690 ( .A1(n19774), .A2(n19765), .A3(n19773), .ZN(n19766) );
  INV_X1 U22691 ( .A(NA), .ZN(n20653) );
  NOR3_X1 U22692 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20653), .ZN(n19781) );
  AOI21_X1 U22693 ( .B1(n19784), .B2(n19766), .A(n19781), .ZN(n19767) );
  OAI221_X1 U22694 ( .B1(n19768), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19768), .C2(n20648), .A(n19767), .ZN(P2_U3209) );
  AOI21_X1 U22695 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20648), .A(n19784), 
        .ZN(n19777) );
  NOR3_X1 U22696 ( .A1(n19777), .A2(n19774), .A3(n19765), .ZN(n19769) );
  NOR2_X1 U22697 ( .A1(n19769), .A2(n19773), .ZN(n19771) );
  OAI211_X1 U22698 ( .C1(n20648), .C2(n19772), .A(n19771), .B(n19770), .ZN(
        P2_U3210) );
  AOI22_X1 U22699 ( .A1(n19775), .A2(n19774), .B1(n19773), .B2(n20653), .ZN(
        n19783) );
  OAI21_X1 U22700 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19782) );
  NOR2_X1 U22701 ( .A1(n19776), .A2(n19784), .ZN(n19779) );
  AOI21_X1 U22702 ( .B1(n19779), .B2(n19778), .A(n19777), .ZN(n19780) );
  OAI22_X1 U22703 ( .A1(n19783), .A2(n19782), .B1(n19781), .B2(n19780), .ZN(
        P2_U3211) );
  OAI222_X1 U22704 ( .A1(n19838), .A2(n19786), .B1(n19785), .B2(n19835), .C1(
        n10419), .C2(n19834), .ZN(P2_U3212) );
  OAI222_X1 U22705 ( .A1(n19838), .A2(n13729), .B1(n19787), .B2(n19835), .C1(
        n19786), .C2(n19834), .ZN(P2_U3213) );
  INV_X1 U22706 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19789) );
  OAI222_X1 U22707 ( .A1(n19838), .A2(n19789), .B1(n19788), .B2(n19835), .C1(
        n13729), .C2(n19834), .ZN(P2_U3214) );
  OAI222_X1 U22708 ( .A1(n19838), .A2(n13863), .B1(n19790), .B2(n19835), .C1(
        n19789), .C2(n19834), .ZN(P2_U3215) );
  OAI222_X1 U22709 ( .A1(n19838), .A2(n19792), .B1(n19791), .B2(n19835), .C1(
        n13863), .C2(n19834), .ZN(P2_U3216) );
  OAI222_X1 U22710 ( .A1(n19838), .A2(n19794), .B1(n19793), .B2(n19835), .C1(
        n19792), .C2(n19834), .ZN(P2_U3217) );
  OAI222_X1 U22711 ( .A1(n19838), .A2(n19796), .B1(n19795), .B2(n19835), .C1(
        n19794), .C2(n19834), .ZN(P2_U3218) );
  OAI222_X1 U22712 ( .A1(n19838), .A2(n11280), .B1(n19797), .B2(n19835), .C1(
        n19796), .C2(n19834), .ZN(P2_U3219) );
  OAI222_X1 U22713 ( .A1(n19838), .A2(n19799), .B1(n19798), .B2(n19835), .C1(
        n11280), .C2(n19834), .ZN(P2_U3220) );
  OAI222_X1 U22714 ( .A1(n19838), .A2(n11310), .B1(n19800), .B2(n19835), .C1(
        n19799), .C2(n19834), .ZN(P2_U3221) );
  INV_X1 U22715 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19802) );
  OAI222_X1 U22716 ( .A1(n19838), .A2(n19802), .B1(n19801), .B2(n19835), .C1(
        n11310), .C2(n19834), .ZN(P2_U3222) );
  OAI222_X1 U22717 ( .A1(n19838), .A2(n11342), .B1(n19803), .B2(n19835), .C1(
        n19802), .C2(n19834), .ZN(P2_U3223) );
  OAI222_X1 U22718 ( .A1(n19838), .A2(n19805), .B1(n19804), .B2(n19835), .C1(
        n11342), .C2(n19834), .ZN(P2_U3224) );
  OAI222_X1 U22719 ( .A1(n19838), .A2(n15090), .B1(n19806), .B2(n19835), .C1(
        n19805), .C2(n19834), .ZN(P2_U3225) );
  OAI222_X1 U22720 ( .A1(n19838), .A2(n19808), .B1(n19807), .B2(n19835), .C1(
        n15090), .C2(n19834), .ZN(P2_U3226) );
  OAI222_X1 U22721 ( .A1(n19838), .A2(n19810), .B1(n19809), .B2(n19835), .C1(
        n19808), .C2(n19834), .ZN(P2_U3227) );
  OAI222_X1 U22722 ( .A1(n19838), .A2(n15070), .B1(n19811), .B2(n19835), .C1(
        n19810), .C2(n19834), .ZN(P2_U3228) );
  OAI222_X1 U22723 ( .A1(n19838), .A2(n19813), .B1(n19812), .B2(n19835), .C1(
        n15070), .C2(n19834), .ZN(P2_U3229) );
  OAI222_X1 U22724 ( .A1(n19838), .A2(n15043), .B1(n19814), .B2(n19835), .C1(
        n19813), .C2(n19834), .ZN(P2_U3230) );
  OAI222_X1 U22725 ( .A1(n19838), .A2(n19816), .B1(n19815), .B2(n19835), .C1(
        n15043), .C2(n19834), .ZN(P2_U3231) );
  OAI222_X1 U22726 ( .A1(n19838), .A2(n19818), .B1(n19817), .B2(n19835), .C1(
        n19816), .C2(n19834), .ZN(P2_U3232) );
  OAI222_X1 U22727 ( .A1(n19838), .A2(n19820), .B1(n19819), .B2(n19835), .C1(
        n19818), .C2(n19834), .ZN(P2_U3233) );
  INV_X1 U22728 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19822) );
  OAI222_X1 U22729 ( .A1(n19838), .A2(n19822), .B1(n19821), .B2(n19835), .C1(
        n19820), .C2(n19834), .ZN(P2_U3234) );
  OAI222_X1 U22730 ( .A1(n19838), .A2(n19824), .B1(n19823), .B2(n19835), .C1(
        n19822), .C2(n19834), .ZN(P2_U3235) );
  OAI222_X1 U22731 ( .A1(n19838), .A2(n19826), .B1(n19825), .B2(n19835), .C1(
        n19824), .C2(n19834), .ZN(P2_U3236) );
  OAI222_X1 U22732 ( .A1(n19838), .A2(n19829), .B1(n19827), .B2(n19835), .C1(
        n19826), .C2(n19834), .ZN(P2_U3237) );
  INV_X1 U22733 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19830) );
  OAI222_X1 U22734 ( .A1(n19834), .A2(n19829), .B1(n19828), .B2(n19835), .C1(
        n19830), .C2(n19838), .ZN(P2_U3238) );
  OAI222_X1 U22735 ( .A1(n19838), .A2(n19832), .B1(n19831), .B2(n19835), .C1(
        n19830), .C2(n19834), .ZN(P2_U3239) );
  OAI222_X1 U22736 ( .A1(n19838), .A2(n14235), .B1(n19833), .B2(n19835), .C1(
        n19832), .C2(n19834), .ZN(P2_U3240) );
  INV_X1 U22737 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19837) );
  OAI222_X1 U22738 ( .A1(n19838), .A2(n19837), .B1(n19836), .B2(n19835), .C1(
        n14235), .C2(n19834), .ZN(P2_U3241) );
  OAI22_X1 U22739 ( .A1(n19910), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19835), .ZN(n19839) );
  INV_X1 U22740 ( .A(n19839), .ZN(P2_U3585) );
  MUX2_X1 U22741 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19910), .Z(P2_U3586) );
  OAI22_X1 U22742 ( .A1(n19910), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19835), .ZN(n19840) );
  INV_X1 U22743 ( .A(n19840), .ZN(P2_U3587) );
  OAI22_X1 U22744 ( .A1(n19910), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19835), .ZN(n19841) );
  INV_X1 U22745 ( .A(n19841), .ZN(P2_U3588) );
  OAI21_X1 U22746 ( .B1(n19845), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19843), 
        .ZN(n19842) );
  INV_X1 U22747 ( .A(n19842), .ZN(P2_U3591) );
  OAI21_X1 U22748 ( .B1(n19845), .B2(n19844), .A(n19843), .ZN(P2_U3592) );
  INV_X1 U22749 ( .A(n19846), .ZN(n19847) );
  NOR2_X1 U22750 ( .A1(n19848), .A2(n19847), .ZN(n19849) );
  AOI21_X1 U22751 ( .B1(n19851), .B2(n19850), .A(n19849), .ZN(n19852) );
  OAI21_X1 U22752 ( .B1(n19854), .B2(n19853), .A(n19852), .ZN(n19856) );
  OAI22_X1 U22753 ( .A1(n19857), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n19856), .B2(n19855), .ZN(n19858) );
  INV_X1 U22754 ( .A(n19858), .ZN(P2_U3600) );
  INV_X1 U22755 ( .A(n19894), .ZN(n19897) );
  INV_X1 U22756 ( .A(n19859), .ZN(n19860) );
  NAND2_X1 U22757 ( .A1(n19860), .A2(n19876), .ZN(n19870) );
  NAND3_X1 U22758 ( .A1(n19883), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19861), 
        .ZN(n19862) );
  NAND2_X1 U22759 ( .A1(n19862), .A2(n19887), .ZN(n19871) );
  NAND2_X1 U22760 ( .A1(n19870), .A2(n19871), .ZN(n19867) );
  AOI222_X1 U22761 ( .A1(n19867), .A2(n19866), .B1(n19865), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n19864), .C2(n19863), .ZN(n19868) );
  AOI22_X1 U22762 ( .A1(n19897), .A2(n19869), .B1(n19868), .B2(n19894), .ZN(
        P2_U3602) );
  OAI21_X1 U22763 ( .B1(n19872), .B2(n19871), .A(n19870), .ZN(n19873) );
  AOI21_X1 U22764 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19874), .A(n19873), 
        .ZN(n19875) );
  AOI22_X1 U22765 ( .A1(n19897), .A2(n12599), .B1(n19875), .B2(n19894), .ZN(
        P2_U3603) );
  INV_X1 U22766 ( .A(n19876), .ZN(n19882) );
  INV_X1 U22767 ( .A(n19877), .ZN(n19878) );
  NAND3_X1 U22768 ( .A1(n19883), .A2(n19887), .A3(n19878), .ZN(n19881) );
  OR2_X1 U22769 ( .A1(n19879), .A2(n19888), .ZN(n19880) );
  OAI211_X1 U22770 ( .C1(n19883), .C2(n19882), .A(n19881), .B(n19880), .ZN(
        n19884) );
  INV_X1 U22771 ( .A(n19884), .ZN(n19885) );
  AOI22_X1 U22772 ( .A1(n19897), .A2(n19886), .B1(n19885), .B2(n19894), .ZN(
        P2_U3604) );
  INV_X1 U22773 ( .A(n19887), .ZN(n19889) );
  OAI22_X1 U22774 ( .A1(n19890), .A2(n19889), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19888), .ZN(n19891) );
  AOI21_X1 U22775 ( .B1(n19893), .B2(n19892), .A(n19891), .ZN(n19895) );
  AOI22_X1 U22776 ( .A1(n19897), .A2(n19896), .B1(n19895), .B2(n19894), .ZN(
        P2_U3605) );
  INV_X1 U22777 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19898) );
  AOI22_X1 U22778 ( .A1(n19835), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19898), 
        .B2(n19910), .ZN(P2_U3608) );
  INV_X1 U22779 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19909) );
  INV_X1 U22780 ( .A(n19899), .ZN(n19908) );
  INV_X1 U22781 ( .A(n19900), .ZN(n19902) );
  AOI22_X1 U22782 ( .A1(n19904), .A2(n19903), .B1(n19902), .B2(n19901), .ZN(
        n19907) );
  NOR2_X1 U22783 ( .A1(n19908), .A2(n19905), .ZN(n19906) );
  AOI22_X1 U22784 ( .A1(n19909), .A2(n19908), .B1(n19907), .B2(n19906), .ZN(
        P2_U3609) );
  MUX2_X1 U22785 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n19910), .Z(P2_U3611) );
  AOI21_X1 U22786 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20660), .A(n20657), 
        .ZN(n19918) );
  INV_X1 U22787 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19912) );
  NOR2_X2 U22788 ( .A1(n19911), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20732) );
  AOI21_X1 U22789 ( .B1(n19918), .B2(n19912), .A(n20732), .ZN(P1_U2802) );
  OAI21_X1 U22790 ( .B1(n19914), .B2(n19913), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19915) );
  OAI21_X1 U22791 ( .B1(n19916), .B2(n20644), .A(n19915), .ZN(P1_U2803) );
  INV_X2 U22792 ( .A(n20732), .ZN(n20745) );
  NOR2_X1 U22793 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19919) );
  OAI21_X1 U22794 ( .B1(n19919), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20745), .ZN(
        n19917) );
  OAI21_X1 U22795 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20745), .A(n19917), 
        .ZN(P1_U2804) );
  NOR2_X1 U22796 ( .A1(n20732), .A2(n19918), .ZN(n20707) );
  OAI21_X1 U22797 ( .B1(BS16), .B2(n19919), .A(n20707), .ZN(n20705) );
  OAI21_X1 U22798 ( .B1(n20707), .B2(n20535), .A(n20705), .ZN(P1_U2805) );
  OAI21_X1 U22799 ( .B1(n19922), .B2(n19921), .A(n19920), .ZN(P1_U2806) );
  NOR4_X1 U22800 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19926) );
  NOR4_X1 U22801 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19925) );
  NOR4_X1 U22802 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19924) );
  NOR4_X1 U22803 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19923) );
  NAND4_X1 U22804 ( .A1(n19926), .A2(n19925), .A3(n19924), .A4(n19923), .ZN(
        n19932) );
  NOR4_X1 U22805 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19930) );
  AOI211_X1 U22806 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_18__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19929) );
  NOR4_X1 U22807 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19928) );
  NOR4_X1 U22808 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19927) );
  NAND4_X1 U22809 ( .A1(n19930), .A2(n19929), .A3(n19928), .A4(n19927), .ZN(
        n19931) );
  NOR2_X1 U22810 ( .A1(n19932), .A2(n19931), .ZN(n20731) );
  INV_X1 U22811 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19934) );
  NOR3_X1 U22812 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19935) );
  OAI21_X1 U22813 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19935), .A(n20731), .ZN(
        n19933) );
  OAI21_X1 U22814 ( .B1(n20731), .B2(n19934), .A(n19933), .ZN(P1_U2807) );
  INV_X1 U22815 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20706) );
  AOI21_X1 U22816 ( .B1(n20724), .B2(n20706), .A(n19935), .ZN(n19937) );
  INV_X1 U22817 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19936) );
  INV_X1 U22818 ( .A(n20731), .ZN(n20726) );
  AOI22_X1 U22819 ( .A1(n20731), .A2(n19937), .B1(n19936), .B2(n20726), .ZN(
        P1_U2808) );
  OAI22_X1 U22820 ( .A1(n19939), .A2(n19985), .B1(n19984), .B2(n19938), .ZN(
        n19940) );
  AOI211_X1 U22821 ( .C1(n19977), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19955), .B(n19940), .ZN(n19949) );
  NAND2_X1 U22822 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19941) );
  NOR2_X1 U22823 ( .A1(n19941), .A2(n19975), .ZN(n19943) );
  AOI21_X1 U22824 ( .B1(n19941), .B2(n19993), .A(n19969), .ZN(n19962) );
  INV_X1 U22825 ( .A(n19962), .ZN(n19942) );
  MUX2_X1 U22826 ( .A(n19943), .B(n19942), .S(P1_REIP_REG_7__SCAN_IN), .Z(
        n19947) );
  NOR2_X1 U22827 ( .A1(n19945), .A2(n19944), .ZN(n19946) );
  NOR2_X1 U22828 ( .A1(n19947), .A2(n19946), .ZN(n19948) );
  OAI211_X1 U22829 ( .C1(n19950), .C2(n19995), .A(n19949), .B(n19948), .ZN(
        P1_U2833) );
  INV_X1 U22830 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19961) );
  AOI22_X1 U22831 ( .A1(n19994), .A2(n19951), .B1(n19997), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n19952) );
  OAI21_X1 U22832 ( .B1(n19953), .B2(n19995), .A(n19952), .ZN(n19954) );
  AOI211_X1 U22833 ( .C1(n19977), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19955), .B(n19954), .ZN(n19960) );
  NOR2_X1 U22834 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19975), .ZN(n19956) );
  AOI22_X1 U22835 ( .A1(n19958), .A2(n19957), .B1(n19956), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n19959) );
  OAI211_X1 U22836 ( .C1(n19962), .C2(n19961), .A(n19960), .B(n19959), .ZN(
        P1_U2834) );
  OAI21_X1 U22837 ( .B1(n19996), .B2(n19964), .A(n19963), .ZN(n19968) );
  OAI22_X1 U22838 ( .A1(n19966), .A2(n19985), .B1(n19984), .B2(n19965), .ZN(
        n19967) );
  AOI211_X1 U22839 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n19969), .A(n19968), .B(
        n19967), .ZN(n19974) );
  OAI22_X1 U22840 ( .A1(n19971), .A2(n20002), .B1(n19970), .B2(n19995), .ZN(
        n19972) );
  INV_X1 U22841 ( .A(n19972), .ZN(n19973) );
  OAI211_X1 U22842 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n19975), .A(n19974), .B(
        n19973), .ZN(P1_U2835) );
  AOI22_X1 U22843 ( .A1(n19977), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19976), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n19979) );
  OAI211_X1 U22844 ( .C1(n13545), .C2(n19980), .A(n19979), .B(n19978), .ZN(
        n19981) );
  INV_X1 U22845 ( .A(n19981), .ZN(n19991) );
  INV_X1 U22846 ( .A(n19982), .ZN(n19986) );
  OAI22_X1 U22847 ( .A1(n19986), .A2(n19985), .B1(n19984), .B2(n19983), .ZN(
        n19987) );
  AOI21_X1 U22848 ( .B1(n19989), .B2(n19988), .A(n19987), .ZN(n19990) );
  OAI211_X1 U22849 ( .C1(n20002), .C2(n19992), .A(n19991), .B(n19990), .ZN(
        P1_U2839) );
  AOI22_X1 U22850 ( .A1(n19994), .A2(n20088), .B1(P1_REIP_REG_0__SCAN_IN), 
        .B2(n19993), .ZN(n20001) );
  NAND2_X1 U22851 ( .A1(n19996), .A2(n19995), .ZN(n19999) );
  AOI222_X1 U22852 ( .A1(n19999), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19998), .B2(n11689), .C1(P1_EBX_REG_0__SCAN_IN), .C2(n19997), .ZN(
        n20000) );
  OAI211_X1 U22853 ( .C1(n20002), .C2(n20072), .A(n20001), .B(n20000), .ZN(
        P1_U2840) );
  AOI22_X1 U22854 ( .A1(n20005), .A2(n20004), .B1(n20003), .B2(n20073), .ZN(
        n20006) );
  OAI21_X1 U22855 ( .B1(n20008), .B2(n20007), .A(n20006), .ZN(P1_U2870) );
  OAI222_X1 U22856 ( .A1(n20735), .A2(n20012), .B1(n20033), .B2(n20011), .C1(
        n20010), .C2(n20009), .ZN(P1_U2921) );
  AOI22_X1 U22857 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20013) );
  OAI21_X1 U22858 ( .B1(n14050), .B2(n20033), .A(n20013), .ZN(P1_U2922) );
  INV_X1 U22859 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U22860 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20014) );
  OAI21_X1 U22861 ( .B1(n20015), .B2(n20033), .A(n20014), .ZN(P1_U2923) );
  AOI22_X1 U22862 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20016) );
  OAI21_X1 U22863 ( .B1(n14570), .B2(n20033), .A(n20016), .ZN(P1_U2924) );
  AOI22_X1 U22864 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20017) );
  OAI21_X1 U22865 ( .B1(n14054), .B2(n20033), .A(n20017), .ZN(P1_U2925) );
  AOI22_X1 U22866 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22867 ( .B1(n14033), .B2(n20033), .A(n20018), .ZN(P1_U2926) );
  AOI22_X1 U22868 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20019) );
  OAI21_X1 U22869 ( .B1(n13987), .B2(n20033), .A(n20019), .ZN(P1_U2927) );
  AOI22_X1 U22870 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20020) );
  OAI21_X1 U22871 ( .B1(n20021), .B2(n20033), .A(n20020), .ZN(P1_U2928) );
  AOI22_X1 U22872 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20022) );
  OAI21_X1 U22873 ( .B1(n11801), .B2(n20033), .A(n20022), .ZN(P1_U2929) );
  AOI22_X1 U22874 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20023) );
  OAI21_X1 U22875 ( .B1(n11788), .B2(n20033), .A(n20023), .ZN(P1_U2930) );
  AOI22_X1 U22876 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20024) );
  OAI21_X1 U22877 ( .B1(n11771), .B2(n20033), .A(n20024), .ZN(P1_U2931) );
  AOI22_X1 U22878 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20025) );
  OAI21_X1 U22879 ( .B1(n20026), .B2(n20033), .A(n20025), .ZN(P1_U2932) );
  AOI22_X1 U22880 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20027) );
  OAI21_X1 U22881 ( .B1(n11724), .B2(n20033), .A(n20027), .ZN(P1_U2933) );
  AOI22_X1 U22882 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20028) );
  OAI21_X1 U22883 ( .B1(n11676), .B2(n20033), .A(n20028), .ZN(P1_U2934) );
  AOI22_X1 U22884 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20029) );
  OAI21_X1 U22885 ( .B1(n11682), .B2(n20033), .A(n20029), .ZN(P1_U2935) );
  AOI22_X1 U22886 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20031), .B1(n20030), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U22887 ( .B1(n20034), .B2(n20033), .A(n20032), .ZN(P1_U2936) );
  AOI22_X1 U22888 ( .A1(n20061), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20060), .ZN(n20037) );
  INV_X1 U22889 ( .A(n20035), .ZN(n20036) );
  NAND2_X1 U22890 ( .A1(n20048), .A2(n20036), .ZN(n20050) );
  NAND2_X1 U22891 ( .A1(n20037), .A2(n20050), .ZN(P1_U2946) );
  AOI22_X1 U22892 ( .A1(n20061), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20040) );
  INV_X1 U22893 ( .A(n20038), .ZN(n20039) );
  NAND2_X1 U22894 ( .A1(n20048), .A2(n20039), .ZN(n20052) );
  NAND2_X1 U22895 ( .A1(n20040), .A2(n20052), .ZN(P1_U2947) );
  AOI22_X1 U22896 ( .A1(n20061), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20043) );
  INV_X1 U22897 ( .A(n20041), .ZN(n20042) );
  NAND2_X1 U22898 ( .A1(n20048), .A2(n20042), .ZN(n20054) );
  NAND2_X1 U22899 ( .A1(n20043), .A2(n20054), .ZN(P1_U2948) );
  AOI22_X1 U22900 ( .A1(n20061), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20046) );
  INV_X1 U22901 ( .A(n20044), .ZN(n20045) );
  NAND2_X1 U22902 ( .A1(n20048), .A2(n20045), .ZN(n20056) );
  NAND2_X1 U22903 ( .A1(n20046), .A2(n20056), .ZN(P1_U2949) );
  AOI22_X1 U22904 ( .A1(n20061), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20060), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20049) );
  NAND2_X1 U22905 ( .A1(n20048), .A2(n20047), .ZN(n20058) );
  NAND2_X1 U22906 ( .A1(n20049), .A2(n20058), .ZN(P1_U2950) );
  AOI22_X1 U22907 ( .A1(n20061), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20060), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20051) );
  NAND2_X1 U22908 ( .A1(n20051), .A2(n20050), .ZN(P1_U2961) );
  AOI22_X1 U22909 ( .A1(n20061), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20060), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20053) );
  NAND2_X1 U22910 ( .A1(n20053), .A2(n20052), .ZN(P1_U2962) );
  AOI22_X1 U22911 ( .A1(n20061), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20060), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20055) );
  NAND2_X1 U22912 ( .A1(n20055), .A2(n20054), .ZN(P1_U2963) );
  AOI22_X1 U22913 ( .A1(n20061), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20060), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U22914 ( .A1(n20057), .A2(n20056), .ZN(P1_U2964) );
  AOI22_X1 U22915 ( .A1(n20061), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20060), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20059) );
  NAND2_X1 U22916 ( .A1(n20059), .A2(n20058), .ZN(P1_U2965) );
  AOI22_X1 U22917 ( .A1(n20061), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20060), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20063) );
  NAND2_X1 U22918 ( .A1(n20063), .A2(n20062), .ZN(P1_U2966) );
  INV_X1 U22919 ( .A(n20064), .ZN(n20066) );
  AOI21_X1 U22920 ( .B1(n20066), .B2(n20094), .A(n20065), .ZN(n20091) );
  OR2_X1 U22921 ( .A1(n20068), .A2(n20067), .ZN(n20069) );
  AOI22_X1 U22922 ( .A1(n20091), .A2(n20070), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20069), .ZN(n20071) );
  NAND2_X1 U22923 ( .A1(n20074), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20099) );
  OAI211_X1 U22924 ( .C1(n20072), .C2(n20104), .A(n20071), .B(n20099), .ZN(
        P1_U2999) );
  AOI22_X1 U22925 ( .A1(n20074), .A2(P1_REIP_REG_2__SCAN_IN), .B1(n20089), 
        .B2(n20073), .ZN(n20087) );
  NOR2_X1 U22926 ( .A1(n20094), .A2(n12422), .ZN(n20076) );
  OAI221_X1 U22927 ( .B1(n20077), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n20077), .C2(n20076), .A(n20075), .ZN(n20086) );
  OAI21_X1 U22928 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20079), .A(
        n20078), .ZN(n20080) );
  AOI22_X1 U22929 ( .A1(n20081), .A2(n20090), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20080), .ZN(n20085) );
  NAND3_X1 U22930 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20083), .A3(
        n20082), .ZN(n20084) );
  NAND4_X1 U22931 ( .A1(n20087), .A2(n20086), .A3(n20085), .A4(n20084), .ZN(
        P1_U3029) );
  AOI22_X1 U22932 ( .A1(n20091), .A2(n20090), .B1(n20089), .B2(n20088), .ZN(
        n20100) );
  NAND3_X1 U22933 ( .A1(n20094), .A2(n20093), .A3(n20092), .ZN(n20095) );
  OAI21_X1 U22934 ( .B1(n20097), .B2(n20096), .A(n20095), .ZN(n20098) );
  NAND3_X1 U22935 ( .A1(n20100), .A2(n20099), .A3(n20098), .ZN(P1_U3031) );
  NOR2_X1 U22936 ( .A1(n20101), .A2(n20723), .ZN(P1_U3032) );
  NOR2_X2 U22937 ( .A1(n20102), .A2(n20104), .ZN(n20149) );
  AOI22_X1 U22938 ( .A1(DATAI_16_), .A2(n20149), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20105), .ZN(n20595) );
  INV_X1 U22939 ( .A(n9672), .ZN(n20106) );
  NOR2_X2 U22940 ( .A1(n20148), .A2(n20107), .ZN(n20583) );
  NOR3_X1 U22941 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20163) );
  NAND2_X1 U22942 ( .A1(n20504), .A2(n20163), .ZN(n20114) );
  INV_X1 U22943 ( .A(n20114), .ZN(n20151) );
  AOI22_X1 U22944 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20105), .B1(DATAI_24_), 
        .B2(n20149), .ZN(n20546) );
  INV_X1 U22945 ( .A(n20546), .ZN(n20592) );
  AOI22_X1 U22946 ( .A1(n20583), .A2(n20151), .B1(n20150), .B2(n20592), .ZN(
        n20123) );
  INV_X1 U22947 ( .A(n20183), .ZN(n20110) );
  OAI21_X1 U22948 ( .B1(n20110), .B2(n20150), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20111) );
  NAND2_X1 U22949 ( .A1(n20111), .A2(n20718), .ZN(n20121) );
  OR2_X1 U22950 ( .A1(n20711), .A2(n20112), .ZN(n20218) );
  NOR2_X1 U22951 ( .A1(n20218), .A2(n20538), .ZN(n20118) );
  INV_X1 U22952 ( .A(n20415), .ZN(n20113) );
  OR2_X1 U22953 ( .A1(n20113), .A2(n20361), .ZN(n20249) );
  AOI22_X1 U22954 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20249), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20114), .ZN(n20116) );
  NAND2_X1 U22955 ( .A1(n20119), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20532) );
  NAND2_X1 U22956 ( .A1(n20115), .A2(n20532), .ZN(n20187) );
  OAI211_X1 U22957 ( .C1(n20121), .C2(n20118), .A(n20116), .B(n20416), .ZN(
        n20154) );
  NOR2_X2 U22958 ( .A1(n20117), .A2(n20254), .ZN(n20582) );
  INV_X1 U22959 ( .A(n20118), .ZN(n20120) );
  NOR2_X1 U22960 ( .A1(n20119), .A2(n11673), .ZN(n20253) );
  INV_X1 U22961 ( .A(n20253), .ZN(n20420) );
  OAI22_X1 U22962 ( .A1(n20121), .A2(n20120), .B1(n20420), .B2(n20249), .ZN(
        n20153) );
  AOI22_X1 U22963 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20154), .B1(
        n20582), .B2(n20153), .ZN(n20122) );
  OAI211_X1 U22964 ( .C1(n20595), .C2(n20183), .A(n20123), .B(n20122), .ZN(
        P1_U3033) );
  AOI22_X1 U22965 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20105), .B1(DATAI_17_), 
        .B2(n20149), .ZN(n20601) );
  NOR2_X2 U22966 ( .A1(n20148), .A2(n20124), .ZN(n20597) );
  AOI22_X1 U22967 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20105), .B1(DATAI_25_), 
        .B2(n20149), .ZN(n20550) );
  INV_X1 U22968 ( .A(n20550), .ZN(n20598) );
  AOI22_X1 U22969 ( .A1(n20597), .A2(n20151), .B1(n20150), .B2(n20598), .ZN(
        n20127) );
  NOR2_X2 U22970 ( .A1(n20125), .A2(n20254), .ZN(n20596) );
  AOI22_X1 U22971 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20154), .B1(
        n20596), .B2(n20153), .ZN(n20126) );
  OAI211_X1 U22972 ( .C1(n20601), .C2(n20183), .A(n20127), .B(n20126), .ZN(
        P1_U3034) );
  AOI22_X1 U22973 ( .A1(DATAI_18_), .A2(n20149), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20105), .ZN(n20607) );
  NOR2_X2 U22974 ( .A1(n20148), .A2(n13249), .ZN(n20603) );
  AOI22_X1 U22975 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20105), .B1(DATAI_26_), 
        .B2(n20149), .ZN(n20554) );
  INV_X1 U22976 ( .A(n20554), .ZN(n20604) );
  AOI22_X1 U22977 ( .A1(n20603), .A2(n20151), .B1(n20150), .B2(n20604), .ZN(
        n20130) );
  NOR2_X2 U22978 ( .A1(n20128), .A2(n20254), .ZN(n20602) );
  AOI22_X1 U22979 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20154), .B1(
        n20602), .B2(n20153), .ZN(n20129) );
  OAI211_X1 U22980 ( .C1(n20607), .C2(n20183), .A(n20130), .B(n20129), .ZN(
        P1_U3035) );
  AOI22_X1 U22981 ( .A1(DATAI_19_), .A2(n20149), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20105), .ZN(n20613) );
  NOR2_X2 U22982 ( .A1(n20148), .A2(n20131), .ZN(n20609) );
  AOI22_X1 U22983 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20105), .B1(DATAI_27_), 
        .B2(n20149), .ZN(n20558) );
  INV_X1 U22984 ( .A(n20558), .ZN(n20610) );
  AOI22_X1 U22985 ( .A1(n20609), .A2(n20151), .B1(n20150), .B2(n20610), .ZN(
        n20134) );
  NOR2_X2 U22986 ( .A1(n20132), .A2(n20254), .ZN(n20608) );
  AOI22_X1 U22987 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20154), .B1(
        n20608), .B2(n20153), .ZN(n20133) );
  OAI211_X1 U22988 ( .C1(n20613), .C2(n20183), .A(n20134), .B(n20133), .ZN(
        P1_U3036) );
  AOI22_X1 U22989 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20105), .B1(DATAI_20_), 
        .B2(n20149), .ZN(n20619) );
  NOR2_X2 U22990 ( .A1(n20148), .A2(n20135), .ZN(n20615) );
  AOI22_X1 U22991 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20105), .B1(DATAI_28_), 
        .B2(n20149), .ZN(n20562) );
  INV_X1 U22992 ( .A(n20562), .ZN(n20616) );
  AOI22_X1 U22993 ( .A1(n20615), .A2(n20151), .B1(n20150), .B2(n20616), .ZN(
        n20138) );
  NOR2_X2 U22994 ( .A1(n20136), .A2(n20254), .ZN(n20614) );
  AOI22_X1 U22995 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20154), .B1(
        n20614), .B2(n20153), .ZN(n20137) );
  OAI211_X1 U22996 ( .C1(n20619), .C2(n20183), .A(n20138), .B(n20137), .ZN(
        P1_U3037) );
  AOI22_X1 U22997 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20105), .B1(DATAI_21_), 
        .B2(n20149), .ZN(n20625) );
  NOR2_X2 U22998 ( .A1(n20148), .A2(n20139), .ZN(n20621) );
  AOI22_X1 U22999 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20105), .B1(DATAI_29_), 
        .B2(n20149), .ZN(n20566) );
  INV_X1 U23000 ( .A(n20566), .ZN(n20622) );
  AOI22_X1 U23001 ( .A1(n20621), .A2(n20151), .B1(n20150), .B2(n20622), .ZN(
        n20142) );
  NOR2_X2 U23002 ( .A1(n20140), .A2(n20254), .ZN(n20620) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20154), .B1(
        n20620), .B2(n20153), .ZN(n20141) );
  OAI211_X1 U23004 ( .C1(n20625), .C2(n20183), .A(n20142), .B(n20141), .ZN(
        P1_U3038) );
  AOI22_X1 U23005 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20105), .B1(DATAI_22_), 
        .B2(n20149), .ZN(n20631) );
  NOR2_X2 U23006 ( .A1(n20148), .A2(n20143), .ZN(n20627) );
  AOI22_X1 U23007 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20105), .B1(DATAI_30_), 
        .B2(n20149), .ZN(n20570) );
  INV_X1 U23008 ( .A(n20570), .ZN(n20628) );
  AOI22_X1 U23009 ( .A1(n20627), .A2(n20151), .B1(n20150), .B2(n20628), .ZN(
        n20146) );
  NOR2_X2 U23010 ( .A1(n20144), .A2(n20254), .ZN(n20626) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20154), .B1(
        n20626), .B2(n20153), .ZN(n20145) );
  OAI211_X1 U23012 ( .C1(n20631), .C2(n20183), .A(n20146), .B(n20145), .ZN(
        P1_U3039) );
  AOI22_X1 U23013 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20105), .B1(DATAI_23_), 
        .B2(n20149), .ZN(n20642) );
  NOR2_X2 U23014 ( .A1(n20148), .A2(n20147), .ZN(n20635) );
  AOI22_X1 U23015 ( .A1(DATAI_31_), .A2(n20149), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20105), .ZN(n20578) );
  INV_X1 U23016 ( .A(n20578), .ZN(n20636) );
  AOI22_X1 U23017 ( .A1(n20635), .A2(n20151), .B1(n20150), .B2(n20636), .ZN(
        n20156) );
  NOR2_X2 U23018 ( .A1(n20152), .A2(n20254), .ZN(n20633) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20154), .B1(
        n20633), .B2(n20153), .ZN(n20155) );
  OAI211_X1 U23020 ( .C1(n20642), .C2(n20183), .A(n20156), .B(n20155), .ZN(
        P1_U3040) );
  INV_X1 U23021 ( .A(n20163), .ZN(n20160) );
  NOR2_X1 U23022 ( .A1(n20504), .A2(n20160), .ZN(n20179) );
  OR2_X1 U23023 ( .A1(n20218), .A2(n20157), .ZN(n20159) );
  INV_X1 U23024 ( .A(n20179), .ZN(n20158) );
  OAI22_X1 U23025 ( .A1(n20161), .A2(n20590), .B1(n20160), .B2(n11673), .ZN(
        n20178) );
  AOI22_X1 U23026 ( .A1(n20583), .A2(n20179), .B1(n20582), .B2(n20178), .ZN(
        n20165) );
  INV_X1 U23027 ( .A(n20214), .ZN(n20215) );
  OR2_X1 U23028 ( .A1(n20185), .A2(n20535), .ZN(n20508) );
  OAI21_X1 U23029 ( .B1(n20215), .B2(n20508), .A(n20161), .ZN(n20162) );
  OAI221_X1 U23030 ( .B1(n20718), .B2(n20163), .C1(n20590), .C2(n20162), .A(
        n20588), .ZN(n20180) );
  NAND2_X1 U23031 ( .A1(n20214), .A2(n9734), .ZN(n20195) );
  INV_X1 U23032 ( .A(n20595), .ZN(n20543) );
  AOI22_X1 U23033 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20543), .ZN(n20164) );
  OAI211_X1 U23034 ( .C1(n20546), .C2(n20183), .A(n20165), .B(n20164), .ZN(
        P1_U3041) );
  AOI22_X1 U23035 ( .A1(n20597), .A2(n20179), .B1(n20596), .B2(n20178), .ZN(
        n20167) );
  INV_X1 U23036 ( .A(n20601), .ZN(n20547) );
  AOI22_X1 U23037 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20547), .ZN(n20166) );
  OAI211_X1 U23038 ( .C1(n20550), .C2(n20183), .A(n20167), .B(n20166), .ZN(
        P1_U3042) );
  AOI22_X1 U23039 ( .A1(n20603), .A2(n20179), .B1(n20602), .B2(n20178), .ZN(
        n20169) );
  INV_X1 U23040 ( .A(n20607), .ZN(n20551) );
  AOI22_X1 U23041 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20551), .ZN(n20168) );
  OAI211_X1 U23042 ( .C1(n20554), .C2(n20183), .A(n20169), .B(n20168), .ZN(
        P1_U3043) );
  AOI22_X1 U23043 ( .A1(n20609), .A2(n20179), .B1(n20608), .B2(n20178), .ZN(
        n20171) );
  INV_X1 U23044 ( .A(n20613), .ZN(n20555) );
  AOI22_X1 U23045 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20555), .ZN(n20170) );
  OAI211_X1 U23046 ( .C1(n20558), .C2(n20183), .A(n20171), .B(n20170), .ZN(
        P1_U3044) );
  AOI22_X1 U23047 ( .A1(n20615), .A2(n20179), .B1(n20614), .B2(n20178), .ZN(
        n20173) );
  INV_X1 U23048 ( .A(n20619), .ZN(n20559) );
  AOI22_X1 U23049 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20559), .ZN(n20172) );
  OAI211_X1 U23050 ( .C1(n20562), .C2(n20183), .A(n20173), .B(n20172), .ZN(
        P1_U3045) );
  AOI22_X1 U23051 ( .A1(n20621), .A2(n20179), .B1(n20620), .B2(n20178), .ZN(
        n20175) );
  INV_X1 U23052 ( .A(n20625), .ZN(n20563) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20563), .ZN(n20174) );
  OAI211_X1 U23054 ( .C1(n20566), .C2(n20183), .A(n20175), .B(n20174), .ZN(
        P1_U3046) );
  AOI22_X1 U23055 ( .A1(n20627), .A2(n20179), .B1(n20626), .B2(n20178), .ZN(
        n20177) );
  INV_X1 U23056 ( .A(n20631), .ZN(n20567) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20567), .ZN(n20176) );
  OAI211_X1 U23058 ( .C1(n20570), .C2(n20183), .A(n20177), .B(n20176), .ZN(
        P1_U3047) );
  AOI22_X1 U23059 ( .A1(n20635), .A2(n20179), .B1(n20633), .B2(n20178), .ZN(
        n20182) );
  INV_X1 U23060 ( .A(n20642), .ZN(n20573) );
  AOI22_X1 U23061 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20180), .B1(
        n20208), .B2(n20573), .ZN(n20181) );
  OAI211_X1 U23062 ( .C1(n20578), .C2(n20183), .A(n20182), .B(n20181), .ZN(
        P1_U3048) );
  NAND3_X1 U23063 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20722), .A3(
        n20474), .ZN(n20223) );
  NOR2_X1 U23064 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20223), .ZN(
        n20209) );
  INV_X1 U23065 ( .A(n20246), .ZN(n20238) );
  AOI22_X1 U23066 ( .A1(n20583), .A2(n20209), .B1(n20238), .B2(n20543), .ZN(
        n20194) );
  OAI21_X1 U23067 ( .B1(n20238), .B2(n20208), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20186) );
  NAND2_X1 U23068 ( .A1(n20186), .A2(n20718), .ZN(n20192) );
  NOR2_X1 U23069 ( .A1(n20218), .A2(n13545), .ZN(n20190) );
  INV_X1 U23070 ( .A(n20209), .ZN(n20188) );
  OR2_X1 U23071 ( .A1(n20415), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20307) );
  AND2_X1 U23072 ( .A1(n20307), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20304) );
  AOI211_X1 U23073 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20188), .A(n20304), 
        .B(n20187), .ZN(n20189) );
  INV_X1 U23074 ( .A(n20190), .ZN(n20191) );
  OAI22_X1 U23075 ( .A1(n20192), .A2(n20191), .B1(n20307), .B2(n20420), .ZN(
        n20210) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20211), .B1(
        n20582), .B2(n20210), .ZN(n20193) );
  OAI211_X1 U23077 ( .C1(n20546), .C2(n20195), .A(n20194), .B(n20193), .ZN(
        P1_U3049) );
  AOI22_X1 U23078 ( .A1(n20597), .A2(n20209), .B1(n20208), .B2(n20598), .ZN(
        n20197) );
  AOI22_X1 U23079 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20211), .B1(
        n20596), .B2(n20210), .ZN(n20196) );
  OAI211_X1 U23080 ( .C1(n20601), .C2(n20246), .A(n20197), .B(n20196), .ZN(
        P1_U3050) );
  AOI22_X1 U23081 ( .A1(n20603), .A2(n20209), .B1(n20208), .B2(n20604), .ZN(
        n20199) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20211), .B1(
        n20602), .B2(n20210), .ZN(n20198) );
  OAI211_X1 U23083 ( .C1(n20607), .C2(n20246), .A(n20199), .B(n20198), .ZN(
        P1_U3051) );
  AOI22_X1 U23084 ( .A1(n20609), .A2(n20209), .B1(n20208), .B2(n20610), .ZN(
        n20201) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20211), .B1(
        n20608), .B2(n20210), .ZN(n20200) );
  OAI211_X1 U23086 ( .C1(n20613), .C2(n20246), .A(n20201), .B(n20200), .ZN(
        P1_U3052) );
  AOI22_X1 U23087 ( .A1(n20615), .A2(n20209), .B1(n20208), .B2(n20616), .ZN(
        n20203) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20211), .B1(
        n20614), .B2(n20210), .ZN(n20202) );
  OAI211_X1 U23089 ( .C1(n20619), .C2(n20246), .A(n20203), .B(n20202), .ZN(
        P1_U3053) );
  AOI22_X1 U23090 ( .A1(n20621), .A2(n20209), .B1(n20208), .B2(n20622), .ZN(
        n20205) );
  AOI22_X1 U23091 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20211), .B1(
        n20620), .B2(n20210), .ZN(n20204) );
  OAI211_X1 U23092 ( .C1(n20625), .C2(n20246), .A(n20205), .B(n20204), .ZN(
        P1_U3054) );
  AOI22_X1 U23093 ( .A1(n20627), .A2(n20209), .B1(n20208), .B2(n20628), .ZN(
        n20207) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20211), .B1(
        n20626), .B2(n20210), .ZN(n20206) );
  OAI211_X1 U23095 ( .C1(n20631), .C2(n20246), .A(n20207), .B(n20206), .ZN(
        P1_U3055) );
  AOI22_X1 U23096 ( .A1(n20635), .A2(n20209), .B1(n20208), .B2(n20636), .ZN(
        n20213) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20211), .B1(
        n20633), .B2(n20210), .ZN(n20212) );
  OAI211_X1 U23098 ( .C1(n20642), .C2(n20246), .A(n20213), .B(n20212), .ZN(
        P1_U3056) );
  NOR2_X1 U23099 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20446), .ZN(
        n20241) );
  AOI22_X1 U23100 ( .A1(n20583), .A2(n20241), .B1(n20273), .B2(n20543), .ZN(
        n20227) );
  OAI21_X1 U23101 ( .B1(n20215), .B2(n20586), .A(n20718), .ZN(n20224) );
  AND2_X1 U23102 ( .A1(n20216), .A2(n11689), .ZN(n20579) );
  INV_X1 U23103 ( .A(n20579), .ZN(n20217) );
  OR2_X1 U23104 ( .A1(n20218), .A2(n20217), .ZN(n20220) );
  INV_X1 U23105 ( .A(n20241), .ZN(n20219) );
  AND2_X1 U23106 ( .A1(n20220), .A2(n20219), .ZN(n20225) );
  INV_X1 U23107 ( .A(n20225), .ZN(n20222) );
  INV_X1 U23108 ( .A(n20588), .ZN(n20333) );
  AOI21_X1 U23109 ( .B1(n20590), .B2(n20223), .A(n20333), .ZN(n20221) );
  OAI21_X1 U23110 ( .B1(n20224), .B2(n20222), .A(n20221), .ZN(n20243) );
  OAI22_X1 U23111 ( .A1(n20225), .A2(n20224), .B1(n11673), .B2(n20223), .ZN(
        n20242) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20243), .B1(
        n20582), .B2(n20242), .ZN(n20226) );
  OAI211_X1 U23113 ( .C1(n20546), .C2(n20246), .A(n20227), .B(n20226), .ZN(
        P1_U3057) );
  AOI22_X1 U23114 ( .A1(n20597), .A2(n20241), .B1(n20273), .B2(n20547), .ZN(
        n20229) );
  AOI22_X1 U23115 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20243), .B1(
        n20596), .B2(n20242), .ZN(n20228) );
  OAI211_X1 U23116 ( .C1(n20550), .C2(n20246), .A(n20229), .B(n20228), .ZN(
        P1_U3058) );
  AOI22_X1 U23117 ( .A1(n20603), .A2(n20241), .B1(n20273), .B2(n20551), .ZN(
        n20231) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20243), .B1(
        n20602), .B2(n20242), .ZN(n20230) );
  OAI211_X1 U23119 ( .C1(n20554), .C2(n20246), .A(n20231), .B(n20230), .ZN(
        P1_U3059) );
  AOI22_X1 U23120 ( .A1(n20609), .A2(n20241), .B1(n20273), .B2(n20555), .ZN(
        n20233) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20243), .B1(
        n20608), .B2(n20242), .ZN(n20232) );
  OAI211_X1 U23122 ( .C1(n20558), .C2(n20246), .A(n20233), .B(n20232), .ZN(
        P1_U3060) );
  AOI22_X1 U23123 ( .A1(n20615), .A2(n20241), .B1(n20273), .B2(n20559), .ZN(
        n20235) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20243), .B1(
        n20614), .B2(n20242), .ZN(n20234) );
  OAI211_X1 U23125 ( .C1(n20562), .C2(n20246), .A(n20235), .B(n20234), .ZN(
        P1_U3061) );
  AOI22_X1 U23126 ( .A1(n20621), .A2(n20241), .B1(n20273), .B2(n20563), .ZN(
        n20237) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20243), .B1(
        n20620), .B2(n20242), .ZN(n20236) );
  OAI211_X1 U23128 ( .C1(n20566), .C2(n20246), .A(n20237), .B(n20236), .ZN(
        P1_U3062) );
  INV_X1 U23129 ( .A(n20273), .ZN(n20258) );
  AOI22_X1 U23130 ( .A1(n20627), .A2(n20241), .B1(n20238), .B2(n20628), .ZN(
        n20240) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20243), .B1(
        n20626), .B2(n20242), .ZN(n20239) );
  OAI211_X1 U23132 ( .C1(n20631), .C2(n20258), .A(n20240), .B(n20239), .ZN(
        P1_U3063) );
  AOI22_X1 U23133 ( .A1(n20635), .A2(n20241), .B1(n20273), .B2(n20573), .ZN(
        n20245) );
  AOI22_X1 U23134 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20243), .B1(
        n20633), .B2(n20242), .ZN(n20244) );
  OAI211_X1 U23135 ( .C1(n20578), .C2(n20246), .A(n20245), .B(n20244), .ZN(
        P1_U3064) );
  NOR3_X1 U23136 ( .A1(n20474), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20281) );
  INV_X1 U23137 ( .A(n20281), .ZN(n20277) );
  NOR2_X1 U23138 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20277), .ZN(
        n20272) );
  NOR2_X1 U23139 ( .A1(n13515), .A2(n20247), .ZN(n20332) );
  NAND3_X1 U23140 ( .A1(n20332), .A2(n20718), .A3(n13545), .ZN(n20248) );
  OAI21_X1 U23141 ( .B1(n20249), .B2(n20532), .A(n20248), .ZN(n20271) );
  AOI22_X1 U23142 ( .A1(n20583), .A2(n20272), .B1(n20582), .B2(n20271), .ZN(
        n20257) );
  AOI21_X1 U23143 ( .B1(n20258), .B2(n20296), .A(n20535), .ZN(n20251) );
  AOI21_X1 U23144 ( .B1(n20332), .B2(n13545), .A(n20251), .ZN(n20252) );
  NOR2_X1 U23145 ( .A1(n20252), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20255) );
  INV_X1 U23146 ( .A(n20296), .ZN(n20299) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20274), .B1(
        n20299), .B2(n20543), .ZN(n20256) );
  OAI211_X1 U23148 ( .C1(n20546), .C2(n20258), .A(n20257), .B(n20256), .ZN(
        P1_U3065) );
  AOI22_X1 U23149 ( .A1(n20597), .A2(n20272), .B1(n20596), .B2(n20271), .ZN(
        n20260) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20598), .ZN(n20259) );
  OAI211_X1 U23151 ( .C1(n20601), .C2(n20296), .A(n20260), .B(n20259), .ZN(
        P1_U3066) );
  AOI22_X1 U23152 ( .A1(n20603), .A2(n20272), .B1(n20602), .B2(n20271), .ZN(
        n20262) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20604), .ZN(n20261) );
  OAI211_X1 U23154 ( .C1(n20607), .C2(n20296), .A(n20262), .B(n20261), .ZN(
        P1_U3067) );
  AOI22_X1 U23155 ( .A1(n20609), .A2(n20272), .B1(n20608), .B2(n20271), .ZN(
        n20264) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20610), .ZN(n20263) );
  OAI211_X1 U23157 ( .C1(n20613), .C2(n20296), .A(n20264), .B(n20263), .ZN(
        P1_U3068) );
  AOI22_X1 U23158 ( .A1(n20615), .A2(n20272), .B1(n20614), .B2(n20271), .ZN(
        n20266) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20616), .ZN(n20265) );
  OAI211_X1 U23160 ( .C1(n20619), .C2(n20296), .A(n20266), .B(n20265), .ZN(
        P1_U3069) );
  AOI22_X1 U23161 ( .A1(n20621), .A2(n20272), .B1(n20620), .B2(n20271), .ZN(
        n20268) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20622), .ZN(n20267) );
  OAI211_X1 U23163 ( .C1(n20625), .C2(n20296), .A(n20268), .B(n20267), .ZN(
        P1_U3070) );
  AOI22_X1 U23164 ( .A1(n20627), .A2(n20272), .B1(n20626), .B2(n20271), .ZN(
        n20270) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20628), .ZN(n20269) );
  OAI211_X1 U23166 ( .C1(n20631), .C2(n20296), .A(n20270), .B(n20269), .ZN(
        P1_U3071) );
  AOI22_X1 U23167 ( .A1(n20635), .A2(n20272), .B1(n20633), .B2(n20271), .ZN(
        n20276) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20274), .B1(
        n20273), .B2(n20636), .ZN(n20275) );
  OAI211_X1 U23169 ( .C1(n20642), .C2(n20296), .A(n20276), .B(n20275), .ZN(
        P1_U3072) );
  NOR2_X1 U23170 ( .A1(n20504), .A2(n20277), .ZN(n20298) );
  INV_X1 U23171 ( .A(n20157), .ZN(n20505) );
  AOI21_X1 U23172 ( .B1(n20332), .B2(n20505), .A(n20298), .ZN(n20278) );
  OAI22_X1 U23173 ( .A1(n20278), .A2(n20590), .B1(n20277), .B2(n11673), .ZN(
        n20297) );
  AOI22_X1 U23174 ( .A1(n20583), .A2(n20298), .B1(n20582), .B2(n20297), .ZN(
        n20283) );
  INV_X1 U23175 ( .A(n20337), .ZN(n20279) );
  OAI21_X1 U23176 ( .B1(n20279), .B2(n20508), .A(n20278), .ZN(n20280) );
  OAI221_X1 U23177 ( .B1(n20718), .B2(n20281), .C1(n20590), .C2(n20280), .A(
        n20588), .ZN(n20300) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20592), .ZN(n20282) );
  OAI211_X1 U23179 ( .C1(n20595), .C2(n20324), .A(n20283), .B(n20282), .ZN(
        P1_U3073) );
  AOI22_X1 U23180 ( .A1(n20597), .A2(n20298), .B1(n20596), .B2(n20297), .ZN(
        n20285) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20300), .B1(
        n20325), .B2(n20547), .ZN(n20284) );
  OAI211_X1 U23182 ( .C1(n20550), .C2(n20296), .A(n20285), .B(n20284), .ZN(
        P1_U3074) );
  AOI22_X1 U23183 ( .A1(n20603), .A2(n20298), .B1(n20602), .B2(n20297), .ZN(
        n20287) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20604), .ZN(n20286) );
  OAI211_X1 U23185 ( .C1(n20607), .C2(n20324), .A(n20287), .B(n20286), .ZN(
        P1_U3075) );
  AOI22_X1 U23186 ( .A1(n20609), .A2(n20298), .B1(n20608), .B2(n20297), .ZN(
        n20289) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20300), .B1(
        n20325), .B2(n20555), .ZN(n20288) );
  OAI211_X1 U23188 ( .C1(n20558), .C2(n20296), .A(n20289), .B(n20288), .ZN(
        P1_U3076) );
  AOI22_X1 U23189 ( .A1(n20615), .A2(n20298), .B1(n20614), .B2(n20297), .ZN(
        n20291) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20300), .B1(
        n20325), .B2(n20559), .ZN(n20290) );
  OAI211_X1 U23191 ( .C1(n20562), .C2(n20296), .A(n20291), .B(n20290), .ZN(
        P1_U3077) );
  AOI22_X1 U23192 ( .A1(n20621), .A2(n20298), .B1(n20620), .B2(n20297), .ZN(
        n20293) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20300), .B1(
        n20325), .B2(n20563), .ZN(n20292) );
  OAI211_X1 U23194 ( .C1(n20566), .C2(n20296), .A(n20293), .B(n20292), .ZN(
        P1_U3078) );
  AOI22_X1 U23195 ( .A1(n20627), .A2(n20298), .B1(n20626), .B2(n20297), .ZN(
        n20295) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20300), .B1(
        n20325), .B2(n20567), .ZN(n20294) );
  OAI211_X1 U23197 ( .C1(n20570), .C2(n20296), .A(n20295), .B(n20294), .ZN(
        P1_U3079) );
  AOI22_X1 U23198 ( .A1(n20635), .A2(n20298), .B1(n20633), .B2(n20297), .ZN(
        n20302) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20636), .ZN(n20301) );
  OAI211_X1 U23200 ( .C1(n20642), .C2(n20324), .A(n20302), .B(n20301), .ZN(
        P1_U3080) );
  NOR2_X1 U23201 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20335), .ZN(
        n20326) );
  AOI22_X1 U23202 ( .A1(n20583), .A2(n20326), .B1(n20349), .B2(n20543), .ZN(
        n20311) );
  OR2_X1 U23203 ( .A1(n20349), .A2(n20325), .ZN(n20303) );
  AOI21_X1 U23204 ( .B1(n20303), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20590), 
        .ZN(n20306) );
  NAND2_X1 U23205 ( .A1(n20332), .A2(n20538), .ZN(n20308) );
  AOI21_X1 U23206 ( .B1(n20306), .B2(n20308), .A(n20304), .ZN(n20305) );
  OAI211_X1 U23207 ( .C1(n20326), .C2(n20479), .A(n20541), .B(n20305), .ZN(
        n20328) );
  INV_X1 U23208 ( .A(n20306), .ZN(n20309) );
  OAI22_X1 U23209 ( .A1(n20309), .A2(n20308), .B1(n20532), .B2(n20307), .ZN(
        n20327) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20328), .B1(
        n20582), .B2(n20327), .ZN(n20310) );
  OAI211_X1 U23211 ( .C1(n20546), .C2(n20324), .A(n20311), .B(n20310), .ZN(
        P1_U3081) );
  AOI22_X1 U23212 ( .A1(n20597), .A2(n20326), .B1(n20349), .B2(n20547), .ZN(
        n20313) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20328), .B1(
        n20596), .B2(n20327), .ZN(n20312) );
  OAI211_X1 U23214 ( .C1(n20550), .C2(n20324), .A(n20313), .B(n20312), .ZN(
        P1_U3082) );
  AOI22_X1 U23215 ( .A1(n20603), .A2(n20326), .B1(n20349), .B2(n20551), .ZN(
        n20315) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20328), .B1(
        n20602), .B2(n20327), .ZN(n20314) );
  OAI211_X1 U23217 ( .C1(n20554), .C2(n20324), .A(n20315), .B(n20314), .ZN(
        P1_U3083) );
  AOI22_X1 U23218 ( .A1(n20609), .A2(n20326), .B1(n20349), .B2(n20555), .ZN(
        n20317) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20328), .B1(
        n20608), .B2(n20327), .ZN(n20316) );
  OAI211_X1 U23220 ( .C1(n20558), .C2(n20324), .A(n20317), .B(n20316), .ZN(
        P1_U3084) );
  AOI22_X1 U23221 ( .A1(n20615), .A2(n20326), .B1(n20349), .B2(n20559), .ZN(
        n20319) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20328), .B1(
        n20614), .B2(n20327), .ZN(n20318) );
  OAI211_X1 U23223 ( .C1(n20562), .C2(n20324), .A(n20319), .B(n20318), .ZN(
        P1_U3085) );
  AOI22_X1 U23224 ( .A1(n20621), .A2(n20326), .B1(n20325), .B2(n20622), .ZN(
        n20321) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20328), .B1(
        n20620), .B2(n20327), .ZN(n20320) );
  OAI211_X1 U23226 ( .C1(n20625), .C2(n20360), .A(n20321), .B(n20320), .ZN(
        P1_U3086) );
  AOI22_X1 U23227 ( .A1(n20627), .A2(n20326), .B1(n20349), .B2(n20567), .ZN(
        n20323) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20328), .B1(
        n20626), .B2(n20327), .ZN(n20322) );
  OAI211_X1 U23229 ( .C1(n20570), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        P1_U3087) );
  AOI22_X1 U23230 ( .A1(n20635), .A2(n20326), .B1(n20325), .B2(n20636), .ZN(
        n20330) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20328), .B1(
        n20633), .B2(n20327), .ZN(n20329) );
  OAI211_X1 U23232 ( .C1(n20642), .C2(n20360), .A(n20330), .B(n20329), .ZN(
        P1_U3088) );
  INV_X1 U23233 ( .A(n20586), .ZN(n20331) );
  NAND2_X1 U23234 ( .A1(n20337), .A2(n20331), .ZN(n20709) );
  AOI21_X1 U23235 ( .B1(n20332), .B2(n20579), .A(n20356), .ZN(n20336) );
  AND2_X1 U23236 ( .A1(n20709), .A2(n20336), .ZN(n20334) );
  AOI221_X1 U23237 ( .B1(n20334), .B2(n20718), .C1(n20335), .C2(n20590), .A(
        n20333), .ZN(n20340) );
  INV_X1 U23238 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n20872) );
  OAI22_X1 U23239 ( .A1(n20336), .A2(n20590), .B1(n20335), .B2(n11673), .ZN(
        n20355) );
  AOI22_X1 U23240 ( .A1(n20583), .A2(n20356), .B1(n20582), .B2(n20355), .ZN(
        n20339) );
  NAND2_X1 U23241 ( .A1(n20337), .A2(n20444), .ZN(n20352) );
  AOI22_X1 U23242 ( .A1(n20382), .A2(n20543), .B1(n20349), .B2(n20592), .ZN(
        n20338) );
  OAI211_X1 U23243 ( .C1(n20340), .C2(n20872), .A(n20339), .B(n20338), .ZN(
        P1_U3089) );
  AOI22_X1 U23244 ( .A1(n20597), .A2(n20356), .B1(n20596), .B2(n20355), .ZN(
        n20342) );
  INV_X1 U23245 ( .A(n20340), .ZN(n20357) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20357), .B1(
        n20349), .B2(n20598), .ZN(n20341) );
  OAI211_X1 U23247 ( .C1(n20601), .C2(n20352), .A(n20342), .B(n20341), .ZN(
        P1_U3090) );
  AOI22_X1 U23248 ( .A1(n20603), .A2(n20356), .B1(n20602), .B2(n20355), .ZN(
        n20344) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20357), .B1(
        n20349), .B2(n20604), .ZN(n20343) );
  OAI211_X1 U23250 ( .C1(n20607), .C2(n20352), .A(n20344), .B(n20343), .ZN(
        P1_U3091) );
  AOI22_X1 U23251 ( .A1(n20609), .A2(n20356), .B1(n20608), .B2(n20355), .ZN(
        n20346) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20357), .B1(
        n20382), .B2(n20555), .ZN(n20345) );
  OAI211_X1 U23253 ( .C1(n20558), .C2(n20360), .A(n20346), .B(n20345), .ZN(
        P1_U3092) );
  AOI22_X1 U23254 ( .A1(n20615), .A2(n20356), .B1(n20614), .B2(n20355), .ZN(
        n20348) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20357), .B1(
        n20382), .B2(n20559), .ZN(n20347) );
  OAI211_X1 U23256 ( .C1(n20562), .C2(n20360), .A(n20348), .B(n20347), .ZN(
        P1_U3093) );
  AOI22_X1 U23257 ( .A1(n20621), .A2(n20356), .B1(n20620), .B2(n20355), .ZN(
        n20351) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20357), .B1(
        n20349), .B2(n20622), .ZN(n20350) );
  OAI211_X1 U23259 ( .C1(n20625), .C2(n20352), .A(n20351), .B(n20350), .ZN(
        P1_U3094) );
  AOI22_X1 U23260 ( .A1(n20627), .A2(n20356), .B1(n20626), .B2(n20355), .ZN(
        n20354) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20357), .B1(
        n20382), .B2(n20567), .ZN(n20353) );
  OAI211_X1 U23262 ( .C1(n20570), .C2(n20360), .A(n20354), .B(n20353), .ZN(
        P1_U3095) );
  AOI22_X1 U23263 ( .A1(n20635), .A2(n20356), .B1(n20633), .B2(n20355), .ZN(
        n20359) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20357), .B1(
        n20382), .B2(n20573), .ZN(n20358) );
  OAI211_X1 U23265 ( .C1(n20578), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        P1_U3096) );
  NOR3_X1 U23266 ( .A1(n20722), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20391) );
  INV_X1 U23267 ( .A(n20391), .ZN(n20388) );
  NOR2_X1 U23268 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20388), .ZN(
        n20381) );
  NAND2_X1 U23269 ( .A1(n20711), .A2(n13515), .ZN(n20414) );
  INV_X1 U23270 ( .A(n20414), .ZN(n20447) );
  AOI21_X1 U23271 ( .B1(n20447), .B2(n13545), .A(n20381), .ZN(n20363) );
  NAND2_X1 U23272 ( .A1(n20361), .A2(n20415), .ZN(n20481) );
  OAI22_X1 U23273 ( .A1(n20363), .A2(n20590), .B1(n20420), .B2(n20481), .ZN(
        n20380) );
  AOI22_X1 U23274 ( .A1(n20583), .A2(n20381), .B1(n20582), .B2(n20380), .ZN(
        n20367) );
  INV_X1 U23275 ( .A(n20411), .ZN(n20362) );
  OAI21_X1 U23276 ( .B1(n20362), .B2(n20382), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20364) );
  NAND2_X1 U23277 ( .A1(n20364), .A2(n20363), .ZN(n20365) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20592), .ZN(n20366) );
  OAI211_X1 U23279 ( .C1(n20595), .C2(n20411), .A(n20367), .B(n20366), .ZN(
        P1_U3097) );
  AOI22_X1 U23280 ( .A1(n20597), .A2(n20381), .B1(n20596), .B2(n20380), .ZN(
        n20369) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20598), .ZN(n20368) );
  OAI211_X1 U23282 ( .C1(n20601), .C2(n20411), .A(n20369), .B(n20368), .ZN(
        P1_U3098) );
  AOI22_X1 U23283 ( .A1(n20603), .A2(n20381), .B1(n20602), .B2(n20380), .ZN(
        n20371) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20604), .ZN(n20370) );
  OAI211_X1 U23285 ( .C1(n20607), .C2(n20411), .A(n20371), .B(n20370), .ZN(
        P1_U3099) );
  AOI22_X1 U23286 ( .A1(n20609), .A2(n20381), .B1(n20608), .B2(n20380), .ZN(
        n20373) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20610), .ZN(n20372) );
  OAI211_X1 U23288 ( .C1(n20613), .C2(n20411), .A(n20373), .B(n20372), .ZN(
        P1_U3100) );
  AOI22_X1 U23289 ( .A1(n20615), .A2(n20381), .B1(n20614), .B2(n20380), .ZN(
        n20375) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20616), .ZN(n20374) );
  OAI211_X1 U23291 ( .C1(n20619), .C2(n20411), .A(n20375), .B(n20374), .ZN(
        P1_U3101) );
  AOI22_X1 U23292 ( .A1(n20621), .A2(n20381), .B1(n20620), .B2(n20380), .ZN(
        n20377) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20622), .ZN(n20376) );
  OAI211_X1 U23294 ( .C1(n20625), .C2(n20411), .A(n20377), .B(n20376), .ZN(
        P1_U3102) );
  AOI22_X1 U23295 ( .A1(n20627), .A2(n20381), .B1(n20626), .B2(n20380), .ZN(
        n20379) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20628), .ZN(n20378) );
  OAI211_X1 U23297 ( .C1(n20631), .C2(n20411), .A(n20379), .B(n20378), .ZN(
        P1_U3103) );
  AOI22_X1 U23298 ( .A1(n20635), .A2(n20381), .B1(n20633), .B2(n20380), .ZN(
        n20385) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20383), .B1(
        n20382), .B2(n20636), .ZN(n20384) );
  OAI211_X1 U23300 ( .C1(n20642), .C2(n20411), .A(n20385), .B(n20384), .ZN(
        P1_U3104) );
  NOR2_X1 U23301 ( .A1(n20504), .A2(n20388), .ZN(n20407) );
  OR2_X1 U23302 ( .A1(n20414), .A2(n20157), .ZN(n20387) );
  INV_X1 U23303 ( .A(n20407), .ZN(n20386) );
  AND2_X1 U23304 ( .A1(n20387), .A2(n20386), .ZN(n20389) );
  OAI22_X1 U23305 ( .A1(n20389), .A2(n20590), .B1(n20388), .B2(n11673), .ZN(
        n20406) );
  AOI22_X1 U23306 ( .A1(n20583), .A2(n20407), .B1(n20582), .B2(n20406), .ZN(
        n20393) );
  OAI21_X1 U23307 ( .B1(n20708), .B2(n20508), .A(n20389), .ZN(n20390) );
  OAI221_X1 U23308 ( .B1(n20718), .B2(n20391), .C1(n20590), .C2(n20390), .A(
        n20588), .ZN(n20408) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20543), .ZN(n20392) );
  OAI211_X1 U23310 ( .C1(n20546), .C2(n20411), .A(n20393), .B(n20392), .ZN(
        P1_U3105) );
  AOI22_X1 U23311 ( .A1(n20597), .A2(n20407), .B1(n20596), .B2(n20406), .ZN(
        n20395) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20547), .ZN(n20394) );
  OAI211_X1 U23313 ( .C1(n20550), .C2(n20411), .A(n20395), .B(n20394), .ZN(
        P1_U3106) );
  AOI22_X1 U23314 ( .A1(n20603), .A2(n20407), .B1(n20602), .B2(n20406), .ZN(
        n20397) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20551), .ZN(n20396) );
  OAI211_X1 U23316 ( .C1(n20554), .C2(n20411), .A(n20397), .B(n20396), .ZN(
        P1_U3107) );
  AOI22_X1 U23317 ( .A1(n20609), .A2(n20407), .B1(n20608), .B2(n20406), .ZN(
        n20399) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20555), .ZN(n20398) );
  OAI211_X1 U23319 ( .C1(n20558), .C2(n20411), .A(n20399), .B(n20398), .ZN(
        P1_U3108) );
  AOI22_X1 U23320 ( .A1(n20615), .A2(n20407), .B1(n20614), .B2(n20406), .ZN(
        n20401) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20559), .ZN(n20400) );
  OAI211_X1 U23322 ( .C1(n20562), .C2(n20411), .A(n20401), .B(n20400), .ZN(
        P1_U3109) );
  AOI22_X1 U23323 ( .A1(n20621), .A2(n20407), .B1(n20620), .B2(n20406), .ZN(
        n20403) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20563), .ZN(n20402) );
  OAI211_X1 U23325 ( .C1(n20566), .C2(n20411), .A(n20403), .B(n20402), .ZN(
        P1_U3110) );
  AOI22_X1 U23326 ( .A1(n20627), .A2(n20407), .B1(n20626), .B2(n20406), .ZN(
        n20405) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20567), .ZN(n20404) );
  OAI211_X1 U23328 ( .C1(n20570), .C2(n20411), .A(n20405), .B(n20404), .ZN(
        P1_U3111) );
  AOI22_X1 U23329 ( .A1(n20635), .A2(n20407), .B1(n20633), .B2(n20406), .ZN(
        n20410) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20408), .B1(
        n20435), .B2(n20573), .ZN(n20409) );
  OAI211_X1 U23331 ( .C1(n20578), .C2(n20411), .A(n20410), .B(n20409), .ZN(
        P1_U3112) );
  NOR3_X1 U23332 ( .A1(n20722), .A2(n20412), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20450) );
  INV_X1 U23333 ( .A(n20450), .ZN(n20448) );
  NOR2_X1 U23334 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20448), .ZN(
        n20438) );
  AOI22_X1 U23335 ( .A1(n20583), .A2(n20438), .B1(n20470), .B2(n20543), .ZN(
        n20424) );
  OAI21_X1 U23336 ( .B1(n20470), .B2(n20435), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20413) );
  NAND2_X1 U23337 ( .A1(n20413), .A2(n20718), .ZN(n20422) );
  NOR2_X1 U23338 ( .A1(n20414), .A2(n13545), .ZN(n20419) );
  OR2_X1 U23339 ( .A1(n20415), .A2(n20722), .ZN(n20533) );
  NAND2_X1 U23340 ( .A1(n20533), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20540) );
  OAI211_X1 U23341 ( .C1(n20479), .C2(n20438), .A(n20540), .B(n20416), .ZN(
        n20417) );
  INV_X1 U23342 ( .A(n20417), .ZN(n20418) );
  INV_X1 U23343 ( .A(n20419), .ZN(n20421) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20440), .B1(
        n20582), .B2(n20439), .ZN(n20423) );
  OAI211_X1 U23345 ( .C1(n20546), .C2(n20443), .A(n20424), .B(n20423), .ZN(
        P1_U3113) );
  AOI22_X1 U23346 ( .A1(n20597), .A2(n20438), .B1(n20470), .B2(n20547), .ZN(
        n20426) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20440), .B1(
        n20596), .B2(n20439), .ZN(n20425) );
  OAI211_X1 U23348 ( .C1(n20550), .C2(n20443), .A(n20426), .B(n20425), .ZN(
        P1_U3114) );
  AOI22_X1 U23349 ( .A1(n20603), .A2(n20438), .B1(n20470), .B2(n20551), .ZN(
        n20428) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20440), .B1(
        n20602), .B2(n20439), .ZN(n20427) );
  OAI211_X1 U23351 ( .C1(n20554), .C2(n20443), .A(n20428), .B(n20427), .ZN(
        P1_U3115) );
  AOI22_X1 U23352 ( .A1(n20609), .A2(n20438), .B1(n20435), .B2(n20610), .ZN(
        n20430) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20440), .B1(
        n20608), .B2(n20439), .ZN(n20429) );
  OAI211_X1 U23354 ( .C1(n20613), .C2(n20467), .A(n20430), .B(n20429), .ZN(
        P1_U3116) );
  AOI22_X1 U23355 ( .A1(n20615), .A2(n20438), .B1(n20435), .B2(n20616), .ZN(
        n20432) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20440), .B1(
        n20614), .B2(n20439), .ZN(n20431) );
  OAI211_X1 U23357 ( .C1(n20619), .C2(n20467), .A(n20432), .B(n20431), .ZN(
        P1_U3117) );
  AOI22_X1 U23358 ( .A1(n20621), .A2(n20438), .B1(n20470), .B2(n20563), .ZN(
        n20434) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20440), .B1(
        n20620), .B2(n20439), .ZN(n20433) );
  OAI211_X1 U23360 ( .C1(n20566), .C2(n20443), .A(n20434), .B(n20433), .ZN(
        P1_U3118) );
  AOI22_X1 U23361 ( .A1(n20627), .A2(n20438), .B1(n20435), .B2(n20628), .ZN(
        n20437) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20440), .B1(
        n20626), .B2(n20439), .ZN(n20436) );
  OAI211_X1 U23363 ( .C1(n20631), .C2(n20467), .A(n20437), .B(n20436), .ZN(
        P1_U3119) );
  AOI22_X1 U23364 ( .A1(n20635), .A2(n20438), .B1(n20470), .B2(n20573), .ZN(
        n20442) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20440), .B1(
        n20633), .B2(n20439), .ZN(n20441) );
  OAI211_X1 U23366 ( .C1(n20578), .C2(n20443), .A(n20442), .B(n20441), .ZN(
        P1_U3120) );
  NOR2_X1 U23367 ( .A1(n20722), .A2(n20446), .ZN(n20469) );
  AOI21_X1 U23368 ( .B1(n20447), .B2(n20579), .A(n20469), .ZN(n20449) );
  OAI22_X1 U23369 ( .A1(n20449), .A2(n20590), .B1(n20448), .B2(n11673), .ZN(
        n20468) );
  AOI22_X1 U23370 ( .A1(n20583), .A2(n20469), .B1(n20582), .B2(n20468), .ZN(
        n20453) );
  NOR3_X1 U23371 ( .A1(n20708), .A2(n20590), .A3(n20586), .ZN(n20451) );
  OAI21_X1 U23372 ( .B1(n20451), .B2(n20450), .A(n20588), .ZN(n20471) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20471), .B1(
        n20470), .B2(n20592), .ZN(n20452) );
  OAI211_X1 U23374 ( .C1(n20595), .C2(n20503), .A(n20453), .B(n20452), .ZN(
        P1_U3121) );
  AOI22_X1 U23375 ( .A1(n20597), .A2(n20469), .B1(n20596), .B2(n20468), .ZN(
        n20455) );
  INV_X1 U23376 ( .A(n20503), .ZN(n20464) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20471), .B1(
        n20464), .B2(n20547), .ZN(n20454) );
  OAI211_X1 U23378 ( .C1(n20550), .C2(n20467), .A(n20455), .B(n20454), .ZN(
        P1_U3122) );
  AOI22_X1 U23379 ( .A1(n20603), .A2(n20469), .B1(n20602), .B2(n20468), .ZN(
        n20457) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20471), .B1(
        n20464), .B2(n20551), .ZN(n20456) );
  OAI211_X1 U23381 ( .C1(n20554), .C2(n20467), .A(n20457), .B(n20456), .ZN(
        P1_U3123) );
  AOI22_X1 U23382 ( .A1(n20609), .A2(n20469), .B1(n20608), .B2(n20468), .ZN(
        n20459) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20471), .B1(
        n20470), .B2(n20610), .ZN(n20458) );
  OAI211_X1 U23384 ( .C1(n20613), .C2(n20503), .A(n20459), .B(n20458), .ZN(
        P1_U3124) );
  AOI22_X1 U23385 ( .A1(n20615), .A2(n20469), .B1(n20614), .B2(n20468), .ZN(
        n20461) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20471), .B1(
        n20464), .B2(n20559), .ZN(n20460) );
  OAI211_X1 U23387 ( .C1(n20562), .C2(n20467), .A(n20461), .B(n20460), .ZN(
        P1_U3125) );
  AOI22_X1 U23388 ( .A1(n20621), .A2(n20469), .B1(n20620), .B2(n20468), .ZN(
        n20463) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20471), .B1(
        n20464), .B2(n20563), .ZN(n20462) );
  OAI211_X1 U23390 ( .C1(n20566), .C2(n20467), .A(n20463), .B(n20462), .ZN(
        P1_U3126) );
  AOI22_X1 U23391 ( .A1(n20627), .A2(n20469), .B1(n20626), .B2(n20468), .ZN(
        n20466) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20471), .B1(
        n20464), .B2(n20567), .ZN(n20465) );
  OAI211_X1 U23393 ( .C1(n20570), .C2(n20467), .A(n20466), .B(n20465), .ZN(
        P1_U3127) );
  AOI22_X1 U23394 ( .A1(n20635), .A2(n20469), .B1(n20633), .B2(n20468), .ZN(
        n20473) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20471), .B1(
        n20470), .B2(n20636), .ZN(n20472) );
  OAI211_X1 U23396 ( .C1(n20642), .C2(n20503), .A(n20473), .B(n20472), .ZN(
        P1_U3128) );
  NOR3_X1 U23397 ( .A1(n20474), .A2(n20722), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20510) );
  INV_X1 U23398 ( .A(n20510), .ZN(n20506) );
  NOR2_X1 U23399 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20506), .ZN(
        n20498) );
  AOI22_X1 U23400 ( .A1(n20583), .A2(n20498), .B1(n20527), .B2(n20543), .ZN(
        n20485) );
  INV_X1 U23401 ( .A(n20527), .ZN(n20475) );
  NAND2_X1 U23402 ( .A1(n20503), .A2(n20475), .ZN(n20476) );
  AOI21_X1 U23403 ( .B1(n20476), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20590), 
        .ZN(n20480) );
  NOR2_X1 U23404 ( .A1(n13515), .A2(n20477), .ZN(n20580) );
  NAND2_X1 U23405 ( .A1(n20580), .A2(n13545), .ZN(n20482) );
  AOI22_X1 U23406 ( .A1(n20480), .A2(n20482), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20481), .ZN(n20478) );
  OAI211_X1 U23407 ( .C1(n20498), .C2(n20479), .A(n20541), .B(n20478), .ZN(
        n20500) );
  INV_X1 U23408 ( .A(n20480), .ZN(n20483) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20500), .B1(
        n20582), .B2(n20499), .ZN(n20484) );
  OAI211_X1 U23410 ( .C1(n20546), .C2(n20503), .A(n20485), .B(n20484), .ZN(
        P1_U3129) );
  AOI22_X1 U23411 ( .A1(n20597), .A2(n20498), .B1(n20527), .B2(n20547), .ZN(
        n20487) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20500), .B1(
        n20596), .B2(n20499), .ZN(n20486) );
  OAI211_X1 U23413 ( .C1(n20550), .C2(n20503), .A(n20487), .B(n20486), .ZN(
        P1_U3130) );
  AOI22_X1 U23414 ( .A1(n20603), .A2(n20498), .B1(n20527), .B2(n20551), .ZN(
        n20489) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20500), .B1(
        n20602), .B2(n20499), .ZN(n20488) );
  OAI211_X1 U23416 ( .C1(n20554), .C2(n20503), .A(n20489), .B(n20488), .ZN(
        P1_U3131) );
  AOI22_X1 U23417 ( .A1(n20609), .A2(n20498), .B1(n20527), .B2(n20555), .ZN(
        n20491) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20500), .B1(
        n20608), .B2(n20499), .ZN(n20490) );
  OAI211_X1 U23419 ( .C1(n20558), .C2(n20503), .A(n20491), .B(n20490), .ZN(
        P1_U3132) );
  AOI22_X1 U23420 ( .A1(n20615), .A2(n20498), .B1(n20527), .B2(n20559), .ZN(
        n20493) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20500), .B1(
        n20614), .B2(n20499), .ZN(n20492) );
  OAI211_X1 U23422 ( .C1(n20562), .C2(n20503), .A(n20493), .B(n20492), .ZN(
        P1_U3133) );
  AOI22_X1 U23423 ( .A1(n20621), .A2(n20498), .B1(n20527), .B2(n20563), .ZN(
        n20495) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20500), .B1(
        n20620), .B2(n20499), .ZN(n20494) );
  OAI211_X1 U23425 ( .C1(n20566), .C2(n20503), .A(n20495), .B(n20494), .ZN(
        P1_U3134) );
  AOI22_X1 U23426 ( .A1(n20627), .A2(n20498), .B1(n20527), .B2(n20567), .ZN(
        n20497) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20500), .B1(
        n20626), .B2(n20499), .ZN(n20496) );
  OAI211_X1 U23428 ( .C1(n20570), .C2(n20503), .A(n20497), .B(n20496), .ZN(
        P1_U3135) );
  AOI22_X1 U23429 ( .A1(n20635), .A2(n20498), .B1(n20527), .B2(n20573), .ZN(
        n20502) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20500), .B1(
        n20633), .B2(n20499), .ZN(n20501) );
  OAI211_X1 U23431 ( .C1(n20578), .C2(n20503), .A(n20502), .B(n20501), .ZN(
        P1_U3136) );
  NOR2_X1 U23432 ( .A1(n20504), .A2(n20506), .ZN(n20526) );
  AOI21_X1 U23433 ( .B1(n20580), .B2(n20505), .A(n20526), .ZN(n20507) );
  OAI22_X1 U23434 ( .A1(n20507), .A2(n20590), .B1(n20506), .B2(n11673), .ZN(
        n20525) );
  AOI22_X1 U23435 ( .A1(n20583), .A2(n20526), .B1(n20582), .B2(n20525), .ZN(
        n20512) );
  NOR2_X1 U23436 ( .A1(n20508), .A2(n20590), .ZN(n20509) );
  AND2_X1 U23437 ( .A1(n20584), .A2(n20509), .ZN(n20715) );
  OAI21_X1 U23438 ( .B1(n20510), .B2(n20715), .A(n20588), .ZN(n20528) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20592), .ZN(n20511) );
  OAI211_X1 U23440 ( .C1(n20595), .C2(n20577), .A(n20512), .B(n20511), .ZN(
        P1_U3137) );
  AOI22_X1 U23441 ( .A1(n20597), .A2(n20526), .B1(n20596), .B2(n20525), .ZN(
        n20514) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20598), .ZN(n20513) );
  OAI211_X1 U23443 ( .C1(n20601), .C2(n20577), .A(n20514), .B(n20513), .ZN(
        P1_U3138) );
  AOI22_X1 U23444 ( .A1(n20603), .A2(n20526), .B1(n20602), .B2(n20525), .ZN(
        n20516) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20604), .ZN(n20515) );
  OAI211_X1 U23446 ( .C1(n20607), .C2(n20577), .A(n20516), .B(n20515), .ZN(
        P1_U3139) );
  AOI22_X1 U23447 ( .A1(n20609), .A2(n20526), .B1(n20608), .B2(n20525), .ZN(
        n20518) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20610), .ZN(n20517) );
  OAI211_X1 U23449 ( .C1(n20613), .C2(n20577), .A(n20518), .B(n20517), .ZN(
        P1_U3140) );
  AOI22_X1 U23450 ( .A1(n20615), .A2(n20526), .B1(n20614), .B2(n20525), .ZN(
        n20520) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20616), .ZN(n20519) );
  OAI211_X1 U23452 ( .C1(n20619), .C2(n20577), .A(n20520), .B(n20519), .ZN(
        P1_U3141) );
  AOI22_X1 U23453 ( .A1(n20621), .A2(n20526), .B1(n20620), .B2(n20525), .ZN(
        n20522) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20622), .ZN(n20521) );
  OAI211_X1 U23455 ( .C1(n20625), .C2(n20577), .A(n20522), .B(n20521), .ZN(
        P1_U3142) );
  AOI22_X1 U23456 ( .A1(n20627), .A2(n20526), .B1(n20626), .B2(n20525), .ZN(
        n20524) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20628), .ZN(n20523) );
  OAI211_X1 U23458 ( .C1(n20631), .C2(n20577), .A(n20524), .B(n20523), .ZN(
        P1_U3143) );
  AOI22_X1 U23459 ( .A1(n20635), .A2(n20526), .B1(n20633), .B2(n20525), .ZN(
        n20530) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20528), .B1(
        n20527), .B2(n20636), .ZN(n20529) );
  OAI211_X1 U23461 ( .C1(n20642), .C2(n20577), .A(n20530), .B(n20529), .ZN(
        P1_U3144) );
  NOR2_X1 U23462 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20581), .ZN(
        n20572) );
  NAND3_X1 U23463 ( .A1(n20580), .A2(n20538), .A3(n20718), .ZN(n20531) );
  OAI21_X1 U23464 ( .B1(n20533), .B2(n20532), .A(n20531), .ZN(n20571) );
  AOI22_X1 U23465 ( .A1(n20583), .A2(n20572), .B1(n20582), .B2(n20571), .ZN(
        n20545) );
  INV_X1 U23466 ( .A(n20637), .ZN(n20536) );
  AOI21_X1 U23467 ( .B1(n20536), .B2(n20577), .A(n20535), .ZN(n20537) );
  AOI21_X1 U23468 ( .B1(n20580), .B2(n20538), .A(n20537), .ZN(n20539) );
  NOR2_X1 U23469 ( .A1(n20539), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20542) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20543), .ZN(n20544) );
  OAI211_X1 U23471 ( .C1(n20546), .C2(n20577), .A(n20545), .B(n20544), .ZN(
        P1_U3145) );
  AOI22_X1 U23472 ( .A1(n20597), .A2(n20572), .B1(n20596), .B2(n20571), .ZN(
        n20549) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20547), .ZN(n20548) );
  OAI211_X1 U23474 ( .C1(n20550), .C2(n20577), .A(n20549), .B(n20548), .ZN(
        P1_U3146) );
  AOI22_X1 U23475 ( .A1(n20603), .A2(n20572), .B1(n20602), .B2(n20571), .ZN(
        n20553) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20551), .ZN(n20552) );
  OAI211_X1 U23477 ( .C1(n20554), .C2(n20577), .A(n20553), .B(n20552), .ZN(
        P1_U3147) );
  AOI22_X1 U23478 ( .A1(n20609), .A2(n20572), .B1(n20608), .B2(n20571), .ZN(
        n20557) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20555), .ZN(n20556) );
  OAI211_X1 U23480 ( .C1(n20558), .C2(n20577), .A(n20557), .B(n20556), .ZN(
        P1_U3148) );
  AOI22_X1 U23481 ( .A1(n20615), .A2(n20572), .B1(n20614), .B2(n20571), .ZN(
        n20561) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20559), .ZN(n20560) );
  OAI211_X1 U23483 ( .C1(n20562), .C2(n20577), .A(n20561), .B(n20560), .ZN(
        P1_U3149) );
  AOI22_X1 U23484 ( .A1(n20621), .A2(n20572), .B1(n20620), .B2(n20571), .ZN(
        n20565) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20563), .ZN(n20564) );
  OAI211_X1 U23486 ( .C1(n20566), .C2(n20577), .A(n20565), .B(n20564), .ZN(
        P1_U3150) );
  AOI22_X1 U23487 ( .A1(n20627), .A2(n20572), .B1(n20626), .B2(n20571), .ZN(
        n20569) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20567), .ZN(n20568) );
  OAI211_X1 U23489 ( .C1(n20570), .C2(n20577), .A(n20569), .B(n20568), .ZN(
        P1_U3151) );
  AOI22_X1 U23490 ( .A1(n20635), .A2(n20572), .B1(n20633), .B2(n20571), .ZN(
        n20576) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20574), .B1(
        n20637), .B2(n20573), .ZN(n20575) );
  OAI211_X1 U23492 ( .C1(n20578), .C2(n20577), .A(n20576), .B(n20575), .ZN(
        P1_U3152) );
  AOI21_X1 U23493 ( .B1(n20580), .B2(n20579), .A(n20634), .ZN(n20585) );
  OAI22_X1 U23494 ( .A1(n20585), .A2(n20590), .B1(n20581), .B2(n11673), .ZN(
        n20632) );
  AOI22_X1 U23495 ( .A1(n20583), .A2(n20634), .B1(n20582), .B2(n20632), .ZN(
        n20594) );
  INV_X1 U23496 ( .A(n20584), .ZN(n20587) );
  OAI21_X1 U23497 ( .B1(n20587), .B2(n20586), .A(n20585), .ZN(n20589) );
  OAI221_X1 U23498 ( .B1(n20718), .B2(n20591), .C1(n20590), .C2(n20589), .A(
        n20588), .ZN(n20638) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20592), .ZN(n20593) );
  OAI211_X1 U23500 ( .C1(n20595), .C2(n20641), .A(n20594), .B(n20593), .ZN(
        P1_U3153) );
  AOI22_X1 U23501 ( .A1(n20597), .A2(n20634), .B1(n20596), .B2(n20632), .ZN(
        n20600) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20598), .ZN(n20599) );
  OAI211_X1 U23503 ( .C1(n20601), .C2(n20641), .A(n20600), .B(n20599), .ZN(
        P1_U3154) );
  AOI22_X1 U23504 ( .A1(n20603), .A2(n20634), .B1(n20602), .B2(n20632), .ZN(
        n20606) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20604), .ZN(n20605) );
  OAI211_X1 U23506 ( .C1(n20607), .C2(n20641), .A(n20606), .B(n20605), .ZN(
        P1_U3155) );
  AOI22_X1 U23507 ( .A1(n20609), .A2(n20634), .B1(n20608), .B2(n20632), .ZN(
        n20612) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20610), .ZN(n20611) );
  OAI211_X1 U23509 ( .C1(n20613), .C2(n20641), .A(n20612), .B(n20611), .ZN(
        P1_U3156) );
  AOI22_X1 U23510 ( .A1(n20615), .A2(n20634), .B1(n20614), .B2(n20632), .ZN(
        n20618) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20616), .ZN(n20617) );
  OAI211_X1 U23512 ( .C1(n20619), .C2(n20641), .A(n20618), .B(n20617), .ZN(
        P1_U3157) );
  AOI22_X1 U23513 ( .A1(n20621), .A2(n20634), .B1(n20620), .B2(n20632), .ZN(
        n20624) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20622), .ZN(n20623) );
  OAI211_X1 U23515 ( .C1(n20625), .C2(n20641), .A(n20624), .B(n20623), .ZN(
        P1_U3158) );
  AOI22_X1 U23516 ( .A1(n20627), .A2(n20634), .B1(n20626), .B2(n20632), .ZN(
        n20630) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20628), .ZN(n20629) );
  OAI211_X1 U23518 ( .C1(n20631), .C2(n20641), .A(n20630), .B(n20629), .ZN(
        P1_U3159) );
  AOI22_X1 U23519 ( .A1(n20635), .A2(n20634), .B1(n20633), .B2(n20632), .ZN(
        n20640) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20636), .ZN(n20639) );
  OAI211_X1 U23521 ( .C1(n20642), .C2(n20641), .A(n20640), .B(n20639), .ZN(
        P1_U3160) );
  NOR2_X1 U23522 ( .A1(n20644), .A2(n20643), .ZN(n20646) );
  OAI21_X1 U23523 ( .B1(n20646), .B2(n11673), .A(n20645), .ZN(P1_U3163) );
  AND2_X1 U23524 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20647), .ZN(
        P1_U3164) );
  AND2_X1 U23525 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20647), .ZN(
        P1_U3165) );
  AND2_X1 U23526 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20647), .ZN(
        P1_U3166) );
  AND2_X1 U23527 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20647), .ZN(
        P1_U3167) );
  AND2_X1 U23528 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20647), .ZN(
        P1_U3168) );
  AND2_X1 U23529 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20647), .ZN(
        P1_U3169) );
  AND2_X1 U23530 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20647), .ZN(
        P1_U3170) );
  AND2_X1 U23531 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20647), .ZN(
        P1_U3171) );
  AND2_X1 U23532 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20647), .ZN(
        P1_U3172) );
  AND2_X1 U23533 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20647), .ZN(
        P1_U3173) );
  AND2_X1 U23534 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20647), .ZN(
        P1_U3174) );
  AND2_X1 U23535 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20647), .ZN(
        P1_U3175) );
  AND2_X1 U23536 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20647), .ZN(
        P1_U3176) );
  INV_X1 U23537 ( .A(P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20888) );
  NOR2_X1 U23538 ( .A1(n20707), .A2(n20888), .ZN(P1_U3177) );
  AND2_X1 U23539 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20647), .ZN(
        P1_U3178) );
  AND2_X1 U23540 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20647), .ZN(
        P1_U3179) );
  AND2_X1 U23541 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20647), .ZN(
        P1_U3180) );
  AND2_X1 U23542 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20647), .ZN(
        P1_U3181) );
  AND2_X1 U23543 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20647), .ZN(
        P1_U3182) );
  AND2_X1 U23544 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20647), .ZN(
        P1_U3183) );
  AND2_X1 U23545 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20647), .ZN(
        P1_U3184) );
  AND2_X1 U23546 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20647), .ZN(
        P1_U3185) );
  AND2_X1 U23547 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20647), .ZN(P1_U3186) );
  AND2_X1 U23548 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20647), .ZN(P1_U3187) );
  AND2_X1 U23549 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20647), .ZN(P1_U3188) );
  AND2_X1 U23550 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20647), .ZN(P1_U3189) );
  AND2_X1 U23551 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20647), .ZN(P1_U3190) );
  AND2_X1 U23552 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20647), .ZN(P1_U3191) );
  AND2_X1 U23553 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20647), .ZN(P1_U3192) );
  AND2_X1 U23554 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20647), .ZN(P1_U3193) );
  AOI21_X1 U23555 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20736), .A(n20657), 
        .ZN(n20659) );
  OAI22_X1 U23556 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20653), .B1(n20660), 
        .B2(n20648), .ZN(n20649) );
  NOR3_X1 U23557 ( .A1(n20650), .A2(n20743), .A3(n20649), .ZN(n20651) );
  OAI22_X1 U23558 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20659), .B1(n20732), 
        .B2(n20651), .ZN(P1_U3194) );
  AOI222_X1 U23559 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20653), .B1(
        P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_1__SCAN_IN), .C1(n20653), 
        .C2(n20652), .ZN(n20658) );
  OAI211_X1 U23560 ( .C1(NA), .C2(n20654), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20660), .ZN(n20655) );
  OAI211_X1 U23561 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20743), .A(HOLD), .B(
        n20655), .ZN(n20656) );
  OAI22_X1 U23562 ( .A1(n20659), .A2(n20658), .B1(n20657), .B2(n20656), .ZN(
        P1_U3196) );
  NAND2_X1 U23563 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20732), .ZN(n20688) );
  NAND2_X1 U23564 ( .A1(n20660), .A2(n20732), .ZN(n20683) );
  AOI22_X1 U23565 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20933), .ZN(n20661) );
  OAI21_X1 U23566 ( .B1(n20724), .B2(n20688), .A(n20661), .ZN(P1_U3197) );
  INV_X1 U23567 ( .A(n20688), .ZN(n20934) );
  AOI22_X1 U23568 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20934), .ZN(n20662) );
  OAI21_X1 U23569 ( .B1(n13593), .B2(n20683), .A(n20662), .ZN(P1_U3198) );
  INV_X1 U23570 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20758) );
  OAI222_X1 U23571 ( .A1(n20688), .A2(n13593), .B1(n20758), .B2(n20732), .C1(
        n20663), .C2(n20683), .ZN(P1_U3199) );
  AOI222_X1 U23572 ( .A1(n20933), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20934), .ZN(n20664) );
  INV_X1 U23573 ( .A(n20664), .ZN(P1_U3200) );
  AOI222_X1 U23574 ( .A1(n20934), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20933), .ZN(n20665) );
  INV_X1 U23575 ( .A(n20665), .ZN(P1_U3201) );
  AOI222_X1 U23576 ( .A1(n20934), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20933), .ZN(n20666) );
  INV_X1 U23577 ( .A(n20666), .ZN(P1_U3202) );
  AOI222_X1 U23578 ( .A1(n20934), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20933), .ZN(n20667) );
  INV_X1 U23579 ( .A(n20667), .ZN(P1_U3203) );
  AOI22_X1 U23580 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20933), .ZN(n20668) );
  OAI21_X1 U23581 ( .B1(n20669), .B2(n20688), .A(n20668), .ZN(P1_U3204) );
  AOI22_X1 U23582 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20934), .ZN(n20670) );
  OAI21_X1 U23583 ( .B1(n20671), .B2(n20683), .A(n20670), .ZN(P1_U3205) );
  AOI222_X1 U23584 ( .A1(n20934), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20933), .ZN(n20672) );
  INV_X1 U23585 ( .A(n20672), .ZN(P1_U3206) );
  AOI22_X1 U23586 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20933), .ZN(n20673) );
  OAI21_X1 U23587 ( .B1(n20674), .B2(n20688), .A(n20673), .ZN(P1_U3207) );
  AOI22_X1 U23588 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20934), .ZN(n20675) );
  OAI21_X1 U23589 ( .B1(n20676), .B2(n20683), .A(n20675), .ZN(P1_U3208) );
  AOI222_X1 U23590 ( .A1(n20934), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20933), .ZN(n20677) );
  INV_X1 U23591 ( .A(n20677), .ZN(P1_U3209) );
  AOI22_X1 U23592 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20933), .ZN(n20678) );
  OAI21_X1 U23593 ( .B1(n20679), .B2(n20688), .A(n20678), .ZN(P1_U3210) );
  AOI22_X1 U23594 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20933), .ZN(n20680) );
  OAI21_X1 U23595 ( .B1(n20681), .B2(n20688), .A(n20680), .ZN(P1_U3212) );
  AOI22_X1 U23596 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20934), .ZN(n20682) );
  OAI21_X1 U23597 ( .B1(n20685), .B2(n20683), .A(n20682), .ZN(P1_U3213) );
  AOI22_X1 U23598 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20933), .ZN(n20684) );
  OAI21_X1 U23599 ( .B1(n20685), .B2(n20688), .A(n20684), .ZN(P1_U3214) );
  AOI222_X1 U23600 ( .A1(n20933), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20934), .ZN(n20686) );
  INV_X1 U23601 ( .A(n20686), .ZN(P1_U3215) );
  AOI22_X1 U23602 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20745), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20933), .ZN(n20687) );
  OAI21_X1 U23603 ( .B1(n20689), .B2(n20688), .A(n20687), .ZN(P1_U3216) );
  AOI222_X1 U23604 ( .A1(n20934), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20933), .ZN(n20690) );
  INV_X1 U23605 ( .A(n20690), .ZN(P1_U3217) );
  AOI222_X1 U23606 ( .A1(n20934), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20933), .ZN(n20691) );
  INV_X1 U23607 ( .A(n20691), .ZN(P1_U3218) );
  AOI222_X1 U23608 ( .A1(n20934), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20933), .ZN(n20692) );
  INV_X1 U23609 ( .A(n20692), .ZN(P1_U3219) );
  AOI222_X1 U23610 ( .A1(n20934), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20933), .ZN(n20693) );
  INV_X1 U23611 ( .A(n20693), .ZN(P1_U3220) );
  AOI222_X1 U23612 ( .A1(n20934), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20933), .ZN(n20694) );
  INV_X1 U23613 ( .A(n20694), .ZN(P1_U3221) );
  AOI222_X1 U23614 ( .A1(n20934), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20933), .ZN(n20695) );
  INV_X1 U23615 ( .A(n20695), .ZN(P1_U3222) );
  AOI222_X1 U23616 ( .A1(n20934), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20933), .ZN(n20696) );
  INV_X1 U23617 ( .A(n20696), .ZN(P1_U3223) );
  AOI222_X1 U23618 ( .A1(n20934), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20933), .ZN(n20697) );
  INV_X1 U23619 ( .A(n20697), .ZN(P1_U3224) );
  AOI222_X1 U23620 ( .A1(n20934), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20933), .ZN(n20698) );
  INV_X1 U23621 ( .A(n20698), .ZN(P1_U3225) );
  AOI222_X1 U23622 ( .A1(n20934), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20745), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20933), .ZN(n20699) );
  INV_X1 U23623 ( .A(n20699), .ZN(P1_U3226) );
  OAI22_X1 U23624 ( .A1(n20745), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20732), .ZN(n20700) );
  INV_X1 U23625 ( .A(n20700), .ZN(P1_U3458) );
  OAI22_X1 U23626 ( .A1(n20745), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20732), .ZN(n20701) );
  INV_X1 U23627 ( .A(n20701), .ZN(P1_U3459) );
  OAI22_X1 U23628 ( .A1(n20745), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20732), .ZN(n20702) );
  INV_X1 U23629 ( .A(n20702), .ZN(P1_U3460) );
  OAI22_X1 U23630 ( .A1(n20745), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20732), .ZN(n20703) );
  INV_X1 U23631 ( .A(n20703), .ZN(P1_U3461) );
  OAI21_X1 U23632 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20707), .A(n20705), 
        .ZN(n20704) );
  INV_X1 U23633 ( .A(n20704), .ZN(P1_U3464) );
  OAI21_X1 U23634 ( .B1(n20707), .B2(n20706), .A(n20705), .ZN(P1_U3465) );
  OAI211_X1 U23635 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20710), .A(n20709), 
        .B(n20708), .ZN(n20717) );
  INV_X1 U23636 ( .A(n20711), .ZN(n20714) );
  INV_X1 U23637 ( .A(n20712), .ZN(n20713) );
  NOR2_X1 U23638 ( .A1(n20714), .A2(n20713), .ZN(n20716) );
  AOI211_X1 U23639 ( .C1(n20718), .C2(n20717), .A(n20716), .B(n20715), .ZN(
        n20719) );
  OR2_X1 U23640 ( .A1(n20720), .A2(n20719), .ZN(n20721) );
  OAI21_X1 U23641 ( .B1(n20723), .B2(n20722), .A(n20721), .ZN(P1_U3475) );
  AOI21_X1 U23642 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20725) );
  AOI22_X1 U23643 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20725), .B2(n20724), .ZN(n20728) );
  INV_X1 U23644 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20727) );
  AOI22_X1 U23645 ( .A1(n20731), .A2(n20728), .B1(n20727), .B2(n20726), .ZN(
        P1_U3481) );
  INV_X1 U23646 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20730) );
  OAI21_X1 U23647 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20731), .ZN(n20729) );
  OAI21_X1 U23648 ( .B1(n20731), .B2(n20730), .A(n20729), .ZN(P1_U3482) );
  AOI22_X1 U23649 ( .A1(n20732), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20759), 
        .B2(n20745), .ZN(P1_U3483) );
  OAI211_X1 U23650 ( .C1(n20736), .C2(n20735), .A(n20734), .B(n20733), .ZN(
        n20744) );
  NOR2_X1 U23651 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20737), .ZN(n20742) );
  OAI211_X1 U23652 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20739), .A(n20738), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20740) );
  NAND2_X1 U23653 ( .A1(n20744), .A2(n20740), .ZN(n20741) );
  OAI22_X1 U23654 ( .A1(n20744), .A2(n20743), .B1(n20742), .B2(n20741), .ZN(
        P1_U3485) );
  MUX2_X1 U23655 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20745), .Z(P1_U3486) );
  INV_X1 U23656 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20915) );
  INV_X1 U23657 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20906) );
  AOI22_X1 U23658 ( .A1(n20915), .A2(keyinput95), .B1(keyinput126), .B2(n20906), .ZN(n20746) );
  OAI221_X1 U23659 ( .B1(n20915), .B2(keyinput95), .C1(n20906), .C2(
        keyinput126), .A(n20746), .ZN(n20756) );
  INV_X1 U23660 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n20748) );
  AOI22_X1 U23661 ( .A1(n20748), .A2(keyinput76), .B1(keyinput93), .B2(n20898), 
        .ZN(n20747) );
  OAI221_X1 U23662 ( .B1(n20748), .B2(keyinput76), .C1(n20898), .C2(keyinput93), .A(n20747), .ZN(n20755) );
  INV_X1 U23663 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U23664 ( .A1(n20897), .A2(keyinput122), .B1(keyinput83), .B2(n20901), .ZN(n20749) );
  OAI221_X1 U23665 ( .B1(n20897), .B2(keyinput122), .C1(n20901), .C2(
        keyinput83), .A(n20749), .ZN(n20754) );
  XOR2_X1 U23666 ( .A(n20750), .B(keyinput64), .Z(n20752) );
  XNOR2_X1 U23667 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B(keyinput123), .ZN(
        n20751) );
  NAND2_X1 U23668 ( .A1(n20752), .A2(n20751), .ZN(n20753) );
  NOR4_X1 U23669 ( .A1(n20756), .A2(n20755), .A3(n20754), .A4(n20753), .ZN(
        n20794) );
  AOI22_X1 U23670 ( .A1(n20759), .A2(keyinput104), .B1(n20758), .B2(keyinput73), .ZN(n20757) );
  OAI221_X1 U23671 ( .B1(n20759), .B2(keyinput104), .C1(n20758), .C2(
        keyinput73), .A(n20757), .ZN(n20767) );
  AOI22_X1 U23672 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput110), 
        .B1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B2(keyinput99), .ZN(n20760) );
  OAI221_X1 U23673 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput110), 
        .C1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .C2(keyinput99), .A(n20760), .ZN(
        n20766) );
  XNOR2_X1 U23674 ( .A(n20888), .B(keyinput96), .ZN(n20765) );
  XOR2_X1 U23675 ( .A(n14525), .B(keyinput121), .Z(n20763) );
  XNOR2_X1 U23676 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B(keyinput120), .ZN(
        n20762) );
  XNOR2_X1 U23677 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B(keyinput112), .ZN(
        n20761) );
  NAND3_X1 U23678 ( .A1(n20763), .A2(n20762), .A3(n20761), .ZN(n20764) );
  NOR4_X1 U23679 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20793) );
  INV_X1 U23680 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U23681 ( .A1(n20883), .A2(keyinput68), .B1(keyinput69), .B2(n20913), 
        .ZN(n20768) );
  OAI221_X1 U23682 ( .B1(n20883), .B2(keyinput68), .C1(n20913), .C2(keyinput69), .A(n20768), .ZN(n20778) );
  AOI22_X1 U23683 ( .A1(n20884), .A2(keyinput100), .B1(keyinput90), .B2(n20770), .ZN(n20769) );
  OAI221_X1 U23684 ( .B1(n20884), .B2(keyinput100), .C1(n20770), .C2(
        keyinput90), .A(n20769), .ZN(n20777) );
  AOI22_X1 U23685 ( .A1(n10522), .A2(keyinput124), .B1(keyinput101), .B2(
        n20772), .ZN(n20771) );
  OAI221_X1 U23686 ( .B1(n10522), .B2(keyinput124), .C1(n20772), .C2(
        keyinput101), .A(n20771), .ZN(n20776) );
  INV_X1 U23687 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20774) );
  AOI22_X1 U23688 ( .A1(n20774), .A2(keyinput108), .B1(n20871), .B2(keyinput71), .ZN(n20773) );
  OAI221_X1 U23689 ( .B1(n20774), .B2(keyinput108), .C1(n20871), .C2(
        keyinput71), .A(n20773), .ZN(n20775) );
  NOR4_X1 U23690 ( .A1(n20778), .A2(n20777), .A3(n20776), .A4(n20775), .ZN(
        n20792) );
  INV_X1 U23691 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20868) );
  AOI22_X1 U23692 ( .A1(n20780), .A2(keyinput81), .B1(keyinput107), .B2(n20868), .ZN(n20779) );
  OAI221_X1 U23693 ( .B1(n20780), .B2(keyinput81), .C1(n20868), .C2(
        keyinput107), .A(n20779), .ZN(n20790) );
  AOI22_X1 U23694 ( .A1(n20782), .A2(keyinput113), .B1(n20886), .B2(keyinput66), .ZN(n20781) );
  OAI221_X1 U23695 ( .B1(n20782), .B2(keyinput113), .C1(n20886), .C2(
        keyinput66), .A(n20781), .ZN(n20789) );
  INV_X1 U23696 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20784) );
  AOI22_X1 U23697 ( .A1(n20784), .A2(keyinput70), .B1(keyinput82), .B2(n20889), 
        .ZN(n20783) );
  OAI221_X1 U23698 ( .B1(n20784), .B2(keyinput70), .C1(n20889), .C2(keyinput82), .A(n20783), .ZN(n20788) );
  INV_X1 U23699 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20786) );
  INV_X1 U23700 ( .A(DATAI_22_), .ZN(n20891) );
  AOI22_X1 U23701 ( .A1(n20786), .A2(keyinput92), .B1(keyinput109), .B2(n20891), .ZN(n20785) );
  OAI221_X1 U23702 ( .B1(n20786), .B2(keyinput92), .C1(n20891), .C2(
        keyinput109), .A(n20785), .ZN(n20787) );
  NOR4_X1 U23703 ( .A1(n20790), .A2(n20789), .A3(n20788), .A4(n20787), .ZN(
        n20791) );
  AND4_X1 U23704 ( .A1(n20794), .A2(n20793), .A3(n20792), .A4(n20791), .ZN(
        n20932) );
  OAI22_X1 U23705 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(keyinput72), .B1(
        keyinput75), .B2(P3_LWORD_REG_15__SCAN_IN), .ZN(n20795) );
  AOI221_X1 U23706 ( .B1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput72), 
        .C1(P3_LWORD_REG_15__SCAN_IN), .C2(keyinput75), .A(n20795), .ZN(n20802) );
  OAI22_X1 U23707 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(keyinput102), 
        .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput74), .ZN(n20796)
         );
  AOI221_X1 U23708 ( .B1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput102), 
        .C1(keyinput74), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n20796), 
        .ZN(n20801) );
  OAI22_X1 U23709 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput116), .B1(
        keyinput119), .B2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20797) );
  AOI221_X1 U23710 ( .B1(P1_EAX_REG_22__SCAN_IN), .B2(keyinput116), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(keyinput119), .A(n20797), .ZN(
        n20800) );
  OAI22_X1 U23711 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput80), 
        .B1(keyinput84), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20798) );
  AOI221_X1 U23712 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput80), 
        .C1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .C2(keyinput84), .A(n20798), 
        .ZN(n20799) );
  NAND4_X1 U23713 ( .A1(n20802), .A2(n20801), .A3(n20800), .A4(n20799), .ZN(
        n20830) );
  OAI22_X1 U23714 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(keyinput88), 
        .B1(keyinput85), .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n20803) );
  AOI221_X1 U23715 ( .B1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput88), 
        .C1(P1_DATAO_REG_20__SCAN_IN), .C2(keyinput85), .A(n20803), .ZN(n20810) );
  OAI22_X1 U23716 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput98), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(keyinput125), .ZN(n20804) );
  AOI221_X1 U23717 ( .B1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput98), 
        .C1(keyinput125), .C2(P3_UWORD_REG_10__SCAN_IN), .A(n20804), .ZN(
        n20809) );
  OAI22_X1 U23718 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(keyinput86), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(keyinput97), .ZN(n20805) );
  AOI221_X1 U23719 ( .B1(P2_EAX_REG_21__SCAN_IN), .B2(keyinput86), .C1(
        keyinput97), .C2(P1_EBX_REG_29__SCAN_IN), .A(n20805), .ZN(n20808) );
  OAI22_X1 U23720 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(keyinput65), .B1(
        P3_W_R_N_REG_SCAN_IN), .B2(keyinput118), .ZN(n20806) );
  AOI221_X1 U23721 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(keyinput65), .C1(
        keyinput118), .C2(P3_W_R_N_REG_SCAN_IN), .A(n20806), .ZN(n20807) );
  NAND4_X1 U23722 ( .A1(n20810), .A2(n20809), .A3(n20808), .A4(n20807), .ZN(
        n20829) );
  OAI22_X1 U23723 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput111), 
        .B1(keyinput77), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20811) );
  AOI221_X1 U23724 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput111), 
        .C1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .C2(keyinput77), .A(n20811), .ZN(
        n20818) );
  OAI22_X1 U23725 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(keyinput117), .B1(
        keyinput67), .B2(P3_BE_N_REG_3__SCAN_IN), .ZN(n20812) );
  AOI221_X1 U23726 ( .B1(P2_LWORD_REG_3__SCAN_IN), .B2(keyinput117), .C1(
        P3_BE_N_REG_3__SCAN_IN), .C2(keyinput67), .A(n20812), .ZN(n20817) );
  OAI22_X1 U23727 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(keyinput103), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(keyinput106), .ZN(n20813) );
  AOI221_X1 U23728 ( .B1(P2_ADDRESS_REG_2__SCAN_IN), .B2(keyinput103), .C1(
        keyinput106), .C2(P3_ADDRESS_REG_20__SCAN_IN), .A(n20813), .ZN(n20816)
         );
  OAI22_X1 U23729 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(keyinput78), .B1(
        keyinput89), .B2(P3_EAX_REG_29__SCAN_IN), .ZN(n20814) );
  AOI221_X1 U23730 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(keyinput78), .C1(
        P3_EAX_REG_29__SCAN_IN), .C2(keyinput89), .A(n20814), .ZN(n20815) );
  NAND4_X1 U23731 ( .A1(n20818), .A2(n20817), .A3(n20816), .A4(n20815), .ZN(
        n20828) );
  OAI22_X1 U23732 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput105), 
        .B1(P3_DATAO_REG_23__SCAN_IN), .B2(keyinput79), .ZN(n20819) );
  AOI221_X1 U23733 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput105), 
        .C1(keyinput79), .C2(P3_DATAO_REG_23__SCAN_IN), .A(n20819), .ZN(n20826) );
  OAI22_X1 U23734 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(keyinput114), 
        .B1(P1_UWORD_REG_6__SCAN_IN), .B2(keyinput94), .ZN(n20820) );
  AOI221_X1 U23735 ( .B1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(keyinput114), 
        .C1(keyinput94), .C2(P1_UWORD_REG_6__SCAN_IN), .A(n20820), .ZN(n20825)
         );
  OAI22_X1 U23736 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(keyinput87), .B1(
        keyinput115), .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20821) );
  AOI221_X1 U23737 ( .B1(P1_ADDRESS_REG_18__SCAN_IN), .B2(keyinput87), .C1(
        P1_DATAO_REG_15__SCAN_IN), .C2(keyinput115), .A(n20821), .ZN(n20824)
         );
  OAI22_X1 U23738 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(keyinput127), .B1(
        keyinput91), .B2(BUF2_REG_26__SCAN_IN), .ZN(n20822) );
  AOI221_X1 U23739 ( .B1(P2_REIP_REG_11__SCAN_IN), .B2(keyinput127), .C1(
        BUF2_REG_26__SCAN_IN), .C2(keyinput91), .A(n20822), .ZN(n20823) );
  NAND4_X1 U23740 ( .A1(n20826), .A2(n20825), .A3(n20824), .A4(n20823), .ZN(
        n20827) );
  NOR4_X1 U23741 ( .A1(n20830), .A2(n20829), .A3(n20828), .A4(n20827), .ZN(
        n20931) );
  AOI22_X1 U23742 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(keyinput24), 
        .B1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput34), .ZN(n20831) );
  OAI221_X1 U23743 ( .B1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput24), 
        .C1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .C2(keyinput34), .A(n20831), .ZN(
        n20838) );
  AOI22_X1 U23744 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(keyinput14), .B1(
        P2_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput6), .ZN(n20832) );
  OAI221_X1 U23745 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(keyinput14), .C1(
        P2_INSTQUEUE_REG_9__2__SCAN_IN), .C2(keyinput6), .A(n20832), .ZN(
        n20837) );
  AOI22_X1 U23746 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput12), .B1(
        P1_INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput28), .ZN(n20833) );
  OAI221_X1 U23747 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput12), .C1(
        P1_INSTQUEUE_REG_2__0__SCAN_IN), .C2(keyinput28), .A(n20833), .ZN(
        n20836) );
  AOI22_X1 U23748 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(keyinput54), .B1(
        P3_EBX_REG_27__SCAN_IN), .B2(keyinput1), .ZN(n20834) );
  OAI221_X1 U23749 ( .B1(P3_W_R_N_REG_SCAN_IN), .B2(keyinput54), .C1(
        P3_EBX_REG_27__SCAN_IN), .C2(keyinput1), .A(n20834), .ZN(n20835) );
  NOR4_X1 U23750 ( .A1(n20838), .A2(n20837), .A3(n20836), .A4(n20835), .ZN(
        n20866) );
  AOI22_X1 U23751 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput49), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput17), .ZN(n20839) );
  OAI221_X1 U23752 ( .B1(P2_DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput49), .C1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput17), .A(n20839), .ZN(
        n20846) );
  AOI22_X1 U23753 ( .A1(P3_LWORD_REG_15__SCAN_IN), .A2(keyinput11), .B1(
        BUF2_REG_26__SCAN_IN), .B2(keyinput27), .ZN(n20840) );
  OAI221_X1 U23754 ( .B1(P3_LWORD_REG_15__SCAN_IN), .B2(keyinput11), .C1(
        BUF2_REG_26__SCAN_IN), .C2(keyinput27), .A(n20840), .ZN(n20845) );
  AOI22_X1 U23755 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(keyinput39), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(keyinput22), .ZN(n20841) );
  OAI221_X1 U23756 ( .B1(P2_ADDRESS_REG_2__SCAN_IN), .B2(keyinput39), .C1(
        P2_EAX_REG_21__SCAN_IN), .C2(keyinput22), .A(n20841), .ZN(n20844) );
  AOI22_X1 U23757 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput26), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(keyinput63), .ZN(n20842) );
  OAI221_X1 U23758 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput26), .C1(
        P2_REIP_REG_11__SCAN_IN), .C2(keyinput63), .A(n20842), .ZN(n20843) );
  NOR4_X1 U23759 ( .A1(n20846), .A2(n20845), .A3(n20844), .A4(n20843), .ZN(
        n20865) );
  AOI22_X1 U23760 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(keyinput21), .B1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput41), .ZN(n20847) );
  OAI221_X1 U23761 ( .B1(P1_DATAO_REG_20__SCAN_IN), .B2(keyinput21), .C1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput41), .A(n20847), .ZN(
        n20854) );
  AOI22_X1 U23762 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(keyinput30), .B1(
        P3_INSTQUEUE_REG_11__0__SCAN_IN), .B2(keyinput44), .ZN(n20848) );
  OAI221_X1 U23763 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(keyinput30), .C1(
        P3_INSTQUEUE_REG_11__0__SCAN_IN), .C2(keyinput44), .A(n20848), .ZN(
        n20853) );
  AOI22_X1 U23764 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(keyinput53), .B1(
        BUF1_REG_27__SCAN_IN), .B2(keyinput0), .ZN(n20849) );
  OAI221_X1 U23765 ( .B1(P2_LWORD_REG_3__SCAN_IN), .B2(keyinput53), .C1(
        BUF1_REG_27__SCAN_IN), .C2(keyinput0), .A(n20849), .ZN(n20852) );
  AOI22_X1 U23766 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput51), .B1(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput37), .ZN(n20850) );
  OAI221_X1 U23767 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput51), .C1(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .C2(keyinput37), .A(n20850), .ZN(
        n20851) );
  NOR4_X1 U23768 ( .A1(n20854), .A2(n20853), .A3(n20852), .A4(n20851), .ZN(
        n20864) );
  AOI22_X1 U23769 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput57), .B1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(keyinput50), .ZN(n20855) );
  OAI221_X1 U23770 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput57), .C1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .C2(keyinput50), .A(n20855), .ZN(
        n20862) );
  AOI22_X1 U23771 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput40), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput47), .ZN(n20856) );
  OAI221_X1 U23772 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput40), .C1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(keyinput47), .A(n20856), .ZN(
        n20861) );
  AOI22_X1 U23773 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(keyinput23), .B1(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput10), .ZN(n20857) );
  OAI221_X1 U23774 ( .B1(P1_ADDRESS_REG_18__SCAN_IN), .B2(keyinput23), .C1(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(keyinput10), .A(n20857), .ZN(
        n20860) );
  AOI22_X1 U23775 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(keyinput9), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(keyinput33), .ZN(n20858) );
  OAI221_X1 U23776 ( .B1(P1_ADDRESS_REG_2__SCAN_IN), .B2(keyinput9), .C1(
        P1_EBX_REG_29__SCAN_IN), .C2(keyinput33), .A(n20858), .ZN(n20859) );
  NOR4_X1 U23777 ( .A1(n20862), .A2(n20861), .A3(n20860), .A4(n20859), .ZN(
        n20863) );
  NAND4_X1 U23778 ( .A1(n20866), .A2(n20865), .A3(n20864), .A4(n20863), .ZN(
        n20930) );
  AOI22_X1 U23779 ( .A1(n20869), .A2(keyinput20), .B1(n20868), .B2(keyinput43), 
        .ZN(n20867) );
  OAI221_X1 U23780 ( .B1(n20869), .B2(keyinput20), .C1(n20868), .C2(keyinput43), .A(n20867), .ZN(n20881) );
  AOI22_X1 U23781 ( .A1(n20872), .A2(keyinput35), .B1(n20871), .B2(keyinput7), 
        .ZN(n20870) );
  OAI221_X1 U23782 ( .B1(n20872), .B2(keyinput35), .C1(n20871), .C2(keyinput7), 
        .A(n20870), .ZN(n20880) );
  INV_X1 U23783 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U23784 ( .A1(n20874), .A2(keyinput38), .B1(n12880), .B2(keyinput8), 
        .ZN(n20873) );
  OAI221_X1 U23785 ( .B1(n20874), .B2(keyinput38), .C1(n12880), .C2(keyinput8), 
        .A(n20873), .ZN(n20879) );
  INV_X1 U23786 ( .A(P3_UWORD_REG_10__SCAN_IN), .ZN(n20875) );
  XOR2_X1 U23787 ( .A(keyinput61), .B(n20875), .Z(n20877) );
  XNOR2_X1 U23788 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B(keyinput56), .ZN(
        n20876) );
  NAND2_X1 U23789 ( .A1(n20877), .A2(n20876), .ZN(n20878) );
  NOR4_X1 U23790 ( .A1(n20881), .A2(n20880), .A3(n20879), .A4(n20878), .ZN(
        n20928) );
  AOI22_X1 U23791 ( .A1(n20884), .A2(keyinput36), .B1(n20883), .B2(keyinput4), 
        .ZN(n20882) );
  OAI221_X1 U23792 ( .B1(n20884), .B2(keyinput36), .C1(n20883), .C2(keyinput4), 
        .A(n20882), .ZN(n20895) );
  AOI22_X1 U23793 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput46), 
        .B1(n20886), .B2(keyinput2), .ZN(n20885) );
  OAI221_X1 U23794 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput46), 
        .C1(n20886), .C2(keyinput2), .A(n20885), .ZN(n20894) );
  AOI22_X1 U23795 ( .A1(n20889), .A2(keyinput18), .B1(keyinput32), .B2(n20888), 
        .ZN(n20887) );
  OAI221_X1 U23796 ( .B1(n20889), .B2(keyinput18), .C1(n20888), .C2(keyinput32), .A(n20887), .ZN(n20893) );
  AOI22_X1 U23797 ( .A1(n20891), .A2(keyinput45), .B1(n14534), .B2(keyinput52), 
        .ZN(n20890) );
  OAI221_X1 U23798 ( .B1(n20891), .B2(keyinput45), .C1(n14534), .C2(keyinput52), .A(n20890), .ZN(n20892) );
  NOR4_X1 U23799 ( .A1(n20895), .A2(n20894), .A3(n20893), .A4(n20892), .ZN(
        n20927) );
  AOI22_X1 U23800 ( .A1(n20898), .A2(keyinput29), .B1(n20897), .B2(keyinput58), 
        .ZN(n20896) );
  OAI221_X1 U23801 ( .B1(n20898), .B2(keyinput29), .C1(n20897), .C2(keyinput58), .A(n20896), .ZN(n20910) );
  AOI22_X1 U23802 ( .A1(n20901), .A2(keyinput19), .B1(keyinput42), .B2(n20900), 
        .ZN(n20899) );
  OAI221_X1 U23803 ( .B1(n20901), .B2(keyinput19), .C1(n20900), .C2(keyinput42), .A(n20899), .ZN(n20909) );
  INV_X1 U23804 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n20903) );
  AOI22_X1 U23805 ( .A1(n20903), .A2(keyinput15), .B1(n10522), .B2(keyinput60), 
        .ZN(n20902) );
  OAI221_X1 U23806 ( .B1(n20903), .B2(keyinput15), .C1(n10522), .C2(keyinput60), .A(n20902), .ZN(n20908) );
  AOI22_X1 U23807 ( .A1(n20906), .A2(keyinput62), .B1(keyinput25), .B2(n20905), 
        .ZN(n20904) );
  OAI221_X1 U23808 ( .B1(n20906), .B2(keyinput62), .C1(n20905), .C2(keyinput25), .A(n20904), .ZN(n20907) );
  NOR4_X1 U23809 ( .A1(n20910), .A2(n20909), .A3(n20908), .A4(n20907), .ZN(
        n20926) );
  AOI22_X1 U23810 ( .A1(n20913), .A2(keyinput5), .B1(keyinput55), .B2(n20912), 
        .ZN(n20911) );
  OAI221_X1 U23811 ( .B1(n20913), .B2(keyinput5), .C1(n20912), .C2(keyinput55), 
        .A(n20911), .ZN(n20924) );
  INV_X1 U23812 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20916) );
  AOI22_X1 U23813 ( .A1(n20916), .A2(keyinput13), .B1(keyinput31), .B2(n20915), 
        .ZN(n20914) );
  OAI221_X1 U23814 ( .B1(n20916), .B2(keyinput13), .C1(n20915), .C2(keyinput31), .A(n20914), .ZN(n20923) );
  XNOR2_X1 U23815 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B(keyinput59), .ZN(
        n20919) );
  XNOR2_X1 U23816 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B(keyinput48), .ZN(
        n20918) );
  XNOR2_X1 U23817 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B(keyinput16), 
        .ZN(n20917) );
  NAND3_X1 U23818 ( .A1(n20919), .A2(n20918), .A3(n20917), .ZN(n20922) );
  XNOR2_X1 U23819 ( .A(n20920), .B(keyinput3), .ZN(n20921) );
  NOR4_X1 U23820 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n20925) );
  NAND4_X1 U23821 ( .A1(n20928), .A2(n20927), .A3(n20926), .A4(n20925), .ZN(
        n20929) );
  AOI211_X1 U23822 ( .C1(n20932), .C2(n20931), .A(n20930), .B(n20929), .ZN(
        n20936) );
  AOI222_X1 U23823 ( .A1(n20745), .A2(P1_ADDRESS_REG_14__SCAN_IN), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20934), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20933), .ZN(n20935) );
  XNOR2_X1 U23824 ( .A(n20936), .B(n20935), .ZN(P1_U3211) );
  NAND2_X2 U11483 ( .A1(n10281), .A2(n10280), .ZN(n13763) );
  INV_X1 U14521 ( .A(n11548), .ZN(n20139) );
  BUF_X2 U11095 ( .A(n15355), .Z(n17109) );
  CLKBUF_X1 U11154 ( .A(n11643), .Z(n11699) );
  OAI21_X1 U11246 ( .B1(n10353), .B2(n10352), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10354) );
  CLKBUF_X2 U11406 ( .A(n15482), .Z(n17099) );
  CLKBUF_X1 U12302 ( .A(n12063), .Z(n14438) );
  CLKBUF_X2 U12337 ( .A(n14285), .Z(n14295) );
  CLKBUF_X1 U12860 ( .A(n17486), .Z(n17493) );
  CLKBUF_X1 U13217 ( .A(n16496), .Z(n16507) );
endmodule

