

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987;

  NAND2_X1 U3545 ( .A1(n6010), .A2(n5442), .ZN(n5441) );
  CLKBUF_X1 U3546 ( .A(n3704), .Z(n3112) );
  CLKBUF_X2 U3547 ( .A(n3740), .Z(n3837) );
  NAND2_X2 U3548 ( .A1(n4637), .A2(n3111), .ZN(n3750) );
  CLKBUF_X2 U3549 ( .A(n3286), .Z(n4522) );
  CLKBUF_X2 U3550 ( .A(n3303), .Z(n4368) );
  CLKBUF_X2 U3551 ( .A(n3421), .Z(n4361) );
  CLKBUF_X2 U3552 ( .A(n3448), .Z(n3412) );
  CLKBUF_X2 U3553 ( .A(n3285), .Z(n4370) );
  CLKBUF_X2 U3554 ( .A(n3292), .Z(n4187) );
  CLKBUF_X2 U3555 ( .A(n3420), .Z(n4311) );
  CLKBUF_X2 U3556 ( .A(n3387), .Z(n4360) );
  CLKBUF_X2 U3557 ( .A(n3388), .Z(n4369) );
  CLKBUF_X2 U3558 ( .A(n4345), .Z(n4367) );
  CLKBUF_X1 U3559 ( .A(n3317), .Z(n3719) );
  AND4_X1 U3560 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3283)
         );
  AND4_X1 U3561 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3282)
         );
  AND4_X1 U3562 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3281)
         );
  CLKBUF_X2 U3563 ( .A(n3263), .Z(n3736) );
  AND4_X1 U3564 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3310)
         );
  AND4_X1 U3565 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3235)
         );
  AND2_X2 U3566 ( .A1(n4524), .A2(n3165), .ZN(n3387) );
  OR2_X1 U3567 ( .A1(n3735), .A2(n3316), .ZN(n3152) );
  AND2_X1 U3568 ( .A1(n3314), .A2(n4452), .ZN(n3371) );
  AND4_X1 U3569 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n3233)
         );
  AND4_X1 U3570 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3309)
         );
  AND2_X1 U3571 ( .A1(n3704), .A2(n3111), .ZN(n4399) );
  NAND2_X1 U3572 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5204), .ZN(n4938) );
  INV_X1 U3573 ( .A(n3734), .ZN(n4632) );
  NOR2_X1 U3574 ( .A1(n5401), .A2(n5314), .ZN(n5950) );
  INV_X1 U3575 ( .A(n4563), .ZN(n6325) );
  INV_X1 U3576 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6656) );
  INV_X1 U3577 ( .A(n6099), .ZN(n6149) );
  NAND2_X2 U3578 ( .A1(n3367), .A2(n3325), .ZN(n3340) );
  NOR2_X4 U3579 ( .A1(n5497), .A2(n5496), .ZN(n5495) );
  BUF_X1 U3580 ( .A(n3336), .Z(n3900) );
  INV_X2 U3581 ( .A(n4940), .ZN(n5336) );
  AND2_X2 U3582 ( .A1(n3174), .A2(n4524), .ZN(n4345) );
  NOR2_X2 U3583 ( .A1(n6590), .A2(n5445), .ZN(n6070) );
  NAND2_X2 U3584 ( .A1(n3629), .A2(n5698), .ZN(n5688) );
  INV_X1 U3585 ( .A(n5912), .ZN(n5541) );
  NOR2_X1 U3586 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  AND2_X1 U3587 ( .A1(n5455), .A2(n5454), .ZN(n5912) );
  AOI211_X1 U3588 ( .C1(n6258), .C2(n5595), .A(n5594), .B(n5593), .ZN(n5596)
         );
  NAND2_X1 U3589 ( .A1(n3142), .A2(n3119), .ZN(n5746) );
  CLKBUF_X1 U3590 ( .A(n5648), .Z(n5649) );
  NAND2_X1 U3591 ( .A1(n5668), .A2(n5667), .ZN(n5653) );
  AOI211_X1 U3592 ( .C1(n5322), .C2(n6312), .A(n3868), .B(n3867), .ZN(n3884)
         );
  NOR2_X1 U3593 ( .A1(n5367), .A2(n5462), .ZN(n3834) );
  XNOR2_X1 U3594 ( .A(n3622), .B(n5260), .ZN(n5165) );
  INV_X2 U3595 ( .A(n5652), .ZN(n5689) );
  INV_X2 U3597 ( .A(n3625), .ZN(n5652) );
  NAND2_X1 U3598 ( .A1(n3614), .A2(n3617), .ZN(n3625) );
  XNOR2_X1 U3599 ( .A(n3614), .B(n3604), .ZN(n3901) );
  NAND2_X1 U3600 ( .A1(n3595), .A2(n3572), .ZN(n3957) );
  CLKBUF_X1 U3601 ( .A(n4552), .Z(n4553) );
  XNOR2_X1 U3602 ( .A(n3406), .B(n3405), .ZN(n3502) );
  NAND2_X1 U3603 ( .A1(n3524), .A2(n3523), .ZN(n4656) );
  AND2_X2 U3604 ( .A1(n5184), .A2(n3771), .ZN(n5185) );
  NAND2_X1 U3605 ( .A1(n5858), .A2(n6660), .ZN(n3524) );
  NAND2_X1 U3606 ( .A1(n3385), .A2(n3384), .ZN(n4545) );
  AOI21_X1 U3607 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6660), .A(n3698), 
        .ZN(n3699) );
  AOI21_X1 U3608 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3697) );
  INV_X1 U3609 ( .A(n3460), .ZN(n3486) );
  AND2_X1 U3610 ( .A1(n3334), .A2(n3333), .ZN(n3704) );
  NOR2_X1 U3611 ( .A1(n3339), .A2(n3338), .ZN(n3341) );
  BUF_X2 U3612 ( .A(n3366), .Z(n6658) );
  INV_X1 U3613 ( .A(n3679), .ZN(n3695) );
  INV_X1 U3614 ( .A(n3740), .ZN(n3313) );
  INV_X1 U3615 ( .A(n3618), .ZN(n3603) );
  NAND2_X1 U3616 ( .A1(n4632), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3509) );
  OR2_X1 U3617 ( .A1(n3736), .A2(n6660), .ZN(n3510) );
  AND2_X1 U3618 ( .A1(n3323), .A2(n3337), .ZN(n3264) );
  AND2_X2 U3619 ( .A1(n3337), .A2(n3900), .ZN(n3345) );
  OR2_X1 U3620 ( .A1(n3432), .A2(n3431), .ZN(n3618) );
  NOR2_X1 U3621 ( .A1(n3163), .A2(n3162), .ZN(n3183) );
  AND3_X2 U3622 ( .A1(n3262), .A2(n3261), .A3(n3151), .ZN(n3342) );
  AND4_X1 U3623 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3180)
         );
  AND4_X1 U3624 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3261)
         );
  AND4_X1 U3625 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3181)
         );
  AND4_X1 U3626 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n3182)
         );
  AND4_X1 U3627 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3216)
         );
  AND4_X1 U3628 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3236)
         );
  INV_X2 U3629 ( .A(n3395), .ZN(n4359) );
  AND4_X1 U3630 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3234)
         );
  AND4_X1 U3631 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  AND4_X1 U3632 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3214)
         );
  NOR2_X1 U3633 ( .A1(n3389), .A2(n3199), .ZN(n3204) );
  INV_X2 U3634 ( .A(n6667), .ZN(n6651) );
  INV_X1 U3635 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6552) );
  INV_X2 U3636 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U3637 ( .A1(n3754), .A2(n3753), .ZN(n4491) );
  NAND2_X1 U3639 ( .A1(n5489), .A2(n5488), .ZN(n5385) );
  OR2_X2 U3640 ( .A1(n5629), .A2(n5630), .ZN(n5600) );
  AND2_X2 U3641 ( .A1(n5430), .A2(n3794), .ZN(n3154) );
  AND2_X2 U3643 ( .A1(n4485), .A2(n4486), .ZN(n4487) );
  OR2_X4 U3644 ( .A1(n5456), .A2(n5457), .ZN(n5459) );
  OR2_X2 U3645 ( .A1(n3835), .A2(EBX_REG_1__SCAN_IN), .ZN(n3745) );
  OR2_X2 U3646 ( .A1(n3442), .A2(n3441), .ZN(n3443) );
  NAND2_X2 U3647 ( .A1(n5438), .A2(n3129), .ZN(n5412) );
  NOR2_X4 U3648 ( .A1(n5412), .A2(n5415), .ZN(n5413) );
  NOR3_X2 U3649 ( .A1(n5504), .A2(n3806), .A3(n3805), .ZN(n3807) );
  NAND2_X4 U3650 ( .A1(n3444), .A2(n3443), .ZN(n3911) );
  AND2_X4 U3651 ( .A1(n3488), .A2(n3487), .ZN(n4563) );
  NAND2_X1 U3652 ( .A1(n3103), .A2(n3579), .ZN(n3098) );
  NAND2_X1 U3653 ( .A1(n3637), .A2(n3102), .ZN(n3099) );
  AND2_X2 U3654 ( .A1(n3099), .A2(n3100), .ZN(n5661) );
  OR2_X1 U3655 ( .A1(n3101), .A2(n5667), .ZN(n3100) );
  INV_X1 U3656 ( .A(n3638), .ZN(n3101) );
  AND2_X1 U3657 ( .A1(n3636), .A2(n3638), .ZN(n3102) );
  NAND2_X1 U3658 ( .A1(n4694), .A2(n4695), .ZN(n3103) );
  NAND2_X1 U3659 ( .A1(n5688), .A2(n3107), .ZN(n3104) );
  AND2_X2 U3660 ( .A1(n3104), .A2(n3105), .ZN(n5674) );
  OR2_X1 U3661 ( .A1(n3106), .A2(n3117), .ZN(n3105) );
  INV_X1 U3662 ( .A(n3634), .ZN(n3106) );
  AND2_X1 U3663 ( .A1(n3630), .A2(n3634), .ZN(n3107) );
  NAND3_X1 U3665 ( .A1(n3350), .A2(n3349), .A3(n3351), .ZN(n3109) );
  NAND2_X1 U3666 ( .A1(n3580), .A2(n3579), .ZN(n4876) );
  XNOR2_X2 U3667 ( .A(n3578), .B(n3863), .ZN(n4695) );
  NAND3_X1 U3668 ( .A1(n3350), .A2(n3349), .A3(n3351), .ZN(n3375) );
  OAI211_X1 U3669 ( .C1(n3957), .C2(n4084), .A(n3956), .B(n3955), .ZN(n4514)
         );
  INV_X2 U3670 ( .A(n3336), .ZN(n4622) );
  NOR2_X2 U3671 ( .A1(n4513), .A2(n4761), .ZN(n4762) );
  NAND2_X2 U3672 ( .A1(n3725), .A2(n3344), .ZN(n3737) );
  BUF_X1 U3673 ( .A(n5326), .Z(n5348) );
  AOI22_X2 U3674 ( .A1(n5640), .A2(n5598), .B1(n5652), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5636) );
  NAND2_X2 U3675 ( .A1(n5613), .A2(n3641), .ZN(n5640) );
  NOR2_X4 U3676 ( .A1(n3111), .A2(n3735), .ZN(n3344) );
  AND2_X1 U3678 ( .A1(n3174), .A2(n4524), .ZN(n3110) );
  BUF_X4 U3679 ( .A(n3315), .Z(n3735) );
  NAND3_X2 U3680 ( .A1(n3331), .A2(n3330), .A3(n3329), .ZN(n3376) );
  AND2_X2 U3681 ( .A1(n3174), .A2(n4540), .ZN(n3426) );
  AND2_X2 U3682 ( .A1(n3174), .A2(n4523), .ZN(n3420) );
  NAND2_X1 U3683 ( .A1(n3545), .A2(n3544), .ZN(n3571) );
  NAND2_X2 U3684 ( .A1(n3554), .A2(n3553), .ZN(n4694) );
  NAND2_X2 U3685 ( .A1(n3386), .A2(n4545), .ZN(n4451) );
  XNOR2_X1 U3686 ( .A(n3502), .B(n3501), .ZN(n4558) );
  AND2_X2 U3687 ( .A1(n5362), .A2(n5365), .ZN(n5363) );
  NOR2_X2 U3688 ( .A1(n5385), .A2(n3133), .ZN(n5362) );
  AND2_X1 U3689 ( .A1(n3383), .A2(n3109), .ZN(n3385) );
  NAND2_X2 U3690 ( .A1(n3375), .A2(n3355), .ZN(n3407) );
  OAI21_X1 U3691 ( .B1(n4602), .B2(n4084), .A(n3940), .ZN(n4486) );
  AND2_X2 U3692 ( .A1(n3341), .A2(n3340), .ZN(n3725) );
  NAND2_X1 U3693 ( .A1(n3313), .A2(n3359), .ZN(n4452) );
  NOR2_X2 U3694 ( .A1(n5120), .A2(n5243), .ZN(n5219) );
  NAND2_X2 U3695 ( .A1(n3547), .A2(n3527), .ZN(n4602) );
  OAI22_X2 U3696 ( .A1(n5636), .A2(n5635), .B1(n5601), .B2(n5599), .ZN(n5629)
         );
  NOR2_X4 U3697 ( .A1(n5270), .A2(n5560), .ZN(n5438) );
  XNOR2_X2 U3698 ( .A(n5350), .B(n5292), .ZN(n5301) );
  AND2_X2 U3699 ( .A1(n5349), .A2(n4358), .ZN(n5350) );
  AND2_X1 U3700 ( .A1(n5586), .A2(n3115), .ZN(n5564) );
  AND2_X1 U3701 ( .A1(n5839), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U3702 ( .A1(n3471), .A2(n3315), .ZN(n3740) );
  NAND2_X2 U3703 ( .A1(n3664), .A2(n3736), .ZN(n3679) );
  AND3_X1 U3704 ( .A1(n5829), .A2(n6541), .A3(n6543), .ZN(n4932) );
  AND2_X1 U3705 ( .A1(n5601), .A2(n5751), .ZN(n3649) );
  AND2_X1 U3706 ( .A1(n6168), .A2(n3345), .ZN(n6160) );
  AND2_X1 U3707 ( .A1(n6168), .A2(n4587), .ZN(n6164) );
  CLKBUF_X1 U3708 ( .A(n3559), .Z(n4366) );
  AND3_X1 U3709 ( .A1(n3435), .A2(n3445), .A3(n3434), .ZN(n3437) );
  AND2_X2 U3710 ( .A1(n4525), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3174)
         );
  INV_X1 U3711 ( .A(n3710), .ZN(n3671) );
  OAI22_X1 U3712 ( .A1(n3700), .A2(n3592), .B1(n3679), .B2(n3591), .ZN(n3593)
         );
  AOI21_X1 U3713 ( .B1(n3506), .B2(n5006), .A(n3348), .ZN(n3351) );
  AND2_X1 U3714 ( .A1(n3505), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3348)
         );
  AND2_X1 U3715 ( .A1(n4410), .A2(n3337), .ZN(n3240) );
  AOI21_X1 U3716 ( .B1(n3361), .B2(n3344), .A(n3360), .ZN(n3859) );
  CLKBUF_X1 U3717 ( .A(n3358), .Z(n3361) );
  AND2_X1 U3718 ( .A1(n5427), .A2(n5440), .ZN(n3131) );
  AND2_X1 U3719 ( .A1(n3977), .A2(n3123), .ZN(n3143) );
  INV_X1 U3720 ( .A(n4925), .ZN(n3144) );
  OAI22_X1 U3721 ( .A1(n3700), .A2(n3603), .B1(n3602), .B2(n3679), .ZN(n3604)
         );
  INV_X1 U3722 ( .A(n3925), .ZN(n4391) );
  NOR2_X1 U3723 ( .A1(n3900), .A2(n6656), .ZN(n4065) );
  NAND2_X1 U3724 ( .A1(n5487), .A2(n5388), .ZN(n5377) );
  INV_X1 U3725 ( .A(n3342), .ZN(n3855) );
  NAND4_X1 U3726 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3263)
         );
  NAND2_X1 U3727 ( .A1(n3374), .A2(n3444), .ZN(n3384) );
  AND2_X1 U3728 ( .A1(n3734), .A2(n4616), .ZN(n3366) );
  AND3_X1 U3729 ( .A1(n3752), .A2(n3818), .A3(n3751), .ZN(n4475) );
  AND2_X1 U3730 ( .A1(n3748), .A2(n3747), .ZN(n4430) );
  AOI21_X1 U3731 ( .B1(n4390), .B2(n4389), .A(n4388), .ZN(n5292) );
  INV_X1 U3732 ( .A(n5351), .ZN(n4358) );
  OR2_X1 U3733 ( .A1(n3134), .A2(n5479), .ZN(n3133) );
  AND2_X1 U3734 ( .A1(n4202), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4229)
         );
  NOR2_X1 U3735 ( .A1(n5503), .A2(n3128), .ZN(n3126) );
  NAND2_X1 U3736 ( .A1(n4406), .A2(n3929), .ZN(n4494) );
  NAND2_X1 U3737 ( .A1(n3910), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U3738 ( .A1(n3750), .A2(n3837), .ZN(n5337) );
  NOR2_X1 U3739 ( .A1(n5746), .A2(n3645), .ZN(n5748) );
  OAI21_X1 U3740 ( .B1(n3911), .B2(STATE2_REG_0__SCAN_IN), .A(n3486), .ZN(
        n3464) );
  INV_X1 U3741 ( .A(n3315), .ZN(n4616) );
  INV_X1 U3742 ( .A(n4401), .ZN(n4402) );
  INV_X1 U3743 ( .A(n6167), .ZN(n5561) );
  OAI211_X2 U3744 ( .C1(n6034), .C2(n4585), .A(n6251), .B(n4584), .ZN(n6168)
         );
  NAND2_X1 U3745 ( .A1(n6277), .A2(n3890), .ZN(n6266) );
  CLKBUF_X1 U3746 ( .A(n4558), .Z(n4559) );
  OR2_X1 U3747 ( .A1(n3590), .A2(n3589), .ZN(n3606) );
  OR2_X1 U3748 ( .A1(n3565), .A2(n3564), .ZN(n3575) );
  OR2_X1 U3749 ( .A1(n3543), .A2(n3542), .ZN(n3549) );
  OR2_X1 U3750 ( .A1(n3520), .A2(n3519), .ZN(n3529) );
  OR2_X1 U3751 ( .A1(n3418), .A2(n3417), .ZN(n3478) );
  AND2_X1 U3752 ( .A1(n3734), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3664) );
  NOR2_X1 U3753 ( .A1(n3402), .A2(n3401), .ZN(n3470) );
  AOI21_X1 U3754 ( .B1(n3297), .B2(INSTQUEUE_REG_1__3__SCAN_IN), .A(n3241), 
        .ZN(n3245) );
  AND2_X1 U3755 ( .A1(n3298), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U3756 ( .A1(n3421), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U3757 ( .A1(n3303), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U3758 ( .A1(n3672), .A2(n3671), .ZN(n3673) );
  NAND2_X1 U3759 ( .A1(n3690), .A2(n3689), .ZN(n3691) );
  NAND2_X1 U3760 ( .A1(n3683), .A2(n3682), .ZN(n3690) );
  OR3_X1 U3761 ( .A1(n3694), .A2(n6966), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n3713) );
  NAND2_X1 U3762 ( .A1(n4249), .A2(n3135), .ZN(n3134) );
  INV_X1 U3763 ( .A(n5386), .ZN(n3135) );
  INV_X1 U3764 ( .A(n4065), .ZN(n4084) );
  INV_X1 U3765 ( .A(n3140), .ZN(n3139) );
  OAI21_X1 U3766 ( .B1(n3120), .B2(n3141), .A(n3642), .ZN(n3140) );
  NAND2_X1 U3767 ( .A1(n4940), .A2(n3837), .ZN(n5331) );
  NAND2_X1 U3768 ( .A1(n4410), .A2(n3264), .ZN(n3722) );
  INV_X1 U3769 ( .A(n3345), .ZN(n3854) );
  XNOR2_X1 U3770 ( .A(n3475), .B(n3476), .ZN(n4552) );
  INV_X1 U3771 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4887) );
  INV_X1 U3772 ( .A(n4411), .ZN(n3505) );
  OAI21_X1 U3773 ( .B1(n3358), .B2(n3735), .A(n3327), .ZN(n3330) );
  AND2_X1 U3774 ( .A1(n3504), .A2(n4744), .ZN(n5007) );
  OAI21_X1 U3775 ( .B1(n4930), .B2(n6549), .A(n6539), .ZN(n4607) );
  NAND2_X1 U3776 ( .A1(n3695), .A2(n3688), .ZN(n3701) );
  NAND2_X1 U3777 ( .A1(n3661), .A2(n3660), .ZN(n3712) );
  OR2_X1 U3778 ( .A1(n3694), .A2(n3659), .ZN(n3661) );
  AND2_X1 U3779 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6966), .ZN(n3659)
         );
  AND2_X1 U3780 ( .A1(n4520), .A2(n4519), .ZN(n6511) );
  INV_X1 U3781 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6969) );
  NOR2_X2 U3782 ( .A1(n5317), .A2(n5316), .ZN(n5356) );
  NAND2_X1 U3783 ( .A1(n4017), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4021)
         );
  INV_X1 U3784 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5213) );
  AND4_X1 U3785 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n4533), .ZN(n3373)
         );
  XNOR2_X1 U3786 ( .A(n4393), .B(n4392), .ZN(n5326) );
  AOI22_X1 U3787 ( .A1(n3912), .A2(EAX_REG_31__SCAN_IN), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4392) );
  OR2_X1 U3788 ( .A1(n4331), .A2(n4330), .ZN(n4337) );
  INV_X1 U3789 ( .A(n5349), .ZN(n5455) );
  OR2_X1 U3790 ( .A1(n4306), .A2(n4305), .ZN(n4331) );
  AND2_X1 U3791 ( .A1(n5595), .A2(n4931), .ZN(n4287) );
  NOR2_X1 U3792 ( .A1(n4264), .A2(n3895), .ZN(n4286) );
  AND2_X1 U3793 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3894), .ZN(n4202)
         );
  AND2_X1 U3794 ( .A1(n4205), .A2(n4204), .ZN(n5488) );
  NAND2_X1 U3795 ( .A1(n4154), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4184)
         );
  AND2_X1 U3796 ( .A1(n4153), .A2(n4152), .ZN(n5397) );
  NOR2_X1 U3797 ( .A1(n4116), .A2(n5419), .ZN(n4133) );
  CLKBUF_X1 U3798 ( .A(n5413), .Z(n5414) );
  NOR2_X1 U3799 ( .A1(n5526), .A2(n3130), .ZN(n3129) );
  INV_X1 U3800 ( .A(n3131), .ZN(n3130) );
  OR2_X1 U3801 ( .A1(n5444), .A2(n4053), .ZN(n4068) );
  INV_X1 U3802 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6856) );
  NOR2_X1 U3803 ( .A1(n4068), .A2(n6856), .ZN(n4098) );
  NAND2_X1 U3804 ( .A1(n4038), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4053)
         );
  CLKBUF_X1 U3805 ( .A(n5270), .Z(n5271) );
  AND2_X1 U3806 ( .A1(n3992), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4017)
         );
  NOR2_X1 U3807 ( .A1(n5213), .A2(n3973), .ZN(n3988) );
  AND3_X1 U3808 ( .A1(n3976), .A2(n3975), .A3(n3974), .ZN(n5070) );
  NOR2_X1 U3809 ( .A1(n3958), .A2(n3893), .ZN(n3902) );
  INV_X1 U3810 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U3811 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3902), .ZN(n3973)
         );
  OAI21_X1 U3812 ( .B1(n4326), .B2(n3904), .A(n3903), .ZN(n3905) );
  AOI21_X1 U3813 ( .B1(n3962), .B2(n4065), .A(n3961), .ZN(n4761) );
  NAND2_X1 U3814 ( .A1(n3954), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3958)
         );
  AND2_X1 U3815 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3954)
         );
  NAND2_X1 U3816 ( .A1(n3953), .A2(n3952), .ZN(n4566) );
  CLKBUF_X1 U3817 ( .A(n4511), .Z(n4512) );
  NAND2_X1 U3818 ( .A1(n3931), .A2(n3930), .ZN(n3932) );
  NAND2_X1 U3819 ( .A1(n4428), .A2(n3918), .ZN(n4407) );
  NAND2_X1 U3820 ( .A1(n3917), .A2(n3916), .ZN(n4428) );
  INV_X1 U3821 ( .A(n4425), .ZN(n3916) );
  INV_X1 U3822 ( .A(n4426), .ZN(n3917) );
  CLKBUF_X1 U3823 ( .A(n5456), .Z(n5465) );
  CLKBUF_X1 U3824 ( .A(n5367), .Z(n5463) );
  NOR2_X2 U3825 ( .A1(n5377), .A2(n3828), .ZN(n5472) );
  CLKBUF_X1 U3826 ( .A(n5377), .Z(n5476) );
  NAND2_X1 U3827 ( .A1(n5648), .A2(n3120), .ZN(n5613) );
  INV_X1 U3828 ( .A(n5600), .ZN(n5628) );
  INV_X1 U3829 ( .A(n5682), .ZN(n3633) );
  AND2_X1 U3830 ( .A1(n5831), .A2(n3874), .ZN(n5818) );
  NAND2_X1 U3831 ( .A1(n3624), .A2(n3137), .ZN(n3136) );
  AND2_X1 U3832 ( .A1(n3769), .A2(n3768), .ZN(n5182) );
  AND3_X1 U3833 ( .A1(n3765), .A2(n3818), .A3(n3764), .ZN(n4770) );
  AND2_X1 U3834 ( .A1(n5839), .A2(n3853), .ZN(n6522) );
  NAND2_X1 U3835 ( .A1(n3763), .A2(n3762), .ZN(n4771) );
  INV_X1 U3836 ( .A(n4570), .ZN(n3763) );
  INV_X1 U3837 ( .A(n4475), .ZN(n3753) );
  INV_X1 U3838 ( .A(n4476), .ZN(n3754) );
  INV_X1 U3839 ( .A(n4697), .ZN(n5831) );
  NAND2_X1 U3840 ( .A1(n3731), .A2(n6544), .ZN(n3870) );
  NOR2_X1 U3841 ( .A1(n3367), .A2(n3318), .ZN(n5839) );
  NOR2_X1 U3842 ( .A1(n4602), .A2(n4559), .ZN(n6435) );
  INV_X1 U3843 ( .A(n4609), .ZN(n6322) );
  INV_X1 U3844 ( .A(n3719), .ZN(n3318) );
  INV_X1 U3845 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U3846 ( .A1(n6626), .A2(n4607), .ZN(n4648) );
  AND2_X1 U3847 ( .A1(n6552), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4411) );
  INV_X1 U3848 ( .A(n6118), .ZN(n6143) );
  INV_X1 U3849 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6084) );
  AND2_X1 U3850 ( .A1(n4940), .A2(n4939), .ZN(n6119) );
  AND2_X1 U3851 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4944), .ZN(n4939) );
  AND2_X1 U3852 ( .A1(n4950), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4933) );
  INV_X1 U3853 ( .A(n6097), .ZN(n6133) );
  AND2_X1 U3854 ( .A1(n5204), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6097) );
  AND2_X1 U3855 ( .A1(n5204), .A2(n4951), .ZN(n6099) );
  CLKBUF_X1 U3856 ( .A(n5535), .Z(n5528) );
  AND2_X1 U3857 ( .A1(n6156), .A2(n5327), .ZN(n6670) );
  NAND2_X2 U3858 ( .A1(n4417), .A2(n4416), .ZN(n6156) );
  OR2_X1 U3859 ( .A1(n6521), .A2(n4409), .ZN(n4417) );
  INV_X1 U3860 ( .A(n6670), .ZN(n5532) );
  INV_X1 U3861 ( .A(n5923), .ZN(n5544) );
  AND2_X1 U3862 ( .A1(n4589), .A2(n4588), .ZN(n6167) );
  AND2_X1 U3863 ( .A1(n4433), .A2(n6042), .ZN(n6188) );
  INV_X1 U3865 ( .A(n6189), .ZN(n6200) );
  INV_X1 U3866 ( .A(n6254), .ZN(n6249) );
  OR2_X1 U3867 ( .A1(n4431), .A2(n6536), .ZN(n6254) );
  INV_X1 U3868 ( .A(n5695), .ZN(n6262) );
  INV_X1 U3869 ( .A(n6272), .ZN(n6258) );
  XNOR2_X1 U3870 ( .A(n3887), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5713)
         );
  NAND2_X1 U3871 ( .A1(n3886), .A2(n3145), .ZN(n3887) );
  XNOR2_X1 U3872 ( .A(n5582), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5737)
         );
  NOR2_X1 U3873 ( .A1(n6290), .A2(n3875), .ZN(n5812) );
  INV_X1 U3874 ( .A(n6318), .ZN(n6014) );
  INV_X1 U3875 ( .A(n5984), .ZN(n6294) );
  INV_X1 U3876 ( .A(n6276), .ZN(n5829) );
  CLKBUF_X1 U3877 ( .A(n5001), .Z(n5002) );
  INV_X1 U3878 ( .A(n6312), .ZN(n6018) );
  CLKBUF_X1 U3879 ( .A(n4574), .Z(n4575) );
  NOR2_X1 U3880 ( .A1(n6014), .A2(n5817), .ZN(n4699) );
  INV_X1 U3881 ( .A(n3878), .ZN(n5792) );
  NAND2_X1 U3882 ( .A1(n3486), .A2(n3485), .ZN(n3487) );
  INV_X1 U3883 ( .A(n3484), .ZN(n3485) );
  INV_X1 U3884 ( .A(n4553), .ZN(n4885) );
  INV_X1 U3885 ( .A(n4554), .ZN(n5843) );
  INV_X1 U3886 ( .A(n6639), .ZN(n6642) );
  INV_X1 U3887 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6966) );
  CLKBUF_X1 U3888 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n5854) );
  OR2_X1 U3889 ( .A1(n4779), .A2(n4563), .ZN(n4829) );
  OR2_X1 U3890 ( .A1(n4779), .A2(n6325), .ZN(n4806) );
  AND2_X1 U3891 ( .A1(n6408), .A2(n6356), .ZN(n6427) );
  NOR2_X1 U3892 ( .A1(n4648), .A2(n5327), .ZN(n6492) );
  INV_X1 U3893 ( .A(n6374), .ZN(n6460) );
  INV_X1 U3894 ( .A(n6377), .ZN(n6466) );
  INV_X1 U3895 ( .A(n6381), .ZN(n6472) );
  INV_X1 U3896 ( .A(n6388), .ZN(n6484) );
  INV_X1 U3897 ( .A(n6392), .ZN(n6490) );
  INV_X1 U3898 ( .A(n6397), .ZN(n6500) );
  AND2_X1 U3899 ( .A1(n4411), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6544) );
  AND2_X1 U3900 ( .A1(n4549), .A2(n6530), .ZN(n6532) );
  NAND2_X1 U3901 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6521), .ZN(n6539) );
  INV_X1 U3902 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U3903 ( .B1(n5319), .B2(n6272), .A(n5296), .ZN(n5297) );
  AND2_X1 U3904 ( .A1(n3144), .A2(n3977), .ZN(n3113) );
  INV_X1 U3905 ( .A(n3298), .ZN(n3389) );
  NAND2_X1 U3906 ( .A1(n3909), .A2(n3736), .ZN(n3367) );
  OR2_X1 U3907 ( .A1(n3097), .A2(n5386), .ZN(n3114) );
  INV_X1 U3908 ( .A(n3132), .ZN(n5375) );
  AND2_X1 U3909 ( .A1(n5588), .A2(n3146), .ZN(n3115) );
  NAND2_X1 U3910 ( .A1(n6411), .A2(n4394), .ZN(n6283) );
  NAND2_X1 U3911 ( .A1(n5601), .A2(n5264), .ZN(n3116) );
  NAND2_X1 U3912 ( .A1(n5413), .A2(n3126), .ZN(n5493) );
  AND2_X1 U3913 ( .A1(n5438), .A2(n5440), .ZN(n5426) );
  NOR2_X1 U3914 ( .A1(n5748), .A2(n3649), .ZN(n5586) );
  AND2_X1 U3915 ( .A1(n3323), .A2(n3317), .ZN(n3359) );
  AND2_X1 U3916 ( .A1(n3633), .A2(n3631), .ZN(n3117) );
  NAND2_X1 U3917 ( .A1(n4622), .A2(n3317), .ZN(n3328) );
  NAND2_X1 U3918 ( .A1(n5572), .A2(n3646), .ZN(n5574) );
  INV_X1 U3919 ( .A(n3263), .ZN(n3323) );
  NOR2_X1 U3920 ( .A1(n3097), .A2(n3134), .ZN(n3132) );
  AND2_X1 U3921 ( .A1(n5413), .A2(n5513), .ZN(n5396) );
  NAND2_X1 U3922 ( .A1(n3328), .A2(n3471), .ZN(n3335) );
  AND2_X1 U3923 ( .A1(n5748), .A2(n5587), .ZN(n5572) );
  AND2_X1 U3924 ( .A1(n3116), .A2(n3626), .ZN(n3118) );
  CLKBUF_X3 U3925 ( .A(n3287), .Z(n3559) );
  INV_X1 U3926 ( .A(n3912), .ZN(n4326) );
  NAND2_X1 U3927 ( .A1(n5438), .A2(n3131), .ZN(n5425) );
  OR2_X1 U3928 ( .A1(n5689), .A2(n3644), .ZN(n3119) );
  NAND2_X1 U3929 ( .A1(n5601), .A2(n3852), .ZN(n3120) );
  AND2_X1 U3930 ( .A1(n3735), .A2(n3719), .ZN(n3688) );
  NAND2_X1 U3931 ( .A1(n5413), .A2(n3127), .ZN(n5395) );
  NAND2_X1 U3932 ( .A1(n3136), .A2(n3626), .ZN(n5253) );
  AND2_X1 U3933 ( .A1(n4622), .A2(n3337), .ZN(n3909) );
  INV_X1 U3934 ( .A(n3332), .ZN(n3479) );
  NOR2_X1 U3935 ( .A1(n3362), .A2(n3332), .ZN(n3720) );
  NAND2_X1 U3936 ( .A1(n3632), .A2(n3117), .ZN(n5680) );
  NAND2_X1 U3937 ( .A1(n3632), .A2(n3631), .ZN(n5681) );
  INV_X1 U3938 ( .A(n3128), .ZN(n3127) );
  NAND2_X1 U3939 ( .A1(n5397), .A2(n5513), .ZN(n3128) );
  AND2_X1 U3940 ( .A1(n3568), .A2(n3593), .ZN(n3121) );
  OR2_X1 U3941 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4357) );
  NOR2_X1 U3942 ( .A1(n5223), .A2(n6009), .ZN(n3122) );
  NAND2_X1 U3943 ( .A1(n3933), .A2(n3932), .ZN(n4485) );
  NOR2_X2 U3944 ( .A1(n4491), .A2(n4492), .ZN(n4490) );
  AND2_X1 U3945 ( .A1(n3500), .A2(n4472), .ZN(n4573) );
  NAND3_X1 U3946 ( .A1(n3991), .A2(n3990), .A3(n3989), .ZN(n3123) );
  INV_X1 U3947 ( .A(n3882), .ZN(n3146) );
  INV_X1 U3948 ( .A(n6624), .ZN(n3124) );
  INV_X1 U3949 ( .A(n3124), .ZN(n3125) );
  AOI221_X1 U3950 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6031), .C2(STATE_REG_0__SCAN_IN), .A(n6667), .ZN(n6624) );
  NOR4_X2 U3951 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n6649)
         );
  NAND2_X1 U3952 ( .A1(n3136), .A2(n3118), .ZN(n3628) );
  NAND2_X1 U3953 ( .A1(n3624), .A2(n3623), .ZN(n5246) );
  NOR2_X1 U3954 ( .A1(n3627), .A2(n3138), .ZN(n3137) );
  INV_X1 U3955 ( .A(n3623), .ZN(n3138) );
  OAI21_X1 U3956 ( .B1(n5648), .B2(n3141), .A(n3139), .ZN(n3142) );
  INV_X1 U3957 ( .A(n3641), .ZN(n3141) );
  NAND2_X1 U3958 ( .A1(n3144), .A2(n3143), .ZN(n5120) );
  NAND2_X1 U3959 ( .A1(n5586), .A2(n5588), .ZN(n5580) );
  NAND2_X1 U3960 ( .A1(n5564), .A2(n3155), .ZN(n3145) );
  NAND2_X1 U3961 ( .A1(n3569), .A2(n3568), .ZN(n3595) );
  NAND2_X1 U3962 ( .A1(n3569), .A2(n3121), .ZN(n3614) );
  AND2_X2 U3963 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4540) );
  INV_X1 U3964 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3157) );
  INV_X1 U3965 ( .A(n3497), .ZN(n3499) );
  NAND2_X1 U3966 ( .A1(n3376), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3350) );
  INV_X1 U3967 ( .A(n5649), .ZN(n5650) );
  INV_X1 U3968 ( .A(n5574), .ZN(n3648) );
  INV_X1 U3969 ( .A(n6169), .ZN(n6161) );
  NOR2_X1 U3970 ( .A1(n5229), .A2(n5399), .ZN(n3147) );
  AND2_X1 U3971 ( .A1(n3647), .A2(n5709), .ZN(n3148) );
  OR2_X1 U3972 ( .A1(n3352), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3149)
         );
  AND2_X1 U3973 ( .A1(n4345), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3150) );
  AND3_X1 U3974 ( .A1(n3260), .A2(n3259), .A3(n3258), .ZN(n3151) );
  NAND3_X1 U3975 ( .A1(n3773), .A2(n3818), .A3(n3772), .ZN(n3153) );
  AND2_X1 U3976 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3155) );
  INV_X1 U3977 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3498) );
  NOR2_X1 U3978 ( .A1(n5400), .A2(n5399), .ZN(n3156) );
  INV_X1 U3979 ( .A(n5024), .ZN(n6630) );
  INV_X1 U3980 ( .A(n6630), .ZN(n6411) );
  INV_X1 U3981 ( .A(n4559), .ZN(n4658) );
  NAND2_X1 U3982 ( .A1(n3152), .A2(n3318), .ZN(n3319) );
  INV_X1 U3983 ( .A(n3700), .ZN(n3678) );
  INV_X1 U3984 ( .A(n3701), .ZN(n3672) );
  NAND2_X1 U3985 ( .A1(n3688), .A2(n3687), .ZN(n3689) );
  AND2_X1 U3986 ( .A1(n6362), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3663)
         );
  AND2_X1 U3987 ( .A1(n5601), .A2(n6850), .ZN(n3639) );
  INV_X1 U3988 ( .A(n3549), .ZN(n3573) );
  AND2_X1 U3989 ( .A1(n4345), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3163) );
  OR2_X1 U3990 ( .A1(n3458), .A2(n3457), .ZN(n3491) );
  INV_X1 U3991 ( .A(n5376), .ZN(n4249) );
  INV_X1 U3992 ( .A(n5273), .ZN(n4036) );
  INV_X1 U3993 ( .A(n5070), .ZN(n3977) );
  AOI22_X1 U3994 ( .A1(n4345), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3286), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3243) );
  AND2_X1 U3995 ( .A1(n4940), .A2(n3841), .ZN(n3842) );
  INV_X1 U3996 ( .A(n4337), .ZN(n3896) );
  INV_X1 U3997 ( .A(n4184), .ZN(n3894) );
  NOR2_X1 U3998 ( .A1(n4151), .A2(n5404), .ZN(n4154) );
  INV_X1 U3999 ( .A(n4383), .ZN(n4354) );
  INV_X1 U4000 ( .A(n3905), .ZN(n3906) );
  NAND2_X1 U4001 ( .A1(n3488), .A2(n3616), .ZN(n3476) );
  INV_X1 U4002 ( .A(n5750), .ZN(n3645) );
  NAND2_X1 U4003 ( .A1(n4563), .A2(n3688), .ZN(n3494) );
  AND2_X1 U4004 ( .A1(n4941), .A2(n6533), .ZN(n4944) );
  INV_X1 U4005 ( .A(n5523), .ZN(n3794) );
  INV_X1 U4006 ( .A(n4516), .ZN(n3762) );
  NAND2_X1 U4007 ( .A1(n3896), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4387)
         );
  AND2_X1 U4008 ( .A1(n4136), .A2(n4135), .ZN(n5513) );
  NOR2_X1 U4009 ( .A1(n4021), .A2(n6084), .ZN(n4038) );
  INV_X1 U4010 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3647) );
  OR2_X1 U4011 ( .A1(n5601), .A2(n3640), .ZN(n3641) );
  AND2_X1 U4012 ( .A1(n4890), .A2(n5024), .ZN(n4892) );
  NAND2_X1 U4013 ( .A1(n3508), .A2(n3507), .ZN(n6359) );
  AND2_X1 U4014 ( .A1(n4537), .A2(n4536), .ZN(n6513) );
  OR2_X1 U4015 ( .A1(n3701), .A2(n3712), .ZN(n3702) );
  NAND2_X1 U4016 ( .A1(n6070), .A2(n5313), .ZN(n5401) );
  NAND2_X1 U4017 ( .A1(n6075), .A2(REIP_REG_13__SCAN_IN), .ZN(n5445) );
  AND2_X1 U4018 ( .A1(n3988), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3992)
         );
  AND3_X1 U4019 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .A3(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n3934) );
  NAND2_X1 U4020 ( .A1(n4229), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4264)
         );
  NAND2_X1 U4021 ( .A1(n4098), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4116)
         );
  NAND2_X1 U4022 ( .A1(n3862), .A2(n6522), .ZN(n4697) );
  OR2_X1 U4023 ( .A1(n5821), .A2(n6014), .ZN(n3878) );
  OR2_X1 U4024 ( .A1(n6516), .A2(n4616), .ZN(n6503) );
  OR2_X1 U4025 ( .A1(n5105), .A2(n4563), .ZN(n5149) );
  AND2_X1 U4026 ( .A1(n4559), .A2(n4774), .ZN(n6408) );
  INV_X1 U4027 ( .A(n6495), .ZN(n5900) );
  INV_X1 U4028 ( .A(n5073), .ZN(n5097) );
  AOI21_X1 U4029 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6362), .A(n5013), .ZN(
        n6448) );
  OR3_X1 U4030 ( .A1(n6516), .A2(n4398), .A3(n6036), .ZN(n4401) );
  NOR2_X1 U4031 ( .A1(n6600), .A2(n5942), .ZN(n5392) );
  OR2_X1 U4032 ( .A1(n5343), .A2(n4947), .ZN(n6118) );
  NOR2_X1 U4033 ( .A1(n6111), .A2(n5226), .ZN(n6102) );
  INV_X1 U4034 ( .A(n5905), .ZN(n6114) );
  INV_X1 U4035 ( .A(n6121), .ZN(n6135) );
  INV_X1 U4036 ( .A(n6156), .ZN(n6671) );
  INV_X1 U4037 ( .A(n6168), .ZN(n6163) );
  INV_X1 U4038 ( .A(n6200), .ZN(n6191) );
  INV_X1 U4039 ( .A(n6202), .ZN(n6243) );
  NAND2_X1 U4040 ( .A1(n4133), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4151)
         );
  NAND2_X1 U4041 ( .A1(n6521), .A2(n6544), .ZN(n4431) );
  INV_X1 U4042 ( .A(n6266), .ZN(n6280) );
  NAND2_X1 U4043 ( .A1(n5580), .A2(n5581), .ZN(n5582) );
  INV_X1 U4044 ( .A(n3870), .ZN(n3862) );
  NAND2_X1 U4045 ( .A1(n6660), .A2(n4607), .ZN(n5013) );
  NOR2_X1 U4046 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6545) );
  INV_X1 U4047 ( .A(n5149), .ZN(n4691) );
  AND2_X1 U4048 ( .A1(n4559), .A2(n4657), .ZN(n4719) );
  INV_X1 U4049 ( .A(n4849), .ZN(n5152) );
  OAI21_X1 U4050 ( .B1(n4816), .B2(n4817), .A(n6364), .ZN(n4842) );
  INV_X1 U4051 ( .A(n4829), .ZN(n4846) );
  INV_X1 U4052 ( .A(n4806), .ZN(n4652) );
  NOR2_X1 U4053 ( .A1(n6326), .A2(n4563), .ZN(n6349) );
  INV_X1 U4054 ( .A(n6357), .ZN(n6399) );
  AND2_X1 U4055 ( .A1(n6408), .A2(n5022), .ZN(n6429) );
  NOR2_X2 U4056 ( .A1(n4895), .A2(n6325), .ZN(n5902) );
  NOR2_X1 U4057 ( .A1(n5856), .A2(n6355), .ZN(n6495) );
  AND2_X1 U4058 ( .A1(n6435), .A2(n5022), .ZN(n6494) );
  NOR2_X1 U4059 ( .A1(n4856), .A2(n4563), .ZN(n5014) );
  INV_X1 U4060 ( .A(n4973), .ZN(n4996) );
  NOR2_X1 U4061 ( .A1(n6220), .A2(n5013), .ZN(n6371) );
  INV_X1 U4062 ( .A(n4720), .ZN(n4746) );
  NOR2_X1 U4063 ( .A1(n4403), .A2(n4402), .ZN(n6662) );
  INV_X1 U4064 ( .A(n6119), .ZN(n6132) );
  NAND2_X1 U4065 ( .A1(n5204), .A2(n4933), .ZN(n5905) );
  INV_X1 U4066 ( .A(n5646), .ZN(n5554) );
  NOR2_X1 U4067 ( .A1(n6188), .A2(n6184), .ZN(n6189) );
  INV_X1 U4068 ( .A(n6188), .ZN(n6199) );
  INV_X1 U4069 ( .A(n6246), .ZN(n6202) );
  OR2_X2 U4070 ( .A1(n4431), .A2(n4420), .ZN(n6251) );
  INV_X1 U4071 ( .A(n6262), .ZN(n6277) );
  OR2_X1 U4072 ( .A1(n4431), .A2(n3888), .ZN(n5695) );
  NOR2_X1 U4073 ( .A1(n5818), .A2(n5830), .ZN(n6290) );
  INV_X1 U4074 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6641) );
  INV_X1 U4075 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U4076 ( .A1(n4719), .A2(n4563), .ZN(n4720) );
  OR2_X1 U4077 ( .A1(n5105), .A2(n6325), .ZN(n4849) );
  INV_X1 U4078 ( .A(n6349), .ZN(n4655) );
  AOI21_X1 U4079 ( .B1(n6630), .B2(n6327), .A(n6324), .ZN(n6354) );
  NOR2_X1 U4080 ( .A1(n6367), .A2(n6366), .ZN(n6403) );
  NAND2_X1 U4081 ( .A1(n4886), .A2(n6325), .ZN(n5066) );
  AOI22_X1 U4082 ( .A1(n5864), .A2(n6437), .B1(n5861), .B2(n5860), .ZN(n5904)
         );
  INV_X1 U4083 ( .A(n6385), .ZN(n6478) );
  INV_X1 U4084 ( .A(n5014), .ZN(n5104) );
  NAND2_X1 U4085 ( .A1(n4850), .A2(n4563), .ZN(n4973) );
  INV_X1 U4086 ( .A(n6371), .ZN(n6454) );
  INV_X1 U4087 ( .A(n4976), .ZN(n4999) );
  INV_X1 U4088 ( .A(n6609), .ZN(n6617) );
  AND2_X4 U4089 ( .A1(n3157), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4524)
         );
  INV_X1 U4090 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3158) );
  AND2_X2 U4091 ( .A1(n3158), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3165)
         );
  NOR2_X4 U4092 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3175) );
  AND2_X2 U4093 ( .A1(n3165), .A2(n3175), .ZN(n3304) );
  NAND2_X1 U4094 ( .A1(n3304), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3161) );
  AND2_X2 U4095 ( .A1(n3165), .A2(n4540), .ZN(n3303) );
  NAND2_X1 U4096 ( .A1(n3303), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3160)
         );
  AND2_X4 U4097 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4459) );
  AND2_X4 U4098 ( .A1(n4524), .A2(n4459), .ZN(n3286) );
  NAND2_X1 U4099 ( .A1(n3286), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3159) );
  NAND3_X1 U4100 ( .A1(n3161), .A2(n3160), .A3(n3159), .ZN(n3162) );
  AND2_X2 U4101 ( .A1(n4540), .A2(n4459), .ZN(n3390) );
  NAND2_X1 U4102 ( .A1(n3390), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3169)
         );
  NAND2_X1 U4103 ( .A1(n3387), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3168) );
  INV_X1 U4104 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3164) );
  AND2_X4 U4105 ( .A1(n3164), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4523)
         );
  NOR2_X4 U4106 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4543) );
  AND2_X4 U4107 ( .A1(n4523), .A2(n4543), .ZN(n3292) );
  NAND2_X1 U4108 ( .A1(n3292), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3167) );
  AND2_X2 U4109 ( .A1(n4523), .A2(n3165), .ZN(n3388) );
  NAND2_X1 U4110 ( .A1(n3388), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3166)
         );
  AND2_X2 U4111 ( .A1(n3174), .A2(n3175), .ZN(n3297) );
  NAND2_X1 U4112 ( .A1(n3297), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U4113 ( .A1(n3420), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3172) );
  AND2_X4 U4114 ( .A1(n4524), .A2(n4543), .ZN(n3421) );
  NAND2_X1 U4115 ( .A1(n3421), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3171) );
  AND2_X2 U4116 ( .A1(n3175), .A2(n4459), .ZN(n3298) );
  NAND2_X1 U4117 ( .A1(n3298), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3170) );
  AND2_X4 U4118 ( .A1(n4459), .A2(n4523), .ZN(n3287) );
  NAND2_X1 U4119 ( .A1(n3287), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3179)
         );
  NAND2_X1 U4120 ( .A1(n3426), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3178)
         );
  AND2_X4 U4121 ( .A1(n4543), .A2(n3175), .ZN(n3448) );
  NAND2_X1 U4122 ( .A1(n3448), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3177) );
  AND2_X4 U4123 ( .A1(n4543), .A2(n4540), .ZN(n3285) );
  NAND2_X1 U4124 ( .A1(n3285), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3176)
         );
  INV_X1 U4126 ( .A(n3317), .ZN(n3194) );
  AOI22_X1 U4127 ( .A1(n3387), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4128 ( .A1(n3420), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4129 ( .A1(n3298), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3184) );
  AND4_X2 U4130 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3193)
         );
  AOI22_X1 U4131 ( .A1(n4345), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4132 ( .A1(n3426), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4133 ( .A1(n3286), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3188) );
  AND4_X2 U4134 ( .A1(n3191), .A2(n3190), .A3(n3189), .A4(n3188), .ZN(n3192)
         );
  NAND2_X2 U4135 ( .A1(n3193), .A2(n3192), .ZN(n3336) );
  NAND2_X2 U4136 ( .A1(n3194), .A2(n3336), .ZN(n4410) );
  NAND2_X1 U4137 ( .A1(n4345), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4138 ( .A1(n3426), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4139 ( .A1(n3448), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4140 ( .A1(n3285), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3195)
         );
  INV_X1 U4141 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4142 ( .A1(n3292), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4143 ( .A1(n3421), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4144 ( .A1(n3388), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3200)
         );
  NAND3_X1 U4145 ( .A1(n3202), .A2(n3201), .A3(n3200), .ZN(n3203) );
  NOR2_X2 U4146 ( .A1(n3204), .A2(n3203), .ZN(n3215) );
  NAND2_X1 U4147 ( .A1(n3387), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4148 ( .A1(n3420), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4149 ( .A1(n3297), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4150 ( .A1(n3390), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4151 ( .A1(n3286), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4152 ( .A1(n3287), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3211)
         );
  NAND2_X1 U4153 ( .A1(n3303), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3210)
         );
  NAND2_X1 U4154 ( .A1(n3304), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3209) );
  NAND4_X4 U4155 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3337)
         );
  INV_X1 U4156 ( .A(n3328), .ZN(n3238) );
  NAND2_X1 U4157 ( .A1(n3390), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4158 ( .A1(n3297), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4159 ( .A1(n3421), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4160 ( .A1(n3298), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4161 ( .A1(n3420), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4162 ( .A1(n3387), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4163 ( .A1(n3388), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3222)
         );
  NAND2_X1 U4164 ( .A1(n3292), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4165 ( .A1(n3426), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4166 ( .A1(n3303), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3227)
         );
  NAND2_X1 U4167 ( .A1(n3304), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4168 ( .A1(n3448), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4169 ( .A1(n3110), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4170 ( .A1(n3287), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3231)
         );
  NAND2_X1 U4171 ( .A1(n3286), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4172 ( .A1(n3285), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3229)
         );
  INV_X1 U4173 ( .A(n3736), .ZN(n3237) );
  NAND2_X1 U4174 ( .A1(n3238), .A2(n3237), .ZN(n3239) );
  NAND2_X1 U4175 ( .A1(n3240), .A2(n3239), .ZN(n3362) );
  AOI22_X1 U4176 ( .A1(n3426), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4177 ( .A1(n3420), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3387), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3242) );
  NAND4_X1 U4178 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3251)
         );
  AOI22_X1 U4179 ( .A1(n3388), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4180 ( .A1(n3303), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4181 ( .A1(n3287), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4182 ( .A1(n3421), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4183 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  OR2_X2 U4184 ( .A1(n3251), .A2(n3250), .ZN(n3471) );
  NAND2_X1 U4185 ( .A1(n3286), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4186 ( .A1(n3285), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3252)
         );
  AND2_X1 U4187 ( .A1(n3253), .A2(n3252), .ZN(n3262) );
  AOI22_X1 U4188 ( .A1(n3420), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4189 ( .A1(n3387), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4190 ( .A1(n3421), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4191 ( .A1(n3298), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4192 ( .A1(n4345), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4193 ( .A1(n3426), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4194 ( .A1(n3303), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3258) );
  NAND2_X1 U4195 ( .A1(n3471), .A2(n3342), .ZN(n3332) );
  NAND2_X1 U4196 ( .A1(n4345), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4197 ( .A1(n3559), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3267)
         );
  NAND2_X1 U4198 ( .A1(n3286), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4199 ( .A1(n3285), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3265)
         );
  AND4_X2 U4200 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3284)
         );
  NAND2_X1 U4201 ( .A1(n3420), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4202 ( .A1(n3387), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4203 ( .A1(n3388), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3270)
         );
  NAND2_X1 U4204 ( .A1(n3292), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4205 ( .A1(n3426), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3276)
         );
  NAND2_X1 U4206 ( .A1(n3303), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3275)
         );
  NAND2_X1 U4207 ( .A1(n3304), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4208 ( .A1(n3448), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3273) );
  NAND2_X1 U4209 ( .A1(n3421), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4210 ( .A1(n3297), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4211 ( .A1(n3390), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3278)
         );
  NAND2_X1 U4212 ( .A1(n3298), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3277) );
  NAND4_X4 U4213 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3734)
         );
  NAND2_X1 U4214 ( .A1(n3285), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3290)
         );
  NAND2_X1 U4215 ( .A1(n3286), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4216 ( .A1(n3287), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3288)
         );
  NAND3_X1 U4217 ( .A1(n3290), .A2(n3289), .A3(n3288), .ZN(n3291) );
  NOR2_X1 U4218 ( .A1(n3150), .A2(n3291), .ZN(n3312) );
  NAND2_X1 U4219 ( .A1(n3420), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3296) );
  NAND2_X1 U4220 ( .A1(n3387), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4221 ( .A1(n3388), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3294)
         );
  NAND2_X1 U4222 ( .A1(n3292), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3293) );
  AND4_X2 U4223 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3311)
         );
  NAND2_X1 U4224 ( .A1(n3390), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3302)
         );
  NAND2_X1 U4225 ( .A1(n3297), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4226 ( .A1(n3421), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U4227 ( .A1(n3298), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4228 ( .A1(n3426), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3308)
         );
  NAND2_X1 U4229 ( .A1(n3303), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U4230 ( .A1(n3304), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4231 ( .A1(n3448), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3305) );
  NAND4_X2 U4232 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3315)
         );
  NAND2_X1 U4233 ( .A1(n3722), .A2(n3366), .ZN(n3314) );
  NAND2_X1 U4234 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6568) );
  OAI21_X1 U4235 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6568), .ZN(n3705) );
  INV_X1 U4236 ( .A(n3705), .ZN(n3316) );
  NAND3_X1 U4237 ( .A1(n3720), .A2(n3371), .A3(n3319), .ZN(n3320) );
  NAND2_X1 U4238 ( .A1(n3320), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3331) );
  INV_X1 U4239 ( .A(n3909), .ZN(n3321) );
  NAND3_X1 U4240 ( .A1(n3321), .A2(n3323), .A3(n4410), .ZN(n3322) );
  NAND2_X1 U4241 ( .A1(n3322), .A2(n3855), .ZN(n3326) );
  NAND2_X1 U4242 ( .A1(n4410), .A2(n3342), .ZN(n3324) );
  NAND2_X1 U4243 ( .A1(n3324), .A2(n3337), .ZN(n3325) );
  NAND3_X1 U4244 ( .A1(n3326), .A2(n3340), .A3(n3335), .ZN(n3358) );
  INV_X1 U4245 ( .A(n3509), .ZN(n3327) );
  INV_X1 U4246 ( .A(n3238), .ZN(n3363) );
  NAND2_X1 U4247 ( .A1(n3695), .A2(n3363), .ZN(n3329) );
  INV_X1 U4248 ( .A(n3722), .ZN(n3334) );
  NOR2_X1 U4249 ( .A1(n3332), .A2(n3719), .ZN(n3333) );
  NAND2_X1 U4250 ( .A1(n4399), .A2(n3152), .ZN(n3347) );
  INV_X1 U4251 ( .A(n3335), .ZN(n3339) );
  NAND2_X1 U4252 ( .A1(n3359), .A2(n3345), .ZN(n3338) );
  NOR2_X1 U4253 ( .A1(n3719), .A2(n3471), .ZN(n3343) );
  NAND3_X1 U4254 ( .A1(n3344), .A2(n3342), .A3(n3343), .ZN(n4453) );
  NOR2_X2 U4255 ( .A1(n4453), .A2(n3854), .ZN(n3733) );
  INV_X1 U4256 ( .A(n3733), .ZN(n3346) );
  NAND3_X1 U4257 ( .A1(n3347), .A2(n3737), .A3(n3346), .ZN(n3354) );
  NAND2_X1 U4258 ( .A1(n3354), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4259 ( .A1(n6545), .A2(n6660), .ZN(n3889) );
  INV_X1 U4260 ( .A(n3889), .ZN(n3506) );
  XNOR2_X1 U4261 ( .A(n6362), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5006)
         );
  INV_X1 U4262 ( .A(n3351), .ZN(n3352) );
  AND2_X1 U4263 ( .A1(n3149), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4264 ( .A1(n3354), .A2(n3353), .ZN(n3355) );
  INV_X1 U4265 ( .A(n3407), .ZN(n3374) );
  NAND2_X1 U4266 ( .A1(n3376), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3357) );
  MUX2_X1 U4267 ( .A(n3889), .B(n4411), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3356) );
  NAND2_X1 U4268 ( .A1(n3357), .A2(n3356), .ZN(n3442) );
  NAND2_X1 U4269 ( .A1(n4632), .A2(n3735), .ZN(n4936) );
  OAI22_X1 U4270 ( .A1(n3359), .A2(n4936), .B1(n4632), .B2(n3342), .ZN(n3360)
         );
  NAND2_X1 U4271 ( .A1(n3363), .A2(n3736), .ZN(n3364) );
  NAND2_X1 U4272 ( .A1(n3364), .A2(n3471), .ZN(n3365) );
  OAI21_X1 U4273 ( .B1(n3362), .B2(n3365), .A(n3735), .ZN(n3372) );
  NAND2_X1 U4274 ( .A1(n6545), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6039) );
  AOI21_X1 U4275 ( .B1(n6658), .B2(n3335), .A(n6039), .ZN(n3370) );
  INV_X1 U4276 ( .A(n3367), .ZN(n3369) );
  INV_X1 U4277 ( .A(n3471), .ZN(n4637) );
  AND3_X1 U4278 ( .A1(n3342), .A2(n4637), .A3(n4632), .ZN(n3368) );
  NAND2_X1 U4279 ( .A1(n3369), .A2(n3368), .ZN(n4533) );
  NAND2_X1 U4280 ( .A1(n3859), .A2(n3373), .ZN(n3441) );
  NAND2_X2 U4281 ( .A1(n3442), .A2(n3441), .ZN(n3444) );
  NAND2_X1 U4282 ( .A1(n3384), .A2(n3109), .ZN(n3382) );
  NAND2_X1 U4283 ( .A1(n3376), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4284 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3377) );
  NAND2_X1 U4285 ( .A1(n3377), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3378) );
  NOR2_X1 U4286 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6969), .ZN(n5862)
         );
  NAND2_X1 U4287 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5862), .ZN(n6438) );
  NAND2_X1 U4288 ( .A1(n3378), .A2(n6438), .ZN(n4610) );
  AOI22_X1 U4289 ( .A1(n3506), .A2(n4610), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3505), .ZN(n3379) );
  NAND2_X1 U4290 ( .A1(n3380), .A2(n3379), .ZN(n3383) );
  INV_X1 U4291 ( .A(n3383), .ZN(n3381) );
  NAND2_X1 U4292 ( .A1(n3382), .A2(n3381), .ZN(n3386) );
  AOI22_X1 U4293 ( .A1(n4311), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4294 ( .A1(n4360), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3393) );
  CLKBUF_X2 U4295 ( .A(n3297), .Z(n3447) );
  AOI22_X1 U4296 ( .A1(n4361), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3392) );
  INV_X2 U4297 ( .A(n3389), .ZN(n4372) );
  INV_X1 U4298 ( .A(n3390), .ZN(n4521) );
  INV_X2 U4299 ( .A(n4521), .ZN(n4371) );
  AOI22_X1 U4300 ( .A1(n4372), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4301 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3402)
         );
  INV_X1 U4302 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6933) );
  AOI22_X1 U4303 ( .A1(n4367), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3559), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3400) );
  INV_X1 U4304 ( .A(n3304), .ZN(n3395) );
  AOI22_X1 U4305 ( .A1(n4368), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3399) );
  INV_X1 U4306 ( .A(n3426), .ZN(n3396) );
  INV_X2 U4307 ( .A(n3396), .ZN(n3446) );
  AOI22_X1 U4308 ( .A1(n3446), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4309 ( .A1(n4522), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4310 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  INV_X1 U4312 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3403) );
  OAI22_X1 U4313 ( .A1(n3679), .A2(n3403), .B1(n3509), .B2(n3470), .ZN(n3404)
         );
  INV_X1 U4314 ( .A(n3404), .ZN(n3405) );
  XNOR2_X2 U4315 ( .A(n3444), .B(n3407), .ZN(n4554) );
  INV_X1 U4316 ( .A(n3510), .ZN(n4413) );
  AOI22_X1 U4317 ( .A1(n4369), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4318 ( .A1(n4360), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4319 ( .A1(n4522), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4320 ( .A1(n4361), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3408) );
  NAND4_X1 U4321 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3418)
         );
  AOI22_X1 U4322 ( .A1(n4367), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3559), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4323 ( .A1(n4311), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4324 ( .A1(n4359), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4325 ( .A1(n4187), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3413) );
  NAND4_X1 U4326 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3417)
         );
  NAND2_X1 U4327 ( .A1(n4413), .A2(n3478), .ZN(n3419) );
  OAI21_X2 U4328 ( .B1(n4554), .B2(STATE2_REG_0__SCAN_IN), .A(n3419), .ZN(
        n3439) );
  INV_X1 U4329 ( .A(n3439), .ZN(n3436) );
  NAND2_X1 U4330 ( .A1(n3695), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4331 ( .A1(n4311), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4332 ( .A1(n4360), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4333 ( .A1(n4361), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4334 ( .A1(n4372), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3422) );
  NAND4_X1 U4335 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3432)
         );
  AOI22_X1 U4336 ( .A1(n4367), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3559), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4337 ( .A1(n3303), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4338 ( .A1(n3446), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4339 ( .A1(n3286), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U4340 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3431)
         );
  NAND2_X1 U4341 ( .A1(n4413), .A2(n3603), .ZN(n3445) );
  INV_X1 U4342 ( .A(n3478), .ZN(n3433) );
  OR2_X1 U4343 ( .A1(n3509), .A2(n3433), .ZN(n3434) );
  NAND2_X1 U4344 ( .A1(n3436), .A2(n3437), .ZN(n3468) );
  INV_X1 U4345 ( .A(n3437), .ZN(n3438) );
  NAND2_X1 U4346 ( .A1(n3439), .A2(n3438), .ZN(n3440) );
  NAND2_X1 U4347 ( .A1(n3468), .A2(n3440), .ZN(n3475) );
  INV_X1 U4348 ( .A(n3475), .ZN(n3467) );
  NOR2_X1 U4349 ( .A1(n3603), .A2(n3510), .ZN(n3465) );
  INV_X1 U4350 ( .A(n3445), .ZN(n3459) );
  AOI22_X1 U4351 ( .A1(n4367), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4352 ( .A1(n4369), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4353 ( .A1(n4360), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4354 ( .A1(n4359), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3449) );
  NAND4_X1 U4355 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3458)
         );
  AOI22_X1 U4356 ( .A1(n3286), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4357 ( .A1(n4311), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4361), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4358 ( .A1(n3559), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4359 ( .A1(n4372), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4360 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  MUX2_X1 U4361 ( .A(n3465), .B(n3459), .S(n3491), .Z(n3460) );
  INV_X1 U4362 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3463) );
  AOI21_X1 U4363 ( .B1(n3237), .B2(n3618), .A(n6660), .ZN(n3462) );
  NAND2_X1 U4364 ( .A1(n4632), .A2(n3491), .ZN(n3461) );
  OAI211_X1 U4365 ( .C1(n3679), .C2(n3463), .A(n3462), .B(n3461), .ZN(n3484)
         );
  NAND2_X1 U4366 ( .A1(n3464), .A2(n3484), .ZN(n3488) );
  INV_X1 U4367 ( .A(n3465), .ZN(n3616) );
  INV_X1 U4368 ( .A(n3476), .ZN(n3466) );
  NAND2_X1 U4369 ( .A1(n3467), .A2(n3466), .ZN(n3469) );
  NAND2_X1 U4370 ( .A1(n3469), .A2(n3108), .ZN(n3501) );
  NAND2_X1 U4371 ( .A1(n4558), .A2(n3688), .ZN(n3474) );
  NAND2_X1 U4372 ( .A1(n3491), .A2(n3478), .ZN(n3477) );
  NAND2_X1 U4373 ( .A1(n3477), .A2(n3470), .ZN(n3528) );
  OAI21_X1 U4374 ( .B1(n3470), .B2(n3477), .A(n3528), .ZN(n3472) );
  AND2_X1 U4375 ( .A1(n4632), .A2(n3471), .ZN(n3489) );
  AOI21_X1 U4376 ( .B1(n3472), .B2(n6658), .A(n3489), .ZN(n3473) );
  NAND2_X1 U4377 ( .A1(n3474), .A2(n3473), .ZN(n3497) );
  NAND2_X1 U4378 ( .A1(n3497), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4471)
         );
  NAND2_X1 U4379 ( .A1(n4552), .A2(n3688), .ZN(n3483) );
  OAI21_X1 U4380 ( .B1(n3491), .B2(n3478), .A(n3477), .ZN(n3480) );
  INV_X1 U4381 ( .A(n6658), .ZN(n3723) );
  OAI211_X1 U4382 ( .C1(n3480), .C2(n3723), .A(n3479), .B(n3719), .ZN(n3481)
         );
  INV_X1 U4383 ( .A(n3481), .ZN(n3482) );
  NAND2_X1 U4384 ( .A1(n3483), .A2(n3482), .ZN(n4705) );
  INV_X1 U4385 ( .A(n3489), .ZN(n3490) );
  OAI21_X1 U4386 ( .B1(n3723), .B2(n3491), .A(n3490), .ZN(n3492) );
  INV_X1 U4387 ( .A(n3492), .ZN(n3493) );
  NAND2_X1 U4388 ( .A1(n3494), .A2(n3493), .ZN(n6275) );
  NAND2_X1 U4389 ( .A1(n6275), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6274)
         );
  XNOR2_X1 U4390 ( .A(n6274), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4704)
         );
  NAND2_X1 U4391 ( .A1(n4705), .A2(n4704), .ZN(n4707) );
  INV_X1 U4392 ( .A(n6274), .ZN(n3495) );
  NAND2_X1 U4393 ( .A1(n3495), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3496)
         );
  AND2_X1 U4394 ( .A1(n4707), .A2(n3496), .ZN(n4474) );
  NAND2_X1 U4395 ( .A1(n4471), .A2(n4474), .ZN(n3500) );
  NAND2_X1 U4396 ( .A1(n3499), .A2(n3498), .ZN(n4472) );
  INV_X1 U4397 ( .A(n3501), .ZN(n3503) );
  NAND2_X1 U4398 ( .A1(n3503), .A2(n3502), .ZN(n3526) );
  INV_X1 U4399 ( .A(n3526), .ZN(n3525) );
  NAND2_X1 U4400 ( .A1(n3376), .A2(n5854), .ZN(n3508) );
  NOR3_X1 U4401 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4887), .A3(n6969), 
        .ZN(n6412) );
  NAND2_X1 U4402 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6412), .ZN(n6404) );
  NAND2_X1 U4403 ( .A1(n6641), .A2(n6404), .ZN(n3504) );
  NAND3_X1 U4404 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4956) );
  INV_X1 U4405 ( .A(n4956), .ZN(n4714) );
  NAND2_X1 U4406 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4714), .ZN(n4744) );
  AOI22_X1 U4407 ( .A1(n3506), .A2(n5007), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3505), .ZN(n3507) );
  XNOR2_X2 U4408 ( .A(n4545), .B(n6359), .ZN(n5858) );
  AND2_X4 U4409 ( .A1(n3510), .A2(n3509), .ZN(n3700) );
  AOI22_X1 U4410 ( .A1(n4311), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4411 ( .A1(n4360), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4412 ( .A1(n4361), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3512) );
  INV_X1 U4413 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6935) );
  AOI22_X1 U4414 ( .A1(n4372), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4415 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3520)
         );
  AOI22_X1 U4416 ( .A1(n4367), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3559), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4417 ( .A1(n4368), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4418 ( .A1(n3446), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4419 ( .A1(n4522), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3515) );
  NAND4_X1 U4420 ( .A1(n3518), .A2(n3517), .A3(n3516), .A4(n3515), .ZN(n3519)
         );
  INV_X1 U4421 ( .A(n3529), .ZN(n3521) );
  OAI22_X1 U4422 ( .A1(n3700), .A2(n3521), .B1(n6935), .B2(n3679), .ZN(n3522)
         );
  INV_X1 U4423 ( .A(n3522), .ZN(n3523) );
  NAND2_X2 U4424 ( .A1(n3525), .A2(n4656), .ZN(n3547) );
  INV_X1 U4425 ( .A(n4656), .ZN(n4774) );
  NAND2_X1 U4426 ( .A1(n3526), .A2(n4774), .ZN(n3527) );
  INV_X1 U4427 ( .A(n3688), .ZN(n3615) );
  NAND2_X1 U4428 ( .A1(n3528), .A2(n3529), .ZN(n3574) );
  OAI211_X1 U4429 ( .C1(n3529), .C2(n3528), .A(n3574), .B(n6658), .ZN(n3530)
         );
  OAI21_X2 U4430 ( .B1(n4602), .B2(n3615), .A(n3530), .ZN(n3531) );
  INV_X1 U4431 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4580) );
  XNOR2_X1 U4432 ( .A(n3531), .B(n4580), .ZN(n4574) );
  NAND2_X1 U4433 ( .A1(n4573), .A2(n4574), .ZN(n3533) );
  NAND2_X1 U4434 ( .A1(n3531), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3532)
         );
  NAND2_X1 U4435 ( .A1(n3533), .A2(n3532), .ZN(n4592) );
  INV_X1 U4436 ( .A(n3547), .ZN(n3545) );
  AOI22_X1 U4437 ( .A1(n4367), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4438 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4369), .B1(n4359), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4439 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4360), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4440 ( .A1(n4372), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3534) );
  NAND4_X1 U4441 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(n3543)
         );
  AOI22_X1 U4442 ( .A1(n4311), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4443 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4361), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4444 ( .A1(n4522), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4445 ( .A1(n4366), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4446 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3542)
         );
  INV_X1 U4447 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6929) );
  OAI22_X1 U4448 ( .A1(n3700), .A2(n3573), .B1(n6929), .B2(n3679), .ZN(n3544)
         );
  INV_X1 U4449 ( .A(n3544), .ZN(n3546) );
  NAND2_X1 U4450 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  NAND2_X1 U4451 ( .A1(n3571), .A2(n3548), .ZN(n3941) );
  XNOR2_X1 U4452 ( .A(n3574), .B(n3549), .ZN(n3550) );
  NAND2_X1 U4453 ( .A1(n3550), .A2(n6658), .ZN(n3551) );
  OAI21_X2 U4454 ( .B1(n3941), .B2(n3615), .A(n3551), .ZN(n3552) );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3756) );
  XNOR2_X1 U4456 ( .A(n3552), .B(n3756), .ZN(n4593) );
  NAND2_X1 U4457 ( .A1(n4592), .A2(n4593), .ZN(n3554) );
  NAND2_X1 U4458 ( .A1(n3552), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3553)
         );
  INV_X1 U4459 ( .A(n3571), .ZN(n3569) );
  AOI22_X1 U4460 ( .A1(n4311), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3558) );
  INV_X1 U4461 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6932) );
  AOI22_X1 U4462 ( .A1(n4360), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4463 ( .A1(n4361), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4464 ( .A1(n4372), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3555) );
  NAND4_X1 U4465 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3565)
         );
  AOI22_X1 U4466 ( .A1(n4367), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4467 ( .A1(n4368), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4468 ( .A1(n3446), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4469 ( .A1(n4522), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4470 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3564)
         );
  INV_X1 U4471 ( .A(n3575), .ZN(n3567) );
  INV_X1 U4472 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3566) );
  OAI22_X1 U4473 ( .A1(n3700), .A2(n3567), .B1(n3566), .B2(n3679), .ZN(n3568)
         );
  INV_X1 U4474 ( .A(n3568), .ZN(n3570) );
  NAND2_X1 U4475 ( .A1(n3571), .A2(n3570), .ZN(n3572) );
  NOR2_X1 U4476 ( .A1(n3574), .A2(n3573), .ZN(n3576) );
  NAND2_X1 U4477 ( .A1(n3576), .A2(n3575), .ZN(n3605) );
  OAI211_X1 U4478 ( .C1(n3576), .C2(n3575), .A(n3605), .B(n6658), .ZN(n3577)
         );
  OAI21_X2 U4479 ( .B1(n3957), .B2(n3615), .A(n3577), .ZN(n3578) );
  INV_X1 U4480 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4481 ( .A1(n4694), .A2(n4695), .ZN(n3580) );
  NAND2_X1 U4482 ( .A1(n3578), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3579)
         );
  AOI22_X1 U4483 ( .A1(n4368), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4484 ( .A1(n4369), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4485 ( .A1(n4366), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4486 ( .A1(n4361), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3581) );
  NAND4_X1 U4487 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3590)
         );
  AOI22_X1 U4488 ( .A1(n4367), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4522), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4489 ( .A1(n4311), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4490 ( .A1(n3446), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4491 ( .A1(n4360), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4492 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3589)
         );
  INV_X1 U4493 ( .A(n3606), .ZN(n3592) );
  INV_X1 U4494 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3591) );
  INV_X1 U4495 ( .A(n3593), .ZN(n3594) );
  NAND2_X1 U4496 ( .A1(n3595), .A2(n3594), .ZN(n3962) );
  NAND3_X1 U4497 ( .A1(n3614), .A2(n3688), .A3(n3962), .ZN(n3598) );
  XNOR2_X1 U4498 ( .A(n3605), .B(n3606), .ZN(n3596) );
  NAND2_X1 U4499 ( .A1(n3596), .A2(n6658), .ZN(n3597) );
  NAND2_X1 U4500 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  INV_X1 U4501 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4878) );
  XNOR2_X1 U4502 ( .A(n3599), .B(n4878), .ZN(n4877) );
  NAND2_X1 U4503 ( .A1(n4876), .A2(n4877), .ZN(n3601) );
  NAND2_X1 U4504 ( .A1(n3599), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3600)
         );
  NAND2_X1 U4505 ( .A1(n3601), .A2(n3600), .ZN(n5001) );
  INV_X1 U4506 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4507 ( .A1(n3901), .A2(n3688), .ZN(n3610) );
  INV_X1 U4508 ( .A(n3605), .ZN(n3607) );
  NAND2_X1 U4509 ( .A1(n3607), .A2(n3606), .ZN(n3620) );
  XNOR2_X1 U4510 ( .A(n3620), .B(n3618), .ZN(n3608) );
  NAND2_X1 U4511 ( .A1(n3608), .A2(n6658), .ZN(n3609) );
  NAND2_X1 U4512 ( .A1(n3610), .A2(n3609), .ZN(n3611) );
  INV_X1 U4513 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6299) );
  XNOR2_X1 U4514 ( .A(n3611), .B(n6299), .ZN(n5000) );
  NAND2_X1 U4515 ( .A1(n5001), .A2(n5000), .ZN(n3613) );
  NAND2_X1 U4516 ( .A1(n3611), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3612)
         );
  NAND2_X1 U4517 ( .A1(n3613), .A2(n3612), .ZN(n5164) );
  NOR2_X1 U4518 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  NAND2_X1 U4519 ( .A1(n6658), .A2(n3618), .ZN(n3619) );
  OR2_X1 U4520 ( .A1(n3620), .A2(n3619), .ZN(n3621) );
  NAND2_X1 U4521 ( .A1(n3625), .A2(n3621), .ZN(n3622) );
  INV_X1 U4522 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U4523 ( .A1(n5164), .A2(n5165), .ZN(n3624) );
  NAND2_X1 U4524 ( .A1(n3622), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3623)
         );
  INV_X1 U4525 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6724) );
  NOR2_X1 U4526 ( .A1(n5601), .A2(n6724), .ZN(n3627) );
  NAND2_X1 U4527 ( .A1(n5601), .A2(n6724), .ZN(n3626) );
  INV_X1 U4528 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5264) );
  OR2_X1 U4529 ( .A1(n5601), .A2(n5264), .ZN(n5254) );
  NAND2_X1 U4530 ( .A1(n3628), .A2(n5254), .ZN(n5696) );
  INV_X1 U4531 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U4532 ( .A1(n5689), .A2(n6954), .ZN(n5697) );
  NAND2_X1 U4533 ( .A1(n5696), .A2(n5697), .ZN(n3629) );
  OR2_X1 U4534 ( .A1(n5601), .A2(n6954), .ZN(n5698) );
  INV_X1 U4535 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U4536 ( .A1(n5689), .A2(n6752), .ZN(n3630) );
  NAND2_X1 U4537 ( .A1(n5688), .A2(n3630), .ZN(n3632) );
  OR2_X1 U4538 ( .A1(n5601), .A2(n6752), .ZN(n3631) );
  INV_X1 U4539 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6023) );
  XNOR2_X1 U4540 ( .A(n5689), .B(n6023), .ZN(n5682) );
  NAND2_X1 U4541 ( .A1(n5689), .A2(n6023), .ZN(n3634) );
  INV_X1 U4542 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5822) );
  OR2_X1 U4543 ( .A1(n5601), .A2(n5822), .ZN(n3635) );
  NAND2_X1 U4544 ( .A1(n5689), .A2(n5822), .ZN(n3636) );
  NAND2_X1 U4545 ( .A1(n3637), .A2(n3636), .ZN(n5668) );
  XNOR2_X1 U4546 ( .A(n5689), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5667)
         );
  INV_X1 U4547 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U4548 ( .A1(n5689), .A2(n6898), .ZN(n3638) );
  INV_X1 U4549 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6850) );
  NOR2_X2 U4550 ( .A1(n5661), .A2(n3639), .ZN(n5648) );
  NAND2_X1 U4551 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3852) );
  INV_X1 U4552 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6811) );
  INV_X1 U4553 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6883) );
  AND3_X1 U4554 ( .A1(n6850), .A2(n6811), .A3(n6883), .ZN(n3640) );
  AND2_X1 U4555 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5795) );
  AND2_X1 U4556 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U4557 ( .A1(n5795), .A2(n3879), .ZN(n5609) );
  NAND2_X1 U4558 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3880) );
  OAI21_X1 U4559 ( .B1(n5609), .B2(n3880), .A(n5689), .ZN(n3642) );
  NOR2_X1 U4560 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5794) );
  NOR2_X1 U4561 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3643) );
  INV_X1 U4562 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5765) );
  INV_X1 U4563 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3822) );
  AND4_X1 U4564 ( .A1(n5794), .A2(n3643), .A3(n5765), .A4(n3822), .ZN(n3644)
         );
  XNOR2_X1 U4565 ( .A(n5689), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5750)
         );
  NOR2_X1 U4566 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5587)
         );
  NOR2_X1 U4567 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4568 ( .A1(n3648), .A2(n3647), .ZN(n3651) );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5751) );
  INV_X1 U4570 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U4571 ( .A1(n5652), .A2(n6684), .ZN(n5588) );
  NAND2_X1 U4572 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4573 ( .A1(n5564), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4574 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  XNOR2_X1 U4575 ( .A(n3652), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5300)
         );
  XNOR2_X1 U4576 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3662) );
  NAND2_X1 U4577 ( .A1(n3663), .A2(n3662), .ZN(n3654) );
  NAND2_X1 U4578 ( .A1(n6969), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U4579 ( .A1(n3654), .A2(n3653), .ZN(n3676) );
  XNOR2_X1 U4580 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4581 ( .A1(n3676), .A2(n3677), .ZN(n3656) );
  NAND2_X1 U4582 ( .A1(n4887), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4583 ( .A1(n3656), .A2(n3655), .ZN(n3686) );
  XNOR2_X1 U4584 ( .A(n5854), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3684)
         );
  NAND2_X1 U4585 ( .A1(n3686), .A2(n3684), .ZN(n3658) );
  NAND2_X1 U4586 ( .A1(n6641), .A2(n5854), .ZN(n3657) );
  NAND2_X1 U4587 ( .A1(n3658), .A2(n3657), .ZN(n3694) );
  NAND2_X1 U4588 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6029), .ZN(n3660) );
  XOR2_X1 U4589 ( .A(n3662), .B(n3663), .Z(n3710) );
  OAI21_X1 U4590 ( .B1(n3700), .B2(n4616), .A(n3719), .ZN(n3670) );
  AOI21_X1 U4591 ( .B1(n4616), .B2(n3719), .A(n3344), .ZN(n3680) );
  INV_X1 U4592 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6502) );
  AOI21_X1 U4593 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6502), .A(n3663), 
        .ZN(n3666) );
  INV_X1 U4594 ( .A(n3666), .ZN(n3665) );
  OAI21_X1 U4595 ( .B1(n3359), .B2(n3665), .A(n3664), .ZN(n3668) );
  NAND2_X1 U4596 ( .A1(n3678), .A2(n3666), .ZN(n3667) );
  AOI22_X1 U4597 ( .A1(n3680), .A2(n3668), .B1(n3667), .B2(n3701), .ZN(n3669)
         );
  OAI21_X1 U4598 ( .B1(n3710), .B2(n3670), .A(n3669), .ZN(n3675) );
  NAND3_X1 U4599 ( .A1(n3670), .A2(STATE2_REG_0__SCAN_IN), .A3(n3710), .ZN(
        n3674) );
  NAND3_X1 U4600 ( .A1(n3675), .A2(n3674), .A3(n3673), .ZN(n3693) );
  XOR2_X1 U4601 ( .A(n3677), .B(n3676), .Z(n3709) );
  NAND2_X1 U4602 ( .A1(n3678), .A2(n3709), .ZN(n3681) );
  OAI211_X1 U4603 ( .C1(n3709), .C2(n3679), .A(n3681), .B(n3680), .ZN(n3692)
         );
  INV_X1 U4604 ( .A(n3680), .ZN(n3683) );
  INV_X1 U4605 ( .A(n3681), .ZN(n3682) );
  INV_X1 U4606 ( .A(n3684), .ZN(n3685) );
  XNOR2_X1 U4607 ( .A(n3686), .B(n3685), .ZN(n3708) );
  INV_X1 U4608 ( .A(n3708), .ZN(n3687) );
  AOI21_X1 U4609 ( .B1(n3708), .B2(n3713), .A(n3695), .ZN(n3696) );
  OAI22_X1 U4610 ( .A1(n3697), .A2(n3696), .B1(n3701), .B2(n3713), .ZN(n3698)
         );
  OAI21_X1 U4611 ( .B1(n3712), .B2(n3700), .A(n3699), .ZN(n3703) );
  NAND2_X4 U4612 ( .A1(n3703), .A2(n3702), .ZN(n6521) );
  OR2_X1 U4613 ( .A1(n3705), .A2(STATE_REG_0__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U4614 ( .A1(n4616), .A2(n6563), .ZN(n4934) );
  INV_X1 U4615 ( .A(READY_N), .ZN(n4438) );
  NAND3_X1 U4616 ( .A1(n3112), .A2(n4934), .A3(n4438), .ZN(n3706) );
  NAND3_X1 U4617 ( .A1(n3706), .A2(n3111), .A3(n3854), .ZN(n3707) );
  NAND2_X1 U4618 ( .A1(n6521), .A2(n3707), .ZN(n3718) );
  NAND2_X1 U4619 ( .A1(n3735), .A2(n6563), .ZN(n3716) );
  NAND3_X1 U4620 ( .A1(n3710), .A2(n3709), .A3(n3708), .ZN(n3711) );
  NAND2_X1 U4621 ( .A1(n3712), .A2(n3711), .ZN(n3714) );
  NAND2_X1 U4622 ( .A1(n3714), .A2(n3713), .ZN(n6515) );
  NAND2_X1 U4623 ( .A1(n4438), .A2(n6515), .ZN(n4446) );
  INV_X1 U4624 ( .A(n4446), .ZN(n3715) );
  NAND2_X1 U4625 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  MUX2_X1 U4626 ( .A(n3718), .B(n3717), .S(n3855), .Z(n3730) );
  NAND2_X1 U4627 ( .A1(n5839), .A2(n3735), .ZN(n3727) );
  OR2_X1 U4628 ( .A1(n5839), .A2(n3734), .ZN(n3721) );
  NAND2_X1 U4629 ( .A1(n3720), .A2(n3721), .ZN(n3732) );
  NAND2_X1 U4630 ( .A1(n3722), .A2(n3734), .ZN(n3724) );
  MUX2_X1 U4631 ( .A(n3724), .B(n3723), .S(n3238), .Z(n4454) );
  INV_X1 U4632 ( .A(n4454), .ZN(n3726) );
  NAND2_X1 U4633 ( .A1(n3725), .A2(n4632), .ZN(n6516) );
  OAI21_X1 U4634 ( .B1(n3732), .B2(n3726), .A(n6516), .ZN(n4441) );
  OAI21_X1 U4635 ( .B1(n6521), .B2(n3727), .A(n4441), .ZN(n3728) );
  INV_X1 U4636 ( .A(n3728), .ZN(n3729) );
  NAND2_X1 U4637 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  INV_X1 U4638 ( .A(n3344), .ZN(n6034) );
  NOR2_X1 U4639 ( .A1(n3732), .A2(n6034), .ZN(n4460) );
  NAND4_X1 U4640 ( .A1(n3345), .A2(n3359), .A3(n3479), .A4(n3734), .ZN(n3888)
         );
  INV_X1 U4641 ( .A(n3888), .ZN(n6526) );
  NOR2_X1 U4642 ( .A1(n4460), .A2(n6526), .ZN(n6518) );
  AND2_X4 U4643 ( .A1(n3735), .A2(n3734), .ZN(n4940) );
  AOI22_X1 U4644 ( .A1(n3733), .A2(n3736), .B1(n3112), .B2(n4940), .ZN(n3738)
         );
  NAND3_X1 U4645 ( .A1(n6518), .A2(n3738), .A3(n3737), .ZN(n3739) );
  NAND2_X2 U4646 ( .A1(n3862), .A2(n3739), .ZN(n5984) );
  NAND2_X2 U4647 ( .A1(n3313), .A2(n4940), .ZN(n3835) );
  INV_X1 U4648 ( .A(n3750), .ZN(n3746) );
  INV_X1 U4649 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4650 ( .A1(n3750), .A2(n3741), .ZN(n3743) );
  INV_X1 U4651 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U4652 ( .A1(n4940), .A2(n5189), .ZN(n3742) );
  NAND3_X1 U4653 ( .A1(n3743), .A2(n3837), .A3(n3742), .ZN(n3744) );
  NAND2_X2 U4654 ( .A1(n3745), .A2(n3744), .ZN(n3749) );
  NAND2_X1 U4655 ( .A1(n3750), .A2(EBX_REG_0__SCAN_IN), .ZN(n3748) );
  INV_X1 U4656 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U4657 ( .A1(n3837), .A2(n6821), .ZN(n3747) );
  XNOR2_X2 U4658 ( .A(n3749), .B(n4430), .ZN(n4418) );
  OAI22_X1 U4659 ( .A1(n4418), .A2(n5336), .B1(n4430), .B2(n3749), .ZN(n4476)
         );
  MUX2_X1 U4660 ( .A(n3835), .B(n3750), .S(EBX_REG_2__SCAN_IN), .Z(n3752) );
  NAND2_X1 U4661 ( .A1(n3746), .A2(n5336), .ZN(n3818) );
  NAND2_X1 U4662 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5336), .ZN(n3751)
         );
  MUX2_X1 U4663 ( .A(n5331), .B(n3837), .S(EBX_REG_3__SCAN_IN), .Z(n3755) );
  OAI21_X1 U4664 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5337), .A(n3755), 
        .ZN(n4492) );
  OR2_X1 U4665 ( .A1(n3835), .A2(EBX_REG_4__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4666 ( .A1(n3750), .A2(n3756), .ZN(n3758) );
  INV_X1 U4667 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U4668 ( .A1(n4940), .A2(n6144), .ZN(n3757) );
  NAND3_X1 U4669 ( .A1(n3758), .A2(n3837), .A3(n3757), .ZN(n3759) );
  NAND2_X1 U4670 ( .A1(n3760), .A2(n3759), .ZN(n4568) );
  NAND2_X1 U4671 ( .A1(n4490), .A2(n4568), .ZN(n4570) );
  MUX2_X1 U4672 ( .A(n5331), .B(n3837), .S(EBX_REG_5__SCAN_IN), .Z(n3761) );
  OAI21_X1 U4673 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5337), .A(n3761), 
        .ZN(n4516) );
  MUX2_X1 U4674 ( .A(n3835), .B(n3750), .S(EBX_REG_6__SCAN_IN), .Z(n3765) );
  NAND2_X1 U4675 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3764)
         );
  OR2_X2 U4676 ( .A1(n4771), .A2(n4770), .ZN(n4923) );
  MUX2_X1 U4677 ( .A(n5331), .B(n3837), .S(EBX_REG_7__SCAN_IN), .Z(n3766) );
  OAI21_X1 U4678 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5337), .A(n3766), 
        .ZN(n4922) );
  NOR2_X4 U4679 ( .A1(n4923), .A2(n4922), .ZN(n5184) );
  MUX2_X1 U4680 ( .A(n3835), .B(n3750), .S(EBX_REG_8__SCAN_IN), .Z(n3769) );
  NAND2_X1 U4681 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3767)
         );
  AND2_X1 U4682 ( .A1(n3818), .A2(n3767), .ZN(n3768) );
  MUX2_X1 U4683 ( .A(n5331), .B(n3837), .S(EBX_REG_9__SCAN_IN), .Z(n3770) );
  OAI21_X1 U4684 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5337), .A(n3770), 
        .ZN(n5187) );
  NOR2_X1 U4685 ( .A1(n5182), .A2(n5187), .ZN(n3771) );
  MUX2_X1 U4686 ( .A(n3835), .B(n3750), .S(EBX_REG_10__SCAN_IN), .Z(n3773) );
  NAND2_X1 U4687 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3772) );
  INV_X1 U4689 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U4690 ( .A1(n4940), .A2(n5231), .ZN(n3775) );
  NAND2_X1 U4691 ( .A1(n3837), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3774) );
  NAND3_X1 U4692 ( .A1(n3775), .A2(n3750), .A3(n3774), .ZN(n3776) );
  OAI21_X1 U4693 ( .B1(n5331), .B2(EBX_REG_11__SCAN_IN), .A(n3776), .ZN(n5222)
         );
  NOR2_X4 U4694 ( .A1(n5262), .A2(n5222), .ZN(n6009) );
  INV_X1 U4695 ( .A(n5331), .ZN(n3812) );
  INV_X1 U4696 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U4697 ( .A1(n3812), .A2(n6965), .ZN(n3780) );
  NAND2_X1 U4698 ( .A1(n4940), .A2(n6965), .ZN(n3778) );
  NAND2_X1 U4699 ( .A1(n3837), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3777) );
  NAND3_X1 U4700 ( .A1(n3778), .A2(n3750), .A3(n3777), .ZN(n3779) );
  AND2_X1 U4701 ( .A1(n3780), .A2(n3779), .ZN(n6007) );
  OR2_X1 U4702 ( .A1(n3835), .A2(EBX_REG_12__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4703 ( .A1(n3750), .A2(n6752), .ZN(n3782) );
  INV_X1 U4704 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U4705 ( .A1(n4940), .A2(n6964), .ZN(n3781) );
  NAND3_X1 U4706 ( .A1(n3782), .A2(n3837), .A3(n3781), .ZN(n3783) );
  NAND2_X1 U4707 ( .A1(n3784), .A2(n3783), .ZN(n6008) );
  AND2_X1 U4708 ( .A1(n6007), .A2(n6008), .ZN(n3785) );
  AND2_X2 U4709 ( .A1(n6009), .A2(n3785), .ZN(n6010) );
  NAND2_X1 U4710 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3786) );
  AND2_X1 U4711 ( .A1(n3818), .A2(n3786), .ZN(n3788) );
  MUX2_X1 U4712 ( .A(n3835), .B(n3750), .S(EBX_REG_14__SCAN_IN), .Z(n3787) );
  NAND2_X1 U4713 ( .A1(n3788), .A2(n3787), .ZN(n5442) );
  INV_X1 U4714 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U4715 ( .A1(n4940), .A2(n5531), .ZN(n3790) );
  NAND2_X1 U4716 ( .A1(n3837), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3789) );
  NAND3_X1 U4717 ( .A1(n3790), .A2(n3750), .A3(n3789), .ZN(n3791) );
  OAI21_X1 U4718 ( .B1(n5331), .B2(EBX_REG_15__SCAN_IN), .A(n3791), .ZN(n5431)
         );
  NOR2_X2 U4719 ( .A1(n5441), .A2(n5431), .ZN(n5430) );
  MUX2_X1 U4720 ( .A(n3835), .B(n3750), .S(EBX_REG_16__SCAN_IN), .Z(n3793) );
  NAND2_X1 U4721 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3792) );
  AND3_X1 U4722 ( .A1(n3793), .A2(n3818), .A3(n3792), .ZN(n5523) );
  INV_X1 U4723 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U4724 ( .A1(n3812), .A2(n6766), .ZN(n3798) );
  NAND2_X1 U4725 ( .A1(n4940), .A2(n6766), .ZN(n3796) );
  NAND2_X1 U4726 ( .A1(n3837), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3795) );
  NAND3_X1 U4727 ( .A1(n3796), .A2(n3750), .A3(n3795), .ZN(n3797) );
  AND2_X1 U4728 ( .A1(n3798), .A2(n3797), .ZN(n5417) );
  AND2_X2 U4729 ( .A1(n3154), .A2(n5417), .ZN(n5517) );
  OR2_X1 U4730 ( .A1(n3835), .A2(EBX_REG_19__SCAN_IN), .ZN(n3802) );
  INV_X1 U4731 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U4732 ( .A1(n3750), .A2(n5597), .ZN(n3800) );
  INV_X1 U4733 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U4734 ( .A1(n4940), .A2(n5510), .ZN(n3799) );
  NAND3_X1 U4735 ( .A1(n3800), .A2(n3837), .A3(n3799), .ZN(n3801) );
  NAND2_X1 U4736 ( .A1(n3802), .A2(n3801), .ZN(n5405) );
  NAND2_X1 U4737 ( .A1(n5517), .A2(n5405), .ZN(n5504) );
  INV_X1 U4738 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5508) );
  NOR2_X1 U4739 ( .A1(n3837), .A2(n5508), .ZN(n3806) );
  OAI22_X1 U4740 ( .A1(n5337), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n5336), .B2(EBX_REG_20__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U4741 ( .A1(n5337), .A2(EBX_REG_18__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4742 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4743 ( .A1(n3804), .A2(n3803), .ZN(n5505) );
  MUX2_X1 U4744 ( .A(n3837), .B(n5507), .S(n5505), .Z(n3805) );
  INV_X1 U4745 ( .A(n3807), .ZN(n5497) );
  OR2_X1 U4746 ( .A1(n3835), .A2(EBX_REG_21__SCAN_IN), .ZN(n3811) );
  INV_X1 U4747 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U4748 ( .A1(n3750), .A2(n5779), .ZN(n3809) );
  INV_X1 U4749 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U4750 ( .A1(n4940), .A2(n5944), .ZN(n3808) );
  NAND3_X1 U4751 ( .A1(n3809), .A2(n3837), .A3(n3808), .ZN(n3810) );
  AND2_X1 U4752 ( .A1(n3811), .A2(n3810), .ZN(n5496) );
  INV_X1 U4753 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U4754 ( .A1(n3812), .A2(n5492), .ZN(n3816) );
  NAND2_X1 U4755 ( .A1(n4940), .A2(n5492), .ZN(n3814) );
  NAND2_X1 U4756 ( .A1(n3837), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3813) );
  NAND3_X1 U4757 ( .A1(n3814), .A2(n3750), .A3(n3813), .ZN(n3815) );
  AND2_X1 U4758 ( .A1(n3816), .A2(n3815), .ZN(n5485) );
  AND2_X2 U4759 ( .A1(n5495), .A2(n5485), .ZN(n5487) );
  NAND2_X1 U4760 ( .A1(n5336), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3817) );
  AND2_X1 U4761 ( .A1(n3818), .A2(n3817), .ZN(n3820) );
  MUX2_X1 U4762 ( .A(n3835), .B(n3750), .S(EBX_REG_23__SCAN_IN), .Z(n3819) );
  NAND2_X1 U4763 ( .A1(n3820), .A2(n3819), .ZN(n5388) );
  MUX2_X1 U4764 ( .A(n5331), .B(n3837), .S(EBX_REG_25__SCAN_IN), .Z(n3821) );
  OAI21_X1 U4765 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5337), .A(n3821), 
        .ZN(n5474) );
  INV_X1 U4766 ( .A(n5474), .ZN(n3827) );
  OR2_X1 U4767 ( .A1(n3835), .A2(EBX_REG_24__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4768 ( .A1(n3750), .A2(n3822), .ZN(n3824) );
  INV_X1 U4769 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U4770 ( .A1(n4940), .A2(n5482), .ZN(n3823) );
  NAND3_X1 U4771 ( .A1(n3824), .A2(n3837), .A3(n3823), .ZN(n3825) );
  NAND2_X1 U4772 ( .A1(n3826), .A2(n3825), .ZN(n5473) );
  NAND2_X1 U4773 ( .A1(n3827), .A2(n5473), .ZN(n3828) );
  OR2_X1 U4774 ( .A1(n3835), .A2(EBX_REG_26__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4775 ( .A1(n3750), .A2(n6684), .ZN(n3830) );
  INV_X1 U4776 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U4777 ( .A1(n4940), .A2(n5469), .ZN(n3829) );
  NAND3_X1 U4778 ( .A1(n3830), .A2(n3837), .A3(n3829), .ZN(n3831) );
  NAND2_X1 U4779 ( .A1(n3832), .A2(n3831), .ZN(n5368) );
  NAND2_X1 U4780 ( .A1(n5472), .A2(n5368), .ZN(n5367) );
  MUX2_X1 U4781 ( .A(n5331), .B(n3837), .S(EBX_REG_27__SCAN_IN), .Z(n3833) );
  OAI21_X1 U4782 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5337), .A(n3833), 
        .ZN(n5462) );
  INV_X1 U4783 ( .A(n3834), .ZN(n5456) );
  OR2_X1 U4784 ( .A1(n3835), .A2(EBX_REG_28__SCAN_IN), .ZN(n3840) );
  INV_X1 U4785 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U4786 ( .A1(n3750), .A2(n5724), .ZN(n3838) );
  INV_X1 U4787 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U4788 ( .A1(n4940), .A2(n5906), .ZN(n3836) );
  NAND3_X1 U4789 ( .A1(n3838), .A2(n3837), .A3(n3836), .ZN(n3839) );
  AND2_X1 U4790 ( .A1(n3840), .A2(n3839), .ZN(n5457) );
  INV_X1 U4791 ( .A(n5459), .ZN(n3844) );
  NOR2_X1 U4792 ( .A1(n5337), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5330)
         );
  INV_X1 U4793 ( .A(EBX_REG_29__SCAN_IN), .ZN(n3841) );
  NOR3_X4 U4794 ( .A1(n5459), .A2(n5330), .A3(n3842), .ZN(n3845) );
  INV_X1 U4795 ( .A(n3845), .ZN(n3843) );
  AOI22_X1 U4796 ( .A1(n5337), .A2(EBX_REG_30__SCAN_IN), .B1(n5336), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5335) );
  NOR2_X1 U4797 ( .A1(n3845), .A2(n3313), .ZN(n5334) );
  AOI211_X2 U4798 ( .C1(n3844), .C2(n3843), .A(n5335), .B(n5334), .ZN(n3848)
         );
  INV_X1 U4799 ( .A(n5335), .ZN(n3846) );
  AOI211_X1 U4800 ( .C1(n3313), .C2(n5459), .A(n3846), .B(n3845), .ZN(n3847)
         );
  NOR2_X1 U4801 ( .A1(n3848), .A2(n3847), .ZN(n5322) );
  NAND2_X1 U4802 ( .A1(n3733), .A2(n3323), .ZN(n3849) );
  NAND2_X1 U4803 ( .A1(n3112), .A2(n6658), .ZN(n6536) );
  AND2_X1 U4804 ( .A1(n3849), .A2(n6536), .ZN(n3850) );
  NOR2_X2 U4805 ( .A1(n3870), .A2(n3850), .ZN(n6312) );
  NOR2_X1 U4806 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5024) );
  NOR2_X1 U4807 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n3851) );
  AND2_X2 U4808 ( .A1(n5024), .A2(n3851), .ZN(n6276) );
  NAND2_X1 U4809 ( .A1(n6276), .A2(REIP_REG_30__SCAN_IN), .ZN(n5293) );
  INV_X1 U4810 ( .A(n5293), .ZN(n3868) );
  INV_X1 U4811 ( .A(n3852), .ZN(n3869) );
  AND2_X1 U4812 ( .A1(n3479), .A2(n4940), .ZN(n3853) );
  NAND4_X1 U4813 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4814 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U4815 ( .A1(n3498), .A2(n4478), .ZN(n4576) );
  NAND3_X1 U4816 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n4576), .ZN(n4696) );
  NOR2_X1 U4817 ( .A1(n3863), .A2(n4696), .ZN(n4879) );
  NAND2_X1 U4818 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4879), .ZN(n5170)
         );
  NOR2_X1 U4819 ( .A1(n3864), .A2(n5170), .ZN(n3874) );
  INV_X1 U4820 ( .A(n6503), .ZN(n5285) );
  NAND2_X1 U4821 ( .A1(n3862), .A2(n5285), .ZN(n6318) );
  INV_X1 U4822 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U4823 ( .A1(n3362), .A2(n3313), .B1(n3855), .B2(n3854), .ZN(n3857)
         );
  NOR2_X1 U4824 ( .A1(n4936), .A2(n3855), .ZN(n4439) );
  OAI21_X1 U4825 ( .B1(n4439), .B2(n5337), .A(n3332), .ZN(n3856) );
  AND2_X1 U4826 ( .A1(n3857), .A2(n3856), .ZN(n3858) );
  NAND2_X1 U4827 ( .A1(n3859), .A2(n3858), .ZN(n4458) );
  OAI211_X1 U4828 ( .C1(n4452), .C2(n3111), .A(n4454), .B(n4533), .ZN(n3860)
         );
  OR2_X1 U4829 ( .A1(n4458), .A2(n3860), .ZN(n3861) );
  NAND2_X1 U4830 ( .A1(n3862), .A2(n3861), .ZN(n3871) );
  NOR2_X1 U4831 ( .A1(n6320), .A2(n3871), .ZN(n5817) );
  NAND4_X1 U4832 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4698) );
  OR3_X1 U4833 ( .A1(n4878), .A2(n3863), .A3(n4698), .ZN(n5166) );
  NOR2_X1 U4834 ( .A1(n5166), .A2(n3864), .ZN(n6012) );
  INV_X1 U4835 ( .A(n6012), .ZN(n3872) );
  NOR2_X1 U4836 ( .A1(n4699), .A2(n3872), .ZN(n5830) );
  NAND2_X1 U4837 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5820) );
  NOR2_X1 U4838 ( .A1(n6023), .A2(n5820), .ZN(n5825) );
  NAND2_X1 U4839 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5825), .ZN(n3875) );
  NAND3_X1 U4840 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5812), .ZN(n5997) );
  INV_X1 U4841 ( .A(n5997), .ZN(n3865) );
  NAND2_X1 U4842 ( .A1(n3869), .A2(n3865), .ZN(n5793) );
  NOR2_X1 U4843 ( .A1(n5793), .A2(n5609), .ZN(n5766) );
  INV_X1 U4844 ( .A(n3880), .ZN(n3866) );
  NAND2_X1 U4845 ( .A1(n5766), .A2(n3866), .ZN(n5738) );
  NAND2_X1 U4846 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5739) );
  NOR2_X1 U4847 ( .A1(n5738), .A2(n5739), .ZN(n5731) );
  NAND2_X1 U4848 ( .A1(n5731), .A2(n3146), .ZN(n5715) );
  NOR3_X1 U4849 ( .A1(n5715), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n3647), 
        .ZN(n3867) );
  NAND2_X1 U4850 ( .A1(n4697), .A2(n3871), .ZN(n5821) );
  INV_X1 U4851 ( .A(n5739), .ZN(n3881) );
  NAND2_X1 U4852 ( .A1(n4699), .A2(n4697), .ZN(n5791) );
  NAND2_X1 U4853 ( .A1(n3869), .A2(n5795), .ZN(n3877) );
  NOR2_X1 U4854 ( .A1(n6898), .A2(n6850), .ZN(n3876) );
  NAND2_X1 U4855 ( .A1(n3871), .A2(n6318), .ZN(n5167) );
  NAND2_X1 U4856 ( .A1(n5829), .A2(n3870), .ZN(n6319) );
  OAI21_X1 U4857 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n3871), .A(n6319), 
        .ZN(n5168) );
  AOI21_X1 U4858 ( .B1(n5167), .B2(n3872), .A(n5168), .ZN(n3873) );
  OAI21_X1 U4859 ( .B1(n3874), .B2(n4697), .A(n3873), .ZN(n6286) );
  AOI21_X1 U4860 ( .B1(n3875), .B2(n3878), .A(n6286), .ZN(n6001) );
  OAI21_X1 U4861 ( .B1(n5792), .B2(n3876), .A(n6001), .ZN(n5990) );
  AOI21_X1 U4862 ( .B1(n3878), .B2(n3877), .A(n5990), .ZN(n5778) );
  OAI21_X1 U4863 ( .B1(n3879), .B2(n5792), .A(n5778), .ZN(n5771) );
  AOI21_X1 U4864 ( .B1(n3880), .B2(n5791), .A(n5771), .ZN(n5759) );
  OAI21_X1 U4865 ( .B1(n5792), .B2(n3881), .A(n5759), .ZN(n5735) );
  NOR2_X1 U4866 ( .A1(n5735), .A2(n3882), .ZN(n5718) );
  NAND2_X1 U4867 ( .A1(n5718), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U4868 ( .A1(n5759), .A2(n5792), .ZN(n5716) );
  NAND3_X1 U4869 ( .A1(n5710), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5716), .ZN(n3883) );
  AND2_X1 U4870 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  OAI21_X1 U4871 ( .B1(n5300), .B2(n5984), .A(n3885), .ZN(U2988) );
  INV_X1 U4872 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U4873 ( .A1(n3648), .A2(n3148), .ZN(n3886) );
  AND2_X1 U4874 ( .A1(n6630), .A2(n3889), .ZN(n6663) );
  OR2_X1 U4875 ( .A1(n6663), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4876 ( .A1(n6660), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3892) );
  INV_X1 U4877 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6657) );
  NAND2_X1 U4878 ( .A1(n6657), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3891) );
  NAND2_X1 U4879 ( .A1(n3892), .A2(n3891), .ZN(n6279) );
  NAND2_X2 U4880 ( .A1(n6266), .A2(n6279), .ZN(n6272) );
  INV_X1 U4881 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5444) );
  INV_X1 U4882 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5419) );
  INV_X1 U4883 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U4884 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3895) );
  NAND2_X1 U4885 ( .A1(n4286), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4306)
         );
  INV_X1 U4886 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4305) );
  INV_X1 U4887 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4330) );
  INV_X1 U4888 ( .A(n4387), .ZN(n3897) );
  NAND2_X1 U4889 ( .A1(n3897), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3898)
         );
  XNOR2_X1 U4890 ( .A(n3898), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4950)
         );
  INV_X1 U4891 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U4892 ( .A1(n6276), .A2(REIP_REG_31__SCAN_IN), .ZN(n5705) );
  OAI21_X1 U4893 ( .B1(n6266), .B2(n6754), .A(n5705), .ZN(n3899) );
  AOI21_X1 U4894 ( .B1(n6258), .B2(n4950), .A(n3899), .ZN(n4397) );
  NAND2_X1 U4895 ( .A1(n3901), .A2(n4065), .ZN(n3907) );
  NOR2_X2 U4896 ( .A1(n3337), .A2(n6656), .ZN(n3912) );
  INV_X1 U4897 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3904) );
  INV_X2 U4898 ( .A(n4357), .ZN(n4931) );
  OAI21_X1 U4899 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3902), .A(n3973), 
        .ZN(n6117) );
  NAND2_X1 U4900 ( .A1(n6656), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4901 ( .A1(n4931), .A2(n6117), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3903) );
  NAND2_X1 U4902 ( .A1(n3907), .A2(n3906), .ZN(n4926) );
  NAND2_X1 U4903 ( .A1(n4558), .A2(n4065), .ZN(n3908) );
  NAND2_X1 U4904 ( .A1(n3908), .A2(n3925), .ZN(n4495) );
  NAND2_X1 U4905 ( .A1(n6325), .A2(n3909), .ZN(n3910) );
  INV_X1 U4906 ( .A(n3911), .ZN(n6436) );
  AND2_X1 U4907 ( .A1(n3345), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3923) );
  INV_X1 U4908 ( .A(n3923), .ZN(n3945) );
  NAND2_X1 U4909 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6656), .ZN(n3914)
         );
  NAND2_X1 U4910 ( .A1(n3912), .A2(EAX_REG_0__SCAN_IN), .ZN(n3913) );
  OAI211_X1 U4911 ( .C1(n3945), .C2(n6502), .A(n3914), .B(n3913), .ZN(n3915)
         );
  AOI21_X1 U4912 ( .B1(n6436), .B2(n4065), .A(n3915), .ZN(n4425) );
  NAND2_X1 U4913 ( .A1(n4425), .A2(n4931), .ZN(n3918) );
  NAND2_X1 U4914 ( .A1(n4552), .A2(n4065), .ZN(n3922) );
  NAND2_X1 U4915 ( .A1(n3923), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3920) );
  INV_X1 U4916 ( .A(n4326), .ZN(n4386) );
  AOI22_X1 U4917 ( .A1(n4386), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6656), .ZN(n3919) );
  AND2_X1 U4918 ( .A1(n3920), .A2(n3919), .ZN(n3921) );
  NAND2_X1 U4919 ( .A1(n3922), .A2(n3921), .ZN(n4408) );
  NAND2_X1 U4920 ( .A1(n4407), .A2(n4408), .ZN(n4406) );
  NAND2_X1 U4921 ( .A1(n3923), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3928) );
  INV_X1 U4922 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U4923 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3935) );
  OAI21_X1 U4924 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3935), .ZN(n6273) );
  NAND2_X1 U4925 ( .A1(n6273), .A2(n4931), .ZN(n3924) );
  OAI21_X1 U4926 ( .B1(n6945), .B2(n3925), .A(n3924), .ZN(n3926) );
  AOI21_X1 U4927 ( .B1(n4386), .B2(EAX_REG_2__SCAN_IN), .A(n3926), .ZN(n3927)
         );
  AND2_X1 U4928 ( .A1(n3928), .A2(n3927), .ZN(n3929) );
  NAND2_X1 U4929 ( .A1(n4495), .A2(n4494), .ZN(n3933) );
  INV_X1 U4930 ( .A(n4406), .ZN(n3931) );
  INV_X1 U4931 ( .A(n3929), .ZN(n3930) );
  INV_X1 U4932 ( .A(n3934), .ZN(n3947) );
  INV_X1 U4933 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U4934 ( .A1(n6946), .A2(n3935), .ZN(n3936) );
  NAND2_X1 U4935 ( .A1(n3947), .A2(n3936), .ZN(n5200) );
  AOI22_X1 U4936 ( .A1(n5200), .A2(n4931), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U4937 ( .A1(n4386), .A2(EAX_REG_3__SCAN_IN), .ZN(n3937) );
  OAI211_X1 U4938 ( .C1(n3945), .C2(n3157), .A(n3938), .B(n3937), .ZN(n3939)
         );
  INV_X1 U4939 ( .A(n3939), .ZN(n3940) );
  INV_X1 U4940 ( .A(n3941), .ZN(n3942) );
  NAND2_X1 U4941 ( .A1(n3942), .A2(n4065), .ZN(n3953) );
  NAND2_X1 U4942 ( .A1(n6656), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3944)
         );
  NAND2_X1 U4943 ( .A1(n4386), .A2(EAX_REG_4__SCAN_IN), .ZN(n3943) );
  OAI211_X1 U4944 ( .C1(n3945), .C2(n6029), .A(n3944), .B(n3943), .ZN(n3951)
         );
  INV_X1 U4945 ( .A(n3954), .ZN(n3949) );
  INV_X1 U4946 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4947 ( .A1(n3947), .A2(n3946), .ZN(n3948) );
  NAND2_X1 U4948 ( .A1(n3949), .A2(n3948), .ZN(n6257) );
  AND2_X1 U4949 ( .A1(n6257), .A2(n4931), .ZN(n3950) );
  AOI21_X1 U4950 ( .B1(n3951), .B2(n4357), .A(n3950), .ZN(n3952) );
  AND2_X2 U4951 ( .A1(n4487), .A2(n4566), .ZN(n4511) );
  OAI21_X1 U4952 ( .B1(n3954), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3958), 
        .ZN(n6130) );
  AOI22_X1 U4953 ( .A1(n6130), .A2(n4931), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3956) );
  NAND2_X1 U4954 ( .A1(n4386), .A2(EAX_REG_5__SCAN_IN), .ZN(n3955) );
  NAND2_X1 U4955 ( .A1(n4511), .A2(n4514), .ZN(n4513) );
  NAND2_X1 U4956 ( .A1(n4386), .A2(EAX_REG_6__SCAN_IN), .ZN(n3960) );
  OAI21_X1 U4957 ( .B1(n6657), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6656), 
        .ZN(n3959) );
  XNOR2_X1 U4958 ( .A(n3958), .B(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U4959 ( .A1(n3960), .A2(n3959), .B1(n4931), .B2(n4915), .ZN(n3961)
         );
  NAND2_X1 U4960 ( .A1(n4926), .A2(n4762), .ZN(n4925) );
  AOI22_X1 U4961 ( .A1(n4522), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4962 ( .A1(n4359), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4963 ( .A1(n4367), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4964 ( .A1(n4187), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3963) );
  NAND4_X1 U4965 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3972)
         );
  AOI22_X1 U4966 ( .A1(n4366), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4967 ( .A1(n4311), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4968 ( .A1(n4360), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4969 ( .A1(n4361), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3967) );
  NAND4_X1 U4970 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3971)
         );
  OAI21_X1 U4971 ( .B1(n3972), .B2(n3971), .A(n4065), .ZN(n3976) );
  XOR2_X1 U4972 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3973), .Z(n5212) );
  AOI22_X1 U4973 ( .A1(n4931), .A2(n5212), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3975) );
  NAND2_X1 U4974 ( .A1(n4386), .A2(EAX_REG_8__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4975 ( .A1(n4522), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4976 ( .A1(n4369), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4977 ( .A1(n4360), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4978 ( .A1(n4366), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4979 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3987)
         );
  AOI22_X1 U4980 ( .A1(n4311), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4981 ( .A1(n4187), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4361), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4982 ( .A1(n4367), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4983 ( .A1(n4372), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4984 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  OAI21_X1 U4985 ( .B1(n3987), .B2(n3986), .A(n4065), .ZN(n3991) );
  XNOR2_X1 U4986 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3988), .ZN(n5248) );
  AOI22_X1 U4987 ( .A1(n4931), .A2(n5248), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3990) );
  NAND2_X1 U4988 ( .A1(n3912), .A2(EAX_REG_9__SCAN_IN), .ZN(n3989) );
  XOR2_X1 U4989 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3992), .Z(n6098) );
  INV_X1 U4990 ( .A(n6098), .ZN(n5257) );
  AOI22_X1 U4991 ( .A1(n3446), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4992 ( .A1(n4369), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4993 ( .A1(n4360), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4361), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4994 ( .A1(n4366), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4995 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4002)
         );
  AOI22_X1 U4996 ( .A1(n4367), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4522), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4997 ( .A1(n4311), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4998 ( .A1(n4359), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4999 ( .A1(n4372), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U5000 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  NOR2_X1 U5001 ( .A1(n4002), .A2(n4001), .ZN(n4005) );
  NAND2_X1 U5002 ( .A1(n3912), .A2(EAX_REG_10__SCAN_IN), .ZN(n4004) );
  NAND2_X1 U5003 ( .A1(n4391), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4003)
         );
  OAI211_X1 U5004 ( .C1(n4084), .C2(n4005), .A(n4004), .B(n4003), .ZN(n4006)
         );
  AOI21_X1 U5005 ( .B1(n5257), .B2(n4931), .A(n4006), .ZN(n5243) );
  AOI22_X1 U5006 ( .A1(n4367), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4522), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5007 ( .A1(n3446), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5008 ( .A1(n4311), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4360), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5009 ( .A1(n4361), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U5010 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4016)
         );
  AOI22_X1 U5011 ( .A1(n4369), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5012 ( .A1(n4368), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5013 ( .A1(n4366), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U5014 ( .A1(n4372), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U5015 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  NOR2_X1 U5016 ( .A1(n4016), .A2(n4015), .ZN(n4020) );
  XNOR2_X1 U5017 ( .A(n4017), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5700)
         );
  NAND2_X1 U5018 ( .A1(n5700), .A2(n4931), .ZN(n4019) );
  AOI22_X1 U5019 ( .A1(n3912), .A2(EAX_REG_11__SCAN_IN), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4018) );
  OAI211_X1 U5020 ( .C1(n4020), .C2(n4084), .A(n4019), .B(n4018), .ZN(n5221)
         );
  NAND2_X1 U5021 ( .A1(n5219), .A2(n5221), .ZN(n5220) );
  INV_X1 U5022 ( .A(n5220), .ZN(n4037) );
  XNOR2_X1 U5023 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4021), .ZN(n6090)
         );
  INV_X1 U5024 ( .A(n6090), .ZN(n5692) );
  AOI22_X1 U5025 ( .A1(n4367), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5026 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4369), .B1(n4360), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5027 ( .A1(n4359), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5028 ( .A1(n3446), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U5029 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4031)
         );
  AOI22_X1 U5030 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4311), .B1(n4368), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5031 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4361), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5032 ( .A1(n4522), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5033 ( .A1(n4372), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U5034 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4030)
         );
  NOR2_X1 U5035 ( .A1(n4031), .A2(n4030), .ZN(n4034) );
  NAND2_X1 U5036 ( .A1(n3912), .A2(EAX_REG_12__SCAN_IN), .ZN(n4033) );
  NAND2_X1 U5037 ( .A1(n4391), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4032)
         );
  OAI211_X1 U5038 ( .C1(n4084), .C2(n4034), .A(n4033), .B(n4032), .ZN(n4035)
         );
  AOI21_X1 U5039 ( .B1(n5692), .B2(n4931), .A(n4035), .ZN(n5273) );
  NAND2_X1 U5040 ( .A1(n4037), .A2(n4036), .ZN(n5270) );
  XNOR2_X1 U5041 ( .A(n4038), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6078)
         );
  AOI22_X1 U5042 ( .A1(n4522), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5043 ( .A1(n4360), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5044 ( .A1(n4366), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5045 ( .A1(n4361), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U5046 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4048)
         );
  AOI22_X1 U5047 ( .A1(n4367), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5048 ( .A1(n4311), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5049 ( .A1(n4368), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5050 ( .A1(n4369), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4043) );
  NAND4_X1 U5051 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(n4047)
         );
  NOR2_X1 U5052 ( .A1(n4048), .A2(n4047), .ZN(n4051) );
  NAND2_X1 U5053 ( .A1(n3912), .A2(EAX_REG_13__SCAN_IN), .ZN(n4050) );
  NAND2_X1 U5054 ( .A1(n4391), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4049)
         );
  OAI211_X1 U5055 ( .C1(n4084), .C2(n4051), .A(n4050), .B(n4049), .ZN(n4052)
         );
  AOI21_X1 U5056 ( .B1(n6078), .B2(n4931), .A(n4052), .ZN(n5560) );
  XNOR2_X1 U5057 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4053), .ZN(n5678)
         );
  AOI22_X1 U5058 ( .A1(n4522), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5059 ( .A1(n4311), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5060 ( .A1(n4369), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4361), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5061 ( .A1(n4372), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U5062 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4063)
         );
  AOI22_X1 U5063 ( .A1(n4367), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5064 ( .A1(n4368), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5065 ( .A1(n4360), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5066 ( .A1(n3412), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5067 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4062)
         );
  OR2_X1 U5068 ( .A1(n4063), .A2(n4062), .ZN(n4064) );
  AOI22_X1 U5069 ( .A1(n4065), .A2(n4064), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4067) );
  NAND2_X1 U5070 ( .A1(n3912), .A2(EAX_REG_14__SCAN_IN), .ZN(n4066) );
  OAI211_X1 U5071 ( .C1(n5678), .C2(n4357), .A(n4067), .B(n4066), .ZN(n5440)
         );
  NAND2_X1 U5072 ( .A1(n4068), .A2(n6856), .ZN(n4070) );
  INV_X1 U5073 ( .A(n4098), .ZN(n4069) );
  NAND2_X1 U5074 ( .A1(n4070), .A2(n4069), .ZN(n5669) );
  NAND2_X1 U5075 ( .A1(n5669), .A2(n4931), .ZN(n4087) );
  AOI22_X1 U5076 ( .A1(n4367), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4522), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5077 ( .A1(n4311), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4360), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5078 ( .A1(n4361), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5079 ( .A1(n3446), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U5080 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4080)
         );
  AOI22_X1 U5081 ( .A1(n4368), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5082 ( .A1(n4369), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5083 ( .A1(n4366), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5084 ( .A1(n4372), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5085 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  NOR2_X1 U5086 ( .A1(n4080), .A2(n4079), .ZN(n4083) );
  NAND2_X1 U5087 ( .A1(n3912), .A2(EAX_REG_15__SCAN_IN), .ZN(n4082) );
  NAND2_X1 U5088 ( .A1(n4391), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4081)
         );
  OAI211_X1 U5089 ( .C1(n4084), .C2(n4083), .A(n4082), .B(n4081), .ZN(n4085)
         );
  INV_X1 U5090 ( .A(n4085), .ZN(n4086) );
  NAND2_X1 U5091 ( .A1(n4087), .A2(n4086), .ZN(n5427) );
  AOI22_X1 U5092 ( .A1(n4360), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5093 ( .A1(n4366), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5094 ( .A1(n4311), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5095 ( .A1(n3447), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5096 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4097)
         );
  AOI22_X1 U5097 ( .A1(n4522), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5098 ( .A1(n4368), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5099 ( .A1(n4367), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5100 ( .A1(n4361), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4092) );
  NAND4_X1 U5101 ( .A1(n4095), .A2(n4094), .A3(n4093), .A4(n4092), .ZN(n4096)
         );
  OR2_X1 U5102 ( .A1(n4097), .A2(n4096), .ZN(n4102) );
  INV_X1 U5103 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4100) );
  XOR2_X1 U5104 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4098), .Z(n6065) );
  INV_X1 U5105 ( .A(n6065), .ZN(n5664) );
  AOI22_X1 U5106 ( .A1(n4931), .A2(n5664), .B1(n4391), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4099) );
  OAI21_X1 U5107 ( .B1(n4326), .B2(n4100), .A(n4099), .ZN(n4101) );
  AOI21_X1 U5108 ( .B1(n4383), .B2(n4102), .A(n4101), .ZN(n5526) );
  AOI22_X1 U5109 ( .A1(n4311), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5110 ( .A1(n4360), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5111 ( .A1(n4361), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5112 ( .A1(n4372), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5113 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4112)
         );
  AOI22_X1 U5114 ( .A1(n4367), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5115 ( .A1(n4368), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5116 ( .A1(n3446), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5117 ( .A1(n4522), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U5118 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4111)
         );
  NOR2_X1 U5119 ( .A1(n4112), .A2(n4111), .ZN(n4115) );
  AOI21_X1 U5120 ( .B1(n5419), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4113) );
  AOI21_X1 U5121 ( .B1(n3912), .B2(EAX_REG_17__SCAN_IN), .A(n4113), .ZN(n4114)
         );
  OAI21_X1 U5122 ( .B1(n4354), .B2(n4115), .A(n4114), .ZN(n4118) );
  XNOR2_X1 U5123 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n4116), .ZN(n5657)
         );
  NAND2_X1 U5124 ( .A1(n4931), .A2(n5657), .ZN(n4117) );
  NAND2_X1 U5125 ( .A1(n4118), .A2(n4117), .ZN(n5415) );
  AOI22_X1 U5126 ( .A1(n4367), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5127 ( .A1(n4311), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5128 ( .A1(n4360), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4361), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5129 ( .A1(n3446), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U5130 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4128)
         );
  AOI22_X1 U5131 ( .A1(n4368), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5132 ( .A1(n4187), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5133 ( .A1(n4522), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5134 ( .A1(n4372), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5135 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4127)
         );
  NOR2_X1 U5136 ( .A1(n4128), .A2(n4127), .ZN(n4132) );
  NAND2_X1 U5137 ( .A1(n6656), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4129)
         );
  NAND2_X1 U5138 ( .A1(n4357), .A2(n4129), .ZN(n4130) );
  AOI21_X1 U5139 ( .B1(n3912), .B2(EAX_REG_18__SCAN_IN), .A(n4130), .ZN(n4131)
         );
  OAI21_X1 U5140 ( .B1(n4354), .B2(n4132), .A(n4131), .ZN(n4136) );
  OAI21_X1 U5141 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4133), .A(n4151), 
        .ZN(n6059) );
  INV_X1 U5142 ( .A(n6059), .ZN(n4134) );
  NAND2_X1 U5143 ( .A1(n4134), .A2(n4931), .ZN(n4135) );
  AOI22_X1 U5144 ( .A1(n4522), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5145 ( .A1(n4311), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5146 ( .A1(n4368), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5147 ( .A1(n4361), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U5148 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4146)
         );
  AOI22_X1 U5149 ( .A1(n4367), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5150 ( .A1(n4369), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5151 ( .A1(n4359), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5152 ( .A1(n4360), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4141) );
  NAND4_X1 U5153 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4145)
         );
  NOR2_X1 U5154 ( .A1(n4146), .A2(n4145), .ZN(n4150) );
  NAND2_X1 U5155 ( .A1(n6656), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4147)
         );
  NAND2_X1 U5156 ( .A1(n4357), .A2(n4147), .ZN(n4148) );
  AOI21_X1 U5157 ( .B1(n3912), .B2(EAX_REG_19__SCAN_IN), .A(n4148), .ZN(n4149)
         );
  OAI21_X1 U5158 ( .B1(n4354), .B2(n4150), .A(n4149), .ZN(n4153) );
  XNOR2_X1 U5159 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4151), .ZN(n5642)
         );
  NAND2_X1 U5160 ( .A1(n4931), .A2(n5642), .ZN(n4152) );
  OR2_X1 U5161 ( .A1(n4154), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4155)
         );
  NAND2_X1 U5162 ( .A1(n4155), .A2(n4184), .ZN(n5955) );
  AOI22_X1 U5163 ( .A1(n4522), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5164 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4311), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5165 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4360), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5166 ( .A1(n4361), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4156) );
  NAND4_X1 U5167 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4165)
         );
  AOI22_X1 U5168 ( .A1(n4367), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5169 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3446), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5170 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4359), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5171 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4369), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4160) );
  NAND4_X1 U5172 ( .A1(n4163), .A2(n4162), .A3(n4161), .A4(n4160), .ZN(n4164)
         );
  NOR2_X1 U5173 ( .A1(n4165), .A2(n4164), .ZN(n4166) );
  NOR2_X1 U5174 ( .A1(n4354), .A2(n4166), .ZN(n4170) );
  INV_X1 U5175 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4168) );
  NAND2_X1 U5176 ( .A1(n6656), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4167)
         );
  OAI211_X1 U5177 ( .C1(n4326), .C2(n4168), .A(n4357), .B(n4167), .ZN(n4169)
         );
  OAI22_X1 U5178 ( .A1(n5955), .A2(n4357), .B1(n4170), .B2(n4169), .ZN(n5503)
         );
  AOI22_X1 U5179 ( .A1(n4311), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5180 ( .A1(n4360), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5181 ( .A1(n4361), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5182 ( .A1(n4372), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4171) );
  NAND4_X1 U5183 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4180)
         );
  AOI22_X1 U5184 ( .A1(n4367), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5185 ( .A1(n4368), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5186 ( .A1(n3446), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5187 ( .A1(n4522), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4175) );
  NAND4_X1 U5188 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(n4179)
         );
  NOR2_X1 U5189 ( .A1(n4180), .A2(n4179), .ZN(n4183) );
  INV_X1 U5190 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5945) );
  AOI21_X1 U5191 ( .B1(n5945), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4181) );
  AOI21_X1 U5192 ( .B1(n3912), .B2(EAX_REG_21__SCAN_IN), .A(n4181), .ZN(n4182)
         );
  OAI21_X1 U5193 ( .B1(n4354), .B2(n4183), .A(n4182), .ZN(n4186) );
  XNOR2_X1 U5194 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4184), .ZN(n5947)
         );
  NAND2_X1 U5195 ( .A1(n4931), .A2(n5947), .ZN(n4185) );
  NAND2_X1 U5196 ( .A1(n4186), .A2(n4185), .ZN(n5494) );
  NOR2_X2 U5197 ( .A1(n5493), .A2(n5494), .ZN(n5489) );
  AOI22_X1 U5198 ( .A1(n4367), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5199 ( .A1(n4522), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5200 ( .A1(n4187), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5201 ( .A1(n4372), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4188) );
  NAND4_X1 U5202 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4197)
         );
  AOI22_X1 U5203 ( .A1(n4311), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5204 ( .A1(n4360), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4361), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5205 ( .A1(n4368), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5206 ( .A1(n3446), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4192) );
  NAND4_X1 U5207 ( .A1(n4195), .A2(n4194), .A3(n4193), .A4(n4192), .ZN(n4196)
         );
  NOR2_X1 U5208 ( .A1(n4197), .A2(n4196), .ZN(n4201) );
  OAI21_X1 U5209 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6657), .A(n6656), 
        .ZN(n4198) );
  INV_X1 U5210 ( .A(n4198), .ZN(n4199) );
  AOI21_X1 U5211 ( .B1(n3912), .B2(EAX_REG_22__SCAN_IN), .A(n4199), .ZN(n4200)
         );
  OAI21_X1 U5212 ( .B1(n4354), .B2(n4201), .A(n4200), .ZN(n4205) );
  NOR2_X1 U5213 ( .A1(n4202), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4203)
         );
  NOR2_X1 U5214 ( .A1(n4229), .A2(n4203), .ZN(n5935) );
  NAND2_X1 U5215 ( .A1(n5935), .A2(n4931), .ZN(n4204) );
  AOI22_X1 U5216 ( .A1(n4368), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5217 ( .A1(n4367), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4360), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U5218 ( .A1(n3446), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5219 ( .A1(n4366), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4206) );
  NAND4_X1 U5220 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4215)
         );
  AOI22_X1 U5221 ( .A1(n4311), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U5222 ( .A1(n4522), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U5223 ( .A1(n4361), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5224 ( .A1(n3412), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4210) );
  NAND4_X1 U5225 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(n4214)
         );
  OR2_X1 U5226 ( .A1(n4215), .A2(n4214), .ZN(n4233) );
  AOI22_X1 U5227 ( .A1(n4370), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5228 ( .A1(n3412), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5229 ( .A1(n4369), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5230 ( .A1(n4361), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4216) );
  NAND4_X1 U5231 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4225)
         );
  AOI22_X1 U5232 ( .A1(n4366), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4367), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U5233 ( .A1(n4522), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5234 ( .A1(n4187), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4311), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5235 ( .A1(n4360), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4372), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4220) );
  NAND4_X1 U5236 ( .A1(n4223), .A2(n4222), .A3(n4221), .A4(n4220), .ZN(n4224)
         );
  OR2_X1 U5237 ( .A1(n4225), .A2(n4224), .ZN(n4232) );
  XNOR2_X1 U5238 ( .A(n4233), .B(n4232), .ZN(n4228) );
  INV_X1 U5239 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5615) );
  AOI21_X1 U5240 ( .B1(n5615), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4226) );
  AOI21_X1 U5241 ( .B1(n3912), .B2(EAX_REG_23__SCAN_IN), .A(n4226), .ZN(n4227)
         );
  OAI21_X1 U5242 ( .B1(n4354), .B2(n4228), .A(n4227), .ZN(n4231) );
  XNOR2_X1 U5243 ( .A(n4229), .B(n5615), .ZN(n5619) );
  NAND2_X1 U5244 ( .A1(n5619), .A2(n4931), .ZN(n4230) );
  NAND2_X1 U5245 ( .A1(n4231), .A2(n4230), .ZN(n5386) );
  AND2_X1 U5246 ( .A1(n4233), .A2(n4232), .ZN(n4282) );
  AOI22_X1 U5247 ( .A1(n4311), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5248 ( .A1(n4360), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5249 ( .A1(n4361), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5250 ( .A1(n4372), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4234) );
  NAND4_X1 U5251 ( .A1(n4237), .A2(n4236), .A3(n4235), .A4(n4234), .ZN(n4243)
         );
  AOI22_X1 U5252 ( .A1(n4367), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5253 ( .A1(n4368), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U5254 ( .A1(n3446), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5255 ( .A1(n4522), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4238) );
  NAND4_X1 U5256 ( .A1(n4241), .A2(n4240), .A3(n4239), .A4(n4238), .ZN(n4242)
         );
  OR2_X1 U5257 ( .A1(n4243), .A2(n4242), .ZN(n4281) );
  INV_X1 U5258 ( .A(n4281), .ZN(n4244) );
  XNOR2_X1 U5259 ( .A(n4282), .B(n4244), .ZN(n4248) );
  NAND2_X1 U5260 ( .A1(n4391), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4246)
         );
  INV_X1 U5261 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U5262 ( .A(n4264), .B(n5378), .ZN(n5605) );
  NAND2_X1 U5263 ( .A1(n5605), .A2(n4931), .ZN(n4245) );
  OAI211_X1 U5264 ( .C1(n4326), .C2(n6892), .A(n4246), .B(n4245), .ZN(n4247)
         );
  AOI21_X1 U5265 ( .B1(n4383), .B2(n4248), .A(n4247), .ZN(n5376) );
  AOI22_X1 U5266 ( .A1(n4311), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5267 ( .A1(n4360), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U5268 ( .A1(n4361), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U5269 ( .A1(n4372), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4250) );
  NAND4_X1 U5270 ( .A1(n4253), .A2(n4252), .A3(n4251), .A4(n4250), .ZN(n4259)
         );
  AOI22_X1 U5271 ( .A1(n4367), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U5272 ( .A1(n4368), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U5273 ( .A1(n3446), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U5274 ( .A1(n4522), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4254) );
  NAND4_X1 U5275 ( .A1(n4257), .A2(n4256), .A3(n4255), .A4(n4254), .ZN(n4258)
         );
  OR2_X1 U5276 ( .A1(n4259), .A2(n4258), .ZN(n4280) );
  AND2_X1 U5277 ( .A1(n4281), .A2(n4282), .ZN(n4260) );
  XNOR2_X1 U5278 ( .A(n4280), .B(n4260), .ZN(n4263) );
  INV_X1 U5279 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6913) );
  OAI21_X1 U5280 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6913), .A(n4357), .ZN(
        n4261) );
  AOI21_X1 U5281 ( .B1(n3912), .B2(EAX_REG_25__SCAN_IN), .A(n4261), .ZN(n4262)
         );
  OAI21_X1 U5282 ( .B1(n4354), .B2(n4263), .A(n4262), .ZN(n4269) );
  NOR2_X1 U5283 ( .A1(n4264), .A2(n5378), .ZN(n4265) );
  NOR2_X1 U5284 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4265), .ZN(n4266)
         );
  OR2_X1 U5285 ( .A1(n4286), .A2(n4266), .ZN(n5978) );
  INV_X1 U5286 ( .A(n5978), .ZN(n4267) );
  NAND2_X1 U5287 ( .A1(n4267), .A2(n4931), .ZN(n4268) );
  NAND2_X1 U5288 ( .A1(n4269), .A2(n4268), .ZN(n5479) );
  AOI22_X1 U5289 ( .A1(n4311), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5290 ( .A1(n4361), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5291 ( .A1(n3412), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5292 ( .A1(n4372), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4270) );
  NAND4_X1 U5293 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4279)
         );
  AOI22_X1 U5294 ( .A1(n4367), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5295 ( .A1(n4522), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5296 ( .A1(n4360), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5297 ( .A1(n4359), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5298 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4278)
         );
  NOR2_X1 U5299 ( .A1(n4279), .A2(n4278), .ZN(n4291) );
  NAND3_X1 U5300 ( .A1(n4282), .A2(n4281), .A3(n4280), .ZN(n4290) );
  XOR2_X1 U5301 ( .A(n4291), .B(n4290), .Z(n4283) );
  NAND2_X1 U5302 ( .A1(n4283), .A2(n4383), .ZN(n4289) );
  NAND2_X1 U5303 ( .A1(n6656), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4284)
         );
  NAND2_X1 U5304 ( .A1(n4357), .A2(n4284), .ZN(n4285) );
  AOI21_X1 U5305 ( .B1(n3912), .B2(EAX_REG_26__SCAN_IN), .A(n4285), .ZN(n4288)
         );
  INV_X1 U5306 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U5307 ( .A(n4286), .B(n5591), .ZN(n5595) );
  AOI21_X1 U5308 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(n5365) );
  NOR2_X1 U5309 ( .A1(n4291), .A2(n4290), .ZN(n4323) );
  AOI22_X1 U5310 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4311), .B1(n3292), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U5311 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4369), .B1(n4360), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U5312 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3447), .B1(n4361), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U5313 ( .A1(n4372), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4292) );
  NAND4_X1 U5314 ( .A1(n4295), .A2(n4294), .A3(n4293), .A4(n4292), .ZN(n4301)
         );
  AOI22_X1 U5315 ( .A1(n4367), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U5316 ( .A1(n4368), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U5317 ( .A1(n3446), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U5318 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4522), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4296) );
  NAND4_X1 U5319 ( .A1(n4299), .A2(n4298), .A3(n4297), .A4(n4296), .ZN(n4300)
         );
  OR2_X1 U5320 ( .A1(n4301), .A2(n4300), .ZN(n4322) );
  INV_X1 U5321 ( .A(n4322), .ZN(n4302) );
  XNOR2_X1 U5322 ( .A(n4323), .B(n4302), .ZN(n4303) );
  NAND2_X1 U5323 ( .A1(n4303), .A2(n4383), .ZN(n4310) );
  AOI21_X1 U5324 ( .B1(n4305), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4304) );
  AOI21_X1 U5325 ( .B1(n4386), .B2(EAX_REG_27__SCAN_IN), .A(n4304), .ZN(n4309)
         );
  NAND2_X1 U5326 ( .A1(n4306), .A2(n4305), .ZN(n4307) );
  NAND2_X1 U5327 ( .A1(n4331), .A2(n4307), .ZN(n5917) );
  NOR2_X1 U5328 ( .A1(n5917), .A2(n4357), .ZN(n4308) );
  AOI21_X1 U5329 ( .B1(n4310), .B2(n4309), .A(n4308), .ZN(n5466) );
  NAND2_X1 U5330 ( .A1(n5363), .A2(n5466), .ZN(n5452) );
  AOI22_X1 U5331 ( .A1(n4367), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4522), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4315) );
  AOI22_X1 U5332 ( .A1(n4368), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U5333 ( .A1(n4311), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U5334 ( .A1(n4372), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4312) );
  NAND4_X1 U5335 ( .A1(n4315), .A2(n4314), .A3(n4313), .A4(n4312), .ZN(n4321)
         );
  AOI22_X1 U5336 ( .A1(n4360), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U5337 ( .A1(n4361), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U5338 ( .A1(n3446), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U5339 ( .A1(n4366), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4316) );
  NAND4_X1 U5340 ( .A1(n4319), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(n4320)
         );
  NOR2_X1 U5341 ( .A1(n4321), .A2(n4320), .ZN(n4340) );
  NAND2_X1 U5342 ( .A1(n4323), .A2(n4322), .ZN(n4339) );
  XOR2_X1 U5343 ( .A(n4340), .B(n4339), .Z(n4328) );
  INV_X1 U5344 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4325) );
  NAND2_X1 U5345 ( .A1(n6656), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4324)
         );
  OAI211_X1 U5346 ( .C1(n4326), .C2(n4325), .A(n4357), .B(n4324), .ZN(n4327)
         );
  AOI21_X1 U5347 ( .B1(n4328), .B2(n4383), .A(n4327), .ZN(n4329) );
  INV_X1 U5348 ( .A(n4329), .ZN(n4335) );
  NAND2_X1 U5349 ( .A1(n4331), .A2(n4330), .ZN(n4332) );
  NAND2_X1 U5350 ( .A1(n4337), .A2(n4332), .ZN(n5907) );
  INV_X1 U5351 ( .A(n5907), .ZN(n4333) );
  NAND2_X1 U5352 ( .A1(n4333), .A2(n4931), .ZN(n4334) );
  NAND2_X1 U5353 ( .A1(n4335), .A2(n4334), .ZN(n5453) );
  NOR2_X2 U5354 ( .A1(n5452), .A2(n5453), .ZN(n5349) );
  INV_X1 U5355 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4336) );
  NAND2_X1 U5356 ( .A1(n4337), .A2(n4336), .ZN(n4338) );
  NAND2_X1 U5357 ( .A1(n4387), .A2(n4338), .ZN(n5568) );
  NOR2_X1 U5358 ( .A1(n4340), .A2(n4339), .ZN(n4380) );
  AOI22_X1 U5359 ( .A1(n4311), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U5360 ( .A1(n4360), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4369), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U5361 ( .A1(n4361), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U5362 ( .A1(n4372), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4341) );
  NAND4_X1 U5363 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), .ZN(n4351)
         );
  AOI22_X1 U5364 ( .A1(n4367), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U5365 ( .A1(n4368), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U5366 ( .A1(n3446), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U5367 ( .A1(n4522), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4346) );
  NAND4_X1 U5368 ( .A1(n4349), .A2(n4348), .A3(n4347), .A4(n4346), .ZN(n4350)
         );
  OR2_X1 U5369 ( .A1(n4351), .A2(n4350), .ZN(n4379) );
  XNOR2_X1 U5370 ( .A(n4380), .B(n4379), .ZN(n4355) );
  AOI21_X1 U5371 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6656), .A(n4931), 
        .ZN(n4353) );
  NAND2_X1 U5372 ( .A1(n3912), .A2(EAX_REG_29__SCAN_IN), .ZN(n4352) );
  OAI211_X1 U5373 ( .C1(n4355), .C2(n4354), .A(n4353), .B(n4352), .ZN(n4356)
         );
  OAI21_X1 U5374 ( .B1(n4357), .B2(n5568), .A(n4356), .ZN(n5351) );
  AOI22_X1 U5375 ( .A1(n4311), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U5376 ( .A1(n4360), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U5377 ( .A1(n4361), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U5378 ( .A1(n3446), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4362) );
  NAND4_X1 U5379 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4378)
         );
  AOI22_X1 U5380 ( .A1(n4367), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U5381 ( .A1(n4369), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4368), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U5382 ( .A1(n4522), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4370), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U5383 ( .A1(n4372), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4371), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4373) );
  NAND4_X1 U5384 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(n4377)
         );
  NOR2_X1 U5385 ( .A1(n4378), .A2(n4377), .ZN(n4382) );
  NAND2_X1 U5386 ( .A1(n4380), .A2(n4379), .ZN(n4381) );
  XOR2_X1 U5387 ( .A(n4382), .B(n4381), .Z(n4384) );
  NAND2_X1 U5388 ( .A1(n4384), .A2(n4383), .ZN(n4390) );
  INV_X1 U5389 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5294) );
  AOI21_X1 U5390 ( .B1(n5294), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4385) );
  AOI21_X1 U5391 ( .B1(n4386), .B2(EAX_REG_30__SCAN_IN), .A(n4385), .ZN(n4389)
         );
  XNOR2_X1 U5392 ( .A(n4387), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5311)
         );
  AND2_X1 U5393 ( .A1(n5311), .A2(n4931), .ZN(n4388) );
  NAND2_X1 U5394 ( .A1(n5350), .A2(n5292), .ZN(n4393) );
  INV_X1 U5395 ( .A(n5326), .ZN(n4395) );
  NAND3_X1 U5396 ( .A1(n6660), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6556) );
  INV_X1 U5397 ( .A(n6556), .ZN(n4394) );
  NAND2_X1 U5398 ( .A1(n4395), .A2(n6260), .ZN(n4396) );
  OAI211_X1 U5399 ( .C1(n5713), .C2(n6277), .A(n4397), .B(n4396), .ZN(U2955)
         );
  INV_X1 U5400 ( .A(n6515), .ZN(n4398) );
  INV_X1 U5401 ( .A(n6544), .ZN(n6036) );
  AND2_X1 U5402 ( .A1(n5024), .A2(n6552), .ZN(n5157) );
  INV_X1 U5403 ( .A(n4399), .ZN(n6517) );
  NOR2_X2 U5404 ( .A1(n4431), .A2(n6517), .ZN(n4403) );
  AOI211_X1 U5405 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4401), .A(n5157), .B(
        n4403), .ZN(n4400) );
  INV_X1 U5406 ( .A(n4400), .ZN(U2788) );
  NAND2_X1 U5407 ( .A1(n6034), .A2(n5336), .ZN(n6043) );
  INV_X1 U5408 ( .A(n6043), .ZN(n4405) );
  OAI21_X1 U5409 ( .B1(n5157), .B2(READREQUEST_REG_SCAN_IN), .A(n6662), .ZN(
        n4404) );
  OAI21_X1 U5410 ( .B1(n6662), .B2(n4405), .A(n4404), .ZN(U3474) );
  OAI21_X1 U5411 ( .B1(n4408), .B2(n4407), .A(n4406), .ZN(n5196) );
  NAND2_X1 U5412 ( .A1(n6522), .A2(n6544), .ZN(n4409) );
  INV_X1 U5413 ( .A(n4410), .ZN(n4414) );
  INV_X1 U5414 ( .A(n3337), .ZN(n5327) );
  AND4_X1 U5415 ( .A1(n3342), .A2(n4637), .A3(n5327), .A4(n4411), .ZN(n4412)
         );
  NAND3_X1 U5416 ( .A1(n4414), .A2(n4413), .A3(n4412), .ZN(n4585) );
  INV_X1 U5417 ( .A(n4585), .ZN(n4415) );
  NAND2_X1 U5418 ( .A1(n4415), .A2(n4940), .ZN(n4416) );
  NAND2_X1 U5419 ( .A1(n6156), .A2(n3337), .ZN(n5535) );
  XNOR2_X1 U5420 ( .A(n4418), .B(n5336), .ZN(n4708) );
  AOI22_X1 U5421 ( .A1(n6670), .A2(n4708), .B1(n6671), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4419) );
  OAI21_X1 U5422 ( .B1(n5196), .B2(n5535), .A(n4419), .ZN(U2858) );
  OAI21_X1 U5423 ( .B1(n6658), .B2(n4438), .A(n4403), .ZN(n6246) );
  INV_X1 U5424 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6721) );
  NAND3_X1 U5425 ( .A1(n3112), .A2(n4940), .A3(n4438), .ZN(n4420) );
  INV_X1 U5426 ( .A(DATAI_11_), .ZN(n4421) );
  NOR2_X1 U5427 ( .A1(n6251), .A2(n4421), .ZN(n6240) );
  AOI21_X1 U5428 ( .B1(n6249), .B2(EAX_REG_27__SCAN_IN), .A(n6240), .ZN(n4422)
         );
  OAI21_X1 U5429 ( .B1(n6202), .B2(n6721), .A(n4422), .ZN(U2935) );
  INV_X1 U5430 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6694) );
  INV_X1 U5431 ( .A(DATAI_9_), .ZN(n4423) );
  NOR2_X1 U5432 ( .A1(n6251), .A2(n4423), .ZN(n6234) );
  AOI21_X1 U5433 ( .B1(n6249), .B2(EAX_REG_25__SCAN_IN), .A(n6234), .ZN(n4424)
         );
  OAI21_X1 U5434 ( .B1(n6202), .B2(n6694), .A(n4424), .ZN(U2933) );
  NAND2_X1 U5435 ( .A1(n4426), .A2(n4425), .ZN(n4427) );
  NAND2_X1 U5436 ( .A1(n4428), .A2(n4427), .ZN(n6284) );
  NOR2_X1 U5437 ( .A1(n5337), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4429)
         );
  OR2_X1 U5438 ( .A1(n4430), .A2(n4429), .ZN(n4937) );
  OAI222_X1 U5439 ( .A1(n6284), .A2(n5535), .B1(n6156), .B2(n6821), .C1(n4937), 
        .C2(n5532), .ZN(U2859) );
  OR2_X1 U5440 ( .A1(n4431), .A2(n6503), .ZN(n4432) );
  NAND2_X1 U5441 ( .A1(n6254), .A2(n4432), .ZN(n4433) );
  INV_X1 U5442 ( .A(n6563), .ZN(n6042) );
  NOR2_X1 U5443 ( .A1(n6552), .A2(n6656), .ZN(n6549) );
  NAND2_X1 U5444 ( .A1(n6549), .A2(n6660), .ZN(n6664) );
  INV_X1 U5445 ( .A(n6664), .ZN(n6184) );
  INV_X1 U5446 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U5447 ( .A1(n6188), .A2(n3111), .ZN(n6170) );
  INV_X1 U5448 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6709) );
  INV_X1 U5449 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4434) );
  OAI222_X1 U5450 ( .A1(n6200), .A2(n6897), .B1(n6170), .B2(n6709), .C1(n4434), 
        .C2(n6664), .ZN(U2900) );
  INV_X1 U5451 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6745) );
  INV_X1 U5452 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6795) );
  INV_X1 U5453 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n4435) );
  OAI222_X1 U5454 ( .A1(n6200), .A2(n6745), .B1(n6170), .B2(n6795), .C1(n4435), 
        .C2(n6664), .ZN(U2893) );
  INV_X1 U5455 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6365) );
  NOR2_X1 U5456 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6365), .ZN(n6626) );
  INV_X1 U5457 ( .A(n6522), .ZN(n4444) );
  OAI21_X1 U5458 ( .B1(n6042), .B2(n4940), .A(n3112), .ZN(n4436) );
  OAI21_X1 U5459 ( .B1(n6503), .B2(n6563), .A(n4436), .ZN(n4437) );
  NAND3_X1 U5460 ( .A1(n6521), .A2(n4438), .A3(n4437), .ZN(n4443) );
  INV_X1 U5461 ( .A(n4439), .ZN(n4440) );
  AND2_X1 U5462 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  OAI211_X1 U5463 ( .C1(n6521), .C2(n4444), .A(n4443), .B(n4442), .ZN(n4445)
         );
  INV_X1 U5464 ( .A(n4445), .ZN(n4450) );
  NAND2_X1 U5465 ( .A1(n6521), .A2(n4460), .ZN(n4448) );
  OR2_X1 U5466 ( .A1(n3737), .A2(n4446), .ZN(n4447) );
  NAND2_X1 U5467 ( .A1(n4448), .A2(n4447), .ZN(n4583) );
  INV_X1 U5468 ( .A(n4583), .ZN(n4449) );
  NAND2_X1 U5469 ( .A1(n4450), .A2(n4449), .ZN(n4535) );
  INV_X1 U5470 ( .A(n4535), .ZN(n6508) );
  INV_X1 U5471 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6524) );
  NAND2_X1 U5472 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6549), .ZN(n6553) );
  OAI22_X1 U5473 ( .A1(n6508), .A2(n6036), .B1(n6524), .B2(n6553), .ZN(n6027)
         );
  NOR2_X1 U5474 ( .A1(n6626), .A2(n6027), .ZN(n6025) );
  AND2_X1 U5475 ( .A1(n4453), .A2(n4452), .ZN(n4456) );
  INV_X1 U5476 ( .A(n3112), .ZN(n4455) );
  NAND4_X1 U5477 ( .A1(n3737), .A2(n4456), .A3(n4455), .A4(n4454), .ZN(n4457)
         );
  OR2_X1 U5478 ( .A1(n4458), .A2(n4457), .ZN(n5842) );
  INV_X1 U5479 ( .A(n5842), .ZN(n5286) );
  XNOR2_X1 U5480 ( .A(n4459), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4464)
         );
  OR2_X1 U5481 ( .A1(n4460), .A2(n6522), .ZN(n4530) );
  NAND2_X1 U5482 ( .A1(n4530), .A2(n4464), .ZN(n4463) );
  XNOR2_X1 U5483 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4461) );
  OR2_X1 U5484 ( .A1(n6503), .A2(n4461), .ZN(n4462) );
  OAI211_X1 U5485 ( .C1(n4533), .C2(n4464), .A(n4463), .B(n4462), .ZN(n4465)
         );
  INV_X1 U5486 ( .A(n4465), .ZN(n4466) );
  OAI21_X1 U5487 ( .B1(n4451), .B2(n5286), .A(n4466), .ZN(n4518) );
  INV_X1 U5488 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6714) );
  AOI22_X1 U5489 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n6714), .B2(n3741), .ZN(n5844)
         );
  NOR2_X1 U5490 ( .A1(n6552), .A2(n6320), .ZN(n5845) );
  AND2_X1 U5491 ( .A1(n5844), .A2(n5845), .ZN(n4468) );
  INV_X1 U5492 ( .A(n4459), .ZN(n5838) );
  NOR3_X1 U5493 ( .A1(n5838), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6539), 
        .ZN(n4467) );
  AOI211_X1 U5494 ( .C1(n4518), .C2(n6545), .A(n4468), .B(n4467), .ZN(n4470)
         );
  NOR2_X1 U5495 ( .A1(n4459), .A2(n6539), .ZN(n5848) );
  OAI21_X1 U5496 ( .B1(n6025), .B2(n5848), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4469) );
  OAI21_X1 U5497 ( .B1(n6025), .B2(n4470), .A(n4469), .ZN(U3459) );
  NAND2_X1 U5498 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4577) );
  AOI21_X1 U5499 ( .B1(n5167), .B2(n4577), .A(n5168), .ZN(n4700) );
  NOR2_X1 U5500 ( .A1(n4700), .A2(n3498), .ZN(n4484) );
  NOR3_X1 U5501 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4699), .A3(n3741), 
        .ZN(n4483) );
  NAND2_X1 U5502 ( .A1(n4472), .A2(n4471), .ZN(n4473) );
  XNOR2_X1 U5503 ( .A(n4474), .B(n4473), .ZN(n6268) );
  NAND2_X1 U5504 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  AND2_X1 U5505 ( .A1(n4491), .A2(n4477), .ZN(n5275) );
  AOI22_X1 U5506 ( .A1(n6312), .A2(n5275), .B1(n6276), .B2(REIP_REG_2__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U5507 ( .B1(n4478), .B2(n3498), .A(n4576), .ZN(n4479) );
  NAND2_X1 U5508 ( .A1(n5831), .A2(n4479), .ZN(n4480) );
  OAI211_X1 U5509 ( .C1(n6268), .C2(n5984), .A(n4481), .B(n4480), .ZN(n4482)
         );
  OR3_X1 U5510 ( .A1(n4484), .A2(n4483), .A3(n4482), .ZN(U3016) );
  INV_X1 U5511 ( .A(n4485), .ZN(n4489) );
  INV_X1 U5512 ( .A(n4486), .ZN(n4488) );
  AOI21_X1 U5513 ( .B1(n4489), .B2(n4488), .A(n4487), .ZN(n4752) );
  INV_X1 U5514 ( .A(n4752), .ZN(n5208) );
  AOI21_X1 U5515 ( .B1(n4492), .B2(n4491), .A(n4490), .ZN(n5197) );
  AOI22_X1 U5516 ( .A1(n6670), .A2(n5197), .B1(n6671), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4493) );
  OAI21_X1 U5517 ( .B1(n5208), .B2(n5528), .A(n4493), .ZN(U2856) );
  INV_X1 U5518 ( .A(n5275), .ZN(n4497) );
  INV_X1 U5519 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6952) );
  NOR2_X1 U5520 ( .A1(n4495), .A2(n4494), .ZN(n4496) );
  OR2_X1 U5521 ( .A1(n4485), .A2(n4496), .ZN(n6267) );
  OAI222_X1 U5522 ( .A1(n4497), .A2(n5532), .B1(n6156), .B2(n6952), .C1(n5528), 
        .C2(n6267), .ZN(U2857) );
  INV_X1 U5523 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5524 ( .A1(n6192), .A2(UWORD_REG_6__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4498) );
  OAI21_X1 U5525 ( .B1(n4499), .B2(n6170), .A(n4498), .ZN(U2901) );
  INV_X1 U5526 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6213) );
  AOI22_X1 U5527 ( .A1(n6192), .A2(UWORD_REG_10__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4500) );
  OAI21_X1 U5528 ( .B1(n6213), .B2(n6170), .A(n4500), .ZN(U2897) );
  AOI22_X1 U5529 ( .A1(n6192), .A2(UWORD_REG_0__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4501) );
  OAI21_X1 U5530 ( .B1(n4100), .B2(n6170), .A(n4501), .ZN(U2907) );
  INV_X1 U5531 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6217) );
  AOI22_X1 U5532 ( .A1(n6192), .A2(UWORD_REG_13__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5533 ( .B1(n6217), .B2(n6170), .A(n4502), .ZN(U2894) );
  INV_X1 U5534 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5535 ( .A1(n6192), .A2(UWORD_REG_2__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4503) );
  OAI21_X1 U5536 ( .B1(n4504), .B2(n6170), .A(n4503), .ZN(U2905) );
  AOI22_X1 U5537 ( .A1(n6192), .A2(UWORD_REG_12__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4505) );
  OAI21_X1 U5538 ( .B1(n4325), .B2(n6170), .A(n4505), .ZN(U2895) );
  INV_X1 U5539 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U5540 ( .A1(n6192), .A2(UWORD_REG_5__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4506) );
  OAI21_X1 U5541 ( .B1(n6696), .B2(n6170), .A(n4506), .ZN(U2902) );
  INV_X1 U5542 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6892) );
  AOI22_X1 U5543 ( .A1(n6192), .A2(UWORD_REG_8__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4507) );
  OAI21_X1 U5544 ( .B1(n6892), .B2(n6170), .A(n4507), .ZN(U2899) );
  INV_X1 U5545 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U5546 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6192), .B1(n6191), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4508) );
  OAI21_X1 U5547 ( .B1(n6706), .B2(n6170), .A(n4508), .ZN(U2896) );
  INV_X1 U5548 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6712) );
  AOI22_X1 U5549 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6192), .B1(n6191), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4509) );
  OAI21_X1 U5550 ( .B1(n6712), .B2(n6170), .A(n4509), .ZN(U2898) );
  INV_X1 U5551 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U5552 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6192), .B1(n6191), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4510) );
  OAI21_X1 U5553 ( .B1(n6763), .B2(n6170), .A(n4510), .ZN(U2906) );
  OAI21_X1 U5554 ( .B1(n4512), .B2(n4514), .A(n4513), .ZN(n4755) );
  INV_X1 U5555 ( .A(n4771), .ZN(n4515) );
  AOI21_X1 U5556 ( .B1(n4516), .B2(n4570), .A(n4515), .ZN(n6120) );
  AOI22_X1 U5557 ( .A1(n6670), .A2(n6120), .B1(n6671), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4517) );
  OAI21_X1 U5558 ( .B1(n4755), .B2(n5535), .A(n4517), .ZN(U2854) );
  OR2_X1 U5559 ( .A1(n4535), .A2(n3164), .ZN(n4520) );
  NAND2_X1 U5560 ( .A1(n4535), .A2(n4518), .ZN(n4519) );
  INV_X1 U5561 ( .A(n6511), .ZN(n4538) );
  OR2_X1 U5562 ( .A1(n4535), .A2(n5854), .ZN(n4537) );
  OAI21_X1 U5563 ( .B1(n4522), .B2(n5854), .A(n4521), .ZN(n5851) );
  MUX2_X1 U5564 ( .A(n4524), .B(n5854), .S(n4525), .Z(n4526) );
  OAI21_X1 U5565 ( .B1(n4523), .B2(n4526), .A(n5285), .ZN(n4532) );
  INV_X1 U5566 ( .A(n4523), .ZN(n4528) );
  INV_X1 U5567 ( .A(n4524), .ZN(n4527) );
  OAI211_X1 U5568 ( .C1(n4459), .C2(n4528), .A(n3389), .B(n4527), .ZN(n4529)
         );
  NAND2_X1 U5569 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  OAI211_X1 U5570 ( .C1(n4533), .C2(n5851), .A(n4532), .B(n4531), .ZN(n4534)
         );
  AOI21_X1 U5571 ( .B1(n5858), .B2(n5842), .A(n4534), .ZN(n5853) );
  NAND2_X1 U5572 ( .A1(n4535), .A2(n5853), .ZN(n4536) );
  NAND3_X1 U5573 ( .A1(n4538), .A2(n6513), .A3(n6552), .ZN(n4542) );
  AND2_X1 U5574 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6524), .ZN(n4539) );
  NAND2_X1 U5575 ( .A1(n4540), .A2(n4539), .ZN(n4541) );
  NAND2_X1 U5576 ( .A1(n4542), .A2(n4541), .ZN(n6528) );
  INV_X1 U5577 ( .A(n4543), .ZN(n5847) );
  NAND2_X1 U5578 ( .A1(n6528), .A2(n5847), .ZN(n4549) );
  MUX2_X1 U5579 ( .A(n6524), .B(n6508), .S(n6552), .Z(n4548) );
  INV_X1 U5580 ( .A(n6359), .ZN(n4544) );
  NOR2_X1 U5581 ( .A1(n4545), .A2(n4544), .ZN(n4546) );
  XNOR2_X1 U5582 ( .A(n4546), .B(n6029), .ZN(n6138) );
  NOR2_X1 U5583 ( .A1(n3737), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4547) );
  AND2_X1 U5584 ( .A1(n6138), .A2(n4547), .ZN(n6026) );
  AOI21_X1 U5585 ( .B1(n4548), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n6026), 
        .ZN(n6530) );
  NAND2_X1 U5586 ( .A1(n6532), .A2(n6524), .ZN(n4550) );
  INV_X1 U5587 ( .A(n6553), .ZN(n6625) );
  NAND2_X1 U5588 ( .A1(n4550), .A2(n6625), .ZN(n4551) );
  NAND2_X1 U5589 ( .A1(n6552), .A2(n6656), .ZN(n6659) );
  INV_X1 U5590 ( .A(n6659), .ZN(n4930) );
  NAND2_X1 U5591 ( .A1(n4551), .A2(n5013), .ZN(n6639) );
  AOI21_X1 U5592 ( .B1(n4885), .B2(n6657), .A(n6630), .ZN(n4555) );
  NAND2_X1 U5593 ( .A1(n4553), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6407) );
  NAND2_X1 U5594 ( .A1(n6365), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6633) );
  AOI22_X1 U5595 ( .A1(n4555), .A2(n6407), .B1(n5843), .B2(n6633), .ZN(n4557)
         );
  NAND2_X1 U5596 ( .A1(n6642), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4556) );
  OAI21_X1 U5597 ( .B1(n6642), .B2(n4557), .A(n4556), .ZN(U3464) );
  XNOR2_X1 U5598 ( .A(n4559), .B(n6407), .ZN(n4560) );
  INV_X1 U5599 ( .A(n4451), .ZN(n5276) );
  AOI22_X1 U5600 ( .A1(n4560), .A2(n6411), .B1(n5276), .B2(n6633), .ZN(n4562)
         );
  NAND2_X1 U5601 ( .A1(n6642), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4561) );
  OAI21_X1 U5602 ( .B1(n6642), .B2(n4562), .A(n4561), .ZN(U3463) );
  AOI222_X1 U5603 ( .A1(n4563), .A2(n6411), .B1(n6532), .B2(n6549), .C1(n6436), 
        .C2(n6633), .ZN(n4565) );
  NAND2_X1 U5604 ( .A1(n6642), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U5605 ( .B1(n4565), .B2(n6642), .A(n4564), .ZN(U3465) );
  NOR2_X1 U5606 ( .A1(n4487), .A2(n4566), .ZN(n4567) );
  NOR2_X1 U5607 ( .A1(n4512), .A2(n4567), .ZN(n6261) );
  INV_X1 U5608 ( .A(n6261), .ZN(n4591) );
  OR2_X1 U5609 ( .A1(n4490), .A2(n4568), .ZN(n4569) );
  NAND2_X1 U5610 ( .A1(n4570), .A2(n4569), .ZN(n6131) );
  INV_X1 U5611 ( .A(n6131), .ZN(n4571) );
  AOI22_X1 U5612 ( .A1(n6670), .A2(n4571), .B1(n6671), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4572) );
  OAI21_X1 U5613 ( .B1(n4591), .B2(n5528), .A(n4572), .ZN(U2855) );
  XNOR2_X1 U5614 ( .A(n4573), .B(n4575), .ZN(n4754) );
  OAI21_X1 U5615 ( .B1(n4697), .B2(n4576), .A(n4700), .ZN(n4598) );
  INV_X1 U5616 ( .A(n4576), .ZN(n4579) );
  OAI21_X1 U5617 ( .B1(n4577), .B2(n4699), .A(n4697), .ZN(n4578) );
  INV_X1 U5618 ( .A(n4578), .ZN(n5171) );
  NOR2_X1 U5619 ( .A1(n4579), .A2(n5171), .ZN(n4595) );
  AOI22_X1 U5620 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4598), .B1(n4595), 
        .B2(n4580), .ZN(n4582) );
  INV_X1 U5621 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6681) );
  NOR2_X1 U5622 ( .A1(n5829), .A2(n6681), .ZN(n4749) );
  AOI21_X1 U5623 ( .B1(n6312), .B2(n5197), .A(n4749), .ZN(n4581) );
  OAI211_X1 U5624 ( .C1(n4754), .C2(n5984), .A(n4582), .B(n4581), .ZN(U3015)
         );
  NAND2_X1 U5625 ( .A1(n4583), .A2(n6544), .ZN(n4584) );
  AND2_X1 U5626 ( .A1(n3318), .A2(n3337), .ZN(n4587) );
  NOR2_X1 U5627 ( .A1(n4587), .A2(n3345), .ZN(n4586) );
  NAND2_X2 U5628 ( .A1(n6168), .A2(n4586), .ZN(n6169) );
  INV_X1 U5629 ( .A(n6160), .ZN(n4589) );
  INV_X1 U5630 ( .A(n6164), .ZN(n4588) );
  INV_X1 U5631 ( .A(DATAI_4_), .ZN(n6839) );
  INV_X1 U5632 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4590) );
  OAI222_X1 U5633 ( .A1(n4591), .A2(n6169), .B1(n6167), .B2(n6839), .C1(n6168), 
        .C2(n4590), .ZN(U2887) );
  INV_X1 U5634 ( .A(DATAI_3_), .ZN(n6225) );
  INV_X1 U5635 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6194) );
  OAI222_X1 U5636 ( .A1(n5208), .A2(n6169), .B1(n6167), .B2(n6225), .C1(n6168), 
        .C2(n6194), .ZN(U2888) );
  INV_X1 U5637 ( .A(DATAI_2_), .ZN(n6878) );
  INV_X1 U5638 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6967) );
  OAI222_X1 U5639 ( .A1(n6267), .A2(n6169), .B1(n6167), .B2(n6878), .C1(n6168), 
        .C2(n6967), .ZN(U2889) );
  INV_X1 U5640 ( .A(DATAI_1_), .ZN(n6222) );
  INV_X1 U5641 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6825) );
  OAI222_X1 U5642 ( .A1(n5196), .A2(n6169), .B1(n6167), .B2(n6222), .C1(n6168), 
        .C2(n6825), .ZN(U2890) );
  XNOR2_X1 U5643 ( .A(n4592), .B(n4593), .ZN(n6256) );
  NAND2_X1 U5644 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4594) );
  OAI211_X1 U5645 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4595), .B(n4594), .ZN(n4600) );
  NAND2_X1 U5646 ( .A1(n6276), .A2(REIP_REG_4__SCAN_IN), .ZN(n6264) );
  INV_X1 U5647 ( .A(n6264), .ZN(n4597) );
  NOR2_X1 U5648 ( .A1(n6018), .A2(n6131), .ZN(n4596) );
  AOI211_X1 U5649 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4598), .A(n4597), 
        .B(n4596), .ZN(n4599) );
  OAI211_X1 U5650 ( .C1(n5984), .C2(n6256), .A(n4600), .B(n4599), .ZN(U3014)
         );
  INV_X1 U5651 ( .A(DATAI_5_), .ZN(n6228) );
  INV_X1 U5652 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6852) );
  OAI222_X1 U5653 ( .A1(n4755), .A2(n6169), .B1(n6167), .B2(n6228), .C1(n6168), 
        .C2(n6852), .ZN(U2886) );
  NAND2_X1 U5654 ( .A1(n6408), .A2(n4885), .ZN(n6326) );
  INV_X1 U5655 ( .A(DATAI_20_), .ZN(n4601) );
  OR2_X1 U5656 ( .A1(n6283), .A2(n4601), .ZN(n5885) );
  NAND3_X1 U5657 ( .A1(n4602), .A2(n4658), .A3(n4553), .ZN(n4779) );
  NAND2_X1 U5658 ( .A1(n6411), .A2(n6657), .ZN(n6636) );
  INV_X1 U5659 ( .A(n6636), .ZN(n4954) );
  OR2_X1 U5660 ( .A1(n4451), .A2(n5843), .ZN(n4609) );
  OAI22_X1 U5661 ( .A1(n4806), .A2(n4954), .B1(n6359), .B2(n4609), .ZN(n4605)
         );
  OAI21_X1 U5662 ( .B1(n6326), .B2(n6657), .A(n6411), .ZN(n6329) );
  NAND3_X1 U5663 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6641), .A3(n6969), .ZN(n6327) );
  NOR2_X1 U5664 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6327), .ZN(n4608)
         );
  OR2_X1 U5665 ( .A1(n5007), .A2(n5006), .ZN(n4611) );
  AOI21_X1 U5666 ( .B1(n4611), .B2(STATE2_REG_2__SCAN_IN), .A(n5013), .ZN(
        n4659) );
  OAI21_X1 U5667 ( .B1(n6365), .B2(n4608), .A(n4659), .ZN(n4603) );
  INV_X1 U5668 ( .A(n4603), .ZN(n4604) );
  OR2_X1 U5669 ( .A1(n4610), .A2(n6656), .ZN(n6363) );
  OAI211_X1 U5670 ( .C1(n4605), .C2(n6329), .A(n4604), .B(n6363), .ZN(n4646)
         );
  NAND2_X1 U5671 ( .A1(n4646), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4614) );
  INV_X1 U5672 ( .A(DATAI_28_), .ZN(n4606) );
  OR2_X1 U5673 ( .A1(n6283), .A2(n4606), .ZN(n5143) );
  INV_X1 U5674 ( .A(n5143), .ZN(n6475) );
  NOR2_X1 U5675 ( .A1(n4648), .A2(n3237), .ZN(n6473) );
  INV_X1 U5676 ( .A(n6473), .ZN(n4961) );
  INV_X1 U5677 ( .A(n4608), .ZN(n4650) );
  NOR2_X1 U5678 ( .A1(n5858), .A2(n6630), .ZN(n4819) );
  NAND2_X1 U5679 ( .A1(n4610), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6368) );
  INV_X1 U5680 ( .A(n6368), .ZN(n5010) );
  INV_X1 U5681 ( .A(n4611), .ZN(n4665) );
  AOI22_X1 U5682 ( .A1(n4819), .A2(n6322), .B1(n5010), .B2(n4665), .ZN(n4649)
         );
  NOR2_X1 U5683 ( .A1(n6839), .A2(n5013), .ZN(n6385) );
  OAI22_X1 U5684 ( .A1(n4961), .A2(n4650), .B1(n4649), .B2(n6478), .ZN(n4612)
         );
  AOI21_X1 U5685 ( .B1(n6475), .B2(n4652), .A(n4612), .ZN(n4613) );
  OAI211_X1 U5686 ( .C1(n4655), .C2(n5885), .A(n4614), .B(n4613), .ZN(U3056)
         );
  INV_X1 U5687 ( .A(DATAI_17_), .ZN(n4615) );
  OR2_X1 U5688 ( .A1(n6283), .A2(n4615), .ZN(n5873) );
  NAND2_X1 U5689 ( .A1(n4646), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4619) );
  INV_X1 U5690 ( .A(DATAI_25_), .ZN(n6808) );
  OR2_X1 U5691 ( .A1(n6283), .A2(n6808), .ZN(n5150) );
  INV_X1 U5692 ( .A(n5150), .ZN(n6457) );
  NOR2_X1 U5693 ( .A1(n4648), .A2(n4616), .ZN(n6455) );
  INV_X1 U5694 ( .A(n6455), .ZN(n4969) );
  NOR2_X1 U5695 ( .A1(n6222), .A2(n5013), .ZN(n6374) );
  OAI22_X1 U5696 ( .A1(n4969), .A2(n4650), .B1(n4649), .B2(n6460), .ZN(n4617)
         );
  AOI21_X1 U5697 ( .B1(n6457), .B2(n4652), .A(n4617), .ZN(n4618) );
  OAI211_X1 U5698 ( .C1(n4655), .C2(n5873), .A(n4619), .B(n4618), .ZN(U3053)
         );
  INV_X1 U5699 ( .A(DATAI_22_), .ZN(n4620) );
  OR2_X1 U5700 ( .A1(n6283), .A2(n4620), .ZN(n5893) );
  NAND2_X1 U5701 ( .A1(n4646), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4625) );
  INV_X1 U5702 ( .A(DATAI_30_), .ZN(n4621) );
  OR2_X1 U5703 ( .A1(n6283), .A2(n4621), .ZN(n5135) );
  INV_X1 U5704 ( .A(n5135), .ZN(n6486) );
  NOR2_X1 U5705 ( .A1(n4648), .A2(n4622), .ZN(n6485) );
  INV_X1 U5706 ( .A(n6485), .ZN(n4987) );
  INV_X1 U5707 ( .A(DATAI_6_), .ZN(n6230) );
  NOR2_X1 U5708 ( .A1(n6230), .A2(n5013), .ZN(n6392) );
  OAI22_X1 U5709 ( .A1(n4987), .A2(n4650), .B1(n4649), .B2(n6490), .ZN(n4623)
         );
  AOI21_X1 U5710 ( .B1(n6486), .B2(n4652), .A(n4623), .ZN(n4624) );
  OAI211_X1 U5711 ( .C1(n4655), .C2(n5893), .A(n4625), .B(n4624), .ZN(U3058)
         );
  INV_X1 U5712 ( .A(DATAI_23_), .ZN(n4626) );
  OR2_X1 U5713 ( .A1(n6283), .A2(n4626), .ZN(n5899) );
  NAND2_X1 U5714 ( .A1(n4646), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4630) );
  INV_X1 U5715 ( .A(DATAI_31_), .ZN(n4627) );
  OR2_X1 U5716 ( .A1(n6283), .A2(n4627), .ZN(n5131) );
  INV_X1 U5717 ( .A(n5131), .ZN(n6496) );
  INV_X1 U5718 ( .A(n6492), .ZN(n4983) );
  INV_X1 U5719 ( .A(DATAI_7_), .ZN(n6232) );
  NOR2_X1 U5720 ( .A1(n6232), .A2(n5013), .ZN(n6397) );
  OAI22_X1 U5721 ( .A1(n4983), .A2(n4650), .B1(n4649), .B2(n6500), .ZN(n4628)
         );
  AOI21_X1 U5722 ( .B1(n6496), .B2(n4652), .A(n4628), .ZN(n4629) );
  OAI211_X1 U5723 ( .C1(n4655), .C2(n5899), .A(n4630), .B(n4629), .ZN(U3059)
         );
  INV_X1 U5724 ( .A(DATAI_0_), .ZN(n6220) );
  NAND2_X1 U5725 ( .A1(n4646), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4635) );
  INV_X1 U5726 ( .A(DATAI_16_), .ZN(n4631) );
  OR2_X1 U5727 ( .A1(n6283), .A2(n4631), .ZN(n5869) );
  INV_X1 U5728 ( .A(n5869), .ZN(n6451) );
  NOR2_X1 U5729 ( .A1(n4648), .A2(n4632), .ZN(n6443) );
  INV_X1 U5730 ( .A(n6443), .ZN(n4974) );
  INV_X1 U5731 ( .A(DATAI_24_), .ZN(n6730) );
  OR2_X1 U5732 ( .A1(n6283), .A2(n6730), .ZN(n5117) );
  OAI22_X1 U5733 ( .A1(n4974), .A2(n4650), .B1(n4806), .B2(n5117), .ZN(n4633)
         );
  AOI21_X1 U5734 ( .B1(n6451), .B2(n6349), .A(n4633), .ZN(n4634) );
  OAI211_X1 U5735 ( .C1(n4649), .C2(n6454), .A(n4635), .B(n4634), .ZN(U3052)
         );
  INV_X1 U5736 ( .A(DATAI_19_), .ZN(n4636) );
  OR2_X1 U5737 ( .A1(n6283), .A2(n4636), .ZN(n5881) );
  NAND2_X1 U5738 ( .A1(n4646), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4640) );
  INV_X1 U5739 ( .A(DATAI_27_), .ZN(n6690) );
  OR2_X1 U5740 ( .A1(n6283), .A2(n6690), .ZN(n5127) );
  INV_X1 U5741 ( .A(n5127), .ZN(n6469) );
  NOR2_X1 U5742 ( .A1(n4648), .A2(n4637), .ZN(n6467) );
  INV_X1 U5743 ( .A(n6467), .ZN(n4979) );
  NOR2_X1 U5744 ( .A1(n6225), .A2(n5013), .ZN(n6381) );
  OAI22_X1 U5745 ( .A1(n4979), .A2(n4650), .B1(n4649), .B2(n6472), .ZN(n4638)
         );
  AOI21_X1 U5746 ( .B1(n6469), .B2(n4652), .A(n4638), .ZN(n4639) );
  OAI211_X1 U5747 ( .C1(n4655), .C2(n5881), .A(n4640), .B(n4639), .ZN(U3055)
         );
  INV_X1 U5748 ( .A(DATAI_21_), .ZN(n4641) );
  OR2_X1 U5749 ( .A1(n6283), .A2(n4641), .ZN(n5889) );
  NAND2_X1 U5750 ( .A1(n4646), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4644) );
  INV_X1 U5751 ( .A(DATAI_29_), .ZN(n6691) );
  OR2_X1 U5752 ( .A1(n6283), .A2(n6691), .ZN(n5123) );
  INV_X1 U5753 ( .A(n5123), .ZN(n6481) );
  NOR2_X1 U5754 ( .A1(n4648), .A2(n3318), .ZN(n6479) );
  INV_X1 U5755 ( .A(n6479), .ZN(n4994) );
  NOR2_X1 U5756 ( .A1(n6228), .A2(n5013), .ZN(n6388) );
  OAI22_X1 U5757 ( .A1(n4994), .A2(n4650), .B1(n4649), .B2(n6484), .ZN(n4642)
         );
  AOI21_X1 U5758 ( .B1(n6481), .B2(n4652), .A(n4642), .ZN(n4643) );
  OAI211_X1 U5759 ( .C1(n4655), .C2(n5889), .A(n4644), .B(n4643), .ZN(U3057)
         );
  INV_X1 U5760 ( .A(DATAI_18_), .ZN(n4645) );
  OR2_X1 U5761 ( .A1(n6283), .A2(n4645), .ZN(n5877) );
  NAND2_X1 U5762 ( .A1(n4646), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4654) );
  INV_X1 U5763 ( .A(DATAI_26_), .ZN(n4647) );
  OR2_X1 U5764 ( .A1(n6283), .A2(n4647), .ZN(n5139) );
  INV_X1 U5765 ( .A(n5139), .ZN(n6463) );
  NOR2_X1 U5766 ( .A1(n4648), .A2(n3342), .ZN(n6461) );
  INV_X1 U5767 ( .A(n6461), .ZN(n4965) );
  NOR2_X1 U5768 ( .A1(n6878), .A2(n5013), .ZN(n6377) );
  OAI22_X1 U5769 ( .A1(n4965), .A2(n4650), .B1(n4649), .B2(n6466), .ZN(n4651)
         );
  AOI21_X1 U5770 ( .B1(n6463), .B2(n4652), .A(n4651), .ZN(n4653) );
  OAI211_X1 U5771 ( .C1(n4655), .C2(n5877), .A(n4654), .B(n4653), .ZN(U3054)
         );
  AND2_X1 U5772 ( .A1(n4553), .A2(n4656), .ZN(n4657) );
  NAND3_X1 U5773 ( .A1(n4602), .A2(n4885), .A3(n4658), .ZN(n5105) );
  AOI21_X1 U5774 ( .B1(n5149), .B2(n4720), .A(n6657), .ZN(n4663) );
  NAND2_X1 U5775 ( .A1(n4451), .A2(n4554), .ZN(n5108) );
  OAI21_X1 U5776 ( .B1(n5858), .B2(n5108), .A(n6411), .ZN(n4662) );
  NAND3_X1 U5777 ( .A1(n6641), .A2(n4887), .A3(n6969), .ZN(n5112) );
  NOR2_X1 U5778 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5112), .ZN(n4664)
         );
  OAI21_X1 U5779 ( .B1(n6365), .B2(n4664), .A(n4659), .ZN(n4660) );
  INV_X1 U5780 ( .A(n4660), .ZN(n4661) );
  OAI211_X1 U5781 ( .C1(n4663), .C2(n4662), .A(n4661), .B(n6368), .ZN(n4687)
         );
  NAND2_X1 U5782 ( .A1(n4687), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4668) );
  INV_X1 U5783 ( .A(n5893), .ZN(n6487) );
  INV_X1 U5784 ( .A(n4664), .ZN(n4689) );
  INV_X1 U5785 ( .A(n5108), .ZN(n4888) );
  INV_X1 U5786 ( .A(n6363), .ZN(n5861) );
  AOI22_X1 U5787 ( .A1(n4819), .A2(n4888), .B1(n5861), .B2(n4665), .ZN(n4688)
         );
  OAI22_X1 U5788 ( .A1(n4987), .A2(n4689), .B1(n4688), .B2(n6490), .ZN(n4666)
         );
  AOI21_X1 U5789 ( .B1(n6487), .B2(n4691), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5790 ( .C1(n4720), .C2(n5135), .A(n4668), .B(n4667), .ZN(U3026)
         );
  NAND2_X1 U5791 ( .A1(n4687), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4671) );
  INV_X1 U5792 ( .A(n5117), .ZN(n6444) );
  OAI22_X1 U5793 ( .A1(n4974), .A2(n4689), .B1(n5149), .B2(n5869), .ZN(n4669)
         );
  AOI21_X1 U5794 ( .B1(n6444), .B2(n4746), .A(n4669), .ZN(n4670) );
  OAI211_X1 U5795 ( .C1(n4688), .C2(n6454), .A(n4671), .B(n4670), .ZN(U3020)
         );
  NAND2_X1 U5796 ( .A1(n4687), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4674) );
  INV_X1 U5797 ( .A(n5877), .ZN(n6462) );
  OAI22_X1 U5798 ( .A1(n4965), .A2(n4689), .B1(n4688), .B2(n6466), .ZN(n4672)
         );
  AOI21_X1 U5799 ( .B1(n6462), .B2(n4691), .A(n4672), .ZN(n4673) );
  OAI211_X1 U5800 ( .C1(n4720), .C2(n5139), .A(n4674), .B(n4673), .ZN(U3022)
         );
  NAND2_X1 U5801 ( .A1(n4687), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4677) );
  INV_X1 U5802 ( .A(n5899), .ZN(n6493) );
  OAI22_X1 U5803 ( .A1(n4983), .A2(n4689), .B1(n4688), .B2(n6500), .ZN(n4675)
         );
  AOI21_X1 U5804 ( .B1(n6493), .B2(n4691), .A(n4675), .ZN(n4676) );
  OAI211_X1 U5805 ( .C1(n4720), .C2(n5131), .A(n4677), .B(n4676), .ZN(U3027)
         );
  NAND2_X1 U5806 ( .A1(n4687), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4680) );
  INV_X1 U5807 ( .A(n5873), .ZN(n6456) );
  OAI22_X1 U5808 ( .A1(n4969), .A2(n4689), .B1(n4688), .B2(n6460), .ZN(n4678)
         );
  AOI21_X1 U5809 ( .B1(n6456), .B2(n4691), .A(n4678), .ZN(n4679) );
  OAI211_X1 U5810 ( .C1(n4720), .C2(n5150), .A(n4680), .B(n4679), .ZN(U3021)
         );
  NAND2_X1 U5811 ( .A1(n4687), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4683) );
  INV_X1 U5812 ( .A(n5885), .ZN(n6474) );
  OAI22_X1 U5813 ( .A1(n4961), .A2(n4689), .B1(n4688), .B2(n6478), .ZN(n4681)
         );
  AOI21_X1 U5814 ( .B1(n6474), .B2(n4691), .A(n4681), .ZN(n4682) );
  OAI211_X1 U5815 ( .C1(n4720), .C2(n5143), .A(n4683), .B(n4682), .ZN(U3024)
         );
  NAND2_X1 U5816 ( .A1(n4687), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4686) );
  INV_X1 U5817 ( .A(n5889), .ZN(n6480) );
  OAI22_X1 U5818 ( .A1(n4994), .A2(n4689), .B1(n4688), .B2(n6484), .ZN(n4684)
         );
  AOI21_X1 U5819 ( .B1(n6480), .B2(n4691), .A(n4684), .ZN(n4685) );
  OAI211_X1 U5820 ( .C1(n4720), .C2(n5123), .A(n4686), .B(n4685), .ZN(U3025)
         );
  NAND2_X1 U5821 ( .A1(n4687), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4693) );
  INV_X1 U5822 ( .A(n5881), .ZN(n6468) );
  OAI22_X1 U5823 ( .A1(n4979), .A2(n4689), .B1(n4688), .B2(n6472), .ZN(n4690)
         );
  AOI21_X1 U5824 ( .B1(n6468), .B2(n4691), .A(n4690), .ZN(n4692) );
  OAI211_X1 U5825 ( .C1(n4720), .C2(n5127), .A(n4693), .B(n4692), .ZN(U3023)
         );
  XNOR2_X1 U5826 ( .A(n4694), .B(n4695), .ZN(n4760) );
  OAI22_X1 U5827 ( .A1(n4699), .A2(n4698), .B1(n4697), .B2(n4696), .ZN(n4701)
         );
  OAI21_X1 U5828 ( .B1(n4879), .B2(n5792), .A(n4700), .ZN(n4883) );
  OAI21_X1 U5829 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4701), .A(n4883), 
        .ZN(n4703) );
  AND2_X1 U5830 ( .A1(n6276), .A2(REIP_REG_5__SCAN_IN), .ZN(n4756) );
  AOI21_X1 U5831 ( .B1(n6312), .B2(n6120), .A(n4756), .ZN(n4702) );
  OAI211_X1 U5832 ( .C1(n4760), .C2(n5984), .A(n4703), .B(n4702), .ZN(U3013)
         );
  NAND2_X1 U5833 ( .A1(n6320), .A2(n5821), .ZN(n6309) );
  AOI21_X1 U5834 ( .B1(n6319), .B2(n6309), .A(n3741), .ZN(n4712) );
  AOI211_X1 U5835 ( .C1(n6320), .C2(n6318), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n5792), .ZN(n4711) );
  OR2_X1 U5836 ( .A1(n4705), .A2(n4704), .ZN(n4706) );
  NAND2_X1 U5837 ( .A1(n4707), .A2(n4706), .ZN(n4765) );
  NAND2_X1 U5838 ( .A1(n6312), .A2(n4708), .ZN(n4709) );
  NAND2_X1 U5839 ( .A1(n6276), .A2(REIP_REG_1__SCAN_IN), .ZN(n4764) );
  OAI211_X1 U5840 ( .C1(n5984), .C2(n4765), .A(n4709), .B(n4764), .ZN(n4710)
         );
  OR3_X1 U5841 ( .A1(n4712), .A2(n4711), .A3(n4710), .ZN(U3017) );
  INV_X1 U5842 ( .A(n5858), .ZN(n6635) );
  NOR2_X1 U5843 ( .A1(n6635), .A2(n3911), .ZN(n4889) );
  NOR2_X1 U5844 ( .A1(n4451), .A2(n4554), .ZN(n4960) );
  INV_X1 U5845 ( .A(n4744), .ZN(n4713) );
  AOI21_X1 U5846 ( .B1(n4889), .B2(n4960), .A(n4713), .ZN(n4717) );
  INV_X1 U5847 ( .A(n4717), .ZN(n4715) );
  AOI22_X1 U5848 ( .A1(n4715), .A2(n6411), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4714), .ZN(n4743) );
  OAI21_X1 U5849 ( .B1(n4719), .B2(n6283), .A(n6636), .ZN(n4716) );
  AOI22_X1 U5850 ( .A1(n4717), .A2(n4716), .B1(n6630), .B2(n4956), .ZN(n4718)
         );
  NAND2_X1 U5851 ( .A1(n6448), .A2(n4718), .ZN(n4742) );
  NAND2_X1 U5852 ( .A1(n4742), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4723)
         );
  AND2_X1 U5853 ( .A1(n4719), .A2(n6325), .ZN(n4976) );
  OAI22_X1 U5854 ( .A1(n4974), .A2(n4744), .B1(n5869), .B2(n4720), .ZN(n4721)
         );
  AOI21_X1 U5855 ( .B1(n6444), .B2(n4976), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5856 ( .C1(n4743), .C2(n6454), .A(n4723), .B(n4722), .ZN(U3140)
         );
  NAND2_X1 U5857 ( .A1(n4742), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4726)
         );
  OAI22_X1 U5858 ( .A1(n4965), .A2(n4744), .B1(n4743), .B2(n6466), .ZN(n4724)
         );
  AOI21_X1 U5859 ( .B1(n6462), .B2(n4746), .A(n4724), .ZN(n4725) );
  OAI211_X1 U5860 ( .C1(n4999), .C2(n5139), .A(n4726), .B(n4725), .ZN(U3142)
         );
  NAND2_X1 U5861 ( .A1(n4742), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4729)
         );
  OAI22_X1 U5862 ( .A1(n4969), .A2(n4744), .B1(n4743), .B2(n6460), .ZN(n4727)
         );
  AOI21_X1 U5863 ( .B1(n6456), .B2(n4746), .A(n4727), .ZN(n4728) );
  OAI211_X1 U5864 ( .C1(n4999), .C2(n5150), .A(n4729), .B(n4728), .ZN(U3141)
         );
  NAND2_X1 U5865 ( .A1(n4742), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4732)
         );
  OAI22_X1 U5866 ( .A1(n4987), .A2(n4744), .B1(n4743), .B2(n6490), .ZN(n4730)
         );
  AOI21_X1 U5867 ( .B1(n6487), .B2(n4746), .A(n4730), .ZN(n4731) );
  OAI211_X1 U5868 ( .C1(n4999), .C2(n5135), .A(n4732), .B(n4731), .ZN(U3146)
         );
  NAND2_X1 U5869 ( .A1(n4742), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4735)
         );
  OAI22_X1 U5870 ( .A1(n4961), .A2(n4744), .B1(n4743), .B2(n6478), .ZN(n4733)
         );
  AOI21_X1 U5871 ( .B1(n6474), .B2(n4746), .A(n4733), .ZN(n4734) );
  OAI211_X1 U5872 ( .C1(n4999), .C2(n5143), .A(n4735), .B(n4734), .ZN(U3144)
         );
  NAND2_X1 U5873 ( .A1(n4742), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4738)
         );
  OAI22_X1 U5874 ( .A1(n4983), .A2(n4744), .B1(n4743), .B2(n6500), .ZN(n4736)
         );
  AOI21_X1 U5875 ( .B1(n6493), .B2(n4746), .A(n4736), .ZN(n4737) );
  OAI211_X1 U5876 ( .C1(n4999), .C2(n5131), .A(n4738), .B(n4737), .ZN(U3147)
         );
  NAND2_X1 U5877 ( .A1(n4742), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4741)
         );
  OAI22_X1 U5878 ( .A1(n4994), .A2(n4744), .B1(n4743), .B2(n6484), .ZN(n4739)
         );
  AOI21_X1 U5879 ( .B1(n6480), .B2(n4746), .A(n4739), .ZN(n4740) );
  OAI211_X1 U5880 ( .C1(n4999), .C2(n5123), .A(n4741), .B(n4740), .ZN(U3145)
         );
  NAND2_X1 U5881 ( .A1(n4742), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4748)
         );
  OAI22_X1 U5882 ( .A1(n4979), .A2(n4744), .B1(n4743), .B2(n6472), .ZN(n4745)
         );
  AOI21_X1 U5883 ( .B1(n6468), .B2(n4746), .A(n4745), .ZN(n4747) );
  OAI211_X1 U5884 ( .C1(n4999), .C2(n5127), .A(n4748), .B(n4747), .ZN(U3143)
         );
  INV_X1 U5885 ( .A(n6283), .ZN(n6260) );
  AOI21_X1 U5886 ( .B1(n6280), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4749), 
        .ZN(n4750) );
  OAI21_X1 U5887 ( .B1(n5200), .B2(n6272), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5888 ( .B1(n4752), .B2(n6260), .A(n4751), .ZN(n4753) );
  OAI21_X1 U5889 ( .B1(n4754), .B2(n5695), .A(n4753), .ZN(U2983) );
  INV_X1 U5890 ( .A(n4755), .ZN(n6128) );
  AOI21_X1 U5891 ( .B1(n6280), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4756), 
        .ZN(n4757) );
  OAI21_X1 U5892 ( .B1(n6130), .B2(n6272), .A(n4757), .ZN(n4758) );
  AOI21_X1 U5893 ( .B1(n6128), .B2(n6260), .A(n4758), .ZN(n4759) );
  OAI21_X1 U5894 ( .B1(n4760), .B2(n5695), .A(n4759), .ZN(U2981) );
  AND2_X1 U5895 ( .A1(n4513), .A2(n4761), .ZN(n4763) );
  OR2_X1 U5896 ( .A1(n4763), .A2(n4762), .ZN(n5161) );
  INV_X1 U5897 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6186) );
  OAI222_X1 U5898 ( .A1(n5161), .A2(n6169), .B1(n6167), .B2(n6230), .C1(n6168), 
        .C2(n6186), .ZN(U2885) );
  INV_X1 U5899 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4768) );
  OAI21_X1 U5900 ( .B1(n6266), .B2(n4768), .A(n4764), .ZN(n4767) );
  NOR2_X1 U5901 ( .A1(n4765), .A2(n6277), .ZN(n4766) );
  AOI211_X1 U5902 ( .C1(n6258), .C2(n4768), .A(n4767), .B(n4766), .ZN(n4769)
         );
  OAI21_X1 U5903 ( .B1(n6283), .B2(n5196), .A(n4769), .ZN(U2985) );
  NAND2_X1 U5904 ( .A1(n4771), .A2(n4770), .ZN(n4772) );
  NAND2_X1 U5905 ( .A1(n4923), .A2(n4772), .ZN(n5156) );
  INV_X1 U5906 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4773) );
  OAI222_X1 U5907 ( .A1(n5156), .A2(n5532), .B1(n6156), .B2(n4773), .C1(n5528), 
        .C2(n5161), .ZN(U2853) );
  INV_X1 U5908 ( .A(n6435), .ZN(n5856) );
  NOR2_X1 U5909 ( .A1(n4553), .A2(n4774), .ZN(n4775) );
  NAND2_X1 U5910 ( .A1(n4559), .A2(n4775), .ZN(n4856) );
  INV_X1 U5911 ( .A(n4856), .ZN(n4850) );
  NAND2_X1 U5912 ( .A1(n4850), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5913 ( .A1(n5856), .A2(n4853), .ZN(n6629) );
  NOR3_X1 U5914 ( .A1(n6629), .A2(n4559), .A3(n6407), .ZN(n4776) );
  NOR2_X1 U5915 ( .A1(n4776), .A2(n6630), .ZN(n4783) );
  OR2_X1 U5916 ( .A1(n5858), .A2(n3911), .ZN(n5109) );
  INV_X1 U5917 ( .A(n5109), .ZN(n4777) );
  AND2_X1 U5918 ( .A1(n4451), .A2(n5843), .ZN(n5859) );
  NOR2_X1 U5919 ( .A1(n6438), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4780)
         );
  AOI21_X1 U5920 ( .B1(n4777), .B2(n5859), .A(n4780), .ZN(n4782) );
  INV_X1 U5921 ( .A(n4782), .ZN(n4778) );
  NAND2_X1 U5922 ( .A1(n5862), .A2(n6641), .ZN(n4815) );
  INV_X1 U5923 ( .A(n4815), .ZN(n4785) );
  AOI22_X1 U5924 ( .A1(n4783), .A2(n4778), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4785), .ZN(n4812) );
  INV_X1 U5925 ( .A(n4780), .ZN(n4807) );
  OAI22_X1 U5926 ( .A1(n4969), .A2(n4807), .B1(n4806), .B2(n5873), .ZN(n4781)
         );
  AOI21_X1 U5927 ( .B1(n6457), .B2(n4846), .A(n4781), .ZN(n4787) );
  NAND2_X1 U5928 ( .A1(n4783), .A2(n4782), .ZN(n4784) );
  OAI211_X1 U5929 ( .C1(n6411), .C2(n4785), .A(n4784), .B(n6448), .ZN(n4809)
         );
  NAND2_X1 U5930 ( .A1(n4809), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4786) );
  OAI211_X1 U5931 ( .C1(n4812), .C2(n6460), .A(n4787), .B(n4786), .ZN(U3045)
         );
  OAI22_X1 U5932 ( .A1(n4974), .A2(n4807), .B1(n4806), .B2(n5869), .ZN(n4788)
         );
  AOI21_X1 U5933 ( .B1(n6444), .B2(n4846), .A(n4788), .ZN(n4790) );
  NAND2_X1 U5934 ( .A1(n4809), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4789) );
  OAI211_X1 U5935 ( .C1(n4812), .C2(n6454), .A(n4790), .B(n4789), .ZN(U3044)
         );
  OAI22_X1 U5936 ( .A1(n4983), .A2(n4807), .B1(n4806), .B2(n5899), .ZN(n4791)
         );
  AOI21_X1 U5937 ( .B1(n6496), .B2(n4846), .A(n4791), .ZN(n4793) );
  NAND2_X1 U5938 ( .A1(n4809), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4792) );
  OAI211_X1 U5939 ( .C1(n4812), .C2(n6500), .A(n4793), .B(n4792), .ZN(U3051)
         );
  OAI22_X1 U5940 ( .A1(n4987), .A2(n4807), .B1(n4806), .B2(n5893), .ZN(n4794)
         );
  AOI21_X1 U5941 ( .B1(n6486), .B2(n4846), .A(n4794), .ZN(n4796) );
  NAND2_X1 U5942 ( .A1(n4809), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4795) );
  OAI211_X1 U5943 ( .C1(n4812), .C2(n6490), .A(n4796), .B(n4795), .ZN(U3050)
         );
  OAI22_X1 U5944 ( .A1(n4994), .A2(n4807), .B1(n4806), .B2(n5889), .ZN(n4797)
         );
  AOI21_X1 U5945 ( .B1(n6481), .B2(n4846), .A(n4797), .ZN(n4799) );
  NAND2_X1 U5946 ( .A1(n4809), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4798) );
  OAI211_X1 U5947 ( .C1(n4812), .C2(n6484), .A(n4799), .B(n4798), .ZN(U3049)
         );
  OAI22_X1 U5948 ( .A1(n4961), .A2(n4807), .B1(n4806), .B2(n5885), .ZN(n4800)
         );
  AOI21_X1 U5949 ( .B1(n6475), .B2(n4846), .A(n4800), .ZN(n4802) );
  NAND2_X1 U5950 ( .A1(n4809), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4801) );
  OAI211_X1 U5951 ( .C1(n4812), .C2(n6478), .A(n4802), .B(n4801), .ZN(U3048)
         );
  OAI22_X1 U5952 ( .A1(n4965), .A2(n4807), .B1(n4806), .B2(n5877), .ZN(n4803)
         );
  AOI21_X1 U5953 ( .B1(n6463), .B2(n4846), .A(n4803), .ZN(n4805) );
  NAND2_X1 U5954 ( .A1(n4809), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4804) );
  OAI211_X1 U5955 ( .C1(n4812), .C2(n6466), .A(n4805), .B(n4804), .ZN(U3046)
         );
  OAI22_X1 U5956 ( .A1(n4979), .A2(n4807), .B1(n4806), .B2(n5881), .ZN(n4808)
         );
  AOI21_X1 U5957 ( .B1(n6469), .B2(n4846), .A(n4808), .ZN(n4811) );
  NAND2_X1 U5958 ( .A1(n4809), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4810) );
  OAI211_X1 U5959 ( .C1(n4812), .C2(n6472), .A(n4811), .B(n4810), .ZN(U3047)
         );
  NAND2_X1 U5960 ( .A1(n4849), .A2(n4829), .ZN(n4813) );
  AOI22_X1 U5961 ( .A1(n4813), .A2(n6636), .B1(n6635), .B2(n5859), .ZN(n4814)
         );
  NOR2_X1 U5962 ( .A1(n4814), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4816) );
  NOR2_X1 U5963 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4815), .ZN(n4817)
         );
  NAND2_X1 U5964 ( .A1(n5006), .A2(n6641), .ZN(n6369) );
  AOI21_X1 U5965 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6369), .A(n5013), .ZN(
        n6364) );
  NAND2_X1 U5966 ( .A1(n4842), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4822) );
  INV_X1 U5967 ( .A(n4817), .ZN(n4844) );
  INV_X1 U5968 ( .A(n6369), .ZN(n4818) );
  AOI22_X1 U5969 ( .A1(n4819), .A2(n5859), .B1(n5861), .B2(n4818), .ZN(n4843)
         );
  OAI22_X1 U5970 ( .A1(n4987), .A2(n4844), .B1(n4843), .B2(n6490), .ZN(n4820)
         );
  AOI21_X1 U5971 ( .B1(n6487), .B2(n4846), .A(n4820), .ZN(n4821) );
  OAI211_X1 U5972 ( .C1(n4849), .C2(n5135), .A(n4822), .B(n4821), .ZN(U3042)
         );
  NAND2_X1 U5973 ( .A1(n4842), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4825) );
  OAI22_X1 U5974 ( .A1(n4983), .A2(n4844), .B1(n4843), .B2(n6500), .ZN(n4823)
         );
  AOI21_X1 U5975 ( .B1(n6493), .B2(n4846), .A(n4823), .ZN(n4824) );
  OAI211_X1 U5976 ( .C1(n4849), .C2(n5131), .A(n4825), .B(n4824), .ZN(U3043)
         );
  NAND2_X1 U5977 ( .A1(n4842), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4828) );
  OAI22_X1 U5978 ( .A1(n4979), .A2(n4844), .B1(n4843), .B2(n6472), .ZN(n4826)
         );
  AOI21_X1 U5979 ( .B1(n6468), .B2(n4846), .A(n4826), .ZN(n4827) );
  OAI211_X1 U5980 ( .C1(n4849), .C2(n5127), .A(n4828), .B(n4827), .ZN(U3039)
         );
  NAND2_X1 U5981 ( .A1(n4842), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4832) );
  OAI22_X1 U5982 ( .A1(n4974), .A2(n4844), .B1(n4829), .B2(n5869), .ZN(n4830)
         );
  AOI21_X1 U5983 ( .B1(n6444), .B2(n5152), .A(n4830), .ZN(n4831) );
  OAI211_X1 U5984 ( .C1(n4843), .C2(n6454), .A(n4832), .B(n4831), .ZN(U3036)
         );
  NAND2_X1 U5985 ( .A1(n4842), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4835) );
  OAI22_X1 U5986 ( .A1(n4969), .A2(n4844), .B1(n4843), .B2(n6460), .ZN(n4833)
         );
  AOI21_X1 U5987 ( .B1(n6456), .B2(n4846), .A(n4833), .ZN(n4834) );
  OAI211_X1 U5988 ( .C1(n4849), .C2(n5150), .A(n4835), .B(n4834), .ZN(U3037)
         );
  NAND2_X1 U5989 ( .A1(n4842), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4838) );
  OAI22_X1 U5990 ( .A1(n4965), .A2(n4844), .B1(n4843), .B2(n6466), .ZN(n4836)
         );
  AOI21_X1 U5991 ( .B1(n6462), .B2(n4846), .A(n4836), .ZN(n4837) );
  OAI211_X1 U5992 ( .C1(n4849), .C2(n5139), .A(n4838), .B(n4837), .ZN(U3038)
         );
  NAND2_X1 U5993 ( .A1(n4842), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4841) );
  OAI22_X1 U5994 ( .A1(n4961), .A2(n4844), .B1(n4843), .B2(n6478), .ZN(n4839)
         );
  AOI21_X1 U5995 ( .B1(n6474), .B2(n4846), .A(n4839), .ZN(n4840) );
  OAI211_X1 U5996 ( .C1(n4849), .C2(n5143), .A(n4841), .B(n4840), .ZN(U3040)
         );
  NAND2_X1 U5997 ( .A1(n4842), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4848) );
  OAI22_X1 U5998 ( .A1(n4994), .A2(n4844), .B1(n4843), .B2(n6484), .ZN(n4845)
         );
  AOI21_X1 U5999 ( .B1(n6480), .B2(n4846), .A(n4845), .ZN(n4847) );
  OAI211_X1 U6000 ( .C1(n4849), .C2(n5123), .A(n4848), .B(n4847), .ZN(U3041)
         );
  NAND3_X1 U6001 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6969), .ZN(n5012) );
  INV_X1 U6002 ( .A(n5012), .ZN(n4852) );
  NOR2_X1 U6003 ( .A1(n6362), .A2(n5012), .ZN(n4873) );
  AOI21_X1 U6004 ( .B1(n4889), .B2(n6322), .A(n4873), .ZN(n4855) );
  NAND3_X1 U6005 ( .A1(n6411), .A2(n4855), .A3(n4853), .ZN(n4851) );
  OAI211_X1 U6006 ( .C1(n6411), .C2(n4852), .A(n6448), .B(n4851), .ZN(n4872)
         );
  NAND2_X1 U6007 ( .A1(n6411), .A2(n4853), .ZN(n4854) );
  OAI22_X1 U6008 ( .A1(n4855), .A2(n4854), .B1(n6656), .B2(n5012), .ZN(n4871)
         );
  AOI22_X1 U6009 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4872), .B1(n6374), 
        .B2(n4871), .ZN(n4858) );
  AOI22_X1 U6010 ( .A1(n6455), .A2(n4873), .B1(n5014), .B2(n6457), .ZN(n4857)
         );
  OAI211_X1 U6011 ( .C1(n5873), .C2(n4973), .A(n4858), .B(n4857), .ZN(U3125)
         );
  AOI22_X1 U6012 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4872), .B1(n6371), 
        .B2(n4871), .ZN(n4860) );
  AOI22_X1 U6013 ( .A1(n6443), .A2(n4873), .B1(n5014), .B2(n6444), .ZN(n4859)
         );
  OAI211_X1 U6014 ( .C1(n5869), .C2(n4973), .A(n4860), .B(n4859), .ZN(U3124)
         );
  AOI22_X1 U6015 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4872), .B1(n6377), 
        .B2(n4871), .ZN(n4862) );
  AOI22_X1 U6016 ( .A1(n6461), .A2(n4873), .B1(n5014), .B2(n6463), .ZN(n4861)
         );
  OAI211_X1 U6017 ( .C1(n5877), .C2(n4973), .A(n4862), .B(n4861), .ZN(U3126)
         );
  AOI22_X1 U6018 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4872), .B1(n6397), 
        .B2(n4871), .ZN(n4864) );
  AOI22_X1 U6019 ( .A1(n6492), .A2(n4873), .B1(n5014), .B2(n6496), .ZN(n4863)
         );
  OAI211_X1 U6020 ( .C1(n5899), .C2(n4973), .A(n4864), .B(n4863), .ZN(U3131)
         );
  AOI22_X1 U6021 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4872), .B1(n6392), 
        .B2(n4871), .ZN(n4866) );
  AOI22_X1 U6022 ( .A1(n6485), .A2(n4873), .B1(n5014), .B2(n6486), .ZN(n4865)
         );
  OAI211_X1 U6023 ( .C1(n5893), .C2(n4973), .A(n4866), .B(n4865), .ZN(U3130)
         );
  AOI22_X1 U6024 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4872), .B1(n6388), 
        .B2(n4871), .ZN(n4868) );
  AOI22_X1 U6025 ( .A1(n6479), .A2(n4873), .B1(n5014), .B2(n6481), .ZN(n4867)
         );
  OAI211_X1 U6026 ( .C1(n5889), .C2(n4973), .A(n4868), .B(n4867), .ZN(U3129)
         );
  AOI22_X1 U6027 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4872), .B1(n6385), 
        .B2(n4871), .ZN(n4870) );
  AOI22_X1 U6028 ( .A1(n6473), .A2(n4873), .B1(n5014), .B2(n6475), .ZN(n4869)
         );
  OAI211_X1 U6029 ( .C1(n5885), .C2(n4973), .A(n4870), .B(n4869), .ZN(U3128)
         );
  AOI22_X1 U6030 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4872), .B1(n6381), 
        .B2(n4871), .ZN(n4875) );
  AOI22_X1 U6031 ( .A1(n6467), .A2(n4873), .B1(n5014), .B2(n6469), .ZN(n4874)
         );
  OAI211_X1 U6032 ( .C1(n5881), .C2(n4973), .A(n4875), .B(n4874), .ZN(U3127)
         );
  XNOR2_X1 U6033 ( .A(n4877), .B(n3098), .ZN(n4921) );
  NAND2_X1 U6034 ( .A1(n6276), .A2(REIP_REG_6__SCAN_IN), .ZN(n4917) );
  OAI21_X1 U6035 ( .B1(n6018), .B2(n5156), .A(n4917), .ZN(n4882) );
  NAND2_X1 U6036 ( .A1(n4879), .A2(n4878), .ZN(n4880) );
  NOR2_X1 U6037 ( .A1(n5171), .A2(n4880), .ZN(n4881) );
  AOI211_X1 U6038 ( .C1(n4883), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4882), 
        .B(n4881), .ZN(n4884) );
  OAI21_X1 U6039 ( .B1(n5984), .B2(n4921), .A(n4884), .ZN(U3012) );
  NAND2_X1 U6040 ( .A1(n6435), .A2(n4885), .ZN(n4895) );
  INV_X1 U6041 ( .A(n4895), .ZN(n4886) );
  NAND3_X1 U6042 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4887), .A3(n6969), .ZN(n5026) );
  NOR2_X1 U6043 ( .A1(n6362), .A2(n5026), .ZN(n4912) );
  AOI21_X1 U6044 ( .B1(n4889), .B2(n4888), .A(n4912), .ZN(n4893) );
  OR2_X1 U6045 ( .A1(n4895), .A2(n6657), .ZN(n4890) );
  AOI22_X1 U6046 ( .A1(n4893), .A2(n4892), .B1(n6630), .B2(n5026), .ZN(n4891)
         );
  NAND2_X1 U6047 ( .A1(n6448), .A2(n4891), .ZN(n4911) );
  INV_X1 U6048 ( .A(n4892), .ZN(n4894) );
  OAI22_X1 U6049 ( .A1(n4894), .A2(n4893), .B1(n6656), .B2(n5026), .ZN(n4910)
         );
  AOI22_X1 U6050 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4911), .B1(n6397), 
        .B2(n4910), .ZN(n4897) );
  AOI22_X1 U6051 ( .A1(n5902), .A2(n6493), .B1(n4912), .B2(n6492), .ZN(n4896)
         );
  OAI211_X1 U6052 ( .C1(n5066), .C2(n5131), .A(n4897), .B(n4896), .ZN(U3099)
         );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4911), .B1(n6392), 
        .B2(n4910), .ZN(n4899) );
  AOI22_X1 U6054 ( .A1(n5902), .A2(n6487), .B1(n4912), .B2(n6485), .ZN(n4898)
         );
  OAI211_X1 U6055 ( .C1(n5066), .C2(n5135), .A(n4899), .B(n4898), .ZN(U3098)
         );
  AOI22_X1 U6056 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4911), .B1(n6381), 
        .B2(n4910), .ZN(n4901) );
  AOI22_X1 U6057 ( .A1(n5902), .A2(n6468), .B1(n4912), .B2(n6467), .ZN(n4900)
         );
  OAI211_X1 U6058 ( .C1(n5066), .C2(n5127), .A(n4901), .B(n4900), .ZN(U3095)
         );
  AOI22_X1 U6059 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4911), .B1(n6374), 
        .B2(n4910), .ZN(n4903) );
  AOI22_X1 U6060 ( .A1(n5902), .A2(n6456), .B1(n4912), .B2(n6455), .ZN(n4902)
         );
  OAI211_X1 U6061 ( .C1(n5066), .C2(n5150), .A(n4903), .B(n4902), .ZN(U3093)
         );
  AOI22_X1 U6062 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4911), .B1(n6371), 
        .B2(n4910), .ZN(n4905) );
  AOI22_X1 U6063 ( .A1(n5902), .A2(n6451), .B1(n6443), .B2(n4912), .ZN(n4904)
         );
  OAI211_X1 U6064 ( .C1(n5117), .C2(n5066), .A(n4905), .B(n4904), .ZN(U3092)
         );
  AOI22_X1 U6065 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4911), .B1(n6385), 
        .B2(n4910), .ZN(n4907) );
  AOI22_X1 U6066 ( .A1(n5902), .A2(n6474), .B1(n4912), .B2(n6473), .ZN(n4906)
         );
  OAI211_X1 U6067 ( .C1(n5066), .C2(n5143), .A(n4907), .B(n4906), .ZN(U3096)
         );
  AOI22_X1 U6068 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4911), .B1(n6377), 
        .B2(n4910), .ZN(n4909) );
  AOI22_X1 U6069 ( .A1(n5902), .A2(n6462), .B1(n4912), .B2(n6461), .ZN(n4908)
         );
  OAI211_X1 U6070 ( .C1(n5066), .C2(n5139), .A(n4909), .B(n4908), .ZN(U3094)
         );
  AOI22_X1 U6071 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4911), .B1(n6388), 
        .B2(n4910), .ZN(n4914) );
  AOI22_X1 U6072 ( .A1(n5902), .A2(n6480), .B1(n4912), .B2(n6479), .ZN(n4913)
         );
  OAI211_X1 U6073 ( .C1(n5066), .C2(n5123), .A(n4914), .B(n4913), .ZN(U3097)
         );
  INV_X1 U6074 ( .A(n5161), .ZN(n4919) );
  INV_X1 U6075 ( .A(n4915), .ZN(n5160) );
  NAND2_X1 U6076 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4916)
         );
  OAI211_X1 U6077 ( .C1(n6272), .C2(n5160), .A(n4917), .B(n4916), .ZN(n4918)
         );
  AOI21_X1 U6078 ( .B1(n4919), .B2(n6260), .A(n4918), .ZN(n4920) );
  OAI21_X1 U6079 ( .B1(n4921), .B2(n5695), .A(n4920), .ZN(U2980) );
  AND2_X1 U6080 ( .A1(n4923), .A2(n4922), .ZN(n4924) );
  NOR2_X1 U6081 ( .A1(n5184), .A2(n4924), .ZN(n6302) );
  INV_X1 U6082 ( .A(n6302), .ZN(n4928) );
  INV_X1 U6083 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6953) );
  OR2_X1 U6084 ( .A1(n4762), .A2(n4926), .ZN(n4927) );
  AND2_X1 U6085 ( .A1(n4925), .A2(n4927), .ZN(n6115) );
  INV_X1 U6086 ( .A(n6115), .ZN(n4929) );
  OAI222_X1 U6087 ( .A1(n4928), .A2(n5532), .B1(n6156), .B2(n6953), .C1(n5528), 
        .C2(n4929), .ZN(U2852) );
  OAI222_X1 U6088 ( .A1(n4929), .A2(n6169), .B1(n6167), .B2(n6232), .C1(n6168), 
        .C2(n3904), .ZN(U2884) );
  NAND3_X1 U6089 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n4930), .ZN(n6541) );
  NAND3_X1 U6090 ( .A1(n6660), .A2(STATE2_REG_1__SCAN_IN), .A3(n4931), .ZN(
        n6543) );
  NAND2_X4 U6091 ( .A1(n6662), .A2(n4932), .ZN(n5204) );
  OAI21_X1 U6092 ( .B1(n4938), .B2(n6034), .A(n5905), .ZN(n6146) );
  INV_X1 U6093 ( .A(n6146), .ZN(n5284) );
  NAND2_X1 U6094 ( .A1(n4438), .A2(n6657), .ZN(n6533) );
  NOR2_X1 U6095 ( .A1(n4938), .A2(n6533), .ZN(n4935) );
  NAND3_X1 U6096 ( .A1(n4935), .A2(n3734), .A3(n4934), .ZN(n6140) );
  NAND2_X1 U6097 ( .A1(n5204), .A2(n6140), .ZN(n6086) );
  NOR2_X1 U6098 ( .A1(n4936), .A2(n4938), .ZN(n6137) );
  INV_X1 U6099 ( .A(n6137), .ZN(n5199) );
  INV_X1 U6100 ( .A(n4937), .ZN(n6311) );
  INV_X1 U6101 ( .A(n4938), .ZN(n4941) );
  OAI21_X1 U6102 ( .B1(n6563), .B2(n6533), .A(n4941), .ZN(n4942) );
  INV_X1 U6103 ( .A(n4942), .ZN(n4943) );
  AND2_X1 U6104 ( .A1(n6658), .A2(n4943), .ZN(n5343) );
  INV_X1 U6105 ( .A(n4944), .ZN(n4945) );
  NOR2_X1 U6106 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4945), .ZN(n4946) );
  AND2_X1 U6107 ( .A1(n3734), .A2(n4946), .ZN(n4947) );
  AOI22_X1 U6108 ( .A1(n6311), .A2(n6119), .B1(EBX_REG_0__SCAN_IN), .B2(n6118), 
        .ZN(n4948) );
  OAI21_X1 U6109 ( .B1(n3911), .B2(n5199), .A(n4948), .ZN(n4949) );
  AOI21_X1 U6110 ( .B1(n6086), .B2(REIP_REG_0__SCAN_IN), .A(n4949), .ZN(n4953)
         );
  NOR2_X1 U6111 ( .A1(n4950), .A2(n6552), .ZN(n4951) );
  OAI21_X1 U6112 ( .B1(n6097), .B2(n6099), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4952) );
  OAI211_X1 U6113 ( .C1(n5284), .C2(n6284), .A(n4953), .B(n4952), .ZN(U2827)
         );
  NOR3_X1 U6114 ( .A1(n4996), .A2(n4976), .A3(n6630), .ZN(n4955) );
  INV_X1 U6115 ( .A(n4960), .ZN(n6360) );
  OAI22_X1 U6116 ( .A1(n4955), .A2(n4954), .B1(n6635), .B2(n6360), .ZN(n4958)
         );
  NAND2_X1 U6117 ( .A1(n5006), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4959) );
  AOI21_X1 U6118 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4959), .A(n5013), .ZN(
        n5867) );
  OR2_X1 U6119 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4956), .ZN(n4993)
         );
  NAND2_X1 U6120 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4993), .ZN(n4957) );
  NAND4_X1 U6121 ( .A1(n4958), .A2(n5867), .A3(n6363), .A4(n4957), .ZN(n4991)
         );
  NAND2_X1 U6122 ( .A1(n4991), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4964)
         );
  NAND2_X1 U6123 ( .A1(n5858), .A2(n6411), .ZN(n5030) );
  INV_X1 U6124 ( .A(n5030), .ZN(n5011) );
  INV_X1 U6125 ( .A(n4959), .ZN(n5860) );
  AOI22_X1 U6126 ( .A1(n5011), .A2(n4960), .B1(n5860), .B2(n5010), .ZN(n4992)
         );
  OAI22_X1 U6127 ( .A1(n4961), .A2(n4993), .B1(n4992), .B2(n6478), .ZN(n4962)
         );
  AOI21_X1 U6128 ( .B1(n6475), .B2(n4996), .A(n4962), .ZN(n4963) );
  OAI211_X1 U6129 ( .C1(n4999), .C2(n5885), .A(n4964), .B(n4963), .ZN(U3136)
         );
  NAND2_X1 U6130 ( .A1(n4991), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4968)
         );
  OAI22_X1 U6131 ( .A1(n4965), .A2(n4993), .B1(n4992), .B2(n6466), .ZN(n4966)
         );
  AOI21_X1 U6132 ( .B1(n6463), .B2(n4996), .A(n4966), .ZN(n4967) );
  OAI211_X1 U6133 ( .C1(n4999), .C2(n5877), .A(n4968), .B(n4967), .ZN(U3134)
         );
  NAND2_X1 U6134 ( .A1(n4991), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4972)
         );
  OAI22_X1 U6135 ( .A1(n4969), .A2(n4993), .B1(n4992), .B2(n6460), .ZN(n4970)
         );
  AOI21_X1 U6136 ( .B1(n6457), .B2(n4996), .A(n4970), .ZN(n4971) );
  OAI211_X1 U6137 ( .C1(n4999), .C2(n5873), .A(n4972), .B(n4971), .ZN(U3133)
         );
  NAND2_X1 U6138 ( .A1(n4991), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4978)
         );
  OAI22_X1 U6139 ( .A1(n4974), .A2(n4993), .B1(n5117), .B2(n4973), .ZN(n4975)
         );
  AOI21_X1 U6140 ( .B1(n6451), .B2(n4976), .A(n4975), .ZN(n4977) );
  OAI211_X1 U6141 ( .C1(n4992), .C2(n6454), .A(n4978), .B(n4977), .ZN(U3132)
         );
  NAND2_X1 U6142 ( .A1(n4991), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4982)
         );
  OAI22_X1 U6143 ( .A1(n4979), .A2(n4993), .B1(n4992), .B2(n6472), .ZN(n4980)
         );
  AOI21_X1 U6144 ( .B1(n6469), .B2(n4996), .A(n4980), .ZN(n4981) );
  OAI211_X1 U6145 ( .C1(n4999), .C2(n5881), .A(n4982), .B(n4981), .ZN(U3135)
         );
  NAND2_X1 U6146 ( .A1(n4991), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4986)
         );
  OAI22_X1 U6147 ( .A1(n4983), .A2(n4993), .B1(n4992), .B2(n6500), .ZN(n4984)
         );
  AOI21_X1 U6148 ( .B1(n6496), .B2(n4996), .A(n4984), .ZN(n4985) );
  OAI211_X1 U6149 ( .C1(n4999), .C2(n5899), .A(n4986), .B(n4985), .ZN(U3139)
         );
  NAND2_X1 U6150 ( .A1(n4991), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4990)
         );
  OAI22_X1 U6151 ( .A1(n4987), .A2(n4993), .B1(n4992), .B2(n6490), .ZN(n4988)
         );
  AOI21_X1 U6152 ( .B1(n6486), .B2(n4996), .A(n4988), .ZN(n4989) );
  OAI211_X1 U6153 ( .C1(n4999), .C2(n5893), .A(n4990), .B(n4989), .ZN(U3138)
         );
  NAND2_X1 U6154 ( .A1(n4991), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4998)
         );
  OAI22_X1 U6155 ( .A1(n4994), .A2(n4993), .B1(n4992), .B2(n6484), .ZN(n4995)
         );
  AOI21_X1 U6156 ( .B1(n6481), .B2(n4996), .A(n4995), .ZN(n4997) );
  OAI211_X1 U6157 ( .C1(n4999), .C2(n5889), .A(n4998), .B(n4997), .ZN(U3137)
         );
  XNOR2_X1 U6158 ( .A(n5000), .B(n5002), .ZN(n6305) );
  AND2_X1 U6159 ( .A1(n6276), .A2(REIP_REG_7__SCAN_IN), .ZN(n6301) );
  AOI21_X1 U6160 ( .B1(n6280), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6301), 
        .ZN(n5003) );
  OAI21_X1 U6161 ( .B1(n6117), .B2(n6272), .A(n5003), .ZN(n5004) );
  AOI21_X1 U6162 ( .B1(n6115), .B2(n6260), .A(n5004), .ZN(n5005) );
  OAI21_X1 U6163 ( .B1(n6305), .B2(n5695), .A(n5005), .ZN(U2979) );
  INV_X1 U6164 ( .A(n5006), .ZN(n5008) );
  NAND2_X1 U6165 ( .A1(n5008), .A2(n5007), .ZN(n5031) );
  INV_X1 U6166 ( .A(n5031), .ZN(n5009) );
  AOI22_X1 U6167 ( .A1(n5011), .A2(n6322), .B1(n5010), .B2(n5009), .ZN(n5099)
         );
  AND2_X1 U6168 ( .A1(n4553), .A2(n4563), .ZN(n5022) );
  NOR2_X1 U6169 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5012), .ZN(n5101)
         );
  AOI21_X1 U6170 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5031), .A(n5013), .ZN(
        n5027) );
  INV_X1 U6171 ( .A(n5101), .ZN(n5017) );
  AOI21_X1 U6172 ( .B1(n6322), .B2(n6359), .A(n6630), .ZN(n5016) );
  OAI21_X1 U6173 ( .B1(n5014), .B2(n6494), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5015) );
  AOI22_X1 U6174 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5017), .B1(n5016), .B2(
        n5015), .ZN(n5018) );
  NAND3_X1 U6175 ( .A1(n5027), .A2(n5018), .A3(n6363), .ZN(n5073) );
  AOI22_X1 U6176 ( .A1(n6443), .A2(n5101), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n5073), .ZN(n5019) );
  OAI21_X1 U6177 ( .B1(n5869), .B2(n5104), .A(n5019), .ZN(n5020) );
  AOI21_X1 U6178 ( .B1(n6444), .B2(n6494), .A(n5020), .ZN(n5021) );
  OAI21_X1 U6179 ( .B1(n5099), .B2(n6454), .A(n5021), .ZN(U3116) );
  INV_X1 U6180 ( .A(n5066), .ZN(n5023) );
  OAI21_X1 U6181 ( .B1(n5023), .B2(n6429), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5025) );
  OAI211_X1 U6182 ( .C1(n6635), .C2(n5108), .A(n5025), .B(n5024), .ZN(n5029)
         );
  NOR2_X1 U6183 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5026), .ZN(n5063)
         );
  OR2_X1 U6184 ( .A1(n6365), .A2(n5063), .ZN(n5028) );
  NAND4_X1 U6185 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n6368), .ZN(n5068)
         );
  AOI22_X1 U6186 ( .A1(n6443), .A2(n5063), .B1(n6429), .B2(n6444), .ZN(n5035)
         );
  OR2_X1 U6187 ( .A1(n5030), .A2(n5108), .ZN(n5033) );
  OR2_X1 U6188 ( .A1(n6363), .A2(n5031), .ZN(n5032) );
  NAND2_X1 U6189 ( .A1(n5033), .A2(n5032), .ZN(n5062) );
  NAND2_X1 U6190 ( .A1(n6371), .A2(n5062), .ZN(n5034) );
  OAI211_X1 U6191 ( .C1(n5066), .C2(n5869), .A(n5035), .B(n5034), .ZN(n5036)
         );
  AOI21_X1 U6192 ( .B1(n5068), .B2(INSTQUEUE_REG_8__0__SCAN_IN), .A(n5036), 
        .ZN(n5037) );
  INV_X1 U6193 ( .A(n5037), .ZN(U3084) );
  AOI22_X1 U6194 ( .A1(n6461), .A2(n5063), .B1(n6377), .B2(n5062), .ZN(n5039)
         );
  NAND2_X1 U6195 ( .A1(n6429), .A2(n6463), .ZN(n5038) );
  OAI211_X1 U6196 ( .C1(n5066), .C2(n5877), .A(n5039), .B(n5038), .ZN(n5040)
         );
  AOI21_X1 U6197 ( .B1(n5068), .B2(INSTQUEUE_REG_8__2__SCAN_IN), .A(n5040), 
        .ZN(n5041) );
  INV_X1 U6198 ( .A(n5041), .ZN(U3086) );
  AOI22_X1 U6199 ( .A1(n6473), .A2(n5063), .B1(n6385), .B2(n5062), .ZN(n5043)
         );
  NAND2_X1 U6200 ( .A1(n6429), .A2(n6475), .ZN(n5042) );
  OAI211_X1 U6201 ( .C1(n5066), .C2(n5885), .A(n5043), .B(n5042), .ZN(n5044)
         );
  AOI21_X1 U6202 ( .B1(n5068), .B2(INSTQUEUE_REG_8__4__SCAN_IN), .A(n5044), 
        .ZN(n5045) );
  INV_X1 U6203 ( .A(n5045), .ZN(U3088) );
  AOI22_X1 U6204 ( .A1(n6485), .A2(n5063), .B1(n6392), .B2(n5062), .ZN(n5047)
         );
  NAND2_X1 U6205 ( .A1(n6429), .A2(n6486), .ZN(n5046) );
  OAI211_X1 U6206 ( .C1(n5066), .C2(n5893), .A(n5047), .B(n5046), .ZN(n5048)
         );
  AOI21_X1 U6207 ( .B1(n5068), .B2(INSTQUEUE_REG_8__6__SCAN_IN), .A(n5048), 
        .ZN(n5049) );
  INV_X1 U6208 ( .A(n5049), .ZN(U3090) );
  AOI22_X1 U6209 ( .A1(n6492), .A2(n5063), .B1(n6397), .B2(n5062), .ZN(n5051)
         );
  NAND2_X1 U6210 ( .A1(n6429), .A2(n6496), .ZN(n5050) );
  OAI211_X1 U6211 ( .C1(n5066), .C2(n5899), .A(n5051), .B(n5050), .ZN(n5052)
         );
  AOI21_X1 U6212 ( .B1(n5068), .B2(INSTQUEUE_REG_8__7__SCAN_IN), .A(n5052), 
        .ZN(n5053) );
  INV_X1 U6213 ( .A(n5053), .ZN(U3091) );
  AOI22_X1 U6214 ( .A1(n6455), .A2(n5063), .B1(n6374), .B2(n5062), .ZN(n5055)
         );
  NAND2_X1 U6215 ( .A1(n6429), .A2(n6457), .ZN(n5054) );
  OAI211_X1 U6216 ( .C1(n5066), .C2(n5873), .A(n5055), .B(n5054), .ZN(n5056)
         );
  AOI21_X1 U6217 ( .B1(n5068), .B2(INSTQUEUE_REG_8__1__SCAN_IN), .A(n5056), 
        .ZN(n5057) );
  INV_X1 U6218 ( .A(n5057), .ZN(U3085) );
  AOI22_X1 U6219 ( .A1(n6467), .A2(n5063), .B1(n6381), .B2(n5062), .ZN(n5059)
         );
  NAND2_X1 U6220 ( .A1(n6429), .A2(n6469), .ZN(n5058) );
  OAI211_X1 U6221 ( .C1(n5066), .C2(n5881), .A(n5059), .B(n5058), .ZN(n5060)
         );
  AOI21_X1 U6222 ( .B1(n5068), .B2(INSTQUEUE_REG_8__3__SCAN_IN), .A(n5060), 
        .ZN(n5061) );
  INV_X1 U6223 ( .A(n5061), .ZN(U3087) );
  AOI22_X1 U6224 ( .A1(n6479), .A2(n5063), .B1(n6388), .B2(n5062), .ZN(n5065)
         );
  NAND2_X1 U6225 ( .A1(n6429), .A2(n6481), .ZN(n5064) );
  OAI211_X1 U6226 ( .C1(n5066), .C2(n5889), .A(n5065), .B(n5064), .ZN(n5067)
         );
  AOI21_X1 U6227 ( .B1(n5068), .B2(INSTQUEUE_REG_8__5__SCAN_IN), .A(n5067), 
        .ZN(n5069) );
  INV_X1 U6228 ( .A(n5069), .ZN(U3089) );
  AOI21_X1 U6229 ( .B1(n5070), .B2(n4925), .A(n3113), .ZN(n5179) );
  INV_X1 U6230 ( .A(n5179), .ZN(n5218) );
  INV_X1 U6231 ( .A(DATAI_8_), .ZN(n6832) );
  INV_X1 U6232 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6968) );
  OAI222_X1 U6233 ( .A1(n5218), .A2(n6169), .B1(n6167), .B2(n6832), .C1(n6168), 
        .C2(n6968), .ZN(U2883) );
  XNOR2_X1 U6234 ( .A(n5184), .B(n5182), .ZN(n5210) );
  INV_X1 U6235 ( .A(n5210), .ZN(n5072) );
  INV_X1 U6236 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5071) );
  OAI222_X1 U6237 ( .A1(n5218), .A2(n5528), .B1(n5532), .B2(n5072), .C1(n6156), 
        .C2(n5071), .ZN(U2851) );
  NAND2_X1 U6238 ( .A1(n6494), .A2(n6486), .ZN(n5077) );
  INV_X1 U6239 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5074) );
  OAI22_X1 U6240 ( .A1(n5099), .A2(n6490), .B1(n5074), .B2(n5097), .ZN(n5075)
         );
  AOI21_X1 U6241 ( .B1(n6485), .B2(n5101), .A(n5075), .ZN(n5076) );
  OAI211_X1 U6242 ( .C1(n5104), .C2(n5893), .A(n5077), .B(n5076), .ZN(U3122)
         );
  NAND2_X1 U6243 ( .A1(n6494), .A2(n6457), .ZN(n5081) );
  INV_X1 U6244 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5078) );
  OAI22_X1 U6245 ( .A1(n5099), .A2(n6460), .B1(n5078), .B2(n5097), .ZN(n5079)
         );
  AOI21_X1 U6246 ( .B1(n6455), .B2(n5101), .A(n5079), .ZN(n5080) );
  OAI211_X1 U6247 ( .C1(n5104), .C2(n5873), .A(n5081), .B(n5080), .ZN(U3117)
         );
  NAND2_X1 U6248 ( .A1(n6494), .A2(n6463), .ZN(n5084) );
  OAI22_X1 U6249 ( .A1(n5099), .A2(n6466), .B1(n6933), .B2(n5097), .ZN(n5082)
         );
  AOI21_X1 U6250 ( .B1(n6461), .B2(n5101), .A(n5082), .ZN(n5083) );
  OAI211_X1 U6251 ( .C1(n5104), .C2(n5877), .A(n5084), .B(n5083), .ZN(U3118)
         );
  NAND2_X1 U6252 ( .A1(n6494), .A2(n6496), .ZN(n5088) );
  INV_X1 U6253 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5085) );
  OAI22_X1 U6254 ( .A1(n5099), .A2(n6500), .B1(n5085), .B2(n5097), .ZN(n5086)
         );
  AOI21_X1 U6255 ( .B1(n6492), .B2(n5101), .A(n5086), .ZN(n5087) );
  OAI211_X1 U6256 ( .C1(n5104), .C2(n5899), .A(n5088), .B(n5087), .ZN(U3123)
         );
  NAND2_X1 U6257 ( .A1(n6494), .A2(n6475), .ZN(n5092) );
  INV_X1 U6258 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5089) );
  OAI22_X1 U6259 ( .A1(n5099), .A2(n6478), .B1(n5089), .B2(n5097), .ZN(n5090)
         );
  AOI21_X1 U6260 ( .B1(n6473), .B2(n5101), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6261 ( .C1(n5104), .C2(n5885), .A(n5092), .B(n5091), .ZN(U3120)
         );
  NAND2_X1 U6262 ( .A1(n6494), .A2(n6469), .ZN(n5096) );
  INV_X1 U6263 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5093) );
  OAI22_X1 U6264 ( .A1(n5099), .A2(n6472), .B1(n5093), .B2(n5097), .ZN(n5094)
         );
  AOI21_X1 U6265 ( .B1(n6467), .B2(n5101), .A(n5094), .ZN(n5095) );
  OAI211_X1 U6266 ( .C1(n5104), .C2(n5881), .A(n5096), .B(n5095), .ZN(U3119)
         );
  NAND2_X1 U6267 ( .A1(n6494), .A2(n6481), .ZN(n5103) );
  INV_X1 U6268 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5098) );
  OAI22_X1 U6269 ( .A1(n5099), .A2(n6484), .B1(n5098), .B2(n5097), .ZN(n5100)
         );
  AOI21_X1 U6270 ( .B1(n6479), .B2(n5101), .A(n5100), .ZN(n5102) );
  OAI211_X1 U6271 ( .C1(n5104), .C2(n5889), .A(n5103), .B(n5102), .ZN(U3121)
         );
  INV_X1 U6272 ( .A(n5105), .ZN(n5106) );
  OAI21_X1 U6273 ( .B1(n5106), .B2(n6630), .A(n6636), .ZN(n5113) );
  NOR2_X1 U6274 ( .A1(n6362), .A2(n5112), .ZN(n5147) );
  INV_X1 U6275 ( .A(n5147), .ZN(n5107) );
  OAI21_X1 U6276 ( .B1(n5109), .B2(n5108), .A(n5107), .ZN(n5111) );
  INV_X1 U6277 ( .A(n5112), .ZN(n5110) );
  AOI22_X1 U6278 ( .A1(n5113), .A2(n5111), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5110), .ZN(n5154) );
  INV_X1 U6279 ( .A(n5111), .ZN(n5114) );
  AOI22_X1 U6280 ( .A1(n5114), .A2(n5113), .B1(n5112), .B2(n6630), .ZN(n5115)
         );
  NAND2_X1 U6281 ( .A1(n6448), .A2(n5115), .ZN(n5146) );
  AOI22_X1 U6282 ( .A1(n6443), .A2(n5147), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5146), .ZN(n5116) );
  OAI21_X1 U6283 ( .B1(n5117), .B2(n5149), .A(n5116), .ZN(n5118) );
  AOI21_X1 U6284 ( .B1(n6451), .B2(n5152), .A(n5118), .ZN(n5119) );
  OAI21_X1 U6285 ( .B1(n5154), .B2(n6454), .A(n5119), .ZN(U3028) );
  OAI21_X1 U6286 ( .B1(n3113), .B2(n3123), .A(n5120), .ZN(n5252) );
  AOI22_X1 U6287 ( .A1(n5561), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6163), .ZN(n5121) );
  OAI21_X1 U6288 ( .B1(n5252), .B2(n6169), .A(n5121), .ZN(U2882) );
  AOI22_X1 U6289 ( .A1(n6479), .A2(n5147), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5146), .ZN(n5122) );
  OAI21_X1 U6290 ( .B1(n5123), .B2(n5149), .A(n5122), .ZN(n5124) );
  AOI21_X1 U6291 ( .B1(n6480), .B2(n5152), .A(n5124), .ZN(n5125) );
  OAI21_X1 U6292 ( .B1(n5154), .B2(n6484), .A(n5125), .ZN(U3033) );
  AOI22_X1 U6293 ( .A1(n6467), .A2(n5147), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5146), .ZN(n5126) );
  OAI21_X1 U6294 ( .B1(n5127), .B2(n5149), .A(n5126), .ZN(n5128) );
  AOI21_X1 U6295 ( .B1(n6468), .B2(n5152), .A(n5128), .ZN(n5129) );
  OAI21_X1 U6296 ( .B1(n5154), .B2(n6472), .A(n5129), .ZN(U3031) );
  AOI22_X1 U6297 ( .A1(n6492), .A2(n5147), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5146), .ZN(n5130) );
  OAI21_X1 U6298 ( .B1(n5131), .B2(n5149), .A(n5130), .ZN(n5132) );
  AOI21_X1 U6299 ( .B1(n6493), .B2(n5152), .A(n5132), .ZN(n5133) );
  OAI21_X1 U6300 ( .B1(n5154), .B2(n6500), .A(n5133), .ZN(U3035) );
  AOI22_X1 U6301 ( .A1(n6485), .A2(n5147), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5146), .ZN(n5134) );
  OAI21_X1 U6302 ( .B1(n5135), .B2(n5149), .A(n5134), .ZN(n5136) );
  AOI21_X1 U6303 ( .B1(n6487), .B2(n5152), .A(n5136), .ZN(n5137) );
  OAI21_X1 U6304 ( .B1(n5154), .B2(n6490), .A(n5137), .ZN(U3034) );
  AOI22_X1 U6305 ( .A1(n6461), .A2(n5147), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5146), .ZN(n5138) );
  OAI21_X1 U6306 ( .B1(n5139), .B2(n5149), .A(n5138), .ZN(n5140) );
  AOI21_X1 U6307 ( .B1(n6462), .B2(n5152), .A(n5140), .ZN(n5141) );
  OAI21_X1 U6308 ( .B1(n5154), .B2(n6466), .A(n5141), .ZN(U3030) );
  AOI22_X1 U6309 ( .A1(n6473), .A2(n5147), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5146), .ZN(n5142) );
  OAI21_X1 U6310 ( .B1(n5143), .B2(n5149), .A(n5142), .ZN(n5144) );
  AOI21_X1 U6311 ( .B1(n6474), .B2(n5152), .A(n5144), .ZN(n5145) );
  OAI21_X1 U6312 ( .B1(n5154), .B2(n6478), .A(n5145), .ZN(U3032) );
  AOI22_X1 U6313 ( .A1(n6455), .A2(n5147), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5146), .ZN(n5148) );
  OAI21_X1 U6314 ( .B1(n5150), .B2(n5149), .A(n5148), .ZN(n5151) );
  AOI21_X1 U6315 ( .B1(n6456), .B2(n5152), .A(n5151), .ZN(n5153) );
  OAI21_X1 U6316 ( .B1(n5154), .B2(n6460), .A(n5153), .ZN(U3029) );
  INV_X1 U6317 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6580) );
  INV_X2 U6318 ( .A(n6140), .ZN(n5308) );
  INV_X1 U6319 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6879) );
  INV_X1 U6320 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6575) );
  INV_X1 U6321 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6577) );
  NOR3_X1 U6322 ( .A1(n6681), .A2(n6575), .A3(n6577), .ZN(n5205) );
  INV_X1 U6323 ( .A(n5205), .ZN(n6139) );
  NOR2_X1 U6324 ( .A1(n6879), .A2(n6139), .ZN(n5155) );
  NAND2_X1 U6325 ( .A1(n5308), .A2(n5155), .ZN(n6125) );
  OR2_X2 U6326 ( .A1(n6580), .A2(n6125), .ZN(n6111) );
  INV_X1 U6327 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6581) );
  NAND3_X1 U6328 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5155), .A3(n5204), .ZN(n5209) );
  NAND2_X1 U6329 ( .A1(n6086), .A2(n5209), .ZN(n6124) );
  OAI22_X1 U6330 ( .A1(n5156), .A2(n6132), .B1(n6143), .B2(n4773), .ZN(n5158)
         );
  NAND2_X1 U6331 ( .A1(n5204), .A2(n5157), .ZN(n6121) );
  AOI211_X1 U6332 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5158), 
        .B(n6135), .ZN(n5159) );
  OAI221_X1 U6333 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6111), .C1(n6581), .C2(
        n6124), .A(n5159), .ZN(n5163) );
  OAI22_X1 U6334 ( .A1(n5161), .A2(n5905), .B1(n5160), .B2(n6149), .ZN(n5162)
         );
  OR2_X1 U6335 ( .A1(n5163), .A2(n5162), .ZN(U2821) );
  XNOR2_X1 U6336 ( .A(n5164), .B(n5165), .ZN(n5181) );
  AND2_X1 U6337 ( .A1(n5167), .A2(n5166), .ZN(n5169) );
  AOI211_X1 U6338 ( .C1(n5831), .C2(n5170), .A(n5169), .B(n5168), .ZN(n6300)
         );
  NOR2_X1 U6339 ( .A1(n5171), .A2(n5170), .ZN(n5263) );
  NAND2_X1 U6340 ( .A1(n5263), .A2(n6299), .ZN(n6307) );
  AOI21_X1 U6341 ( .B1(n6300), .B2(n6307), .A(n5260), .ZN(n5175) );
  INV_X1 U6342 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6765) );
  NAND3_X1 U6343 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5263), .A3(n5260), 
        .ZN(n5173) );
  NAND2_X1 U6344 ( .A1(n6312), .A2(n5210), .ZN(n5172) );
  OAI211_X1 U6345 ( .C1(n6765), .C2(n5829), .A(n5173), .B(n5172), .ZN(n5174)
         );
  NOR2_X1 U6346 ( .A1(n5175), .A2(n5174), .ZN(n5176) );
  OAI21_X1 U6347 ( .B1(n5181), .B2(n5984), .A(n5176), .ZN(U3010) );
  AOI22_X1 U6348 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6276), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5177) );
  OAI21_X1 U6349 ( .B1(n6272), .B2(n5212), .A(n5177), .ZN(n5178) );
  AOI21_X1 U6350 ( .B1(n5179), .B2(n6260), .A(n5178), .ZN(n5180) );
  OAI21_X1 U6351 ( .B1(n6277), .B2(n5181), .A(n5180), .ZN(U2978) );
  INV_X1 U6352 ( .A(n5182), .ZN(n5183) );
  NAND2_X1 U6353 ( .A1(n5184), .A2(n5183), .ZN(n5186) );
  AOI21_X1 U6354 ( .B1(n5187), .B2(n5186), .A(n5185), .ZN(n6292) );
  INV_X1 U6355 ( .A(n6292), .ZN(n5188) );
  INV_X1 U6356 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5237) );
  OAI222_X1 U6357 ( .A1(n5188), .A2(n5532), .B1(n5237), .B2(n6156), .C1(n5528), 
        .C2(n5252), .ZN(U2850) );
  OAI22_X1 U6358 ( .A1(n4418), .A2(n6132), .B1(n5204), .B2(n6575), .ZN(n5191)
         );
  NOR2_X1 U6359 ( .A1(n6143), .A2(n5189), .ZN(n5190) );
  AOI211_X1 U6360 ( .C1(n6575), .C2(n5308), .A(n5191), .B(n5190), .ZN(n5192)
         );
  OAI21_X1 U6361 ( .B1(n4554), .B2(n5199), .A(n5192), .ZN(n5194) );
  NOR2_X1 U6362 ( .A1(n6149), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5193)
         );
  AOI211_X1 U6363 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5194), 
        .B(n5193), .ZN(n5195) );
  OAI21_X1 U6364 ( .B1(n5284), .B2(n5196), .A(n5195), .ZN(U2826) );
  AOI22_X1 U6365 ( .A1(n5197), .A2(n6119), .B1(EBX_REG_3__SCAN_IN), .B2(n6118), 
        .ZN(n5198) );
  OAI21_X1 U6366 ( .B1(n6635), .B2(n5199), .A(n5198), .ZN(n5202) );
  NOR2_X1 U6367 ( .A1(n6149), .A2(n5200), .ZN(n5201) );
  AOI211_X1 U6368 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5202), 
        .B(n5201), .ZN(n5207) );
  INV_X1 U6369 ( .A(n6086), .ZN(n5399) );
  AOI21_X1 U6370 ( .B1(n5204), .B2(REIP_REG_1__SCAN_IN), .A(n5399), .ZN(n5203)
         );
  NOR2_X1 U6371 ( .A1(n5203), .A2(n6577), .ZN(n5279) );
  OAI21_X1 U6372 ( .B1(n5205), .B2(n6140), .A(n5204), .ZN(n6136) );
  OAI21_X1 U6373 ( .B1(n5279), .B2(REIP_REG_3__SCAN_IN), .A(n6136), .ZN(n5206)
         );
  OAI211_X1 U6374 ( .C1(n5284), .C2(n5208), .A(n5207), .B(n5206), .ZN(U2824)
         );
  NAND2_X1 U6375 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6109) );
  OAI21_X1 U6376 ( .B1(n6111), .B2(n6109), .A(n6765), .ZN(n5216) );
  NAND3_X1 U6377 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U6378 ( .A1(n5226), .A2(n5209), .ZN(n5229) );
  AOI22_X1 U6379 ( .A1(n5210), .A2(n6119), .B1(EBX_REG_8__SCAN_IN), .B2(n6118), 
        .ZN(n5211) );
  NAND2_X1 U6380 ( .A1(n6121), .A2(n5211), .ZN(n5215) );
  OAI22_X1 U6381 ( .A1(n5213), .A2(n6133), .B1(n6149), .B2(n5212), .ZN(n5214)
         );
  AOI211_X1 U6382 ( .C1(n5216), .C2(n3147), .A(n5215), .B(n5214), .ZN(n5217)
         );
  OAI21_X1 U6383 ( .B1(n5218), .B2(n5905), .A(n5217), .ZN(U2819) );
  OAI21_X1 U6384 ( .B1(n5219), .B2(n5221), .A(n5220), .ZN(n5704) );
  AND2_X1 U6385 ( .A1(n5262), .A2(n5222), .ZN(n5223) );
  AOI22_X1 U6386 ( .A1(n3122), .A2(n6670), .B1(n6671), .B2(EBX_REG_11__SCAN_IN), .ZN(n5224) );
  OAI21_X1 U6387 ( .B1(n5704), .B2(n5528), .A(n5224), .ZN(U2848) );
  AOI22_X1 U6388 ( .A1(n5561), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6163), .ZN(n5225) );
  OAI21_X1 U6389 ( .B1(n5704), .B2(n6169), .A(n5225), .ZN(U2880) );
  AOI22_X1 U6390 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6097), .B1(n6119), 
        .B2(n3122), .ZN(n5228) );
  INV_X1 U6391 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6862) );
  NAND4_X1 U6392 ( .A1(n6102), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n6862), .ZN(n5227) );
  NAND3_X1 U6393 ( .A1(n5228), .A2(n6121), .A3(n5227), .ZN(n5234) );
  NAND4_X1 U6394 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n5229), .ZN(n6085) );
  INV_X1 U6395 ( .A(n6085), .ZN(n5230) );
  NOR3_X1 U6396 ( .A1(n5399), .A2(n6862), .A3(n5230), .ZN(n5233) );
  OAI22_X1 U6397 ( .A1(n6149), .A2(n5700), .B1(n5231), .B2(n6143), .ZN(n5232)
         );
  NOR3_X1 U6398 ( .A1(n5234), .A2(n5233), .A3(n5232), .ZN(n5235) );
  OAI21_X1 U6399 ( .B1(n5704), .B2(n5905), .A(n5235), .ZN(U2816) );
  INV_X1 U6400 ( .A(n6102), .ZN(n5236) );
  NOR2_X1 U6401 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5236), .ZN(n6101) );
  INV_X1 U6402 ( .A(n6101), .ZN(n5242) );
  OAI22_X1 U6403 ( .A1(n6149), .A2(n5248), .B1(n6143), .B2(n5237), .ZN(n5240)
         );
  AOI22_X1 U6404 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6097), .B1(n6119), 
        .B2(n6292), .ZN(n5238) );
  NAND2_X1 U6405 ( .A1(n5238), .A2(n6121), .ZN(n5239) );
  AOI211_X1 U6406 ( .C1(REIP_REG_9__SCAN_IN), .C2(n3147), .A(n5240), .B(n5239), 
        .ZN(n5241) );
  OAI211_X1 U6407 ( .C1(n5252), .C2(n5905), .A(n5242), .B(n5241), .ZN(U2818)
         );
  AND2_X1 U6408 ( .A1(n5120), .A2(n5243), .ZN(n5244) );
  NOR2_X1 U6409 ( .A1(n5219), .A2(n5244), .ZN(n6100) );
  INV_X1 U6410 ( .A(n6100), .ZN(n5269) );
  AOI22_X1 U6411 ( .A1(n5561), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6163), .ZN(n5245) );
  OAI21_X1 U6412 ( .B1(n5269), .B2(n6169), .A(n5245), .ZN(U2881) );
  XNOR2_X1 U6413 ( .A(n5689), .B(n6724), .ZN(n5247) );
  XNOR2_X1 U6414 ( .A(n5246), .B(n5247), .ZN(n6295) );
  NAND2_X1 U6415 ( .A1(n6295), .A2(n6262), .ZN(n5251) );
  AND2_X1 U6416 ( .A1(n6276), .A2(REIP_REG_9__SCAN_IN), .ZN(n6291) );
  NOR2_X1 U6417 ( .A1(n6272), .A2(n5248), .ZN(n5249) );
  AOI211_X1 U6418 ( .C1(n6280), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6291), 
        .B(n5249), .ZN(n5250) );
  OAI211_X1 U6419 ( .C1(n6283), .C2(n5252), .A(n5251), .B(n5250), .ZN(U2977)
         );
  NAND2_X1 U6420 ( .A1(n3116), .A2(n5254), .ZN(n5255) );
  XNOR2_X1 U6421 ( .A(n5253), .B(n5255), .ZN(n5268) );
  AOI22_X1 U6422 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6276), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5256) );
  OAI21_X1 U6423 ( .B1(n6272), .B2(n5257), .A(n5256), .ZN(n5258) );
  AOI21_X1 U6424 ( .B1(n6100), .B2(n6260), .A(n5258), .ZN(n5259) );
  OAI21_X1 U6425 ( .B1(n5268), .B2(n5695), .A(n5259), .ZN(U2976) );
  NOR2_X1 U6426 ( .A1(n5260), .A2(n6299), .ZN(n5261) );
  OAI21_X1 U6427 ( .B1(n5792), .B2(n5261), .A(n6300), .ZN(n6293) );
  OAI21_X1 U6428 ( .B1(n5185), .B2(n3153), .A(n5262), .ZN(n6095) );
  INV_X1 U6429 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6797) );
  OAI22_X1 U6430 ( .A1(n6018), .A2(n6095), .B1(n6797), .B2(n5829), .ZN(n5266)
         );
  NAND3_X1 U6431 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n5263), .ZN(n6298) );
  AOI221_X1 U6432 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n5264), .C2(n6724), .A(n6298), 
        .ZN(n5265) );
  AOI211_X1 U6433 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6293), .A(n5266), .B(n5265), .ZN(n5267) );
  OAI21_X1 U6434 ( .B1(n5984), .B2(n5268), .A(n5267), .ZN(U3008) );
  INV_X1 U6435 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6094) );
  OAI222_X1 U6436 ( .A1(n6095), .A2(n5532), .B1(n6156), .B2(n6094), .C1(n5528), 
        .C2(n5269), .ZN(U2849) );
  INV_X1 U6437 ( .A(n5271), .ZN(n5272) );
  AOI21_X1 U6438 ( .B1(n5273), .B2(n5220), .A(n5272), .ZN(n6154) );
  INV_X1 U6439 ( .A(n6154), .ZN(n5274) );
  INV_X1 U6440 ( .A(DATAI_12_), .ZN(n6783) );
  INV_X1 U6441 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6178) );
  OAI222_X1 U6442 ( .A1(n5274), .A2(n6169), .B1(n6167), .B2(n6783), .C1(n6168), 
        .C2(n6178), .ZN(U2879) );
  AOI22_X1 U6443 ( .A1(n5275), .A2(n6119), .B1(EBX_REG_2__SCAN_IN), .B2(n6118), 
        .ZN(n5278) );
  NAND2_X1 U6444 ( .A1(n5276), .A2(n6137), .ZN(n5277) );
  OAI211_X1 U6445 ( .C1(n6149), .C2(n6273), .A(n5278), .B(n5277), .ZN(n5282)
         );
  NAND2_X1 U6446 ( .A1(n5308), .A2(REIP_REG_1__SCAN_IN), .ZN(n5280) );
  AOI21_X1 U6447 ( .B1(n6577), .B2(n5280), .A(n5279), .ZN(n5281) );
  AOI211_X1 U6448 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5282), 
        .B(n5281), .ZN(n5283) );
  OAI21_X1 U6449 ( .B1(n5284), .B2(n6267), .A(n5283), .ZN(U2825) );
  AOI21_X1 U6450 ( .B1(n5285), .B2(n6545), .A(n6025), .ZN(n5291) );
  OR2_X1 U6451 ( .A1(n3911), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U6452 ( .A1(n5839), .A2(n6502), .ZN(n5287) );
  NAND2_X1 U6453 ( .A1(n5288), .A2(n5287), .ZN(n6505) );
  OAI22_X1 U6454 ( .A1(n6552), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6539), .ZN(n5289) );
  AOI21_X1 U6455 ( .B1(n6505), .B2(n6545), .A(n5289), .ZN(n5290) );
  OAI22_X1 U6456 ( .A1(n5291), .A2(n6502), .B1(n6025), .B2(n5290), .ZN(U3461)
         );
  NOR2_X1 U6457 ( .A1(n5301), .A2(n6283), .ZN(n5298) );
  OAI21_X1 U6458 ( .B1(n6266), .B2(n5294), .A(n5293), .ZN(n5295) );
  INV_X1 U6459 ( .A(n5295), .ZN(n5296) );
  OAI21_X1 U6460 ( .B1(n5300), .B2(n5695), .A(n5299), .ZN(U2956) );
  AOI22_X1 U6461 ( .A1(n5322), .A2(n6670), .B1(EBX_REG_30__SCAN_IN), .B2(n6671), .ZN(n5302) );
  OAI21_X1 U6462 ( .B1(n5301), .B2(n5535), .A(n5302), .ZN(U2829) );
  NAND3_X1 U6463 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5312) );
  INV_X1 U6464 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6875) );
  INV_X1 U6465 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6587) );
  NOR3_X1 U6466 ( .A1(n6875), .A2(n6587), .A3(n6085), .ZN(n6083) );
  NAND2_X1 U6467 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6083), .ZN(n5429) );
  NOR2_X1 U6468 ( .A1(n5312), .A2(n5429), .ZN(n5400) );
  NAND4_X1 U6469 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5400), .ZN(n5943) );
  INV_X1 U6470 ( .A(n5943), .ZN(n5304) );
  AND3_X1 U6471 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6472 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U6473 ( .A1(n6086), .A2(n5305), .ZN(n5929) );
  NAND2_X1 U6474 ( .A1(n5929), .A2(n6140), .ZN(n5340) );
  NAND2_X1 U6475 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n5317) );
  NAND3_X1 U6476 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5315) );
  INV_X1 U6477 ( .A(n5315), .ZN(n5307) );
  INV_X1 U6478 ( .A(n5340), .ZN(n5306) );
  AOI21_X1 U6479 ( .B1(n5929), .B2(n5307), .A(n5306), .ZN(n5919) );
  AOI21_X1 U6480 ( .B1(n5308), .B2(n5317), .A(n5919), .ZN(n5910) );
  NAND2_X1 U6481 ( .A1(n5910), .A2(REIP_REG_29__SCAN_IN), .ZN(n5341) );
  NAND3_X1 U6482 ( .A1(n5340), .A2(REIP_REG_30__SCAN_IN), .A3(n5341), .ZN(
        n5310) );
  AOI22_X1 U6483 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n6118), .ZN(n5309) );
  NAND2_X1 U6484 ( .A1(n5310), .A2(n5309), .ZN(n5321) );
  INV_X1 U6485 ( .A(n5311), .ZN(n5319) );
  INV_X1 U6486 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6600) );
  INV_X1 U6487 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6590) );
  NAND4_X1 U6488 ( .A1(n6102), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n6093) );
  NOR2_X2 U6489 ( .A1(n6093), .A2(n6587), .ZN(n6075) );
  INV_X1 U6490 ( .A(n5312), .ZN(n5313) );
  NAND3_X1 U6491 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6492 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5950), .ZN(n5942) );
  NAND2_X1 U6493 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5392), .ZN(n5930) );
  NOR2_X2 U6494 ( .A1(n5315), .A2(n5930), .ZN(n5920) );
  INV_X1 U6495 ( .A(n5920), .ZN(n5316) );
  INV_X1 U6496 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6614) );
  NAND3_X1 U6497 ( .A1(n5356), .A2(REIP_REG_29__SCAN_IN), .A3(n6614), .ZN(
        n5318) );
  OAI21_X1 U6498 ( .B1(n6149), .B2(n5319), .A(n5318), .ZN(n5320) );
  AOI211_X1 U6499 ( .C1(n5322), .C2(n6119), .A(n5321), .B(n5320), .ZN(n5323)
         );
  OAI21_X1 U6500 ( .B1(n5301), .B2(n5905), .A(n5323), .ZN(U2797) );
  AOI22_X1 U6501 ( .A1(n6160), .A2(DATAI_30_), .B1(n6163), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6502 ( .A1(n6164), .A2(DATAI_14_), .ZN(n5324) );
  OAI211_X1 U6503 ( .C1(n5301), .C2(n6169), .A(n5325), .B(n5324), .ZN(U2861)
         );
  NAND2_X1 U6504 ( .A1(n6168), .A2(n5327), .ZN(n5329) );
  AOI22_X1 U6505 ( .A1(n6160), .A2(DATAI_31_), .B1(n6163), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5328) );
  OAI21_X1 U6506 ( .B1(n5348), .B2(n5329), .A(n5328), .ZN(U2860) );
  MUX2_X1 U6507 ( .A(EBX_REG_29__SCAN_IN), .B(n5330), .S(n3837), .Z(n5333) );
  NOR2_X1 U6508 ( .A1(n5331), .A2(EBX_REG_29__SCAN_IN), .ZN(n5332) );
  OR2_X1 U6509 ( .A1(n5333), .A2(n5332), .ZN(n5352) );
  NOR2_X1 U6510 ( .A1(n5459), .A2(n5352), .ZN(n5354) );
  AOI21_X1 U6511 ( .B1(n5335), .B2(n5354), .A(n5334), .ZN(n5339) );
  OAI22_X1 U6512 ( .A1(n5337), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5336), .B2(EBX_REG_31__SCAN_IN), .ZN(n5338) );
  XNOR2_X1 U6513 ( .A(n5339), .B(n5338), .ZN(n5708) );
  OAI211_X1 U6514 ( .C1(n5341), .C2(n6614), .A(REIP_REG_31__SCAN_IN), .B(n5340), .ZN(n5345) );
  INV_X1 U6515 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5355) );
  NOR3_X1 U6516 ( .A1(n6614), .A2(n5355), .A3(REIP_REG_31__SCAN_IN), .ZN(n5342) );
  AOI22_X1 U6517 ( .A1(n5343), .A2(EBX_REG_31__SCAN_IN), .B1(n5356), .B2(n5342), .ZN(n5344) );
  OAI211_X1 U6518 ( .C1(n6754), .C2(n6133), .A(n5345), .B(n5344), .ZN(n5346)
         );
  AOI21_X1 U6519 ( .B1(n5708), .B2(n6119), .A(n5346), .ZN(n5347) );
  OAI21_X1 U6520 ( .B1(n5348), .B2(n5905), .A(n5347), .ZN(U2796) );
  AOI21_X1 U6521 ( .B1(n5351), .B2(n5455), .A(n5350), .ZN(n5570) );
  INV_X1 U6522 ( .A(n5570), .ZN(n5538) );
  AND2_X1 U6523 ( .A1(n5459), .A2(n5352), .ZN(n5353) );
  NOR2_X1 U6524 ( .A1(n5354), .A2(n5353), .ZN(n5721) );
  NOR2_X1 U6525 ( .A1(n5910), .A2(n5355), .ZN(n5360) );
  AOI22_X1 U6526 ( .A1(n6118), .A2(EBX_REG_29__SCAN_IN), .B1(n5356), .B2(n5355), .ZN(n5358) );
  NAND2_X1 U6527 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5357)
         );
  OAI211_X1 U6528 ( .C1(n6149), .C2(n5568), .A(n5358), .B(n5357), .ZN(n5359)
         );
  AOI211_X1 U6529 ( .C1(n5721), .C2(n6119), .A(n5360), .B(n5359), .ZN(n5361)
         );
  OAI21_X1 U6530 ( .B1(n5538), .B2(n5905), .A(n5361), .ZN(U2798) );
  INV_X1 U6531 ( .A(n5363), .ZN(n5364) );
  OAI21_X1 U6532 ( .B1(n5365), .B2(n5362), .A(n5364), .ZN(n5592) );
  NAND2_X1 U6533 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5366) );
  INV_X1 U6534 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6605) );
  OAI21_X1 U6535 ( .B1(n5930), .B2(n5366), .A(n6605), .ZN(n5373) );
  OR2_X1 U6536 ( .A1(n5472), .A2(n5368), .ZN(n5369) );
  NAND2_X1 U6537 ( .A1(n5463), .A2(n5369), .ZN(n5742) );
  OAI22_X1 U6538 ( .A1(n6133), .A2(n5591), .B1(n5469), .B2(n6143), .ZN(n5370)
         );
  AOI21_X1 U6539 ( .B1(n5595), .B2(n6099), .A(n5370), .ZN(n5371) );
  OAI21_X1 U6540 ( .B1(n5742), .B2(n6132), .A(n5371), .ZN(n5372) );
  AOI21_X1 U6541 ( .B1(n5373), .B2(n5919), .A(n5372), .ZN(n5374) );
  OAI21_X1 U6542 ( .B1(n5592), .B2(n5905), .A(n5374), .ZN(U2801) );
  AOI21_X1 U6543 ( .B1(n5376), .B2(n3114), .A(n3132), .ZN(n5607) );
  INV_X1 U6544 ( .A(n5607), .ZN(n5549) );
  XNOR2_X1 U6545 ( .A(n5476), .B(n5473), .ZN(n5762) );
  INV_X1 U6546 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6601) );
  NOR2_X1 U6547 ( .A1(n5929), .A2(n6601), .ZN(n5383) );
  OR2_X1 U6548 ( .A1(n5930), .A2(REIP_REG_24__SCAN_IN), .ZN(n5381) );
  OAI22_X1 U6549 ( .A1(n5378), .A2(n6133), .B1(n5605), .B2(n6149), .ZN(n5379)
         );
  INV_X1 U6550 ( .A(n5379), .ZN(n5380) );
  OAI211_X1 U6551 ( .C1(n6143), .C2(n5482), .A(n5381), .B(n5380), .ZN(n5382)
         );
  AOI211_X1 U6552 ( .C1(n5762), .C2(n6119), .A(n5383), .B(n5382), .ZN(n5384)
         );
  OAI21_X1 U6553 ( .B1(n5549), .B2(n5905), .A(n5384), .ZN(U2803) );
  NAND2_X1 U6554 ( .A1(n3097), .A2(n5386), .ZN(n5387) );
  NAND2_X1 U6555 ( .A1(n3114), .A2(n5387), .ZN(n5616) );
  INV_X1 U6556 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6683) );
  OAI22_X1 U6557 ( .A1(n6133), .A2(n5615), .B1(n6143), .B2(n6683), .ZN(n5390)
         );
  OAI21_X1 U6558 ( .B1(n5487), .B2(n5388), .A(n5476), .ZN(n5769) );
  NOR2_X1 U6559 ( .A1(n5769), .A2(n6132), .ZN(n5389) );
  AOI211_X1 U6560 ( .C1(n6099), .C2(n5619), .A(n5390), .B(n5389), .ZN(n5394)
         );
  INV_X1 U6561 ( .A(n5929), .ZN(n5391) );
  OAI21_X1 U6562 ( .B1(n5392), .B2(REIP_REG_23__SCAN_IN), .A(n5391), .ZN(n5393) );
  OAI211_X1 U6563 ( .C1(n5616), .C2(n5905), .A(n5394), .B(n5393), .ZN(U2804)
         );
  OR2_X1 U6564 ( .A1(n5396), .A2(n5397), .ZN(n5398) );
  AND2_X1 U6565 ( .A1(n5395), .A2(n5398), .ZN(n5646) );
  INV_X1 U6566 ( .A(n5401), .ZN(n6061) );
  INV_X1 U6567 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6594) );
  XNOR2_X1 U6568 ( .A(REIP_REG_19__SCAN_IN), .B(n6594), .ZN(n5402) );
  AOI22_X1 U6569 ( .A1(REIP_REG_19__SCAN_IN), .A2(n3156), .B1(n6061), .B2(
        n5402), .ZN(n5403) );
  INV_X1 U6570 ( .A(n5403), .ZN(n5410) );
  OAI21_X1 U6571 ( .B1(n6133), .B2(n5404), .A(n6121), .ZN(n5409) );
  XNOR2_X1 U6572 ( .A(n5505), .B(n3837), .ZN(n5516) );
  NAND2_X1 U6573 ( .A1(n5517), .A2(n5516), .ZN(n5519) );
  INV_X1 U6574 ( .A(n5405), .ZN(n5406) );
  XNOR2_X1 U6575 ( .A(n5519), .B(n5406), .ZN(n5805) );
  AOI22_X1 U6576 ( .A1(n6099), .A2(n5642), .B1(EBX_REG_19__SCAN_IN), .B2(n6118), .ZN(n5407) );
  OAI21_X1 U6577 ( .B1(n5805), .B2(n6132), .A(n5407), .ZN(n5408) );
  NOR3_X1 U6578 ( .A1(n5410), .A2(n5409), .A3(n5408), .ZN(n5411) );
  OAI21_X1 U6579 ( .B1(n5554), .B2(n5905), .A(n5411), .ZN(U2808) );
  AOI21_X1 U6580 ( .B1(n5415), .B2(n5412), .A(n5414), .ZN(n5658) );
  INV_X1 U6581 ( .A(n5658), .ZN(n5557) );
  INV_X1 U6582 ( .A(n6070), .ZN(n5416) );
  NAND2_X1 U6583 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6069) );
  INV_X1 U6584 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6867) );
  OAI21_X1 U6585 ( .B1(n5416), .B2(n6069), .A(n6867), .ZN(n5423) );
  NOR2_X1 U6586 ( .A1(n3154), .A2(n5417), .ZN(n5418) );
  OR2_X1 U6587 ( .A1(n5517), .A2(n5418), .ZN(n5992) );
  OAI22_X1 U6588 ( .A1(n5992), .A2(n6132), .B1(n5419), .B2(n6133), .ZN(n5422)
         );
  NAND2_X1 U6589 ( .A1(n6099), .A2(n5657), .ZN(n5420) );
  OAI211_X1 U6590 ( .C1(n6766), .C2(n6143), .A(n5420), .B(n6121), .ZN(n5421)
         );
  AOI211_X1 U6591 ( .C1(n5423), .C2(n3156), .A(n5422), .B(n5421), .ZN(n5424)
         );
  OAI21_X1 U6592 ( .B1(n5557), .B2(n5905), .A(n5424), .ZN(U2810) );
  OR2_X1 U6593 ( .A1(n5426), .A2(n5427), .ZN(n5428) );
  NAND2_X1 U6594 ( .A1(n5425), .A2(n5428), .ZN(n5673) );
  INV_X1 U6595 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U6596 ( .A1(n6086), .A2(n5429), .ZN(n6067) );
  OAI22_X1 U6597 ( .A1(n5669), .A2(n6149), .B1(n6133), .B2(n6856), .ZN(n5434)
         );
  INV_X1 U6598 ( .A(n5430), .ZN(n5524) );
  NAND2_X1 U6599 ( .A1(n5441), .A2(n5431), .ZN(n5432) );
  NAND2_X1 U6600 ( .A1(n5524), .A2(n5432), .ZN(n5998) );
  OAI22_X1 U6601 ( .A1(n5998), .A2(n6132), .B1(n5531), .B2(n6143), .ZN(n5433)
         );
  NOR3_X1 U6602 ( .A1(n5434), .A2(n6135), .A3(n5433), .ZN(n5435) );
  OAI21_X1 U6603 ( .B1(n6067), .B2(n6591), .A(n5435), .ZN(n5436) );
  AOI21_X1 U6604 ( .B1(n6070), .B2(n6591), .A(n5436), .ZN(n5437) );
  OAI21_X1 U6605 ( .B1(n5673), .B2(n5905), .A(n5437), .ZN(U2812) );
  INV_X1 U6606 ( .A(n5426), .ZN(n5439) );
  OAI21_X1 U6607 ( .B1(n5438), .B2(n5440), .A(n5439), .ZN(n6668) );
  OAI21_X1 U6608 ( .B1(n6010), .B2(n5442), .A(n5441), .ZN(n5816) );
  INV_X1 U6609 ( .A(n5816), .ZN(n6669) );
  AOI22_X1 U6610 ( .A1(n6669), .A2(n6119), .B1(EBX_REG_14__SCAN_IN), .B2(n6118), .ZN(n5443) );
  OAI211_X1 U6611 ( .C1(n6133), .C2(n5444), .A(n5443), .B(n6121), .ZN(n5447)
         );
  AOI21_X1 U6612 ( .B1(n6590), .B2(n5445), .A(n6067), .ZN(n5446) );
  AOI211_X1 U6613 ( .C1(n5678), .C2(n6099), .A(n5447), .B(n5446), .ZN(n5448)
         );
  OAI21_X1 U6614 ( .B1(n6668), .B2(n5905), .A(n5448), .ZN(U2813) );
  INV_X1 U6615 ( .A(n5708), .ZN(n5450) );
  INV_X1 U6616 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5449) );
  OAI22_X1 U6617 ( .A1(n5450), .A2(n5532), .B1(n5449), .B2(n6156), .ZN(U2828)
         );
  AOI22_X1 U6618 ( .A1(n5721), .A2(n6670), .B1(n6671), .B2(EBX_REG_29__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U6619 ( .B1(n5538), .B2(n5535), .A(n5451), .ZN(U2830) );
  NAND2_X1 U6620 ( .A1(n5452), .A2(n5453), .ZN(n5454) );
  NAND2_X1 U6621 ( .A1(n5465), .A2(n5457), .ZN(n5458) );
  NAND2_X1 U6622 ( .A1(n5459), .A2(n5458), .ZN(n5915) );
  OAI22_X1 U6623 ( .A1(n5915), .A2(n5532), .B1(n5906), .B2(n6156), .ZN(n5460)
         );
  INV_X1 U6624 ( .A(n5460), .ZN(n5461) );
  OAI21_X1 U6625 ( .B1(n5541), .B2(n5528), .A(n5461), .ZN(U2831) );
  INV_X1 U6626 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6627 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  NAND2_X1 U6628 ( .A1(n5465), .A2(n5464), .ZN(n5921) );
  OR2_X1 U6629 ( .A1(n5363), .A2(n5466), .ZN(n5467) );
  AND2_X1 U6630 ( .A1(n5452), .A2(n5467), .ZN(n5923) );
  OAI222_X1 U6631 ( .A1(n5468), .A2(n6156), .B1(n5532), .B2(n5921), .C1(n5544), 
        .C2(n5528), .ZN(U2832) );
  OAI22_X1 U6632 ( .A1(n5742), .A2(n5532), .B1(n5469), .B2(n6156), .ZN(n5470)
         );
  INV_X1 U6633 ( .A(n5470), .ZN(n5471) );
  OAI21_X1 U6634 ( .B1(n5592), .B2(n5528), .A(n5471), .ZN(U2833) );
  INV_X1 U6635 ( .A(n5472), .ZN(n5478) );
  INV_X1 U6636 ( .A(n5473), .ZN(n5475) );
  OAI21_X1 U6637 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5477) );
  NAND2_X1 U6638 ( .A1(n5478), .A2(n5477), .ZN(n5934) );
  INV_X1 U6639 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5481) );
  AOI21_X1 U6640 ( .B1(n5479), .B2(n5375), .A(n5362), .ZN(n5975) );
  INV_X1 U6641 ( .A(n5975), .ZN(n5480) );
  OAI222_X1 U6642 ( .A1(n5934), .A2(n5532), .B1(n5481), .B2(n6156), .C1(n5480), 
        .C2(n5528), .ZN(U2834) );
  NOR2_X1 U6643 ( .A1(n6156), .A2(n5482), .ZN(n5483) );
  AOI21_X1 U6644 ( .B1(n5762), .B2(n6670), .A(n5483), .ZN(n5484) );
  OAI21_X1 U6645 ( .B1(n5549), .B2(n5528), .A(n5484), .ZN(U2835) );
  OAI222_X1 U6646 ( .A1(n5535), .A2(n5616), .B1(n6156), .B2(n6683), .C1(n5769), 
        .C2(n5532), .ZN(U2836) );
  NOR2_X1 U6647 ( .A1(n5495), .A2(n5485), .ZN(n5486) );
  OR2_X1 U6648 ( .A1(n5487), .A2(n5486), .ZN(n5938) );
  OR2_X1 U6649 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  AND2_X1 U6650 ( .A1(n3097), .A2(n5490), .ZN(n5965) );
  INV_X1 U6651 ( .A(n5965), .ZN(n5491) );
  OAI222_X1 U6652 ( .A1(n5492), .A2(n6156), .B1(n5532), .B2(n5938), .C1(n5491), 
        .C2(n5528), .ZN(U2837) );
  XOR2_X1 U6653 ( .A(n5494), .B(n5493), .Z(n5968) );
  INV_X1 U6654 ( .A(n5535), .ZN(n6672) );
  INV_X1 U6655 ( .A(n5495), .ZN(n5499) );
  NAND2_X1 U6656 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  NAND2_X1 U6657 ( .A1(n5499), .A2(n5498), .ZN(n5953) );
  OAI22_X1 U6658 ( .A1(n5953), .A2(n5532), .B1(n5944), .B2(n6156), .ZN(n5500)
         );
  AOI21_X1 U6659 ( .B1(n5968), .B2(n6672), .A(n5500), .ZN(n5501) );
  INV_X1 U6660 ( .A(n5501), .ZN(U2838) );
  INV_X1 U6661 ( .A(n5493), .ZN(n5502) );
  AOI21_X1 U6662 ( .B1(n5503), .B2(n5395), .A(n5502), .ZN(n5971) );
  INV_X1 U6663 ( .A(n5971), .ZN(n5509) );
  MUX2_X1 U6664 ( .A(n5505), .B(n3313), .S(n5504), .Z(n5506) );
  XOR2_X1 U6665 ( .A(n5507), .B(n5506), .Z(n5957) );
  OAI222_X1 U6666 ( .A1(n5535), .A2(n5509), .B1(n5532), .B2(n5957), .C1(n5508), 
        .C2(n6156), .ZN(U2839) );
  OAI22_X1 U6667 ( .A1(n5805), .A2(n5532), .B1(n5510), .B2(n6156), .ZN(n5511)
         );
  AOI21_X1 U6668 ( .B1(n5646), .B2(n6672), .A(n5511), .ZN(n5512) );
  INV_X1 U6669 ( .A(n5512), .ZN(U2840) );
  INV_X1 U6670 ( .A(n5513), .ZN(n5515) );
  INV_X1 U6671 ( .A(n5414), .ZN(n5514) );
  AOI21_X1 U6672 ( .B1(n5515), .B2(n5514), .A(n5396), .ZN(n6157) );
  INV_X1 U6673 ( .A(n6157), .ZN(n5520) );
  INV_X1 U6674 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6869) );
  OR2_X1 U6675 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  NAND2_X1 U6676 ( .A1(n5519), .A2(n5518), .ZN(n6064) );
  OAI222_X1 U6677 ( .A1(n5520), .A2(n5528), .B1(n6156), .B2(n6869), .C1(n6064), 
        .C2(n5532), .ZN(U2841) );
  OAI22_X1 U6678 ( .A1(n5992), .A2(n5532), .B1(n6766), .B2(n6156), .ZN(n5521)
         );
  AOI21_X1 U6679 ( .B1(n5658), .B2(n6672), .A(n5521), .ZN(n5522) );
  INV_X1 U6680 ( .A(n5522), .ZN(U2842) );
  AND2_X1 U6681 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  OR2_X1 U6682 ( .A1(n5525), .A2(n3154), .ZN(n6066) );
  INV_X1 U6683 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U6684 ( .A1(n5425), .A2(n5526), .ZN(n5527) );
  AND2_X1 U6685 ( .A1(n5412), .A2(n5527), .ZN(n6162) );
  INV_X1 U6686 ( .A(n6162), .ZN(n5529) );
  OAI222_X1 U6687 ( .A1(n6066), .A2(n5532), .B1(n5530), .B2(n6156), .C1(n5529), 
        .C2(n5528), .ZN(U2843) );
  OAI22_X1 U6688 ( .A1(n5998), .A2(n5532), .B1(n5531), .B2(n6156), .ZN(n5533)
         );
  INV_X1 U6689 ( .A(n5533), .ZN(n5534) );
  OAI21_X1 U6690 ( .B1(n5673), .B2(n5535), .A(n5534), .ZN(U2844) );
  AOI22_X1 U6691 ( .A1(n6160), .A2(DATAI_29_), .B1(n6163), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U6692 ( .A1(n6164), .A2(DATAI_13_), .ZN(n5536) );
  OAI211_X1 U6693 ( .C1(n5538), .C2(n6169), .A(n5537), .B(n5536), .ZN(U2862)
         );
  AOI22_X1 U6694 ( .A1(n6164), .A2(DATAI_12_), .B1(n6163), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U6695 ( .A1(n6160), .A2(DATAI_28_), .ZN(n5539) );
  OAI211_X1 U6696 ( .C1(n5541), .C2(n6169), .A(n5540), .B(n5539), .ZN(U2863)
         );
  AOI22_X1 U6697 ( .A1(n6164), .A2(DATAI_11_), .B1(n6163), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U6698 ( .A1(n6160), .A2(DATAI_27_), .ZN(n5542) );
  OAI211_X1 U6699 ( .C1(n5544), .C2(n6169), .A(n5543), .B(n5542), .ZN(U2864)
         );
  AOI22_X1 U6700 ( .A1(n6160), .A2(DATAI_26_), .B1(n6163), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6701 ( .A1(n6164), .A2(DATAI_10_), .ZN(n5545) );
  OAI211_X1 U6702 ( .C1(n5592), .C2(n6169), .A(n5546), .B(n5545), .ZN(U2865)
         );
  AOI22_X1 U6703 ( .A1(n6160), .A2(DATAI_24_), .B1(n6163), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6704 ( .A1(n6164), .A2(DATAI_8_), .ZN(n5547) );
  OAI211_X1 U6705 ( .C1(n5549), .C2(n6169), .A(n5548), .B(n5547), .ZN(U2867)
         );
  AOI22_X1 U6706 ( .A1(n6160), .A2(DATAI_23_), .B1(n6163), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6707 ( .A1(n6164), .A2(DATAI_7_), .ZN(n5550) );
  OAI211_X1 U6708 ( .C1(n5616), .C2(n6169), .A(n5551), .B(n5550), .ZN(U2868)
         );
  AOI22_X1 U6709 ( .A1(n6160), .A2(DATAI_19_), .B1(n6163), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6710 ( .A1(n6164), .A2(DATAI_3_), .ZN(n5552) );
  OAI211_X1 U6711 ( .C1(n5554), .C2(n6169), .A(n5553), .B(n5552), .ZN(U2872)
         );
  AOI22_X1 U6712 ( .A1(n6160), .A2(DATAI_17_), .B1(n6163), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U6713 ( .A1(n6164), .A2(DATAI_1_), .ZN(n5555) );
  OAI211_X1 U6714 ( .C1(n5557), .C2(n6169), .A(n5556), .B(n5555), .ZN(U2874)
         );
  AOI22_X1 U6715 ( .A1(n5561), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6163), .ZN(n5558) );
  OAI21_X1 U6716 ( .B1(n5673), .B2(n6169), .A(n5558), .ZN(U2876) );
  INV_X1 U6717 ( .A(DATAI_14_), .ZN(n6778) );
  INV_X1 U6718 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5559) );
  OAI222_X1 U6719 ( .A1(n6668), .A2(n6169), .B1(n6167), .B2(n6778), .C1(n6168), 
        .C2(n5559), .ZN(U2877) );
  XOR2_X1 U6720 ( .A(n5560), .B(n5271), .Z(n6151) );
  INV_X1 U6721 ( .A(n6151), .ZN(n5563) );
  AOI22_X1 U6722 ( .A1(n5561), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6163), .ZN(n5562) );
  OAI21_X1 U6723 ( .B1(n5563), .B2(n6169), .A(n5562), .ZN(U2878) );
  INV_X1 U6724 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U6725 ( .A1(n5565), .A2(n5574), .ZN(n5566) );
  XNOR2_X1 U6726 ( .A(n5566), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5723)
         );
  NAND2_X1 U6727 ( .A1(n6276), .A2(REIP_REG_29__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6728 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5567)
         );
  OAI211_X1 U6729 ( .C1(n6272), .C2(n5568), .A(n5714), .B(n5567), .ZN(n5569)
         );
  AOI21_X1 U6730 ( .B1(n5570), .B2(n6260), .A(n5569), .ZN(n5571) );
  OAI21_X1 U6731 ( .B1(n5723), .B2(n6277), .A(n5571), .ZN(U2957) );
  NAND2_X1 U6732 ( .A1(n5580), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5573) );
  OAI21_X1 U6733 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5572), .A(n5573), 
        .ZN(n5576) );
  INV_X1 U6734 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6723) );
  NOR3_X1 U6735 ( .A1(n5580), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n6723), 
        .ZN(n5575) );
  AOI211_X1 U6736 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5576), .A(n3648), .B(n5575), .ZN(n5730) );
  NAND2_X1 U6737 ( .A1(n6276), .A2(REIP_REG_28__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U6738 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5577)
         );
  OAI211_X1 U6739 ( .C1(n6272), .C2(n5907), .A(n5727), .B(n5577), .ZN(n5578)
         );
  AOI21_X1 U6740 ( .B1(n5912), .B2(n6260), .A(n5578), .ZN(n5579) );
  OAI21_X1 U6741 ( .B1(n5730), .B2(n5695), .A(n5579), .ZN(U2958) );
  INV_X1 U6742 ( .A(n5572), .ZN(n5581) );
  NAND2_X1 U6743 ( .A1(n6276), .A2(REIP_REG_27__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U6744 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5583)
         );
  OAI211_X1 U6745 ( .C1(n6272), .C2(n5917), .A(n5733), .B(n5583), .ZN(n5584)
         );
  AOI21_X1 U6746 ( .B1(n5923), .B2(n6260), .A(n5584), .ZN(n5585) );
  OAI21_X1 U6747 ( .B1(n5737), .B2(n5695), .A(n5585), .ZN(U2959) );
  INV_X1 U6748 ( .A(n5586), .ZN(n5590) );
  NOR2_X1 U6749 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  XNOR2_X1 U6750 ( .A(n5590), .B(n5589), .ZN(n5745) );
  NAND2_X1 U6751 ( .A1(n6276), .A2(REIP_REG_26__SCAN_IN), .ZN(n5741) );
  OAI21_X1 U6752 ( .B1(n6266), .B2(n5591), .A(n5741), .ZN(n5594) );
  NOR2_X1 U6753 ( .A1(n5592), .A2(n6283), .ZN(n5593) );
  OAI21_X1 U6754 ( .B1(n5745), .B2(n6277), .A(n5596), .ZN(U2960) );
  NAND2_X1 U6755 ( .A1(n5689), .A2(n5597), .ZN(n5598) );
  XNOR2_X1 U6756 ( .A(n5652), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5635)
         );
  INV_X1 U6757 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5599) );
  XNOR2_X1 U6758 ( .A(n5689), .B(n5779), .ZN(n5630) );
  NOR2_X1 U6759 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5621)
         );
  NAND2_X1 U6760 ( .A1(n5628), .A2(n5621), .ZN(n5611) );
  OAI21_X1 U6761 ( .B1(n5652), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5600), 
        .ZN(n5623) );
  NAND3_X1 U6762 ( .A1(n5601), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5602) );
  OAI22_X2 U6763 ( .A1(n5611), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5623), .B2(n5602), .ZN(n5603) );
  XNOR2_X1 U6764 ( .A(n5603), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5764)
         );
  NOR2_X1 U6765 ( .A1(n5829), .A2(n6601), .ZN(n5761) );
  AOI21_X1 U6766 ( .B1(n6280), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5761), 
        .ZN(n5604) );
  OAI21_X1 U6767 ( .B1(n5605), .B2(n6272), .A(n5604), .ZN(n5606) );
  AOI21_X1 U6768 ( .B1(n5607), .B2(n6260), .A(n5606), .ZN(n5608) );
  OAI21_X1 U6769 ( .B1(n5764), .B2(n5695), .A(n5608), .ZN(U2962) );
  INV_X1 U6770 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U6771 ( .A1(n5689), .A2(n5610), .ZN(n5612) );
  OAI21_X1 U6772 ( .B1(n5613), .B2(n5612), .A(n5611), .ZN(n5614) );
  XNOR2_X1 U6773 ( .A(n5614), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5773)
         );
  NAND2_X1 U6774 ( .A1(n6276), .A2(REIP_REG_23__SCAN_IN), .ZN(n5768) );
  OAI21_X1 U6775 ( .B1(n6266), .B2(n5615), .A(n5768), .ZN(n5618) );
  NOR2_X1 U6776 ( .A1(n5616), .A2(n6283), .ZN(n5617) );
  AOI211_X1 U6777 ( .C1(n6258), .C2(n5619), .A(n5618), .B(n5617), .ZN(n5620)
         );
  OAI21_X1 U6778 ( .B1(n5773), .B2(n5695), .A(n5620), .ZN(U2963) );
  AOI21_X1 U6779 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5689), .A(n5621), 
        .ZN(n5622) );
  XNOR2_X1 U6780 ( .A(n5623), .B(n5622), .ZN(n5783) );
  INV_X1 U6781 ( .A(n5935), .ZN(n5625) );
  NOR2_X1 U6782 ( .A1(n5829), .A2(n6600), .ZN(n5776) );
  AOI21_X1 U6783 ( .B1(n6280), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5776), 
        .ZN(n5624) );
  OAI21_X1 U6784 ( .B1(n5625), .B2(n6272), .A(n5624), .ZN(n5626) );
  AOI21_X1 U6785 ( .B1(n5965), .B2(n6260), .A(n5626), .ZN(n5627) );
  OAI21_X1 U6786 ( .B1(n5783), .B2(n5695), .A(n5627), .ZN(U2964) );
  AOI21_X1 U6787 ( .B1(n5630), .B2(n5629), .A(n5628), .ZN(n5790) );
  INV_X1 U6788 ( .A(n5947), .ZN(n5632) );
  INV_X1 U6789 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U6790 ( .A1(n5829), .A2(n6707), .ZN(n5785) );
  AOI21_X1 U6791 ( .B1(n6280), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5785), 
        .ZN(n5631) );
  OAI21_X1 U6792 ( .B1(n5632), .B2(n6272), .A(n5631), .ZN(n5633) );
  AOI21_X1 U6793 ( .B1(n5968), .B2(n6260), .A(n5633), .ZN(n5634) );
  OAI21_X1 U6794 ( .B1(n5790), .B2(n5695), .A(n5634), .ZN(U2965) );
  XNOR2_X1 U6795 ( .A(n5636), .B(n5635), .ZN(n5801) );
  NAND2_X1 U6796 ( .A1(n6276), .A2(REIP_REG_20__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U6797 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5637)
         );
  OAI211_X1 U6798 ( .C1(n6272), .C2(n5955), .A(n5798), .B(n5637), .ZN(n5638)
         );
  AOI21_X1 U6799 ( .B1(n5971), .B2(n6260), .A(n5638), .ZN(n5639) );
  OAI21_X1 U6800 ( .B1(n5801), .B2(n5695), .A(n5639), .ZN(U2966) );
  XNOR2_X1 U6801 ( .A(n5689), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5641)
         );
  XNOR2_X1 U6802 ( .A(n5640), .B(n5641), .ZN(n5809) );
  INV_X1 U6803 ( .A(n5642), .ZN(n5644) );
  NAND2_X1 U6804 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5643)
         );
  NAND2_X1 U6805 ( .A1(n6276), .A2(REIP_REG_19__SCAN_IN), .ZN(n5804) );
  OAI211_X1 U6806 ( .C1(n6272), .C2(n5644), .A(n5643), .B(n5804), .ZN(n5645)
         );
  AOI21_X1 U6807 ( .B1(n5646), .B2(n6260), .A(n5645), .ZN(n5647) );
  OAI21_X1 U6808 ( .B1(n5809), .B2(n5695), .A(n5647), .ZN(U2967) );
  NOR3_X1 U6809 ( .A1(n5649), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5689), 
        .ZN(n5651) );
  OAI22_X1 U6810 ( .A1(n5651), .A2(n6811), .B1(n5652), .B2(n5650), .ZN(n5655)
         );
  NOR3_X1 U6811 ( .A1(n5650), .A2(n5652), .A3(n6811), .ZN(n5980) );
  INV_X1 U6812 ( .A(n5980), .ZN(n5654) );
  NOR4_X1 U6813 ( .A1(n5653), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A4(n5689), .ZN(n5979) );
  AOI21_X1 U6814 ( .B1(n5655), .B2(n5654), .A(n5979), .ZN(n5991) );
  OAI22_X1 U6815 ( .A1(n6266), .A2(n5419), .B1(n5829), .B2(n6867), .ZN(n5656)
         );
  AOI21_X1 U6816 ( .B1(n6258), .B2(n5657), .A(n5656), .ZN(n5660) );
  NAND2_X1 U6817 ( .A1(n5658), .A2(n6260), .ZN(n5659) );
  OAI211_X1 U6818 ( .C1(n5991), .C2(n6277), .A(n5660), .B(n5659), .ZN(U2969)
         );
  XNOR2_X1 U6819 ( .A(n5689), .B(n6850), .ZN(n5662) );
  XNOR2_X1 U6820 ( .A(n5661), .B(n5662), .ZN(n5814) );
  AOI22_X1 U6821 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6276), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5663) );
  OAI21_X1 U6822 ( .B1(n5664), .B2(n6272), .A(n5663), .ZN(n5665) );
  AOI21_X1 U6823 ( .B1(n6162), .B2(n6260), .A(n5665), .ZN(n5666) );
  OAI21_X1 U6824 ( .B1(n5814), .B2(n6277), .A(n5666), .ZN(U2970) );
  OAI21_X1 U6825 ( .B1(n5668), .B2(n5667), .A(n5653), .ZN(n6003) );
  NAND2_X1 U6826 ( .A1(n6003), .A2(n6262), .ZN(n5672) );
  AND2_X1 U6827 ( .A1(n6276), .A2(REIP_REG_15__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U6828 ( .A1(n6272), .A2(n5669), .ZN(n5670) );
  AOI211_X1 U6829 ( .C1(n6280), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5999), 
        .B(n5670), .ZN(n5671) );
  OAI211_X1 U6830 ( .C1(n6283), .C2(n5673), .A(n5672), .B(n5671), .ZN(U2971)
         );
  XNOR2_X1 U6831 ( .A(n5689), .B(n5822), .ZN(n5675) );
  XNOR2_X1 U6832 ( .A(n5674), .B(n5675), .ZN(n5828) );
  NAND2_X1 U6833 ( .A1(n6276), .A2(REIP_REG_14__SCAN_IN), .ZN(n5815) );
  OAI21_X1 U6834 ( .B1(n6266), .B2(n5444), .A(n5815), .ZN(n5677) );
  NOR2_X1 U6835 ( .A1(n6668), .A2(n6283), .ZN(n5676) );
  AOI211_X1 U6836 ( .C1(n6258), .C2(n5678), .A(n5677), .B(n5676), .ZN(n5679)
         );
  OAI21_X1 U6837 ( .B1(n6277), .B2(n5828), .A(n5679), .ZN(U2972) );
  NAND2_X1 U6838 ( .A1(n5681), .A2(n5682), .ZN(n5683) );
  NAND2_X1 U6839 ( .A1(n5680), .A2(n5683), .ZN(n6020) );
  INV_X1 U6840 ( .A(n6020), .ZN(n5687) );
  NAND2_X1 U6841 ( .A1(n6276), .A2(REIP_REG_13__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U6842 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5684)
         );
  OAI211_X1 U6843 ( .C1(n6272), .C2(n6078), .A(n6015), .B(n5684), .ZN(n5685)
         );
  AOI21_X1 U6844 ( .B1(n6151), .B2(n6260), .A(n5685), .ZN(n5686) );
  OAI21_X1 U6845 ( .B1(n5687), .B2(n5695), .A(n5686), .ZN(U2973) );
  XNOR2_X1 U6846 ( .A(n5689), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5690)
         );
  XNOR2_X1 U6847 ( .A(n5688), .B(n5690), .ZN(n5837) );
  AOI22_X1 U6848 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6276), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5691) );
  OAI21_X1 U6849 ( .B1(n6272), .B2(n5692), .A(n5691), .ZN(n5693) );
  AOI21_X1 U6850 ( .B1(n6154), .B2(n6260), .A(n5693), .ZN(n5694) );
  OAI21_X1 U6851 ( .B1(n5837), .B2(n5695), .A(n5694), .ZN(U2974) );
  NAND2_X1 U6852 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  XNOR2_X1 U6853 ( .A(n5696), .B(n5699), .ZN(n6287) );
  NAND2_X1 U6854 ( .A1(n6287), .A2(n6262), .ZN(n5703) );
  AND2_X1 U6855 ( .A1(n6276), .A2(REIP_REG_11__SCAN_IN), .ZN(n6285) );
  NOR2_X1 U6856 ( .A1(n6272), .A2(n5700), .ZN(n5701) );
  AOI211_X1 U6857 ( .C1(n6280), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6285), 
        .B(n5701), .ZN(n5702) );
  OAI211_X1 U6858 ( .C1(n6283), .C2(n5704), .A(n5703), .B(n5702), .ZN(U2975)
         );
  INV_X1 U6859 ( .A(n5705), .ZN(n5707) );
  NOR4_X1 U6860 ( .A1(n5715), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5709), 
        .A4(n3647), .ZN(n5706) );
  AOI211_X1 U6861 ( .C1(n5708), .C2(n6312), .A(n5707), .B(n5706), .ZN(n5712)
         );
  OAI211_X1 U6862 ( .C1(n5710), .C2(n5709), .A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(n5716), .ZN(n5711) );
  OAI211_X1 U6863 ( .C1(n5713), .C2(n5984), .A(n5712), .B(n5711), .ZN(U2987)
         );
  OAI21_X1 U6864 ( .B1(n5715), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5714), 
        .ZN(n5720) );
  INV_X1 U6865 ( .A(n5716), .ZN(n5717) );
  NOR3_X1 U6866 ( .A1(n5718), .A2(n5717), .A3(n3647), .ZN(n5719) );
  AOI211_X1 U6867 ( .C1(n6312), .C2(n5721), .A(n5720), .B(n5719), .ZN(n5722)
         );
  OAI21_X1 U6868 ( .B1(n5723), .B2(n5984), .A(n5722), .ZN(U2989) );
  XNOR2_X1 U6869 ( .A(n5724), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5725)
         );
  NAND2_X1 U6870 ( .A1(n5731), .A2(n5725), .ZN(n5726) );
  OAI211_X1 U6871 ( .C1(n5915), .C2(n6018), .A(n5727), .B(n5726), .ZN(n5728)
         );
  AOI21_X1 U6872 ( .B1(n5735), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5728), 
        .ZN(n5729) );
  OAI21_X1 U6873 ( .B1(n5730), .B2(n5984), .A(n5729), .ZN(U2990) );
  NAND2_X1 U6874 ( .A1(n5731), .A2(n6723), .ZN(n5732) );
  OAI211_X1 U6875 ( .C1(n5921), .C2(n6018), .A(n5733), .B(n5732), .ZN(n5734)
         );
  AOI21_X1 U6876 ( .B1(n5735), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5734), 
        .ZN(n5736) );
  OAI21_X1 U6877 ( .B1(n5737), .B2(n5984), .A(n5736), .ZN(U2991) );
  INV_X1 U6878 ( .A(n5759), .ZN(n5755) );
  INV_X1 U6879 ( .A(n5738), .ZN(n5752) );
  OAI211_X1 U6880 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5752), .B(n5739), .ZN(n5740) );
  OAI211_X1 U6881 ( .C1(n5742), .C2(n6018), .A(n5741), .B(n5740), .ZN(n5743)
         );
  AOI21_X1 U6882 ( .B1(n5755), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5743), 
        .ZN(n5744) );
  OAI21_X1 U6883 ( .B1(n5745), .B2(n5984), .A(n5744), .ZN(U2992) );
  INV_X1 U6884 ( .A(n5746), .ZN(n5747) );
  INV_X1 U6885 ( .A(n5748), .ZN(n5749) );
  OAI21_X1 U6886 ( .B1(n5750), .B2(n5747), .A(n5749), .ZN(n5974) );
  INV_X1 U6887 ( .A(n5974), .ZN(n5757) );
  AOI22_X1 U6888 ( .A1(n5752), .A2(n5751), .B1(REIP_REG_25__SCAN_IN), .B2(
        n6276), .ZN(n5753) );
  OAI21_X1 U6889 ( .B1(n5934), .B2(n6018), .A(n5753), .ZN(n5754) );
  AOI21_X1 U6890 ( .B1(n5755), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5754), 
        .ZN(n5756) );
  OAI21_X1 U6891 ( .B1(n5757), .B2(n5984), .A(n5756), .ZN(U2993) );
  AOI21_X1 U6892 ( .B1(n5766), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5758) );
  NOR2_X1 U6893 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  AOI211_X1 U6894 ( .C1(n6312), .C2(n5762), .A(n5761), .B(n5760), .ZN(n5763)
         );
  OAI21_X1 U6895 ( .B1(n5764), .B2(n5984), .A(n5763), .ZN(U2994) );
  NAND2_X1 U6896 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  OAI211_X1 U6897 ( .C1(n5769), .C2(n6018), .A(n5768), .B(n5767), .ZN(n5770)
         );
  AOI21_X1 U6898 ( .B1(n5771), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5770), 
        .ZN(n5772) );
  OAI21_X1 U6899 ( .B1(n5773), .B2(n5984), .A(n5772), .ZN(U2995) );
  INV_X1 U6900 ( .A(n5938), .ZN(n5777) );
  INV_X1 U6901 ( .A(n5795), .ZN(n5774) );
  NOR4_X1 U6902 ( .A1(n5793), .A2(n5774), .A3(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .A4(n5779), .ZN(n5775) );
  AOI211_X1 U6903 ( .C1(n5777), .C2(n6312), .A(n5776), .B(n5775), .ZN(n5782)
         );
  INV_X1 U6904 ( .A(n5778), .ZN(n5787) );
  NAND2_X1 U6905 ( .A1(n5795), .A2(n5779), .ZN(n5780) );
  NOR2_X1 U6906 ( .A1(n5793), .A2(n5780), .ZN(n5784) );
  OAI21_X1 U6907 ( .B1(n5787), .B2(n5784), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5781) );
  OAI211_X1 U6908 ( .C1(n5783), .C2(n5984), .A(n5782), .B(n5781), .ZN(U2996)
         );
  INV_X1 U6909 ( .A(n5953), .ZN(n5786) );
  AOI211_X1 U6910 ( .C1(n5786), .C2(n6312), .A(n5785), .B(n5784), .ZN(n5789)
         );
  NAND2_X1 U6911 ( .A1(n5787), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5788) );
  OAI211_X1 U6912 ( .C1(n5790), .C2(n5984), .A(n5789), .B(n5788), .ZN(U2997)
         );
  AOI21_X1 U6913 ( .B1(n6811), .B2(n5791), .A(n5990), .ZN(n5985) );
  OAI21_X1 U6914 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5792), .A(n5985), 
        .ZN(n5807) );
  INV_X1 U6915 ( .A(n5793), .ZN(n5802) );
  NOR2_X1 U6916 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U6917 ( .A1(n5802), .A2(n5796), .ZN(n5797) );
  OAI211_X1 U6918 ( .C1(n5957), .C2(n6018), .A(n5798), .B(n5797), .ZN(n5799)
         );
  AOI21_X1 U6919 ( .B1(n5807), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5799), 
        .ZN(n5800) );
  OAI21_X1 U6920 ( .B1(n5801), .B2(n5984), .A(n5800), .ZN(U2998) );
  NAND2_X1 U6921 ( .A1(n5802), .A2(n5597), .ZN(n5803) );
  OAI211_X1 U6922 ( .C1(n5805), .C2(n6018), .A(n5804), .B(n5803), .ZN(n5806)
         );
  AOI21_X1 U6923 ( .B1(n5807), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5806), 
        .ZN(n5808) );
  OAI21_X1 U6924 ( .B1(n5809), .B2(n5984), .A(n5808), .ZN(U2999) );
  NOR2_X1 U6925 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6898), .ZN(n6944)
         );
  INV_X1 U6926 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6592) );
  OAI22_X1 U6927 ( .A1(n6066), .A2(n6018), .B1(n6592), .B2(n5829), .ZN(n5811)
         );
  NAND2_X1 U6928 ( .A1(n5812), .A2(n6898), .ZN(n6004) );
  AOI21_X1 U6929 ( .B1(n6001), .B2(n6004), .A(n6850), .ZN(n5810) );
  AOI211_X1 U6930 ( .C1(n6944), .C2(n5812), .A(n5811), .B(n5810), .ZN(n5813)
         );
  OAI21_X1 U6931 ( .B1(n5814), .B2(n5984), .A(n5813), .ZN(U3002) );
  NOR2_X1 U6932 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6290), .ZN(n5826)
         );
  OAI21_X1 U6933 ( .B1(n6018), .B2(n5816), .A(n5815), .ZN(n5824) );
  NOR2_X1 U6934 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5820), .ZN(n6013)
         );
  OAI221_X1 U6935 ( .B1(n5818), .B2(n6012), .C1(n5818), .C2(n5817), .A(n6013), 
        .ZN(n6022) );
  OAI21_X1 U6936 ( .B1(n5825), .B2(n6318), .A(n6022), .ZN(n5819) );
  AOI211_X1 U6937 ( .C1(n5821), .C2(n5820), .A(n6286), .B(n5819), .ZN(n6024)
         );
  NOR2_X1 U6938 ( .A1(n6024), .A2(n5822), .ZN(n5823) );
  AOI211_X1 U6939 ( .C1(n5826), .C2(n5825), .A(n5824), .B(n5823), .ZN(n5827)
         );
  OAI21_X1 U6940 ( .B1(n5828), .B2(n5984), .A(n5827), .ZN(U3004) );
  XOR2_X1 U6941 ( .A(n6009), .B(n6008), .Z(n6153) );
  NOR2_X1 U6942 ( .A1(n5829), .A2(n6587), .ZN(n5835) );
  AOI221_X1 U6944 ( .B1(n5831), .B2(n6954), .C1(n5830), .C2(n6954), .A(n6286), 
        .ZN(n5832) );
  OAI33_X1 U6945 ( .A1(1'b0), .A2(n5832), .A3(n6752), .B1(
        INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6290), .B3(n6954), .ZN(n5834)
         );
  AOI211_X1 U6946 ( .C1(n6312), .C2(n6153), .A(n5835), .B(n5834), .ZN(n5836)
         );
  OAI21_X1 U6947 ( .B1(n5837), .B2(n5984), .A(n5836), .ZN(U3006) );
  NAND3_X1 U6948 ( .A1(n5839), .A2(n5838), .A3(n5847), .ZN(n5840) );
  OAI21_X1 U6949 ( .B1(n6503), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5840), 
        .ZN(n5841) );
  AOI21_X1 U6950 ( .B1(n5843), .B2(n5842), .A(n5841), .ZN(n6507) );
  INV_X1 U6951 ( .A(n6545), .ZN(n5852) );
  INV_X1 U6952 ( .A(n5844), .ZN(n5846) );
  AOI22_X1 U6953 ( .A1(n5848), .A2(n5847), .B1(n5846), .B2(n5845), .ZN(n5849)
         );
  OAI21_X1 U6954 ( .B1(n6507), .B2(n5852), .A(n5849), .ZN(n5850) );
  MUX2_X1 U6955 ( .A(n5850), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n6025), 
        .Z(U3460) );
  OAI22_X1 U6956 ( .A1(n5853), .A2(n5852), .B1(n6539), .B2(n5851), .ZN(n5855)
         );
  MUX2_X1 U6957 ( .A(n5855), .B(n5854), .S(n6025), .Z(U3456) );
  NAND2_X1 U6958 ( .A1(n4553), .A2(n6325), .ZN(n6355) );
  NAND2_X1 U6959 ( .A1(n5900), .A2(n6411), .ZN(n5857) );
  OAI21_X1 U6960 ( .B1(n5857), .B2(n5902), .A(n6636), .ZN(n5864) );
  AND2_X1 U6961 ( .A1(n5859), .A2(n5858), .ZN(n6437) );
  NAND2_X1 U6962 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5862), .ZN(n6441) );
  NOR2_X1 U6963 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6441), .ZN(n5897)
         );
  INV_X1 U6964 ( .A(n5897), .ZN(n5865) );
  INV_X1 U6965 ( .A(n6437), .ZN(n5863) );
  AOI22_X1 U6966 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5865), .B1(n5864), .B2(
        n5863), .ZN(n5866) );
  NAND3_X1 U6967 ( .A1(n5867), .A2(n5866), .A3(n6368), .ZN(n5896) );
  AOI22_X1 U6968 ( .A1(n6443), .A2(n5897), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5896), .ZN(n5868) );
  OAI21_X1 U6969 ( .B1(n5900), .B2(n5869), .A(n5868), .ZN(n5870) );
  AOI21_X1 U6970 ( .B1(n6444), .B2(n5902), .A(n5870), .ZN(n5871) );
  OAI21_X1 U6971 ( .B1(n5904), .B2(n6454), .A(n5871), .ZN(U3100) );
  AOI22_X1 U6972 ( .A1(n6455), .A2(n5897), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5896), .ZN(n5872) );
  OAI21_X1 U6973 ( .B1(n5900), .B2(n5873), .A(n5872), .ZN(n5874) );
  AOI21_X1 U6974 ( .B1(n5902), .B2(n6457), .A(n5874), .ZN(n5875) );
  OAI21_X1 U6975 ( .B1(n5904), .B2(n6460), .A(n5875), .ZN(U3101) );
  AOI22_X1 U6976 ( .A1(n6461), .A2(n5897), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5896), .ZN(n5876) );
  OAI21_X1 U6977 ( .B1(n5900), .B2(n5877), .A(n5876), .ZN(n5878) );
  AOI21_X1 U6978 ( .B1(n5902), .B2(n6463), .A(n5878), .ZN(n5879) );
  OAI21_X1 U6979 ( .B1(n5904), .B2(n6466), .A(n5879), .ZN(U3102) );
  AOI22_X1 U6980 ( .A1(n6467), .A2(n5897), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5896), .ZN(n5880) );
  OAI21_X1 U6981 ( .B1(n5900), .B2(n5881), .A(n5880), .ZN(n5882) );
  AOI21_X1 U6982 ( .B1(n5902), .B2(n6469), .A(n5882), .ZN(n5883) );
  OAI21_X1 U6983 ( .B1(n5904), .B2(n6472), .A(n5883), .ZN(U3103) );
  AOI22_X1 U6984 ( .A1(n6473), .A2(n5897), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5896), .ZN(n5884) );
  OAI21_X1 U6985 ( .B1(n5900), .B2(n5885), .A(n5884), .ZN(n5886) );
  AOI21_X1 U6986 ( .B1(n5902), .B2(n6475), .A(n5886), .ZN(n5887) );
  OAI21_X1 U6987 ( .B1(n5904), .B2(n6478), .A(n5887), .ZN(U3104) );
  AOI22_X1 U6988 ( .A1(n6479), .A2(n5897), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5896), .ZN(n5888) );
  OAI21_X1 U6989 ( .B1(n5900), .B2(n5889), .A(n5888), .ZN(n5890) );
  AOI21_X1 U6990 ( .B1(n5902), .B2(n6481), .A(n5890), .ZN(n5891) );
  OAI21_X1 U6991 ( .B1(n5904), .B2(n6484), .A(n5891), .ZN(U3105) );
  AOI22_X1 U6992 ( .A1(n6485), .A2(n5897), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5896), .ZN(n5892) );
  OAI21_X1 U6993 ( .B1(n5900), .B2(n5893), .A(n5892), .ZN(n5894) );
  AOI21_X1 U6994 ( .B1(n5902), .B2(n6486), .A(n5894), .ZN(n5895) );
  OAI21_X1 U6995 ( .B1(n5904), .B2(n6490), .A(n5895), .ZN(U3106) );
  AOI22_X1 U6996 ( .A1(n6492), .A2(n5897), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5896), .ZN(n5898) );
  OAI21_X1 U6997 ( .B1(n5900), .B2(n5899), .A(n5898), .ZN(n5901) );
  AOI21_X1 U6998 ( .B1(n5902), .B2(n6496), .A(n5901), .ZN(n5903) );
  OAI21_X1 U6999 ( .B1(n5904), .B2(n6500), .A(n5903), .ZN(U3107) );
  AND2_X1 U7000 ( .A1(n6189), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7001 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6612) );
  OAI22_X1 U7002 ( .A1(n6149), .A2(n5907), .B1(n5906), .B2(n6143), .ZN(n5908)
         );
  AOI21_X1 U7003 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6097), .A(n5908), 
        .ZN(n5909) );
  OAI21_X1 U7004 ( .B1(n5910), .B2(n6612), .A(n5909), .ZN(n5911) );
  AOI21_X1 U7005 ( .B1(n5912), .B2(n6114), .A(n5911), .ZN(n5914) );
  NAND3_X1 U7006 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5920), .A3(n6612), .ZN(
        n5913) );
  OAI211_X1 U7007 ( .C1(n6132), .C2(n5915), .A(n5914), .B(n5913), .ZN(U2799)
         );
  INV_X1 U7008 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6608) );
  AOI22_X1 U7009 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        EBX_REG_27__SCAN_IN), .B2(n6118), .ZN(n5916) );
  OAI21_X1 U7010 ( .B1(n5917), .B2(n6149), .A(n5916), .ZN(n5918) );
  AOI221_X1 U7011 ( .B1(n5920), .B2(n6608), .C1(n5919), .C2(
        REIP_REG_27__SCAN_IN), .A(n5918), .ZN(n5925) );
  NOR2_X1 U7012 ( .A1(n5921), .A2(n6132), .ZN(n5922) );
  AOI21_X1 U7013 ( .B1(n5923), .B2(n6114), .A(n5922), .ZN(n5924) );
  NAND2_X1 U7014 ( .A1(n5925), .A2(n5924), .ZN(U2800) );
  NOR3_X1 U7015 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6601), .A3(n5930), .ZN(n5926) );
  AOI21_X1 U7016 ( .B1(n6118), .B2(EBX_REG_25__SCAN_IN), .A(n5926), .ZN(n5927)
         );
  OAI21_X1 U7017 ( .B1(n6149), .B2(n5978), .A(n5927), .ZN(n5928) );
  AOI21_X1 U7018 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6097), .A(n5928), 
        .ZN(n5933) );
  OAI21_X1 U7019 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5930), .A(n5929), .ZN(n5931) );
  AOI22_X1 U7020 ( .A1(n5975), .A2(n6114), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5931), .ZN(n5932) );
  OAI211_X1 U7021 ( .C1(n5934), .C2(n6132), .A(n5933), .B(n5932), .ZN(U2802)
         );
  AOI22_X1 U7022 ( .A1(n5950), .A2(n6707), .B1(n6086), .B2(n5943), .ZN(n5941)
         );
  AOI22_X1 U7023 ( .A1(n6099), .A2(n5935), .B1(EBX_REG_22__SCAN_IN), .B2(n6118), .ZN(n5937) );
  NAND2_X1 U7024 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5936)
         );
  OAI211_X1 U7025 ( .C1(n5938), .C2(n6132), .A(n5937), .B(n5936), .ZN(n5939)
         );
  AOI21_X1 U7026 ( .B1(n5965), .B2(n6114), .A(n5939), .ZN(n5940) );
  OAI221_X1 U7027 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5942), .C1(n6600), .C2(
        n5941), .A(n5940), .ZN(U2805) );
  NAND2_X1 U7028 ( .A1(n6086), .A2(n5943), .ZN(n5961) );
  OAI22_X1 U7029 ( .A1(n6133), .A2(n5945), .B1(n5944), .B2(n6143), .ZN(n5946)
         );
  AOI21_X1 U7030 ( .B1(n6099), .B2(n5947), .A(n5946), .ZN(n5948) );
  OAI21_X1 U7031 ( .B1(n6707), .B2(n5961), .A(n5948), .ZN(n5949) );
  AOI21_X1 U7032 ( .B1(n5968), .B2(n6114), .A(n5949), .ZN(n5952) );
  NAND2_X1 U7033 ( .A1(n5950), .A2(n6707), .ZN(n5951) );
  OAI211_X1 U7034 ( .C1(n6132), .C2(n5953), .A(n5952), .B(n5951), .ZN(U2806)
         );
  INV_X1 U7035 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6596) );
  NOR2_X1 U7036 ( .A1(n6596), .A2(n6594), .ZN(n5954) );
  AOI21_X1 U7037 ( .B1(n6061), .B2(n5954), .A(REIP_REG_20__SCAN_IN), .ZN(n5962) );
  INV_X1 U7038 ( .A(n5955), .ZN(n5956) );
  AOI222_X1 U7039 ( .A1(n6118), .A2(EBX_REG_20__SCAN_IN), .B1(n5956), .B2(
        n6099), .C1(PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n6097), .ZN(n5960) );
  INV_X1 U7040 ( .A(n5957), .ZN(n5958) );
  AOI22_X1 U7041 ( .A1(n5971), .A2(n6114), .B1(n6119), .B2(n5958), .ZN(n5959)
         );
  OAI211_X1 U7042 ( .C1(n5962), .C2(n5961), .A(n5960), .B(n5959), .ZN(U2807)
         );
  AOI22_X1 U7043 ( .A1(n5975), .A2(n6161), .B1(n6160), .B2(DATAI_25_), .ZN(
        n5964) );
  AOI22_X1 U7044 ( .A1(n6164), .A2(DATAI_9_), .B1(n6163), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7045 ( .A1(n5964), .A2(n5963), .ZN(U2866) );
  AOI22_X1 U7046 ( .A1(n5965), .A2(n6161), .B1(n6160), .B2(DATAI_22_), .ZN(
        n5967) );
  AOI22_X1 U7047 ( .A1(n6164), .A2(DATAI_6_), .B1(n6163), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7048 ( .A1(n5967), .A2(n5966), .ZN(U2869) );
  AOI22_X1 U7049 ( .A1(n5968), .A2(n6161), .B1(n6160), .B2(DATAI_21_), .ZN(
        n5970) );
  AOI22_X1 U7050 ( .A1(n6164), .A2(DATAI_5_), .B1(n6163), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7051 ( .A1(n5970), .A2(n5969), .ZN(U2870) );
  AOI22_X1 U7052 ( .A1(n5971), .A2(n6161), .B1(n6160), .B2(DATAI_20_), .ZN(
        n5973) );
  AOI22_X1 U7053 ( .A1(n6164), .A2(DATAI_4_), .B1(n6163), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7054 ( .A1(n5973), .A2(n5972), .ZN(U2871) );
  AOI22_X1 U7055 ( .A1(n6276), .A2(REIP_REG_25__SCAN_IN), .B1(n6280), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5977) );
  AOI22_X1 U7056 ( .A1(n5975), .A2(n6260), .B1(n6262), .B2(n5974), .ZN(n5976)
         );
  OAI211_X1 U7057 ( .C1(n6272), .C2(n5978), .A(n5977), .B(n5976), .ZN(U2961)
         );
  AOI22_X1 U7058 ( .A1(n6276), .A2(REIP_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6280), .ZN(n5983) );
  NOR2_X1 U7059 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  XNOR2_X1 U7060 ( .A(n5981), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5987)
         );
  AOI22_X1 U7061 ( .A1(n5987), .A2(n6262), .B1(n6260), .B2(n6157), .ZN(n5982)
         );
  OAI211_X1 U7062 ( .C1(n6059), .C2(n6272), .A(n5983), .B(n5982), .ZN(U2968)
         );
  NAND2_X1 U7063 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6883), .ZN(n6951) );
  OAI22_X1 U7064 ( .A1(n5985), .A2(n6883), .B1(n6018), .B2(n6064), .ZN(n5986)
         );
  AOI21_X1 U7065 ( .B1(n5987), .B2(n6294), .A(n5986), .ZN(n5989) );
  NAND2_X1 U7066 ( .A1(n6276), .A2(REIP_REG_18__SCAN_IN), .ZN(n5988) );
  OAI211_X1 U7067 ( .C1(n5997), .C2(n6951), .A(n5989), .B(n5988), .ZN(U3000)
         );
  AOI22_X1 U7068 ( .A1(n6276), .A2(REIP_REG_17__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5990), .ZN(n5996) );
  INV_X1 U7069 ( .A(n5991), .ZN(n5994) );
  INV_X1 U7070 ( .A(n5992), .ZN(n5993) );
  AOI22_X1 U7071 ( .A1(n5994), .A2(n6294), .B1(n6312), .B2(n5993), .ZN(n5995)
         );
  OAI211_X1 U7072 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5997), .A(n5996), .B(n5995), .ZN(U3001) );
  INV_X1 U7073 ( .A(n5998), .ZN(n6000) );
  AOI21_X1 U7074 ( .B1(n6000), .B2(n6312), .A(n5999), .ZN(n6006) );
  INV_X1 U7075 ( .A(n6001), .ZN(n6002) );
  AOI22_X1 U7076 ( .A1(n6003), .A2(n6294), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6002), .ZN(n6005) );
  NAND3_X1 U7077 ( .A1(n6006), .A2(n6005), .A3(n6004), .ZN(U3003) );
  AOI21_X1 U7078 ( .B1(n6009), .B2(n6008), .A(n6007), .ZN(n6011) );
  NOR2_X1 U7079 ( .A1(n6011), .A2(n6010), .ZN(n6150) );
  INV_X1 U7080 ( .A(n6150), .ZN(n6017) );
  NAND3_X1 U7081 ( .A1(n6014), .A2(n6013), .A3(n6012), .ZN(n6016) );
  OAI211_X1 U7082 ( .C1(n6018), .C2(n6017), .A(n6016), .B(n6015), .ZN(n6019)
         );
  AOI21_X1 U7083 ( .B1(n6020), .B2(n6294), .A(n6019), .ZN(n6021) );
  OAI211_X1 U7084 ( .C1(n6024), .C2(n6023), .A(n6022), .B(n6021), .ZN(U3005)
         );
  INV_X1 U7085 ( .A(n6025), .ZN(n6030) );
  NAND3_X1 U7086 ( .A1(n6027), .A2(n6026), .A3(n6365), .ZN(n6028) );
  OAI21_X1 U7087 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(U3455) );
  INV_X1 U7088 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6031) );
  NOR2_X2 U7089 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6031), .ZN(n6667) );
  INV_X1 U7090 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6876) );
  OAI21_X1 U7091 ( .B1(n6667), .B2(n6876), .A(n3124), .ZN(U2789) );
  INV_X1 U7092 ( .A(n6521), .ZN(n6035) );
  INV_X1 U7093 ( .A(n6516), .ZN(n6032) );
  AOI21_X1 U7094 ( .B1(n6032), .B2(n6515), .A(n4399), .ZN(n6033) );
  AOI21_X1 U7095 ( .B1(n6035), .B2(n6034), .A(n6033), .ZN(n6044) );
  INV_X1 U7096 ( .A(n6044), .ZN(n6037) );
  OAI21_X1 U7097 ( .B1(n6037), .B2(n6036), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6038) );
  OAI21_X1 U7098 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6039), .A(n6038), .ZN(
        U2790) );
  NOR2_X1 U7099 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6041) );
  OAI21_X1 U7100 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6041), .A(n6651), .ZN(n6040)
         );
  OAI21_X1 U7101 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6651), .A(n6040), .ZN(
        U2791) );
  OAI21_X1 U7102 ( .B1(BS16_N), .B2(n6041), .A(n3125), .ZN(n6622) );
  OAI21_X1 U7103 ( .B1(n3125), .B2(n6657), .A(n6622), .ZN(U2792) );
  OAI21_X1 U7104 ( .B1(n6043), .B2(n6042), .A(n4438), .ZN(n6655) );
  NAND2_X1 U7105 ( .A1(n6044), .A2(n6655), .ZN(n6523) );
  NAND2_X1 U7106 ( .A1(n6544), .A2(n6523), .ZN(n6652) );
  INV_X1 U7107 ( .A(n6652), .ZN(n6654) );
  OAI21_X1 U7108 ( .B1(n6654), .B2(n6524), .A(n6277), .ZN(U2793) );
  NOR2_X1 U7109 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6943) );
  AOI211_X1 U7110 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_14__SCAN_IN), .B(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6045) );
  INV_X1 U7111 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6697) );
  INV_X1 U7112 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6693) );
  NAND4_X1 U7113 ( .A1(n6943), .A2(n6045), .A3(n6697), .A4(n6693), .ZN(n6053)
         );
  OR4_X1 U7114 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6052) );
  OR4_X1 U7115 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(
        n6051) );
  NOR4_X1 U7116 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6049) );
  NOR4_X1 U7117 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6048) );
  NOR4_X1 U7118 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6047) );
  NOR4_X1 U7119 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6046) );
  NAND4_X1 U7120 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(n6050)
         );
  INV_X1 U7121 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6055) );
  NOR3_X1 U7122 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6056) );
  OAI21_X1 U7123 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6056), .A(n6649), .ZN(n6054)
         );
  OAI21_X1 U7124 ( .B1(n6649), .B2(n6055), .A(n6054), .ZN(U2794) );
  INV_X1 U7125 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6623) );
  AOI21_X1 U7126 ( .B1(n6575), .B2(n6623), .A(n6056), .ZN(n6057) );
  INV_X1 U7127 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6619) );
  INV_X1 U7128 ( .A(n6649), .ZN(n6646) );
  AOI22_X1 U7129 ( .A1(n6649), .A2(n6057), .B1(n6619), .B2(n6646), .ZN(U2795)
         );
  AOI22_X1 U7130 ( .A1(n3156), .A2(REIP_REG_18__SCAN_IN), .B1(
        EBX_REG_18__SCAN_IN), .B2(n6118), .ZN(n6058) );
  OAI21_X1 U7131 ( .B1(n6059), .B2(n6149), .A(n6058), .ZN(n6060) );
  AOI211_X1 U7132 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6135), 
        .B(n6060), .ZN(n6063) );
  AOI22_X1 U7133 ( .A1(n6157), .A2(n6114), .B1(n6594), .B2(n6061), .ZN(n6062)
         );
  OAI211_X1 U7134 ( .C1(n6132), .C2(n6064), .A(n6063), .B(n6062), .ZN(U2809)
         );
  AOI22_X1 U7135 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        EBX_REG_16__SCAN_IN), .B2(n6118), .ZN(n6074) );
  AOI21_X1 U7136 ( .B1(n6099), .B2(n6065), .A(n6135), .ZN(n6073) );
  OAI22_X1 U7137 ( .A1(n6067), .A2(n6592), .B1(n6132), .B2(n6066), .ZN(n6068)
         );
  AOI21_X1 U7138 ( .B1(n6162), .B2(n6114), .A(n6068), .ZN(n6072) );
  OAI211_X1 U7139 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n6070), .B(n6069), .ZN(n6071) );
  NAND4_X1 U7140 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(U2811)
         );
  OAI21_X1 U7141 ( .B1(REIP_REG_13__SCAN_IN), .B2(n6075), .A(n6086), .ZN(n6082) );
  INV_X1 U7142 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6076) );
  OAI22_X1 U7143 ( .A1(n6133), .A2(n6076), .B1(n6965), .B2(n6143), .ZN(n6077)
         );
  AOI211_X1 U7144 ( .C1(n6150), .C2(n6119), .A(n6135), .B(n6077), .ZN(n6081)
         );
  INV_X1 U7145 ( .A(n6078), .ZN(n6079) );
  AOI22_X1 U7146 ( .A1(n6151), .A2(n6114), .B1(n6079), .B2(n6099), .ZN(n6080)
         );
  OAI211_X1 U7147 ( .C1(n6083), .C2(n6082), .A(n6081), .B(n6080), .ZN(U2814)
         );
  OAI21_X1 U7148 ( .B1(n6133), .B2(n6084), .A(n6121), .ZN(n6089) );
  NAND3_X1 U7149 ( .A1(n6086), .A2(n6085), .A3(REIP_REG_12__SCAN_IN), .ZN(
        n6087) );
  OAI21_X1 U7150 ( .B1(n6964), .B2(n6143), .A(n6087), .ZN(n6088) );
  AOI211_X1 U7151 ( .C1(n6119), .C2(n6153), .A(n6089), .B(n6088), .ZN(n6092)
         );
  AOI22_X1 U7152 ( .A1(n6154), .A2(n6114), .B1(n6099), .B2(n6090), .ZN(n6091)
         );
  OAI211_X1 U7153 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6093), .A(n6092), .B(n6091), .ZN(U2815) );
  OAI22_X1 U7154 ( .A1(n6095), .A2(n6132), .B1(n6143), .B2(n6094), .ZN(n6096)
         );
  AOI211_X1 U7155 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6135), 
        .B(n6096), .ZN(n6106) );
  AOI22_X1 U7156 ( .A1(n6100), .A2(n6114), .B1(n6099), .B2(n6098), .ZN(n6105)
         );
  OAI21_X1 U7157 ( .B1(n3147), .B2(n6101), .A(REIP_REG_10__SCAN_IN), .ZN(n6104) );
  NAND3_X1 U7158 ( .A1(n6102), .A2(REIP_REG_9__SCAN_IN), .A3(n6797), .ZN(n6103) );
  NAND4_X1 U7159 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(U2817)
         );
  INV_X1 U7160 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6108) );
  AOI22_X1 U7161 ( .A1(n6302), .A2(n6119), .B1(n6118), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n6107) );
  OAI211_X1 U7162 ( .C1(n6133), .C2(n6108), .A(n6107), .B(n6121), .ZN(n6113)
         );
  OAI21_X1 U7163 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n6109), .ZN(n6110) );
  INV_X1 U7164 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6583) );
  OAI22_X1 U7165 ( .A1(n6111), .A2(n6110), .B1(n6583), .B2(n6124), .ZN(n6112)
         );
  AOI211_X1 U7166 ( .C1(n6115), .C2(n6114), .A(n6113), .B(n6112), .ZN(n6116)
         );
  OAI21_X1 U7167 ( .B1(n6117), .B2(n6149), .A(n6116), .ZN(U2820) );
  INV_X1 U7168 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6123) );
  AOI22_X1 U7169 ( .A1(n6120), .A2(n6119), .B1(EBX_REG_5__SCAN_IN), .B2(n6118), 
        .ZN(n6122) );
  OAI211_X1 U7170 ( .C1(n6133), .C2(n6123), .A(n6122), .B(n6121), .ZN(n6127)
         );
  AOI21_X1 U7171 ( .B1(n6580), .B2(n6125), .A(n6124), .ZN(n6126) );
  AOI211_X1 U7172 ( .C1(n6128), .C2(n6146), .A(n6127), .B(n6126), .ZN(n6129)
         );
  OAI21_X1 U7173 ( .B1(n6130), .B2(n6149), .A(n6129), .ZN(U2822) );
  OAI22_X1 U7174 ( .A1(n3946), .A2(n6133), .B1(n6132), .B2(n6131), .ZN(n6134)
         );
  AOI211_X1 U7175 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6136), .A(n6135), .B(n6134), 
        .ZN(n6148) );
  NAND2_X1 U7176 ( .A1(n6138), .A2(n6137), .ZN(n6142) );
  OR3_X1 U7177 ( .A1(n6140), .A2(REIP_REG_4__SCAN_IN), .A3(n6139), .ZN(n6141)
         );
  OAI211_X1 U7178 ( .C1(n6144), .C2(n6143), .A(n6142), .B(n6141), .ZN(n6145)
         );
  AOI21_X1 U7179 ( .B1(n6261), .B2(n6146), .A(n6145), .ZN(n6147) );
  OAI211_X1 U7180 ( .C1(n6257), .C2(n6149), .A(n6148), .B(n6147), .ZN(U2823)
         );
  AOI22_X1 U7181 ( .A1(n6151), .A2(n6672), .B1(n6670), .B2(n6150), .ZN(n6152)
         );
  OAI21_X1 U7182 ( .B1(n6965), .B2(n6156), .A(n6152), .ZN(U2846) );
  AOI22_X1 U7183 ( .A1(n6154), .A2(n6672), .B1(n6670), .B2(n6153), .ZN(n6155)
         );
  OAI21_X1 U7184 ( .B1(n6964), .B2(n6156), .A(n6155), .ZN(U2847) );
  AOI22_X1 U7185 ( .A1(n6157), .A2(n6161), .B1(n6160), .B2(DATAI_18_), .ZN(
        n6159) );
  AOI22_X1 U7186 ( .A1(n6164), .A2(DATAI_2_), .B1(n6163), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7187 ( .A1(n6159), .A2(n6158), .ZN(U2873) );
  AOI22_X1 U7188 ( .A1(n6162), .A2(n6161), .B1(n6160), .B2(DATAI_16_), .ZN(
        n6166) );
  AOI22_X1 U7189 ( .A1(n6164), .A2(DATAI_0_), .B1(n6163), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7190 ( .A1(n6166), .A2(n6165), .ZN(U2875) );
  INV_X1 U7191 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6198) );
  OAI222_X1 U7192 ( .A1(n6284), .A2(n6169), .B1(n6168), .B2(n6198), .C1(n6167), 
        .C2(n6220), .ZN(U2891) );
  INV_X1 U7193 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6779) );
  INV_X1 U7194 ( .A(n6170), .ZN(n6172) );
  AOI22_X1 U7195 ( .A1(n6191), .A2(DATAO_REG_20__SCAN_IN), .B1(n6172), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6171) );
  OAI21_X1 U7196 ( .B1(n6779), .B2(n6664), .A(n6171), .ZN(U2903) );
  INV_X1 U7197 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6678) );
  AOI22_X1 U7198 ( .A1(n6172), .A2(EAX_REG_19__SCAN_IN), .B1(
        UWORD_REG_3__SCAN_IN), .B2(n6192), .ZN(n6173) );
  OAI21_X1 U7199 ( .B1(n6678), .B2(n6200), .A(n6173), .ZN(U2904) );
  INV_X1 U7200 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6255) );
  AOI22_X1 U7201 ( .A1(n6192), .A2(LWORD_REG_15__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U7202 ( .B1(n6255), .B2(n6199), .A(n6174), .ZN(U2908) );
  AOI222_X1 U7203 ( .A1(n6189), .A2(DATAO_REG_14__SCAN_IN), .B1(n6188), .B2(
        EAX_REG_14__SCAN_IN), .C1(n6192), .C2(LWORD_REG_14__SCAN_IN), .ZN(
        n6175) );
  INV_X1 U7204 ( .A(n6175), .ZN(U2909) );
  INV_X1 U7205 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6248) );
  AOI22_X1 U7206 ( .A1(n6192), .A2(LWORD_REG_13__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7207 ( .B1(n6248), .B2(n6199), .A(n6176), .ZN(U2910) );
  AOI22_X1 U7208 ( .A1(n6192), .A2(LWORD_REG_12__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6177) );
  OAI21_X1 U7209 ( .B1(n6178), .B2(n6199), .A(n6177), .ZN(U2911) );
  INV_X1 U7210 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6242) );
  AOI22_X1 U7211 ( .A1(n6192), .A2(LWORD_REG_11__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6179) );
  OAI21_X1 U7212 ( .B1(n6242), .B2(n6199), .A(n6179), .ZN(U2912) );
  INV_X1 U7213 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6239) );
  AOI22_X1 U7214 ( .A1(n6192), .A2(LWORD_REG_10__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U7215 ( .B1(n6239), .B2(n6199), .A(n6180), .ZN(U2913) );
  INV_X1 U7216 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6236) );
  AOI22_X1 U7217 ( .A1(n6192), .A2(LWORD_REG_9__SCAN_IN), .B1(n6189), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6181) );
  OAI21_X1 U7218 ( .B1(n6236), .B2(n6199), .A(n6181), .ZN(U2914) );
  AOI22_X1 U7219 ( .A1(n6192), .A2(LWORD_REG_8__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6182) );
  OAI21_X1 U7220 ( .B1(n6968), .B2(n6199), .A(n6182), .ZN(U2915) );
  AOI222_X1 U7221 ( .A1(n6189), .A2(DATAO_REG_7__SCAN_IN), .B1(n6188), .B2(
        EAX_REG_7__SCAN_IN), .C1(n6192), .C2(LWORD_REG_7__SCAN_IN), .ZN(n6183)
         );
  INV_X1 U7222 ( .A(n6183), .ZN(U2916) );
  AOI22_X1 U7223 ( .A1(n6184), .A2(LWORD_REG_6__SCAN_IN), .B1(n6191), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6185) );
  OAI21_X1 U7224 ( .B1(n6186), .B2(n6199), .A(n6185), .ZN(U2917) );
  INV_X1 U7225 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6755) );
  INV_X1 U7226 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6187) );
  OAI222_X1 U7227 ( .A1(n6200), .A2(n6755), .B1(n6199), .B2(n6852), .C1(n6664), 
        .C2(n6187), .ZN(U2918) );
  AOI222_X1 U7228 ( .A1(n6189), .A2(DATAO_REG_4__SCAN_IN), .B1(n6188), .B2(
        EAX_REG_4__SCAN_IN), .C1(n6192), .C2(LWORD_REG_4__SCAN_IN), .ZN(n6190)
         );
  INV_X1 U7229 ( .A(n6190), .ZN(U2919) );
  AOI22_X1 U7230 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6192), .B1(n6191), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6193) );
  OAI21_X1 U7231 ( .B1(n6194), .B2(n6199), .A(n6193), .ZN(U2920) );
  INV_X1 U7232 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6810) );
  INV_X1 U7233 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6195) );
  OAI222_X1 U7234 ( .A1(n6200), .A2(n6810), .B1(n6199), .B2(n6967), .C1(n6664), 
        .C2(n6195), .ZN(U2921) );
  INV_X1 U7235 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6731) );
  INV_X1 U7236 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6196) );
  OAI222_X1 U7237 ( .A1(n6200), .A2(n6731), .B1(n6199), .B2(n6825), .C1(n6664), 
        .C2(n6196), .ZN(U2922) );
  INV_X1 U7238 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6725) );
  INV_X1 U7239 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6197) );
  OAI222_X1 U7240 ( .A1(n6200), .A2(n6725), .B1(n6199), .B2(n6198), .C1(n6664), 
        .C2(n6197), .ZN(U2923) );
  AOI22_X1 U7241 ( .A1(n6246), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6249), .ZN(n6201) );
  OAI21_X1 U7242 ( .B1(n6251), .B2(n6220), .A(n6201), .ZN(U2924) );
  AOI22_X1 U7243 ( .A1(n6243), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6249), .ZN(n6203) );
  OAI21_X1 U7244 ( .B1(n6251), .B2(n6222), .A(n6203), .ZN(U2925) );
  AOI22_X1 U7245 ( .A1(n6243), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6249), .ZN(n6204) );
  OAI21_X1 U7246 ( .B1(n6251), .B2(n6878), .A(n6204), .ZN(U2926) );
  AOI22_X1 U7247 ( .A1(n6243), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6249), .ZN(n6205) );
  OAI21_X1 U7248 ( .B1(n6251), .B2(n6225), .A(n6205), .ZN(U2927) );
  AOI22_X1 U7249 ( .A1(n6243), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6249), .ZN(n6206) );
  OAI21_X1 U7250 ( .B1(n6251), .B2(n6839), .A(n6206), .ZN(U2928) );
  AOI22_X1 U7251 ( .A1(n6243), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6249), .ZN(n6207) );
  OAI21_X1 U7252 ( .B1(n6251), .B2(n6228), .A(n6207), .ZN(U2929) );
  AOI22_X1 U7253 ( .A1(n6243), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6249), .ZN(n6208) );
  OAI21_X1 U7254 ( .B1(n6251), .B2(n6230), .A(n6208), .ZN(U2930) );
  AOI22_X1 U7255 ( .A1(n6243), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6249), .ZN(n6209) );
  OAI21_X1 U7256 ( .B1(n6251), .B2(n6232), .A(n6209), .ZN(U2931) );
  AOI22_X1 U7257 ( .A1(n6243), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6249), .ZN(n6210) );
  OAI21_X1 U7258 ( .B1(n6251), .B2(n6832), .A(n6210), .ZN(U2932) );
  INV_X1 U7259 ( .A(DATAI_10_), .ZN(n6211) );
  NOR2_X1 U7260 ( .A1(n6251), .A2(n6211), .ZN(n6237) );
  AOI21_X1 U7261 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6243), .A(n6237), .ZN(
        n6212) );
  OAI21_X1 U7262 ( .B1(n6213), .B2(n6254), .A(n6212), .ZN(U2934) );
  AOI22_X1 U7263 ( .A1(n6243), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6249), .ZN(n6214) );
  OAI21_X1 U7264 ( .B1(n6251), .B2(n6783), .A(n6214), .ZN(U2936) );
  INV_X1 U7265 ( .A(DATAI_13_), .ZN(n6215) );
  NOR2_X1 U7266 ( .A1(n6251), .A2(n6215), .ZN(n6245) );
  AOI21_X1 U7267 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6243), .A(n6245), .ZN(
        n6216) );
  OAI21_X1 U7268 ( .B1(n6217), .B2(n6254), .A(n6216), .ZN(U2937) );
  AOI22_X1 U7269 ( .A1(n6243), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6249), .ZN(n6218) );
  OAI21_X1 U7270 ( .B1(n6251), .B2(n6778), .A(n6218), .ZN(U2938) );
  AOI22_X1 U7271 ( .A1(n6246), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6249), .ZN(n6219) );
  OAI21_X1 U7272 ( .B1(n6251), .B2(n6220), .A(n6219), .ZN(U2939) );
  AOI22_X1 U7273 ( .A1(n6246), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6249), .ZN(n6221) );
  OAI21_X1 U7274 ( .B1(n6251), .B2(n6222), .A(n6221), .ZN(U2940) );
  AOI22_X1 U7275 ( .A1(n6246), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6249), .ZN(n6223) );
  OAI21_X1 U7276 ( .B1(n6251), .B2(n6878), .A(n6223), .ZN(U2941) );
  AOI22_X1 U7277 ( .A1(n6246), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6249), .ZN(n6224) );
  OAI21_X1 U7278 ( .B1(n6251), .B2(n6225), .A(n6224), .ZN(U2942) );
  AOI22_X1 U7279 ( .A1(n6246), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6249), .ZN(n6226) );
  OAI21_X1 U7280 ( .B1(n6251), .B2(n6839), .A(n6226), .ZN(U2943) );
  AOI22_X1 U7281 ( .A1(n6246), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6249), .ZN(n6227) );
  OAI21_X1 U7282 ( .B1(n6251), .B2(n6228), .A(n6227), .ZN(U2944) );
  AOI22_X1 U7283 ( .A1(n6243), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6249), .ZN(n6229) );
  OAI21_X1 U7284 ( .B1(n6251), .B2(n6230), .A(n6229), .ZN(U2945) );
  AOI22_X1 U7285 ( .A1(n6243), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6249), .ZN(n6231) );
  OAI21_X1 U7286 ( .B1(n6251), .B2(n6232), .A(n6231), .ZN(U2946) );
  AOI22_X1 U7287 ( .A1(n6243), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6249), .ZN(n6233) );
  OAI21_X1 U7288 ( .B1(n6251), .B2(n6832), .A(n6233), .ZN(U2947) );
  AOI21_X1 U7289 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6246), .A(n6234), .ZN(n6235) );
  OAI21_X1 U7290 ( .B1(n6236), .B2(n6254), .A(n6235), .ZN(U2948) );
  AOI21_X1 U7291 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6243), .A(n6237), .ZN(
        n6238) );
  OAI21_X1 U7292 ( .B1(n6239), .B2(n6254), .A(n6238), .ZN(U2949) );
  AOI21_X1 U7293 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6246), .A(n6240), .ZN(
        n6241) );
  OAI21_X1 U7294 ( .B1(n6242), .B2(n6254), .A(n6241), .ZN(U2950) );
  AOI22_X1 U7295 ( .A1(n6243), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6249), .ZN(n6244) );
  OAI21_X1 U7296 ( .B1(n6251), .B2(n6783), .A(n6244), .ZN(U2951) );
  AOI21_X1 U7297 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6246), .A(n6245), .ZN(
        n6247) );
  OAI21_X1 U7298 ( .B1(n6248), .B2(n6254), .A(n6247), .ZN(U2952) );
  AOI22_X1 U7299 ( .A1(n6243), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6249), .ZN(n6250) );
  OAI21_X1 U7300 ( .B1(n6251), .B2(n6778), .A(n6250), .ZN(U2953) );
  INV_X1 U7301 ( .A(n6251), .ZN(n6252) );
  AOI22_X1 U7302 ( .A1(n6243), .A2(LWORD_REG_15__SCAN_IN), .B1(n6252), .B2(
        DATAI_15_), .ZN(n6253) );
  OAI21_X1 U7303 ( .B1(n6255), .B2(n6254), .A(n6253), .ZN(U2954) );
  INV_X1 U7304 ( .A(n6256), .ZN(n6263) );
  INV_X1 U7305 ( .A(n6257), .ZN(n6259) );
  AOI222_X1 U7306 ( .A1(n6263), .A2(n6262), .B1(n6261), .B2(n6260), .C1(n6259), 
        .C2(n6258), .ZN(n6265) );
  OAI211_X1 U7307 ( .C1(n6266), .C2(n3946), .A(n6265), .B(n6264), .ZN(U2982)
         );
  AOI22_X1 U7308 ( .A1(n6276), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6280), .ZN(n6271) );
  OAI22_X1 U7309 ( .A1(n6268), .A2(n6277), .B1(n6283), .B2(n6267), .ZN(n6269)
         );
  INV_X1 U7310 ( .A(n6269), .ZN(n6270) );
  OAI211_X1 U7311 ( .C1(n6273), .C2(n6272), .A(n6271), .B(n6270), .ZN(U2984)
         );
  OAI21_X1 U7312 ( .B1(n6275), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6274), 
        .ZN(n6315) );
  NAND2_X1 U7313 ( .A1(n6276), .A2(REIP_REG_0__SCAN_IN), .ZN(n6310) );
  OAI21_X1 U7314 ( .B1(n6277), .B2(n6315), .A(n6310), .ZN(n6278) );
  INV_X1 U7315 ( .A(n6278), .ZN(n6282) );
  OAI21_X1 U7316 ( .B1(n6280), .B2(n6279), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6281) );
  OAI211_X1 U7317 ( .C1(n6284), .C2(n6283), .A(n6282), .B(n6281), .ZN(U2986)
         );
  AOI21_X1 U7318 ( .B1(n6312), .B2(n3122), .A(n6285), .ZN(n6289) );
  AOI22_X1 U7319 ( .A1(n6287), .A2(n6294), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6286), .ZN(n6288) );
  OAI211_X1 U7320 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6290), .A(n6289), .B(n6288), .ZN(U3007) );
  AOI21_X1 U7321 ( .B1(n6312), .B2(n6292), .A(n6291), .ZN(n6297) );
  AOI22_X1 U7322 ( .A1(n6295), .A2(n6294), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6293), .ZN(n6296) );
  OAI211_X1 U7323 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6298), .A(n6297), 
        .B(n6296), .ZN(U3009) );
  OR2_X1 U7324 ( .A1(n6300), .A2(n6299), .ZN(n6304) );
  AOI21_X1 U7325 ( .B1(n6312), .B2(n6302), .A(n6301), .ZN(n6303) );
  OAI211_X1 U7326 ( .C1(n6305), .C2(n5984), .A(n6304), .B(n6303), .ZN(n6306)
         );
  INV_X1 U7327 ( .A(n6306), .ZN(n6308) );
  NAND2_X1 U7328 ( .A1(n6308), .A2(n6307), .ZN(U3011) );
  AND2_X1 U7329 ( .A1(n6310), .A2(n6309), .ZN(n6314) );
  NAND2_X1 U7330 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  OAI211_X1 U7331 ( .C1(n5984), .C2(n6315), .A(n6314), .B(n6313), .ZN(n6316)
         );
  INV_X1 U7332 ( .A(n6316), .ZN(n6317) );
  OAI221_X1 U7333 ( .B1(n6320), .B2(n6319), .C1(n6320), .C2(n6318), .A(n6317), 
        .ZN(U3018) );
  NOR2_X1 U7334 ( .A1(n6966), .A2(n6639), .ZN(U3019) );
  NOR2_X1 U7335 ( .A1(n3911), .A2(n6359), .ZN(n6321) );
  NOR2_X1 U7336 ( .A1(n6362), .A2(n6327), .ZN(n6348) );
  AOI21_X1 U7337 ( .B1(n6322), .B2(n6321), .A(n6348), .ZN(n6328) );
  INV_X1 U7338 ( .A(n6328), .ZN(n6323) );
  OAI21_X1 U7339 ( .B1(n6329), .B2(n6323), .A(n6448), .ZN(n6324) );
  INV_X1 U7340 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6961) );
  OR2_X1 U7341 ( .A1(n6326), .A2(n6325), .ZN(n6357) );
  AOI22_X1 U7342 ( .A1(n6399), .A2(n6451), .B1(n6443), .B2(n6348), .ZN(n6331)
         );
  OAI22_X1 U7343 ( .A1(n6329), .A2(n6328), .B1(n6327), .B2(n6656), .ZN(n6350)
         );
  AOI22_X1 U7344 ( .A1(n6350), .A2(n6371), .B1(n6444), .B2(n6349), .ZN(n6330)
         );
  OAI211_X1 U7345 ( .C1(n6354), .C2(n6961), .A(n6331), .B(n6330), .ZN(U3060)
         );
  INV_X1 U7346 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6836) );
  AOI22_X1 U7347 ( .A1(n6399), .A2(n6456), .B1(n6455), .B2(n6348), .ZN(n6333)
         );
  AOI22_X1 U7348 ( .A1(n6350), .A2(n6374), .B1(n6457), .B2(n6349), .ZN(n6332)
         );
  OAI211_X1 U7349 ( .C1(n6354), .C2(n6836), .A(n6333), .B(n6332), .ZN(U3061)
         );
  INV_X1 U7350 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6336) );
  AOI22_X1 U7351 ( .A1(n6399), .A2(n6462), .B1(n6461), .B2(n6348), .ZN(n6335)
         );
  AOI22_X1 U7352 ( .A1(n6350), .A2(n6377), .B1(n6463), .B2(n6349), .ZN(n6334)
         );
  OAI211_X1 U7353 ( .C1(n6354), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3062)
         );
  INV_X1 U7354 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6339) );
  AOI22_X1 U7355 ( .A1(n6399), .A2(n6468), .B1(n6467), .B2(n6348), .ZN(n6338)
         );
  AOI22_X1 U7356 ( .A1(n6350), .A2(n6381), .B1(n6469), .B2(n6349), .ZN(n6337)
         );
  OAI211_X1 U7357 ( .C1(n6354), .C2(n6339), .A(n6338), .B(n6337), .ZN(U3063)
         );
  INV_X1 U7358 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6700) );
  AOI22_X1 U7359 ( .A1(n6399), .A2(n6474), .B1(n6473), .B2(n6348), .ZN(n6341)
         );
  AOI22_X1 U7360 ( .A1(n6350), .A2(n6385), .B1(n6475), .B2(n6349), .ZN(n6340)
         );
  OAI211_X1 U7361 ( .C1(n6354), .C2(n6700), .A(n6341), .B(n6340), .ZN(U3064)
         );
  INV_X1 U7362 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6344) );
  AOI22_X1 U7363 ( .A1(n6399), .A2(n6480), .B1(n6479), .B2(n6348), .ZN(n6343)
         );
  AOI22_X1 U7364 ( .A1(n6350), .A2(n6388), .B1(n6481), .B2(n6349), .ZN(n6342)
         );
  OAI211_X1 U7365 ( .C1(n6354), .C2(n6344), .A(n6343), .B(n6342), .ZN(U3065)
         );
  INV_X1 U7366 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6347) );
  AOI22_X1 U7367 ( .A1(n6399), .A2(n6487), .B1(n6485), .B2(n6348), .ZN(n6346)
         );
  AOI22_X1 U7368 ( .A1(n6350), .A2(n6392), .B1(n6486), .B2(n6349), .ZN(n6345)
         );
  OAI211_X1 U7369 ( .C1(n6354), .C2(n6347), .A(n6346), .B(n6345), .ZN(U3066)
         );
  INV_X1 U7370 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6353) );
  AOI22_X1 U7371 ( .A1(n6399), .A2(n6493), .B1(n6492), .B2(n6348), .ZN(n6352)
         );
  AOI22_X1 U7372 ( .A1(n6350), .A2(n6397), .B1(n6496), .B2(n6349), .ZN(n6351)
         );
  OAI211_X1 U7373 ( .C1(n6354), .C2(n6353), .A(n6352), .B(n6351), .ZN(U3067)
         );
  INV_X1 U7374 ( .A(n6355), .ZN(n6356) );
  INV_X1 U7375 ( .A(n6427), .ZN(n6358) );
  AOI21_X1 U7376 ( .B1(n6358), .B2(n6357), .A(n6657), .ZN(n6361) );
  NOR2_X1 U7377 ( .A1(n6360), .A2(n6359), .ZN(n6405) );
  NOR3_X1 U7378 ( .A1(n6361), .A2(n6405), .A3(n6630), .ZN(n6367) );
  AND2_X1 U7379 ( .A1(n6362), .A2(n6412), .ZN(n6398) );
  OAI211_X1 U7380 ( .C1(n6398), .C2(n6365), .A(n6364), .B(n6363), .ZN(n6366)
         );
  INV_X1 U7381 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6959) );
  INV_X1 U7382 ( .A(n6405), .ZN(n6370) );
  OAI22_X1 U7383 ( .A1(n6370), .A2(n6630), .B1(n6369), .B2(n6368), .ZN(n6396)
         );
  AOI22_X1 U7384 ( .A1(n6371), .A2(n6396), .B1(n6443), .B2(n6398), .ZN(n6373)
         );
  AOI22_X1 U7385 ( .A1(n6399), .A2(n6444), .B1(n6451), .B2(n6427), .ZN(n6372)
         );
  OAI211_X1 U7386 ( .C1(n6403), .C2(n6959), .A(n6373), .B(n6372), .ZN(U3068)
         );
  INV_X1 U7387 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6781) );
  AOI22_X1 U7388 ( .A1(n6455), .A2(n6398), .B1(n6374), .B2(n6396), .ZN(n6376)
         );
  AOI22_X1 U7389 ( .A1(n6399), .A2(n6457), .B1(n6456), .B2(n6427), .ZN(n6375)
         );
  OAI211_X1 U7390 ( .C1(n6403), .C2(n6781), .A(n6376), .B(n6375), .ZN(U3069)
         );
  INV_X1 U7391 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6380) );
  AOI22_X1 U7392 ( .A1(n6461), .A2(n6398), .B1(n6377), .B2(n6396), .ZN(n6379)
         );
  AOI22_X1 U7393 ( .A1(n6399), .A2(n6463), .B1(n6462), .B2(n6427), .ZN(n6378)
         );
  OAI211_X1 U7394 ( .C1(n6403), .C2(n6380), .A(n6379), .B(n6378), .ZN(U3070)
         );
  INV_X1 U7395 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6384) );
  AOI22_X1 U7396 ( .A1(n6467), .A2(n6398), .B1(n6381), .B2(n6396), .ZN(n6383)
         );
  AOI22_X1 U7397 ( .A1(n6399), .A2(n6469), .B1(n6468), .B2(n6427), .ZN(n6382)
         );
  OAI211_X1 U7398 ( .C1(n6403), .C2(n6384), .A(n6383), .B(n6382), .ZN(U3071)
         );
  INV_X1 U7399 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U7400 ( .A1(n6473), .A2(n6398), .B1(n6385), .B2(n6396), .ZN(n6387)
         );
  AOI22_X1 U7401 ( .A1(n6399), .A2(n6475), .B1(n6474), .B2(n6427), .ZN(n6386)
         );
  OAI211_X1 U7402 ( .C1(n6403), .C2(n6930), .A(n6387), .B(n6386), .ZN(U3072)
         );
  INV_X1 U7403 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6391) );
  AOI22_X1 U7404 ( .A1(n6479), .A2(n6398), .B1(n6388), .B2(n6396), .ZN(n6390)
         );
  AOI22_X1 U7405 ( .A1(n6399), .A2(n6481), .B1(n6480), .B2(n6427), .ZN(n6389)
         );
  OAI211_X1 U7406 ( .C1(n6403), .C2(n6391), .A(n6390), .B(n6389), .ZN(U3073)
         );
  INV_X1 U7407 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6395) );
  AOI22_X1 U7408 ( .A1(n6485), .A2(n6398), .B1(n6392), .B2(n6396), .ZN(n6394)
         );
  AOI22_X1 U7409 ( .A1(n6399), .A2(n6486), .B1(n6487), .B2(n6427), .ZN(n6393)
         );
  OAI211_X1 U7410 ( .C1(n6403), .C2(n6395), .A(n6394), .B(n6393), .ZN(U3074)
         );
  INV_X1 U7411 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6402) );
  AOI22_X1 U7412 ( .A1(n6492), .A2(n6398), .B1(n6397), .B2(n6396), .ZN(n6401)
         );
  AOI22_X1 U7413 ( .A1(n6399), .A2(n6496), .B1(n6493), .B2(n6427), .ZN(n6400)
         );
  OAI211_X1 U7414 ( .C1(n6403), .C2(n6402), .A(n6401), .B(n6400), .ZN(U3075)
         );
  INV_X1 U7415 ( .A(n6404), .ZN(n6428) );
  AOI21_X1 U7416 ( .B1(n6405), .B2(n6436), .A(n6428), .ZN(n6409) );
  NOR2_X1 U7417 ( .A1(n6409), .A2(n6630), .ZN(n6406) );
  AOI21_X1 U7418 ( .B1(n6412), .B2(STATE2_REG_2__SCAN_IN), .A(n6406), .ZN(
        n6433) );
  AOI22_X1 U7419 ( .A1(n6428), .A2(n6443), .B1(n6427), .B2(n6444), .ZN(n6414)
         );
  INV_X1 U7420 ( .A(n6407), .ZN(n6434) );
  NAND2_X1 U7421 ( .A1(n6408), .A2(n6434), .ZN(n6631) );
  NAND3_X1 U7422 ( .A1(n6631), .A2(n6411), .A3(n6409), .ZN(n6410) );
  OAI211_X1 U7423 ( .C1(n6412), .C2(n6411), .A(n6410), .B(n6448), .ZN(n6430)
         );
  AOI22_X1 U7424 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6430), .B1(n6451), 
        .B2(n6429), .ZN(n6413) );
  OAI211_X1 U7425 ( .C1(n6433), .C2(n6454), .A(n6414), .B(n6413), .ZN(U3076)
         );
  AOI22_X1 U7426 ( .A1(n6428), .A2(n6455), .B1(n6427), .B2(n6457), .ZN(n6416)
         );
  AOI22_X1 U7427 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6430), .B1(n6456), 
        .B2(n6429), .ZN(n6415) );
  OAI211_X1 U7428 ( .C1(n6433), .C2(n6460), .A(n6416), .B(n6415), .ZN(U3077)
         );
  AOI22_X1 U7429 ( .A1(n6428), .A2(n6461), .B1(n6429), .B2(n6462), .ZN(n6418)
         );
  AOI22_X1 U7430 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6430), .B1(n6463), 
        .B2(n6427), .ZN(n6417) );
  OAI211_X1 U7431 ( .C1(n6433), .C2(n6466), .A(n6418), .B(n6417), .ZN(U3078)
         );
  AOI22_X1 U7432 ( .A1(n6428), .A2(n6467), .B1(n6429), .B2(n6468), .ZN(n6420)
         );
  AOI22_X1 U7433 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6430), .B1(n6469), 
        .B2(n6427), .ZN(n6419) );
  OAI211_X1 U7434 ( .C1(n6433), .C2(n6472), .A(n6420), .B(n6419), .ZN(U3079)
         );
  AOI22_X1 U7435 ( .A1(n6428), .A2(n6473), .B1(n6429), .B2(n6474), .ZN(n6422)
         );
  AOI22_X1 U7436 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6430), .B1(n6475), 
        .B2(n6427), .ZN(n6421) );
  OAI211_X1 U7437 ( .C1(n6433), .C2(n6478), .A(n6422), .B(n6421), .ZN(U3080)
         );
  AOI22_X1 U7438 ( .A1(n6428), .A2(n6479), .B1(n6427), .B2(n6481), .ZN(n6424)
         );
  AOI22_X1 U7439 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6430), .B1(n6480), 
        .B2(n6429), .ZN(n6423) );
  OAI211_X1 U7440 ( .C1(n6433), .C2(n6484), .A(n6424), .B(n6423), .ZN(U3081)
         );
  AOI22_X1 U7441 ( .A1(n6428), .A2(n6485), .B1(n6429), .B2(n6487), .ZN(n6426)
         );
  AOI22_X1 U7442 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6430), .B1(n6486), 
        .B2(n6427), .ZN(n6425) );
  OAI211_X1 U7443 ( .C1(n6433), .C2(n6490), .A(n6426), .B(n6425), .ZN(U3082)
         );
  AOI22_X1 U7444 ( .A1(n6428), .A2(n6492), .B1(n6427), .B2(n6496), .ZN(n6432)
         );
  AOI22_X1 U7445 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6430), .B1(n6493), 
        .B2(n6429), .ZN(n6431) );
  OAI211_X1 U7446 ( .C1(n6433), .C2(n6500), .A(n6432), .B(n6431), .ZN(U3083)
         );
  AOI21_X1 U7447 ( .B1(n6435), .B2(n6434), .A(n6630), .ZN(n6447) );
  NAND2_X1 U7448 ( .A1(n6437), .A2(n6436), .ZN(n6440) );
  INV_X1 U7449 ( .A(n6438), .ZN(n6439) );
  NAND2_X1 U7450 ( .A1(n6439), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U7451 ( .A1(n6440), .A2(n6442), .ZN(n6445) );
  INV_X1 U7452 ( .A(n6441), .ZN(n6450) );
  AOI22_X1 U7453 ( .A1(n6447), .A2(n6445), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6450), .ZN(n6501) );
  INV_X1 U7454 ( .A(n6442), .ZN(n6491) );
  AOI22_X1 U7455 ( .A1(n6495), .A2(n6444), .B1(n6443), .B2(n6491), .ZN(n6453)
         );
  INV_X1 U7456 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U7457 ( .A1(n6447), .A2(n6446), .ZN(n6449) );
  OAI211_X1 U7458 ( .C1(n6411), .C2(n6450), .A(n6449), .B(n6448), .ZN(n6497)
         );
  AOI22_X1 U7459 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6497), .B1(n6451), 
        .B2(n6494), .ZN(n6452) );
  OAI211_X1 U7460 ( .C1(n6501), .C2(n6454), .A(n6453), .B(n6452), .ZN(U3108)
         );
  AOI22_X1 U7461 ( .A1(n6494), .A2(n6456), .B1(n6455), .B2(n6491), .ZN(n6459)
         );
  AOI22_X1 U7462 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6497), .B1(n6457), 
        .B2(n6495), .ZN(n6458) );
  OAI211_X1 U7463 ( .C1(n6501), .C2(n6460), .A(n6459), .B(n6458), .ZN(U3109)
         );
  AOI22_X1 U7464 ( .A1(n6494), .A2(n6462), .B1(n6461), .B2(n6491), .ZN(n6465)
         );
  AOI22_X1 U7465 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6497), .B1(n6463), 
        .B2(n6495), .ZN(n6464) );
  OAI211_X1 U7466 ( .C1(n6501), .C2(n6466), .A(n6465), .B(n6464), .ZN(U3110)
         );
  AOI22_X1 U7467 ( .A1(n6494), .A2(n6468), .B1(n6467), .B2(n6491), .ZN(n6471)
         );
  AOI22_X1 U7468 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6497), .B1(n6469), 
        .B2(n6495), .ZN(n6470) );
  OAI211_X1 U7469 ( .C1(n6501), .C2(n6472), .A(n6471), .B(n6470), .ZN(U3111)
         );
  AOI22_X1 U7470 ( .A1(n6494), .A2(n6474), .B1(n6473), .B2(n6491), .ZN(n6477)
         );
  AOI22_X1 U7471 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6497), .B1(n6475), 
        .B2(n6495), .ZN(n6476) );
  OAI211_X1 U7472 ( .C1(n6501), .C2(n6478), .A(n6477), .B(n6476), .ZN(U3112)
         );
  AOI22_X1 U7473 ( .A1(n6494), .A2(n6480), .B1(n6479), .B2(n6491), .ZN(n6483)
         );
  AOI22_X1 U7474 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6497), .B1(n6481), 
        .B2(n6495), .ZN(n6482) );
  OAI211_X1 U7475 ( .C1(n6501), .C2(n6484), .A(n6483), .B(n6482), .ZN(U3113)
         );
  AOI22_X1 U7476 ( .A1(n6495), .A2(n6486), .B1(n6485), .B2(n6491), .ZN(n6489)
         );
  AOI22_X1 U7477 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6497), .B1(n6487), 
        .B2(n6494), .ZN(n6488) );
  OAI211_X1 U7478 ( .C1(n6501), .C2(n6490), .A(n6489), .B(n6488), .ZN(U3114)
         );
  AOI22_X1 U7479 ( .A1(n6494), .A2(n6493), .B1(n6492), .B2(n6491), .ZN(n6499)
         );
  AOI22_X1 U7480 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6497), .B1(n6496), 
        .B2(n6495), .ZN(n6498) );
  OAI211_X1 U7481 ( .C1(n6501), .C2(n6500), .A(n6499), .B(n6498), .ZN(U3115)
         );
  OAI21_X1 U7482 ( .B1(n6503), .B2(n6502), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .ZN(n6504) );
  NOR2_X1 U7483 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  INV_X1 U7484 ( .A(n6506), .ZN(n6510) );
  OAI22_X1 U7485 ( .A1(n6508), .A2(n6507), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6506), .ZN(n6509) );
  OAI21_X1 U7486 ( .B1(n6510), .B2(n6969), .A(n6509), .ZN(n6512) );
  AOI222_X1 U7487 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6512), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6511), .C1(n6512), .C2(n6511), 
        .ZN(n6514) );
  AOI222_X1 U7488 ( .A1(n6514), .A2(n6641), .B1(n6514), .B2(n6513), .C1(n6641), 
        .C2(n6513), .ZN(n6531) );
  NOR2_X1 U7489 ( .A1(n6516), .A2(n6515), .ZN(n6520) );
  AOI21_X1 U7490 ( .B1(n6518), .B2(n6517), .A(n6521), .ZN(n6519) );
  AOI211_X1 U7491 ( .C1(n6522), .C2(n6521), .A(n6520), .B(n6519), .ZN(n6653)
         );
  INV_X1 U7492 ( .A(n6653), .ZN(n6527) );
  INV_X1 U7493 ( .A(MORE_REG_SCAN_IN), .ZN(n6794) );
  AOI21_X1 U7494 ( .B1(n6524), .B2(n6794), .A(n6523), .ZN(n6525) );
  NOR4_X1 U7495 ( .A1(n6528), .A2(n6527), .A3(n6526), .A4(n6525), .ZN(n6529)
         );
  OAI211_X1 U7496 ( .C1(n6531), .C2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6530), .B(n6529), .ZN(n6537) );
  AOI22_X1 U7497 ( .A1(n6537), .A2(n6544), .B1(n6532), .B2(n6625), .ZN(n6542)
         );
  OR2_X1 U7498 ( .A1(n6563), .A2(n6533), .ZN(n6535) );
  OAI21_X1 U7499 ( .B1(n6552), .B2(n4438), .A(n6660), .ZN(n6534) );
  OAI211_X1 U7500 ( .C1(n6536), .C2(n6535), .A(STATE2_REG_2__SCAN_IN), .B(
        n6534), .ZN(n6538) );
  AOI221_X1 U7501 ( .B1(STATE2_REG_1__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(n6537), .C2(STATE2_REG_0__SCAN_IN), .A(n6538), .ZN(n6627) );
  OAI221_X1 U7502 ( .B1(n6627), .B2(READY_N), .C1(n6627), .C2(n6656), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6551) );
  OAI211_X1 U7503 ( .C1(n6659), .C2(n6539), .A(n6660), .B(n6538), .ZN(n6540)
         );
  NAND4_X1 U7504 ( .A1(n6542), .A2(n6541), .A3(n6551), .A4(n6540), .ZN(U3148)
         );
  INV_X1 U7505 ( .A(n6543), .ZN(n6548) );
  NOR2_X1 U7506 ( .A1(READY_N), .A2(n6660), .ZN(n6554) );
  AOI21_X1 U7507 ( .B1(n6545), .B2(n6554), .A(n6544), .ZN(n6546) );
  NOR2_X1 U7508 ( .A1(n6546), .A2(n6627), .ZN(n6547) );
  AOI211_X1 U7509 ( .C1(n6627), .C2(n6549), .A(n6548), .B(n6547), .ZN(n6550)
         );
  OAI21_X1 U7510 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(U3149) );
  OAI211_X1 U7511 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6554), .A(n6553), .B(
        n6659), .ZN(n6555) );
  NAND2_X1 U7512 ( .A1(n6556), .A2(n6555), .ZN(U3150) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n3124), .ZN(U3151) );
  AND2_X1 U7514 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n3124), .ZN(U3152) );
  INV_X1 U7515 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6743) );
  NOR2_X1 U7516 ( .A1(n3125), .A2(n6743), .ZN(U3153) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n3124), .ZN(U3154) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n3124), .ZN(U3155) );
  INV_X1 U7519 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6864) );
  NOR2_X1 U7520 ( .A1(n3125), .A2(n6864), .ZN(U3156) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n3124), .ZN(U3157) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n3124), .ZN(U3158) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n3124), .ZN(U3159) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n3124), .ZN(U3160) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n3124), .ZN(U3161) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n3124), .ZN(U3162) );
  AND2_X1 U7527 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n3124), .ZN(U3163) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n3124), .ZN(U3164) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n3124), .ZN(U3165) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n3124), .ZN(U3166) );
  NOR2_X1 U7531 ( .A1(n3125), .A2(n6693), .ZN(U3167) );
  INV_X1 U7532 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6807) );
  NOR2_X1 U7533 ( .A1(n3125), .A2(n6807), .ZN(U3168) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n3124), .ZN(U3169) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n3124), .ZN(U3170) );
  INV_X1 U7536 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6740) );
  NOR2_X1 U7537 ( .A1(n3125), .A2(n6740), .ZN(U3171) );
  AND2_X1 U7538 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n3124), .ZN(U3172) );
  NOR2_X1 U7539 ( .A1(n3125), .A2(n6697), .ZN(U3173) );
  AND2_X1 U7540 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n3124), .ZN(U3174) );
  AND2_X1 U7541 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n3124), .ZN(U3175) );
  AND2_X1 U7542 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n3124), .ZN(U3176) );
  INV_X1 U7543 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U7544 ( .A1(n3125), .A2(n6676), .ZN(U3177) );
  INV_X1 U7545 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U7546 ( .A1(n3125), .A2(n6921), .ZN(U3178) );
  AND2_X1 U7547 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n3124), .ZN(U3179) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n3124), .ZN(U3180) );
  NAND2_X1 U7549 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6561) );
  NAND2_X1 U7550 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6566) );
  NAND2_X1 U7551 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7552 ( .A1(n6566), .A2(n6567), .ZN(n6559) );
  INV_X1 U7553 ( .A(NA_N), .ZN(n6558) );
  INV_X1 U7554 ( .A(n6568), .ZN(n6557) );
  AOI211_X1 U7555 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6558), .A(
        STATE_REG_0__SCAN_IN), .B(n6557), .ZN(n6573) );
  AOI21_X1 U7556 ( .B1(n6568), .B2(n6559), .A(n6573), .ZN(n6560) );
  OAI221_X1 U7557 ( .B1(n6667), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6667), 
        .C2(n6561), .A(n6560), .ZN(U3181) );
  INV_X1 U7558 ( .A(n6566), .ZN(n6565) );
  INV_X1 U7559 ( .A(n6561), .ZN(n6562) );
  AOI21_X1 U7560 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6562), .ZN(n6564) );
  OAI211_X1 U7561 ( .C1(n6565), .C2(n6564), .A(n6563), .B(n6567), .ZN(U3182)
         );
  AOI221_X1 U7562 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4438), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6570) );
  OAI211_X1 U7563 ( .C1(n6568), .C2(n6567), .A(STATE_REG_0__SCAN_IN), .B(n6566), .ZN(n6569) );
  AOI21_X1 U7564 ( .B1(HOLD), .B2(n6570), .A(n6569), .ZN(n6572) );
  NAND4_X1 U7565 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .A3(
        STATE_REG_0__SCAN_IN), .A4(REQUESTPENDING_REG_SCAN_IN), .ZN(n6571) );
  OAI22_X1 U7566 ( .A1(n6573), .A2(n6572), .B1(NA_N), .B2(n6571), .ZN(U3183)
         );
  NAND2_X1 U7567 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6667), .ZN(n6611) );
  NOR2_X2 U7568 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6651), .ZN(n6609) );
  AOI22_X1 U7569 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6651), .ZN(n6574) );
  OAI21_X1 U7570 ( .B1(n6575), .B2(n6611), .A(n6574), .ZN(U3184) );
  AOI22_X1 U7571 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6651), .ZN(n6576) );
  OAI21_X1 U7572 ( .B1(n6577), .B2(n6611), .A(n6576), .ZN(U3185) );
  INV_X1 U7573 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6715) );
  OAI222_X1 U7574 ( .A1(n6611), .A2(n6681), .B1(n6715), .B2(n6667), .C1(n6879), 
        .C2(n6617), .ZN(U3186) );
  AOI22_X1 U7575 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6651), .ZN(n6578) );
  OAI21_X1 U7576 ( .B1(n6879), .B2(n6611), .A(n6578), .ZN(U3187) );
  AOI22_X1 U7577 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6651), .ZN(n6579) );
  OAI21_X1 U7578 ( .B1(n6580), .B2(n6611), .A(n6579), .ZN(U3188) );
  INV_X1 U7579 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6711) );
  OAI222_X1 U7580 ( .A1(n6611), .A2(n6581), .B1(n6711), .B2(n6667), .C1(n6583), 
        .C2(n6617), .ZN(U3189) );
  AOI22_X1 U7581 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6651), .ZN(n6582) );
  OAI21_X1 U7582 ( .B1(n6583), .B2(n6611), .A(n6582), .ZN(U3190) );
  AOI22_X1 U7583 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6651), .ZN(n6584) );
  OAI21_X1 U7584 ( .B1(n6765), .B2(n6611), .A(n6584), .ZN(U3191) );
  INV_X1 U7585 ( .A(n6611), .ZN(n6615) );
  AOI22_X1 U7586 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6651), .ZN(n6585) );
  OAI21_X1 U7587 ( .B1(n6797), .B2(n6617), .A(n6585), .ZN(U3192) );
  INV_X1 U7588 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6769) );
  OAI222_X1 U7589 ( .A1(n6611), .A2(n6797), .B1(n6769), .B2(n6667), .C1(n6862), 
        .C2(n6617), .ZN(U3193) );
  AOI22_X1 U7590 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6651), .ZN(n6586) );
  OAI21_X1 U7591 ( .B1(n6587), .B2(n6617), .A(n6586), .ZN(U3194) );
  AOI22_X1 U7592 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6651), .ZN(n6588) );
  OAI21_X1 U7593 ( .B1(n6875), .B2(n6617), .A(n6588), .ZN(U3195) );
  INV_X1 U7594 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6849) );
  OAI222_X1 U7595 ( .A1(n6611), .A2(n6875), .B1(n6849), .B2(n6667), .C1(n6590), 
        .C2(n6617), .ZN(U3196) );
  AOI22_X1 U7596 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6651), .ZN(n6589) );
  OAI21_X1 U7597 ( .B1(n6590), .B2(n6611), .A(n6589), .ZN(U3197) );
  INV_X1 U7598 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6838) );
  OAI222_X1 U7599 ( .A1(n6611), .A2(n6591), .B1(n6838), .B2(n6667), .C1(n6592), 
        .C2(n6617), .ZN(U3198) );
  INV_X1 U7600 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6894) );
  OAI222_X1 U7601 ( .A1(n6611), .A2(n6592), .B1(n6894), .B2(n6667), .C1(n6867), 
        .C2(n6617), .ZN(U3199) );
  INV_X1 U7602 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6834) );
  OAI222_X1 U7603 ( .A1(n6617), .A2(n6594), .B1(n6834), .B2(n6667), .C1(n6867), 
        .C2(n6611), .ZN(U3200) );
  AOI22_X1 U7604 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6651), .ZN(n6593) );
  OAI21_X1 U7605 ( .B1(n6594), .B2(n6611), .A(n6593), .ZN(U3201) );
  AOI22_X1 U7606 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6651), .ZN(n6595) );
  OAI21_X1 U7607 ( .B1(n6596), .B2(n6611), .A(n6595), .ZN(U3202) );
  INV_X1 U7608 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6597) );
  INV_X1 U7609 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6813) );
  OAI222_X1 U7610 ( .A1(n6611), .A2(n6597), .B1(n6813), .B2(n6667), .C1(n6707), 
        .C2(n6617), .ZN(U3203) );
  AOI22_X1 U7611 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6651), .ZN(n6598) );
  OAI21_X1 U7612 ( .B1(n6600), .B2(n6617), .A(n6598), .ZN(U3204) );
  AOI22_X1 U7613 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6651), .ZN(n6599) );
  OAI21_X1 U7614 ( .B1(n6600), .B2(n6611), .A(n6599), .ZN(U3205) );
  INV_X1 U7615 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6602) );
  INV_X1 U7616 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6884) );
  OAI222_X1 U7617 ( .A1(n6611), .A2(n6602), .B1(n6884), .B2(n6667), .C1(n6601), 
        .C2(n6617), .ZN(U3206) );
  INV_X1 U7618 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6757) );
  AOI22_X1 U7619 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6651), .ZN(n6603) );
  OAI21_X1 U7620 ( .B1(n6757), .B2(n6617), .A(n6603), .ZN(U3207) );
  AOI22_X1 U7621 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6651), .ZN(n6604) );
  OAI21_X1 U7622 ( .B1(n6605), .B2(n6617), .A(n6604), .ZN(U3208) );
  AOI22_X1 U7623 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6651), .ZN(n6606) );
  OAI21_X1 U7624 ( .B1(n6608), .B2(n6617), .A(n6606), .ZN(U3209) );
  AOI22_X1 U7625 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6651), .ZN(n6607) );
  OAI21_X1 U7626 ( .B1(n6608), .B2(n6611), .A(n6607), .ZN(U3210) );
  AOI22_X1 U7627 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6651), .ZN(n6610) );
  OAI21_X1 U7628 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(U3211) );
  AOI22_X1 U7629 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6651), .ZN(n6613) );
  OAI21_X1 U7630 ( .B1(n6614), .B2(n6617), .A(n6613), .ZN(U3212) );
  INV_X1 U7631 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6618) );
  AOI22_X1 U7632 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6615), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6651), .ZN(n6616) );
  OAI21_X1 U7633 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(U3213) );
  INV_X1 U7634 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6823) );
  AOI22_X1 U7635 ( .A1(n6667), .A2(n6619), .B1(n6823), .B2(n6651), .ZN(U3445)
         );
  INV_X1 U7636 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6644) );
  INV_X1 U7637 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U7638 ( .A1(n6667), .A2(n6644), .B1(n6675), .B2(n6651), .ZN(U3446)
         );
  MUX2_X1 U7639 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6667), .Z(U3447) );
  MUX2_X1 U7640 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6667), .Z(U3448) );
  INV_X1 U7641 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6621) );
  INV_X1 U7642 ( .A(n6622), .ZN(n6620) );
  AOI21_X1 U7643 ( .B1(n6621), .B2(n3124), .A(n6620), .ZN(U3451) );
  OAI21_X1 U7644 ( .B1(n3125), .B2(n6623), .A(n6622), .ZN(U3452) );
  AOI211_X1 U7645 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6627), .A(n6626), .B(
        n6625), .ZN(n6628) );
  INV_X1 U7646 ( .A(n6628), .ZN(U3453) );
  INV_X1 U7647 ( .A(n6629), .ZN(n6632) );
  AOI21_X1 U7648 ( .B1(n6632), .B2(n6631), .A(n6630), .ZN(n6638) );
  INV_X1 U7649 ( .A(n6633), .ZN(n6634) );
  OAI22_X1 U7650 ( .A1(n4602), .A2(n6636), .B1(n6635), .B2(n6634), .ZN(n6637)
         );
  NOR2_X1 U7651 ( .A1(n6638), .A2(n6637), .ZN(n6640) );
  AOI22_X1 U7652 ( .A1(n6642), .A2(n6641), .B1(n6640), .B2(n6639), .ZN(U3462)
         );
  AOI211_X1 U7653 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6643) );
  AOI21_X1 U7654 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6643), .ZN(n6645) );
  AOI22_X1 U7655 ( .A1(n6649), .A2(n6645), .B1(n6644), .B2(n6646), .ZN(U3468)
         );
  NOR2_X1 U7656 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6648) );
  INV_X1 U7657 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U7658 ( .A1(n6649), .A2(n6648), .B1(n6647), .B2(n6646), .ZN(U3469)
         );
  NAND2_X1 U7659 ( .A1(n6651), .A2(W_R_N_REG_SCAN_IN), .ZN(n6650) );
  OAI21_X1 U7660 ( .B1(n6651), .B2(READREQUEST_REG_SCAN_IN), .A(n6650), .ZN(
        U3470) );
  AOI22_X1 U7661 ( .A1(n6654), .A2(n6653), .B1(n6794), .B2(n6652), .ZN(U3471)
         );
  AOI211_X1 U7662 ( .C1(n6658), .C2(n6657), .A(n6656), .B(n6655), .ZN(n6661)
         );
  OAI21_X1 U7663 ( .B1(n6661), .B2(n6660), .A(n6659), .ZN(n6666) );
  OAI211_X1 U7664 ( .C1(READY_N), .C2(n6664), .A(n6663), .B(n6662), .ZN(n6665)
         );
  MUX2_X1 U7665 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n6666), .S(n6665), .Z(
        U3472) );
  MUX2_X1 U7666 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6667), .Z(U3473) );
  INV_X1 U7667 ( .A(n6668), .ZN(n6673) );
  AOI222_X1 U7668 ( .A1(n6673), .A2(n6672), .B1(n6671), .B2(
        EBX_REG_14__SCAN_IN), .C1(n6670), .C2(n6669), .ZN(n6912) );
  AOI22_X1 U7669 ( .A1(n6676), .A2(keyinput60), .B1(keyinput103), .B2(n6675), 
        .ZN(n6674) );
  OAI221_X1 U7670 ( .B1(n6676), .B2(keyinput60), .C1(n6675), .C2(keyinput103), 
        .A(n6674), .ZN(n6688) );
  INV_X1 U7671 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6679) );
  AOI22_X1 U7672 ( .A1(n6679), .A2(keyinput4), .B1(keyinput12), .B2(n6678), 
        .ZN(n6677) );
  OAI221_X1 U7673 ( .B1(n6679), .B2(keyinput4), .C1(n6678), .C2(keyinput12), 
        .A(n6677), .ZN(n6687) );
  AOI22_X1 U7674 ( .A1(n6681), .A2(keyinput54), .B1(n5093), .B2(keyinput11), 
        .ZN(n6680) );
  OAI221_X1 U7675 ( .B1(n6681), .B2(keyinput54), .C1(n5093), .C2(keyinput11), 
        .A(n6680), .ZN(n6686) );
  AOI22_X1 U7676 ( .A1(n6684), .A2(keyinput21), .B1(n6683), .B2(keyinput72), 
        .ZN(n6682) );
  OAI221_X1 U7677 ( .B1(n6684), .B2(keyinput21), .C1(n6683), .C2(keyinput72), 
        .A(n6682), .ZN(n6685) );
  NOR4_X1 U7678 ( .A1(n6688), .A2(n6687), .A3(n6686), .A4(n6685), .ZN(n6738)
         );
  AOI22_X1 U7679 ( .A1(n6691), .A2(keyinput112), .B1(keyinput86), .B2(n6690), 
        .ZN(n6689) );
  OAI221_X1 U7680 ( .B1(n6691), .B2(keyinput112), .C1(n6690), .C2(keyinput86), 
        .A(n6689), .ZN(n6704) );
  AOI22_X1 U7681 ( .A1(n6694), .A2(keyinput53), .B1(n6693), .B2(keyinput85), 
        .ZN(n6692) );
  OAI221_X1 U7682 ( .B1(n6694), .B2(keyinput53), .C1(n6693), .C2(keyinput85), 
        .A(n6692), .ZN(n6703) );
  AOI22_X1 U7683 ( .A1(n6697), .A2(keyinput3), .B1(n6696), .B2(keyinput67), 
        .ZN(n6695) );
  OAI221_X1 U7684 ( .B1(n6697), .B2(keyinput3), .C1(n6696), .C2(keyinput67), 
        .A(n6695), .ZN(n6702) );
  INV_X1 U7685 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6699) );
  AOI22_X1 U7686 ( .A1(n6700), .A2(keyinput79), .B1(keyinput120), .B2(n6699), 
        .ZN(n6698) );
  OAI221_X1 U7687 ( .B1(n6700), .B2(keyinput79), .C1(n6699), .C2(keyinput120), 
        .A(n6698), .ZN(n6701) );
  NOR4_X1 U7688 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(n6737)
         );
  AOI22_X1 U7689 ( .A1(n6707), .A2(keyinput9), .B1(n6706), .B2(keyinput70), 
        .ZN(n6705) );
  OAI221_X1 U7690 ( .B1(n6707), .B2(keyinput9), .C1(n6706), .C2(keyinput70), 
        .A(n6705), .ZN(n6719) );
  AOI22_X1 U7691 ( .A1(n4626), .A2(keyinput32), .B1(n6709), .B2(keyinput77), 
        .ZN(n6708) );
  OAI221_X1 U7692 ( .B1(n4626), .B2(keyinput32), .C1(n6709), .C2(keyinput77), 
        .A(n6708), .ZN(n6718) );
  AOI22_X1 U7693 ( .A1(n6712), .A2(keyinput83), .B1(keyinput84), .B2(n6711), 
        .ZN(n6710) );
  OAI221_X1 U7694 ( .B1(n6712), .B2(keyinput83), .C1(n6711), .C2(keyinput84), 
        .A(n6710), .ZN(n6717) );
  AOI22_X1 U7695 ( .A1(n6715), .A2(keyinput28), .B1(n6714), .B2(keyinput109), 
        .ZN(n6713) );
  OAI221_X1 U7696 ( .B1(n6715), .B2(keyinput28), .C1(n6714), .C2(keyinput109), 
        .A(n6713), .ZN(n6716) );
  NOR4_X1 U7697 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6736)
         );
  INV_X1 U7698 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U7699 ( .A1(n6931), .A2(keyinput49), .B1(keyinput80), .B2(n6721), 
        .ZN(n6720) );
  OAI221_X1 U7700 ( .B1(n6931), .B2(keyinput49), .C1(n6721), .C2(keyinput80), 
        .A(n6720), .ZN(n6734) );
  AOI22_X1 U7701 ( .A1(n6724), .A2(keyinput123), .B1(keyinput19), .B2(n6723), 
        .ZN(n6722) );
  OAI221_X1 U7702 ( .B1(n6724), .B2(keyinput123), .C1(n6723), .C2(keyinput19), 
        .A(n6722), .ZN(n6728) );
  XNOR2_X1 U7703 ( .A(n6725), .B(keyinput90), .ZN(n6727) );
  XOR2_X1 U7704 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput95), .Z(n6726)
         );
  OR3_X1 U7705 ( .A1(n6728), .A2(n6727), .A3(n6726), .ZN(n6733) );
  AOI22_X1 U7706 ( .A1(n6731), .A2(keyinput76), .B1(n6730), .B2(keyinput100), 
        .ZN(n6729) );
  OAI221_X1 U7707 ( .B1(n6731), .B2(keyinput76), .C1(n6730), .C2(keyinput100), 
        .A(n6729), .ZN(n6732) );
  NOR3_X1 U7708 ( .A1(n6734), .A2(n6733), .A3(n6732), .ZN(n6735) );
  NAND4_X1 U7709 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .ZN(n6910)
         );
  AOI22_X1 U7710 ( .A1(n6740), .A2(keyinput82), .B1(n4325), .B2(keyinput92), 
        .ZN(n6739) );
  OAI221_X1 U7711 ( .B1(n6740), .B2(keyinput82), .C1(n4325), .C2(keyinput92), 
        .A(n6739), .ZN(n6749) );
  INV_X1 U7712 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7713 ( .A1(n6935), .A2(keyinput17), .B1(n6942), .B2(keyinput64), 
        .ZN(n6741) );
  OAI221_X1 U7714 ( .B1(n6935), .B2(keyinput17), .C1(n6942), .C2(keyinput64), 
        .A(n6741), .ZN(n6748) );
  INV_X1 U7715 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7716 ( .A1(n6960), .A2(keyinput2), .B1(keyinput20), .B2(n6743), 
        .ZN(n6742) );
  OAI221_X1 U7717 ( .B1(n6960), .B2(keyinput2), .C1(n6743), .C2(keyinput20), 
        .A(n6742), .ZN(n6747) );
  AOI22_X1 U7718 ( .A1(n6745), .A2(keyinput110), .B1(n6929), .B2(keyinput42), 
        .ZN(n6744) );
  OAI221_X1 U7719 ( .B1(n6745), .B2(keyinput110), .C1(n6929), .C2(keyinput42), 
        .A(n6744), .ZN(n6746) );
  NOR4_X1 U7720 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n6792)
         );
  AOI22_X1 U7721 ( .A1(n6966), .A2(keyinput43), .B1(keyinput1), .B2(n6933), 
        .ZN(n6750) );
  OAI221_X1 U7722 ( .B1(n6966), .B2(keyinput43), .C1(n6933), .C2(keyinput1), 
        .A(n6750), .ZN(n6761) );
  AOI22_X1 U7723 ( .A1(n6932), .A2(keyinput78), .B1(keyinput35), .B2(n6752), 
        .ZN(n6751) );
  OAI221_X1 U7724 ( .B1(n6932), .B2(keyinput78), .C1(n6752), .C2(keyinput35), 
        .A(n6751), .ZN(n6760) );
  AOI22_X1 U7725 ( .A1(n6755), .A2(keyinput44), .B1(n6754), .B2(keyinput46), 
        .ZN(n6753) );
  OAI221_X1 U7726 ( .B1(n6755), .B2(keyinput44), .C1(n6754), .C2(keyinput46), 
        .A(n6753), .ZN(n6759) );
  AOI22_X1 U7727 ( .A1(n5597), .A2(keyinput124), .B1(keyinput56), .B2(n6757), 
        .ZN(n6756) );
  OAI221_X1 U7728 ( .B1(n5597), .B2(keyinput124), .C1(n6757), .C2(keyinput56), 
        .A(n6756), .ZN(n6758) );
  NOR4_X1 U7729 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6791)
         );
  AOI22_X1 U7730 ( .A1(n6763), .A2(keyinput22), .B1(keyinput59), .B2(n6921), 
        .ZN(n6762) );
  OAI221_X1 U7731 ( .B1(n6763), .B2(keyinput22), .C1(n6921), .C2(keyinput59), 
        .A(n6762), .ZN(n6774) );
  AOI22_X1 U7732 ( .A1(n6766), .A2(keyinput57), .B1(keyinput68), .B2(n6765), 
        .ZN(n6764) );
  OAI221_X1 U7733 ( .B1(n6766), .B2(keyinput57), .C1(n6765), .C2(keyinput68), 
        .A(n6764), .ZN(n6773) );
  AOI22_X1 U7734 ( .A1(n6953), .A2(keyinput75), .B1(keyinput34), .B2(n6967), 
        .ZN(n6767) );
  OAI221_X1 U7735 ( .B1(n6953), .B2(keyinput75), .C1(n6967), .C2(keyinput34), 
        .A(n6767), .ZN(n6772) );
  INV_X1 U7736 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U7737 ( .A1(n6770), .A2(keyinput106), .B1(keyinput40), .B2(n6769), 
        .ZN(n6768) );
  OAI221_X1 U7738 ( .B1(n6770), .B2(keyinput106), .C1(n6769), .C2(keyinput40), 
        .A(n6768), .ZN(n6771) );
  NOR4_X1 U7739 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6790)
         );
  INV_X1 U7740 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6776) );
  AOI22_X1 U7741 ( .A1(n6952), .A2(keyinput37), .B1(keyinput55), .B2(n6776), 
        .ZN(n6775) );
  OAI221_X1 U7742 ( .B1(n6952), .B2(keyinput37), .C1(n6776), .C2(keyinput55), 
        .A(n6775), .ZN(n6788) );
  AOI22_X1 U7743 ( .A1(n6779), .A2(keyinput81), .B1(n6778), .B2(keyinput51), 
        .ZN(n6777) );
  OAI221_X1 U7744 ( .B1(n6779), .B2(keyinput81), .C1(n6778), .C2(keyinput51), 
        .A(n6777), .ZN(n6787) );
  AOI22_X1 U7745 ( .A1(n6946), .A2(keyinput25), .B1(n6781), .B2(keyinput88), 
        .ZN(n6780) );
  OAI221_X1 U7746 ( .B1(n6946), .B2(keyinput25), .C1(n6781), .C2(keyinput88), 
        .A(n6780), .ZN(n6786) );
  INV_X1 U7747 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7748 ( .A1(n6784), .A2(keyinput66), .B1(n6783), .B2(keyinput73), 
        .ZN(n6782) );
  OAI221_X1 U7749 ( .B1(n6784), .B2(keyinput66), .C1(n6783), .C2(keyinput73), 
        .A(n6782), .ZN(n6785) );
  NOR4_X1 U7750 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6789)
         );
  NAND4_X1 U7751 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6909)
         );
  AOI22_X1 U7752 ( .A1(n6795), .A2(keyinput97), .B1(keyinput8), .B2(n6794), 
        .ZN(n6793) );
  OAI221_X1 U7753 ( .B1(n6795), .B2(keyinput97), .C1(n6794), .C2(keyinput8), 
        .A(n6793), .ZN(n6805) );
  INV_X1 U7754 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U7755 ( .A1(n6798), .A2(keyinput121), .B1(keyinput111), .B2(n6797), 
        .ZN(n6796) );
  OAI221_X1 U7756 ( .B1(n6798), .B2(keyinput121), .C1(n6797), .C2(keyinput111), 
        .A(n6796), .ZN(n6804) );
  INV_X1 U7757 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6800) );
  AOI22_X1 U7758 ( .A1(n6964), .A2(keyinput113), .B1(keyinput7), .B2(n6800), 
        .ZN(n6799) );
  OAI221_X1 U7759 ( .B1(n6964), .B2(keyinput113), .C1(n6800), .C2(keyinput7), 
        .A(n6799), .ZN(n6803) );
  AOI22_X1 U7760 ( .A1(n4438), .A2(keyinput118), .B1(keyinput13), .B2(n6945), 
        .ZN(n6801) );
  OAI221_X1 U7761 ( .B1(n4438), .B2(keyinput118), .C1(n6945), .C2(keyinput13), 
        .A(n6801), .ZN(n6802) );
  NOR4_X1 U7762 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6847)
         );
  AOI22_X1 U7763 ( .A1(n6808), .A2(keyinput16), .B1(keyinput38), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7764 ( .B1(n6808), .B2(keyinput16), .C1(n6807), .C2(keyinput38), 
        .A(n6806), .ZN(n6819) );
  AOI22_X1 U7765 ( .A1(n6811), .A2(keyinput47), .B1(keyinput89), .B2(n6810), 
        .ZN(n6809) );
  OAI221_X1 U7766 ( .B1(n6811), .B2(keyinput47), .C1(n6810), .C2(keyinput89), 
        .A(n6809), .ZN(n6818) );
  INV_X1 U7767 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U7768 ( .A1(n6814), .A2(keyinput31), .B1(n6813), .B2(keyinput115), 
        .ZN(n6812) );
  OAI221_X1 U7769 ( .B1(n6814), .B2(keyinput31), .C1(n6813), .C2(keyinput115), 
        .A(n6812), .ZN(n6817) );
  INV_X1 U7770 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6963) );
  INV_X1 U7771 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6941) );
  AOI22_X1 U7772 ( .A1(n6963), .A2(keyinput101), .B1(keyinput30), .B2(n6941), 
        .ZN(n6815) );
  OAI221_X1 U7773 ( .B1(n6963), .B2(keyinput101), .C1(n6941), .C2(keyinput30), 
        .A(n6815), .ZN(n6816) );
  NOR4_X1 U7774 ( .A1(n6819), .A2(n6818), .A3(n6817), .A4(n6816), .ZN(n6846)
         );
  AOI22_X1 U7775 ( .A1(n6821), .A2(keyinput114), .B1(keyinput24), .B2(n4641), 
        .ZN(n6820) );
  OAI221_X1 U7776 ( .B1(n6821), .B2(keyinput114), .C1(n4641), .C2(keyinput24), 
        .A(n6820), .ZN(n6830) );
  AOI22_X1 U7777 ( .A1(n6954), .A2(keyinput102), .B1(keyinput125), .B2(n6823), 
        .ZN(n6822) );
  OAI221_X1 U7778 ( .B1(n6954), .B2(keyinput102), .C1(n6823), .C2(keyinput125), 
        .A(n6822), .ZN(n6829) );
  AOI22_X1 U7779 ( .A1(n6825), .A2(keyinput126), .B1(n3199), .B2(keyinput10), 
        .ZN(n6824) );
  OAI221_X1 U7780 ( .B1(n6825), .B2(keyinput126), .C1(n3199), .C2(keyinput10), 
        .A(n6824), .ZN(n6828) );
  AOI22_X1 U7781 ( .A1(n6968), .A2(keyinput5), .B1(n5078), .B2(keyinput0), 
        .ZN(n6826) );
  OAI221_X1 U7782 ( .B1(n6968), .B2(keyinput5), .C1(n5078), .C2(keyinput0), 
        .A(n6826), .ZN(n6827) );
  NOR4_X1 U7783 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n6845)
         );
  AOI22_X1 U7784 ( .A1(n6832), .A2(keyinput52), .B1(n6961), .B2(keyinput98), 
        .ZN(n6831) );
  OAI221_X1 U7785 ( .B1(n6832), .B2(keyinput52), .C1(n6961), .C2(keyinput98), 
        .A(n6831), .ZN(n6843) );
  AOI22_X1 U7786 ( .A1(n6834), .A2(keyinput26), .B1(n3647), .B2(keyinput69), 
        .ZN(n6833) );
  OAI221_X1 U7787 ( .B1(n6834), .B2(keyinput26), .C1(n3647), .C2(keyinput69), 
        .A(n6833), .ZN(n6842) );
  AOI22_X1 U7788 ( .A1(n6959), .A2(keyinput116), .B1(n6836), .B2(keyinput94), 
        .ZN(n6835) );
  OAI221_X1 U7789 ( .B1(n6959), .B2(keyinput116), .C1(n6836), .C2(keyinput94), 
        .A(n6835), .ZN(n6841) );
  AOI22_X1 U7790 ( .A1(n6839), .A2(keyinput63), .B1(keyinput91), .B2(n6838), 
        .ZN(n6837) );
  OAI221_X1 U7791 ( .B1(n6839), .B2(keyinput63), .C1(n6838), .C2(keyinput91), 
        .A(n6837), .ZN(n6840) );
  NOR4_X1 U7792 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n6844)
         );
  NAND4_X1 U7793 ( .A1(n6847), .A2(n6846), .A3(n6845), .A4(n6844), .ZN(n6908)
         );
  AOI22_X1 U7794 ( .A1(n6850), .A2(keyinput105), .B1(keyinput61), .B2(n6849), 
        .ZN(n6848) );
  OAI221_X1 U7795 ( .B1(n6850), .B2(keyinput105), .C1(n6849), .C2(keyinput61), 
        .A(n6848), .ZN(n6860) );
  AOI22_X1 U7796 ( .A1(n6852), .A2(keyinput99), .B1(n6930), .B2(keyinput33), 
        .ZN(n6851) );
  OAI221_X1 U7797 ( .B1(n6852), .B2(keyinput99), .C1(n6930), .C2(keyinput33), 
        .A(n6851), .ZN(n6859) );
  INV_X1 U7798 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6854) );
  AOI22_X1 U7799 ( .A1(n6854), .A2(keyinput39), .B1(keyinput74), .B2(n6913), 
        .ZN(n6853) );
  OAI221_X1 U7800 ( .B1(n6854), .B2(keyinput39), .C1(n6913), .C2(keyinput74), 
        .A(n6853), .ZN(n6858) );
  INV_X1 U7801 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7802 ( .A1(n6936), .A2(keyinput122), .B1(keyinput107), .B2(n6856), 
        .ZN(n6855) );
  OAI221_X1 U7803 ( .B1(n6936), .B2(keyinput122), .C1(n6856), .C2(keyinput107), 
        .A(n6855), .ZN(n6857) );
  NOR4_X1 U7804 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n6906)
         );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U7806 ( .A1(n6862), .A2(keyinput45), .B1(n6934), .B2(keyinput27), 
        .ZN(n6861) );
  OAI221_X1 U7807 ( .B1(n6862), .B2(keyinput45), .C1(n6934), .C2(keyinput27), 
        .A(n6861), .ZN(n6873) );
  INV_X1 U7808 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U7809 ( .A1(n6865), .A2(keyinput108), .B1(keyinput36), .B2(n6864), 
        .ZN(n6863) );
  OAI221_X1 U7810 ( .B1(n6865), .B2(keyinput108), .C1(n6864), .C2(keyinput36), 
        .A(n6863), .ZN(n6872) );
  AOI22_X1 U7811 ( .A1(n6867), .A2(keyinput117), .B1(n3946), .B2(keyinput71), 
        .ZN(n6866) );
  OAI221_X1 U7812 ( .B1(n6867), .B2(keyinput117), .C1(n3946), .C2(keyinput71), 
        .A(n6866), .ZN(n6871) );
  INV_X1 U7813 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6947) );
  AOI22_X1 U7814 ( .A1(n6869), .A2(keyinput48), .B1(n6947), .B2(keyinput41), 
        .ZN(n6868) );
  OAI221_X1 U7815 ( .B1(n6869), .B2(keyinput48), .C1(n6947), .C2(keyinput41), 
        .A(n6868), .ZN(n6870) );
  NOR4_X1 U7816 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n6905)
         );
  AOI22_X1 U7817 ( .A1(n6876), .A2(keyinput127), .B1(n6875), .B2(keyinput14), 
        .ZN(n6874) );
  OAI221_X1 U7818 ( .B1(n6876), .B2(keyinput127), .C1(n6875), .C2(keyinput14), 
        .A(n6874), .ZN(n6888) );
  AOI22_X1 U7819 ( .A1(n6879), .A2(keyinput87), .B1(keyinput65), .B2(n6878), 
        .ZN(n6877) );
  OAI221_X1 U7820 ( .B1(n6879), .B2(keyinput87), .C1(n6878), .C2(keyinput65), 
        .A(n6877), .ZN(n6887) );
  INV_X1 U7821 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U7822 ( .A1(n6965), .A2(keyinput18), .B1(keyinput96), .B2(n6881), 
        .ZN(n6880) );
  OAI221_X1 U7823 ( .B1(n6965), .B2(keyinput18), .C1(n6881), .C2(keyinput96), 
        .A(n6880), .ZN(n6886) );
  AOI22_X1 U7824 ( .A1(n6884), .A2(keyinput104), .B1(n6883), .B2(keyinput15), 
        .ZN(n6882) );
  OAI221_X1 U7825 ( .B1(n6884), .B2(keyinput104), .C1(n6883), .C2(keyinput15), 
        .A(n6882), .ZN(n6885) );
  NOR4_X1 U7826 ( .A1(n6888), .A2(n6887), .A3(n6886), .A4(n6885), .ZN(n6904)
         );
  INV_X1 U7827 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6890) );
  INV_X1 U7828 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6962) );
  AOI22_X1 U7829 ( .A1(n6890), .A2(keyinput6), .B1(keyinput93), .B2(n6962), 
        .ZN(n6889) );
  OAI221_X1 U7830 ( .B1(n6890), .B2(keyinput6), .C1(n6962), .C2(keyinput93), 
        .A(n6889), .ZN(n6902) );
  AOI22_X1 U7831 ( .A1(n6969), .A2(keyinput29), .B1(keyinput58), .B2(n6892), 
        .ZN(n6891) );
  OAI221_X1 U7832 ( .B1(n6969), .B2(keyinput29), .C1(n6892), .C2(keyinput58), 
        .A(n6891), .ZN(n6901) );
  INV_X1 U7833 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U7834 ( .A1(n6895), .A2(keyinput119), .B1(keyinput23), .B2(n6894), 
        .ZN(n6893) );
  OAI221_X1 U7835 ( .B1(n6895), .B2(keyinput119), .C1(n6894), .C2(keyinput23), 
        .A(n6893), .ZN(n6900) );
  AOI22_X1 U7836 ( .A1(n6898), .A2(keyinput50), .B1(keyinput62), .B2(n6897), 
        .ZN(n6896) );
  OAI221_X1 U7837 ( .B1(n6898), .B2(keyinput50), .C1(n6897), .C2(keyinput62), 
        .A(n6896), .ZN(n6899) );
  NOR4_X1 U7838 ( .A1(n6902), .A2(n6901), .A3(n6900), .A4(n6899), .ZN(n6903)
         );
  NAND4_X1 U7839 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n6907)
         );
  NOR4_X1 U7840 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6911)
         );
  XNOR2_X1 U7841 ( .A(n6912), .B(n6911), .ZN(n6987) );
  NOR4_X1 U7842 ( .A1(EBX_REG_18__SCAN_IN), .A2(DATAWIDTH_REG_29__SCAN_IN), 
        .A3(DATAO_REG_2__SCAN_IN), .A4(MORE_REG_SCAN_IN), .ZN(n6985) );
  NOR4_X1 U7843 ( .A1(ADDRESS_REG_5__SCAN_IN), .A2(DATAO_REG_1__SCAN_IN), .A3(
        DATAO_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6984) );
  NOR4_X1 U7844 ( .A1(EAX_REG_25__SCAN_IN), .A2(EAX_REG_27__SCAN_IN), .A3(
        DATAI_29_), .A4(DATAI_12_), .ZN(n6914) );
  NAND3_X1 U7845 ( .A1(ADS_N_REG_SCAN_IN), .A2(n6914), .A3(n6913), .ZN(n6920)
         );
  NOR4_X1 U7846 ( .A1(REIP_REG_8__SCAN_IN), .A2(DATAO_REG_23__SCAN_IN), .A3(
        UWORD_REG_9__SCAN_IN), .A4(DATAO_REG_30__SCAN_IN), .ZN(n6918) );
  NOR4_X1 U7847 ( .A1(READY_N), .A2(BE_N_REG_3__SCAN_IN), .A3(
        LWORD_REG_3__SCAN_IN), .A4(DATAO_REG_7__SCAN_IN), .ZN(n6917) );
  NOR4_X1 U7848 ( .A1(EAX_REG_21__SCAN_IN), .A2(EAX_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_31__SCAN_IN), .A4(DATAI_24_), .ZN(n6916) );
  NOR4_X1 U7849 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .A4(REIP_REG_10__SCAN_IN), .ZN(n6915) );
  NAND4_X1 U7850 ( .A1(n6918), .A2(n6917), .A3(n6916), .A4(n6915), .ZN(n6919)
         );
  NOR4_X1 U7851 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6921), .A3(n6920), .A4(n6919), 
        .ZN(n6983) );
  NAND4_X1 U7852 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n6981) );
  NAND4_X1 U7853 ( .A1(REIP_REG_21__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        DATAI_14_), .A4(DATAI_27_), .ZN(n6980) );
  NAND4_X1 U7854 ( .A1(EBX_REG_17__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .A4(DATAI_2_), .ZN(n6922) );
  NOR3_X1 U7855 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(ADDRESS_REG_12__SCAN_IN), 
        .A3(n6922), .ZN(n6928) );
  NAND4_X1 U7856 ( .A1(UWORD_REG_4__SCAN_IN), .A2(DATAO_REG_19__SCAN_IN), .A3(
        ADDRESS_REG_22__SCAN_IN), .A4(ADDRESS_REG_19__SCAN_IN), .ZN(n6926) );
  NAND4_X1 U7857 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_14__SCAN_IN), 
        .A3(DATAO_REG_5__SCAN_IN), .A4(ADDRESS_REG_2__SCAN_IN), .ZN(n6925) );
  NAND4_X1 U7858 ( .A1(EAX_REG_17__SCAN_IN), .A2(DATAO_REG_14__SCAN_IN), .A3(
        UWORD_REG_11__SCAN_IN), .A4(UWORD_REG_1__SCAN_IN), .ZN(n6924) );
  NAND4_X1 U7859 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(ADDRESS_REG_16__SCAN_IN), 
        .A3(BE_N_REG_2__SCAN_IN), .A4(DATAO_REG_0__SCAN_IN), .ZN(n6923) );
  NOR4_X1 U7860 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n6927)
         );
  NAND4_X1 U7861 ( .A1(EBX_REG_23__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n6928), .A4(n6927), .ZN(n6979) );
  NAND4_X1 U7862 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(
        INSTQUEUE_REG_5__4__SCAN_IN), .A3(n6929), .A4(n5093), .ZN(n6940) );
  NAND4_X1 U7863 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n6932), .A3(n6931), 
        .A4(n6930), .ZN(n6939) );
  NAND4_X1 U7864 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        INSTQUEUE_REG_8__1__SCAN_IN), .A3(n5078), .A4(n6933), .ZN(n6938) );
  NAND4_X1 U7865 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6936), .A3(n6935), 
        .A4(n6934), .ZN(n6937) );
  NOR4_X1 U7866 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6977)
         );
  NAND4_X1 U7867 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6950)
         );
  NAND4_X1 U7868 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTQUEUE_REG_9__5__SCAN_IN), .A3(n6946), .A4(n6945), .ZN(n6949) );
  NAND4_X1 U7869 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        INSTQUEUE_REG_15__6__SCAN_IN), .A3(INSTQUEUE_REG_14__7__SCAN_IN), .A4(
        n6947), .ZN(n6948) );
  NOR4_X1 U7870 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6976)
         );
  NAND4_X1 U7871 ( .A1(EBX_REG_0__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_11__SCAN_IN), .A4(n6952), .ZN(n6958) );
  NAND4_X1 U7872 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6954), .A4(n6953), .ZN(n6957) );
  NAND4_X1 U7873 ( .A1(EAX_REG_28__SCAN_IN), .A2(DATAI_25_), .A3(DATAI_8_), 
        .A4(DATAI_23_), .ZN(n6956) );
  NAND4_X1 U7874 ( .A1(EAX_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A3(DATAI_21_), .A4(DATAI_4_), .ZN(
        n6955) );
  NOR4_X1 U7875 ( .A1(n6958), .A2(n6957), .A3(n6956), .A4(n6955), .ZN(n6975)
         );
  NAND4_X1 U7876 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6961), .A3(n6960), 
        .A4(n6959), .ZN(n6973) );
  NAND4_X1 U7877 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(
        INSTQUEUE_REG_5__1__SCAN_IN), .A3(n6963), .A4(n6962), .ZN(n6972) );
  NAND4_X1 U7878 ( .A1(EAX_REG_1__SCAN_IN), .A2(n6966), .A3(n6965), .A4(n6964), 
        .ZN(n6971) );
  NAND4_X1 U7879 ( .A1(EAX_REG_5__SCAN_IN), .A2(n6969), .A3(n6968), .A4(n6967), 
        .ZN(n6970) );
  NOR4_X1 U7880 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(n6970), .ZN(n6974)
         );
  NAND4_X1 U7881 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n6978)
         );
  NOR4_X1 U7882 ( .A1(n6981), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n6982)
         );
  NAND4_X1 U7883 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n6986)
         );
  XNOR2_X1 U7884 ( .A(n6987), .B(n6986), .ZN(U2845) );
  OAI22_X1 U4311 ( .A1(n4451), .A2(STATE2_REG_0__SCAN_IN), .B1(n3470), .B2(
        n3510), .ZN(n3406) );
  INV_X1 U3596 ( .A(n5652), .ZN(n5601) );
  NAND2_X1 U3642 ( .A1(n5674), .A2(n3635), .ZN(n3637) );
  CLKBUF_X1 U3638 ( .A(n3468), .Z(n3108) );
  NAND4_X1 U3664 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3317)
         );
  CLKBUF_X1 U3677 ( .A(n5385), .Z(n3097) );
  NAND2_X1 U3864 ( .A1(n5185), .A2(n3153), .ZN(n5262) );
  NAND4_X2 U4125 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3111)
         );
  CLKBUF_X1 U4688 ( .A(n6184), .Z(n6192) );
endmodule

