

module b17_C_gen_AntiSAT_k_256_10 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9800, n9801, n9802, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272;

  OAI21_X1 U11244 ( .B1(n14675), .B2(n14624), .A(n16009), .ZN(n14646) );
  NAND2_X2 U11245 ( .A1(n12688), .A2(n14684), .ZN(n14675) );
  INV_X2 U11246 ( .A(n17001), .ZN(n16975) );
  INV_X1 U11248 ( .A(n10647), .ZN(n10654) );
  INV_X1 U11249 ( .A(n10767), .ZN(n9824) );
  INV_X2 U11250 ( .A(n17161), .ZN(n15694) );
  INV_X1 U11251 ( .A(n9848), .ZN(n17289) );
  INV_X1 U11252 ( .A(n17186), .ZN(n17324) );
  INV_X1 U11253 ( .A(n17304), .ZN(n17327) );
  OR2_X1 U11254 ( .A1(n12917), .A2(n12920), .ZN(n9844) );
  NAND2_X2 U11255 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18828) );
  CLKBUF_X2 U11256 ( .A(n11600), .Z(n12543) );
  CLKBUF_X2 U11257 ( .A(n11583), .Z(n12236) );
  INV_X1 U11258 ( .A(n11616), .ZN(n9812) );
  CLKBUF_X1 U11259 ( .A(n11610), .Z(n11540) );
  AND2_X1 U11260 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15511), .ZN(
        n14255) );
  CLKBUF_X2 U11261 ( .A(n11673), .Z(n12129) );
  AND2_X1 U11262 ( .A1(n13380), .A2(n10005), .ZN(n11599) );
  AND2_X1 U11263 ( .A1(n13382), .A2(n13377), .ZN(n11541) );
  AND2_X1 U11265 ( .A1(n11555), .A2(n12576), .ZN(n10435) );
  INV_X1 U11266 ( .A(n11609), .ZN(n11721) );
  INV_X1 U11267 ( .A(n10767), .ZN(n9823) );
  INV_X1 U11268 ( .A(n14227), .ZN(n11279) );
  INV_X1 U11269 ( .A(n9844), .ZN(n17228) );
  INV_X1 U11270 ( .A(n9850), .ZN(n15735) );
  INV_X2 U11271 ( .A(n9844), .ZN(n17308) );
  INV_X1 U11272 ( .A(n16009), .ZN(n10154) );
  NAND2_X2 U11275 ( .A1(n18999), .A2(n19006), .ZN(n13029) );
  INV_X1 U11276 ( .A(n15607), .ZN(n17287) );
  INV_X1 U11277 ( .A(n12404), .ZN(n13172) );
  NAND3_X1 U11278 ( .A1(n10668), .A2(n10667), .A3(n10666), .ZN(n13278) );
  INV_X1 U11279 ( .A(n17186), .ZN(n17231) );
  INV_X2 U11280 ( .A(n10447), .ZN(n17281) );
  INV_X1 U11281 ( .A(n17968), .ZN(n17988) );
  NOR3_X1 U11282 ( .A1(n16537), .A2(n17902), .A3(n18332), .ZN(n16540) );
  BUF_X1 U11283 ( .A(n13278), .Z(n14305) );
  NOR2_X1 U11284 ( .A1(n17773), .A2(n17808), .ZN(n17968) );
  BUF_X1 U11285 ( .A(n14255), .Z(n9820) );
  AND2_X1 U11287 ( .A1(n10367), .A2(n10775), .ZN(n9800) );
  NAND2_X2 U11288 ( .A1(n12059), .A2(n10437), .ZN(n14377) );
  INV_X2 U11289 ( .A(n14436), .ZN(n12059) );
  NOR2_X2 U11290 ( .A1(n14647), .A2(n12673), .ZN(n13836) );
  NAND2_X2 U11291 ( .A1(n17993), .A2(n17983), .ZN(n17982) );
  NAND2_X1 U11292 ( .A1(n13168), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11095) );
  INV_X2 U11293 ( .A(n9850), .ZN(n17331) );
  NOR2_X2 U11294 ( .A1(n17657), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17656) );
  INV_X2 U11296 ( .A(n10501), .ZN(n9802) );
  INV_X1 U11298 ( .A(n9801), .ZN(n9804) );
  INV_X1 U11299 ( .A(n9801), .ZN(n9805) );
  INV_X1 U11300 ( .A(n9802), .ZN(n9806) );
  INV_X1 U11301 ( .A(n9802), .ZN(n9807) );
  INV_X1 U11302 ( .A(n9802), .ZN(n9808) );
  INV_X1 U11303 ( .A(n9802), .ZN(n9809) );
  AND2_X2 U11304 ( .A1(n10365), .A2(n15503), .ZN(n10501) );
  AOI21_X2 U11305 ( .B1(n13963), .B2(n9994), .A(n9897), .ZN(n9993) );
  XNOR2_X2 U11306 ( .A(n10971), .B(n13973), .ZN(n13963) );
  INV_X1 U11307 ( .A(n14993), .ZN(n9810) );
  OR2_X1 U11308 ( .A1(n17883), .A2(n10113), .ZN(n17850) );
  NAND2_X2 U11309 ( .A1(n13446), .A2(n13484), .ZN(n13483) );
  NOR2_X2 U11310 ( .A1(n18350), .A2(n16651), .ZN(n17986) );
  NOR2_X1 U11311 ( .A1(n15441), .A2(n15440), .ZN(n13647) );
  OR2_X1 U11312 ( .A1(n16384), .A2(n10265), .ZN(n15441) );
  NAND2_X1 U11313 ( .A1(n17909), .A2(n15812), .ZN(n15818) );
  CLKBUF_X1 U11314 ( .A(n13426), .Z(n20586) );
  NAND2_X1 U11315 ( .A1(n11688), .A2(n11687), .ZN(n20364) );
  BUF_X1 U11316 ( .A(n17623), .Z(n17615) );
  OAI21_X1 U11317 ( .B1(n11095), .B2(n10929), .A(n10615), .ZN(n10616) );
  AND2_X1 U11318 ( .A1(n11245), .A2(n13925), .ZN(n9976) );
  INV_X2 U11319 ( .A(n11327), .ZN(n11305) );
  INV_X2 U11320 ( .A(n10184), .ZN(n9816) );
  INV_X4 U11321 ( .A(n19339), .ZN(n11441) );
  NAND2_X1 U11322 ( .A1(n13165), .A2(n11267), .ZN(n10587) );
  OR2_X1 U11323 ( .A1(n12712), .A2(n12327), .ZN(n12737) );
  NAND2_X1 U11324 ( .A1(n13925), .A2(n13291), .ZN(n10366) );
  INV_X1 U11325 ( .A(n11440), .ZN(n19332) );
  INV_X1 U11326 ( .A(n11437), .ZN(n10591) );
  AND2_X2 U11327 ( .A1(n10546), .A2(n10545), .ZN(n14227) );
  OR2_X2 U11328 ( .A1(n11606), .A2(n11605), .ZN(n11616) );
  NAND2_X1 U11329 ( .A1(n11505), .A2(n11504), .ZN(n11610) );
  INV_X2 U11330 ( .A(n17283), .ZN(n15715) );
  BUF_X2 U11331 ( .A(n11592), .Z(n12100) );
  INV_X4 U11332 ( .A(n17317), .ZN(n9811) );
  CLKBUF_X2 U11333 ( .A(n15607), .Z(n9813) );
  INV_X4 U11334 ( .A(n15691), .ZN(n15554) );
  BUF_X2 U11335 ( .A(n11599), .Z(n12083) );
  BUF_X2 U11336 ( .A(n11559), .Z(n12241) );
  BUF_X2 U11337 ( .A(n11541), .Z(n12550) );
  CLKBUF_X2 U11338 ( .A(n11714), .Z(n13379) );
  CLKBUF_X2 U11339 ( .A(n11360), .Z(n14108) );
  CLKBUF_X2 U11340 ( .A(n10715), .Z(n14272) );
  BUF_X2 U11341 ( .A(n10509), .Z(n14264) );
  BUF_X2 U11342 ( .A(n11534), .Z(n12542) );
  INV_X4 U11343 ( .A(n17306), .ZN(n15686) );
  AOI211_X1 U11344 ( .C1(n16043), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14672) );
  OAI21_X1 U11345 ( .B1(n14767), .B2(n20155), .A(n12822), .ZN(n12823) );
  OAI21_X1 U11346 ( .B1(n12442), .B2(n14316), .A(n12255), .ZN(n14629) );
  XNOR2_X1 U11347 ( .A(n12814), .B(n12813), .ZN(n14767) );
  OAI21_X1 U11348 ( .B1(n12814), .B2(n12693), .A(n12692), .ZN(n10012) );
  AOI21_X1 U11349 ( .B1(n12858), .B2(n16391), .A(n12857), .ZN(n12861) );
  NOR2_X1 U11350 ( .A1(n12691), .A2(n12843), .ZN(n12845) );
  OR2_X1 U11351 ( .A1(n12802), .A2(n16356), .ZN(n12810) );
  NAND2_X1 U11352 ( .A1(n12689), .A2(n14769), .ZN(n12691) );
  AND2_X1 U11353 ( .A1(n10127), .A2(n10125), .ZN(n10121) );
  AND2_X1 U11354 ( .A1(n10303), .A2(n10302), .ZN(n10306) );
  NAND2_X1 U11355 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  NAND2_X1 U11356 ( .A1(n14655), .A2(n9961), .ZN(n14635) );
  OR2_X1 U11357 ( .A1(n15422), .A2(n10067), .ZN(n15229) );
  NAND2_X1 U11358 ( .A1(n10039), .A2(n16009), .ZN(n14684) );
  NAND2_X1 U11359 ( .A1(n10145), .A2(n9924), .ZN(n10039) );
  OR2_X1 U11360 ( .A1(n14943), .A2(n10358), .ZN(n14923) );
  NAND2_X1 U11361 ( .A1(n17629), .A2(n17630), .ZN(n17628) );
  AND2_X1 U11362 ( .A1(n10364), .A2(n13868), .ZN(n10859) );
  NOR2_X1 U11363 ( .A1(n13887), .A2(n10417), .ZN(n10416) );
  NAND2_X1 U11364 ( .A1(n10852), .A2(n10334), .ZN(n10961) );
  AND2_X1 U11365 ( .A1(n10863), .A2(n11326), .ZN(n9944) );
  NAND2_X1 U11366 ( .A1(n10827), .A2(n9945), .ZN(n10863) );
  NAND2_X1 U11367 ( .A1(n15008), .A2(n14879), .ZN(n14993) );
  NOR2_X2 U11368 ( .A1(n17689), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17688) );
  NAND2_X1 U11369 ( .A1(n17744), .A2(n10107), .ZN(n17689) );
  NAND2_X1 U11370 ( .A1(n10347), .A2(n10345), .ZN(n13958) );
  NAND2_X1 U11371 ( .A1(n9948), .A2(n10755), .ZN(n10786) );
  XNOR2_X1 U11372 ( .A(n12325), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12892) );
  NAND2_X1 U11373 ( .A1(n12652), .A2(n12602), .ZN(n16008) );
  OR2_X1 U11374 ( .A1(n16265), .A2(n11326), .ZN(n11052) );
  AND3_X1 U11375 ( .A1(n10758), .A2(n9979), .A3(n9978), .ZN(n9980) );
  AND2_X1 U11376 ( .A1(n10150), .A2(n11873), .ZN(n12643) );
  NAND2_X1 U11377 ( .A1(n10025), .A2(n10024), .ZN(n12652) );
  OAI22_X1 U11378 ( .A1(n10692), .A2(n19456), .B1(n19481), .B2(n10691), .ZN(
        n10697) );
  INV_X1 U11379 ( .A(n19419), .ZN(n19422) );
  NAND2_X1 U11380 ( .A1(n13647), .A2(n13648), .ZN(n16367) );
  AND2_X1 U11381 ( .A1(n10705), .A2(n10704), .ZN(n10810) );
  AND2_X1 U11382 ( .A1(n10698), .A2(n10699), .ZN(n10809) );
  AND2_X1 U11383 ( .A1(n10705), .A2(n10693), .ZN(n19606) );
  AND2_X1 U11384 ( .A1(n10703), .A2(n10693), .ZN(n10799) );
  OR2_X1 U11385 ( .A1(n19068), .A2(n11039), .ZN(n15204) );
  AND2_X1 U11386 ( .A1(n10703), .A2(n10704), .ZN(n10803) );
  AND2_X1 U11387 ( .A1(n10698), .A2(n10693), .ZN(n10808) );
  AND2_X1 U11388 ( .A1(n10703), .A2(n10699), .ZN(n10800) );
  AND2_X1 U11389 ( .A1(n10705), .A2(n10702), .ZN(n19663) );
  OAI21_X2 U11390 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19019), .A(n16651), 
        .ZN(n17995) );
  AND2_X1 U11391 ( .A1(n10683), .A2(n10693), .ZN(n19362) );
  AND2_X1 U11392 ( .A1(n10698), .A2(n10704), .ZN(n19511) );
  AND2_X1 U11393 ( .A1(n10703), .A2(n10702), .ZN(n10801) );
  AND2_X1 U11394 ( .A1(n13340), .A2(n14305), .ZN(n10683) );
  NOR2_X1 U11395 ( .A1(n13579), .A2(n14305), .ZN(n10698) );
  NAND2_X1 U11396 ( .A1(n13268), .A2(n13267), .ZN(n16384) );
  NAND2_X1 U11397 ( .A1(n10015), .A2(n11743), .ZN(n11794) );
  NAND2_X1 U11398 ( .A1(n11094), .A2(n11093), .ZN(n10342) );
  NOR2_X2 U11399 ( .A1(n18350), .A2(n18249), .ZN(n18197) );
  CLKBUF_X1 U11400 ( .A(n12593), .Z(n14593) );
  CLKBUF_X1 U11401 ( .A(n14045), .Z(n14595) );
  NAND2_X1 U11402 ( .A1(n13241), .A2(n10454), .ZN(n13268) );
  AND3_X1 U11403 ( .A1(n10017), .A2(n10016), .A3(n10406), .ZN(n10015) );
  OAI211_X1 U11404 ( .C1(n11667), .C2(n10037), .A(n10036), .B(n10034), .ZN(
        n20850) );
  INV_X1 U11405 ( .A(n13164), .ZN(n19208) );
  NAND2_X1 U11406 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  NAND2_X1 U11407 ( .A1(n11091), .A2(n10604), .ZN(n11090) );
  OR2_X1 U11408 ( .A1(n10654), .A2(n10653), .ZN(n10662) );
  AND2_X1 U11409 ( .A1(n11758), .A2(n11760), .ZN(n11686) );
  NOR2_X1 U11410 ( .A1(n11300), .A2(n11299), .ZN(n11309) );
  OAI211_X1 U11411 ( .C1(n10601), .C2(n13577), .A(n10600), .B(n10599), .ZN(
        n10602) );
  NAND2_X1 U11412 ( .A1(n11652), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U11413 ( .A1(n17561), .A2(n14017), .ZN(n16650) );
  AOI21_X1 U11414 ( .B1(n18360), .B2(n13011), .A(n14014), .ZN(n15765) );
  AND4_X1 U11415 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10640) );
  AND2_X2 U11416 ( .A1(n13046), .A2(n13148), .ZN(n13118) );
  AND2_X1 U11417 ( .A1(n10946), .A2(n10945), .ZN(n10958) );
  NAND2_X1 U11418 ( .A1(n15809), .A2(n15808), .ZN(n16533) );
  NOR2_X1 U11419 ( .A1(n15805), .A2(n17501), .ZN(n15809) );
  NAND2_X1 U11420 ( .A1(n11261), .A2(n13150), .ZN(n10638) );
  NOR4_X1 U11421 ( .A1(n18360), .A2(n18365), .A3(n12999), .A4(n15778), .ZN(
        n13012) );
  NAND2_X1 U11422 ( .A1(n10928), .A2(n10927), .ZN(n10953) );
  INV_X1 U11423 ( .A(n9942), .ZN(n9941) );
  NAND2_X1 U11424 ( .A1(n11239), .A2(n9976), .ZN(n11435) );
  AOI21_X1 U11425 ( .B1(n12736), .B2(n13376), .A(n11627), .ZN(n11628) );
  AND2_X1 U11426 ( .A1(n10582), .A2(n11234), .ZN(n11261) );
  NAND2_X1 U11427 ( .A1(n10620), .A2(n12484), .ZN(n16451) );
  NOR2_X1 U11428 ( .A1(n17987), .A2(n16483), .ZN(n16507) );
  NAND2_X1 U11429 ( .A1(n9935), .A2(n9933), .ZN(n15920) );
  CLKBUF_X2 U11430 ( .A(n10587), .Z(n13182) );
  NAND2_X1 U11431 ( .A1(n10493), .A2(n9870), .ZN(n11239) );
  INV_X2 U11432 ( .A(n12717), .ZN(n12718) );
  NOR2_X1 U11433 ( .A1(n11228), .A2(n19863), .ZN(n10624) );
  NAND2_X2 U11434 ( .A1(n10508), .A2(n10507), .ZN(n19339) );
  INV_X2 U11435 ( .A(n14227), .ZN(n14957) );
  INV_X2 U11436 ( .A(n11267), .ZN(n13926) );
  OR2_X1 U11437 ( .A1(n10773), .A2(n10772), .ZN(n11311) );
  NAND2_X2 U11438 ( .A1(n10558), .A2(n10557), .ZN(n16437) );
  INV_X1 U11439 ( .A(n11617), .ZN(n11625) );
  NAND2_X1 U11440 ( .A1(n10570), .A2(n10569), .ZN(n11440) );
  OR2_X2 U11441 ( .A1(n16600), .A2(n16547), .ZN(n16602) );
  INV_X2 U11442 ( .A(U212), .ZN(n16585) );
  NAND2_X1 U11443 ( .A1(n11554), .A2(n11610), .ZN(n11647) );
  AND2_X1 U11444 ( .A1(n11526), .A2(n11522), .ZN(n10413) );
  AND3_X1 U11445 ( .A1(n11524), .A2(n11525), .A3(n11527), .ZN(n10414) );
  AND4_X1 U11446 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11589) );
  AND2_X2 U11447 ( .A1(n9820), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14107) );
  AND4_X1 U11448 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11516) );
  AND4_X1 U11449 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11591) );
  AND4_X1 U11450 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11590) );
  AND4_X1 U11451 ( .A1(n11587), .A2(n11586), .A3(n11585), .A4(n11584), .ZN(
        n11588) );
  AND4_X1 U11452 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11505) );
  AND4_X1 U11453 ( .A1(n11503), .A2(n11502), .A3(n11501), .A4(n11500), .ZN(
        n11504) );
  AND4_X1 U11454 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n9832) );
  AND4_X1 U11455 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(
        n11553) );
  AND4_X1 U11456 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11552) );
  AND4_X1 U11457 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11517) );
  NAND2_X1 U11458 ( .A1(n14276), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10767) );
  INV_X4 U11459 ( .A(n9827), .ZN(n17330) );
  NAND2_X2 U11460 ( .A1(n20005), .A2(n19889), .ZN(n19949) );
  NAND2_X1 U11461 ( .A1(n12912), .A2(n12911), .ZN(n17283) );
  NAND2_X2 U11462 ( .A1(n18966), .A2(n18899), .ZN(n18962) );
  CLKBUF_X1 U11463 ( .A(n13930), .Z(n19313) );
  BUF_X2 U11465 ( .A(n11542), .Z(n12540) );
  AND2_X2 U11466 ( .A1(n12815), .A2(n20703), .ZN(n20149) );
  INV_X2 U11467 ( .A(n16641), .ZN(n16643) );
  AND2_X2 U11468 ( .A1(n14254), .A2(n16411), .ZN(n10734) );
  CLKBUF_X3 U11469 ( .A(n11598), .Z(n12105) );
  OR2_X1 U11470 ( .A1(n12917), .A2(n18828), .ZN(n10447) );
  NAND2_X2 U11471 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12916), .ZN(
        n17161) );
  AND2_X2 U11472 ( .A1(n13334), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11487) );
  AND2_X1 U11473 ( .A1(n11480), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10005) );
  AND2_X2 U11474 ( .A1(n13397), .A2(n11488), .ZN(n11673) );
  AND2_X1 U11475 ( .A1(n18817), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n18824) );
  AND3_X1 U11476 ( .A1(n15503), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10520) );
  AND2_X1 U11477 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11488) );
  NOR2_X2 U11478 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11486) );
  AND2_X2 U11479 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13377) );
  INV_X1 U11480 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13334) );
  CLKBUF_X1 U11481 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15529) );
  INV_X1 U11482 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15503) );
  XOR2_X2 U11483 ( .A(n12722), .B(n12721), .Z(n14504) );
  MUX2_X2 U11484 ( .A(n12865), .B(n13172), .S(n12863), .Z(n12721) );
  OR3_X2 U11485 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n12920), .ZN(n9827) );
  NAND2_X1 U11486 ( .A1(n19006), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12920) );
  AND2_X1 U11487 ( .A1(n10980), .A2(n10978), .ZN(n10976) );
  NOR2_X2 U11488 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  NAND2_X2 U11489 ( .A1(n13594), .A2(n9839), .ZN(n13479) );
  INV_X1 U11490 ( .A(n11138), .ZN(n9814) );
  INV_X1 U11491 ( .A(n9814), .ZN(n9815) );
  INV_X4 U11492 ( .A(n15688), .ZN(n15714) );
  NOR2_X2 U11493 ( .A1(n13808), .A2(n13807), .ZN(n13907) );
  NOR2_X2 U11494 ( .A1(n18985), .A2(n17989), .ZN(n17808) );
  NAND2_X2 U11495 ( .A1(n13955), .A2(n13956), .ZN(n14049) );
  AND2_X2 U11496 ( .A1(n13907), .A2(n13906), .ZN(n13955) );
  AOI21_X2 U11497 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n15027) );
  INV_X2 U11498 ( .A(n10184), .ZN(n12413) );
  NAND2_X4 U11499 ( .A1(n10434), .A2(n11626), .ZN(n10184) );
  XNOR2_X2 U11500 ( .A(n10647), .B(n10653), .ZN(n10669) );
  XNOR2_X2 U11501 ( .A(n14138), .B(n10465), .ZN(n14968) );
  AND2_X1 U11502 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15511), .ZN(
        n9817) );
  AND2_X1 U11503 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15511), .ZN(
        n9818) );
  INV_X1 U11504 ( .A(n14255), .ZN(n9819) );
  INV_X1 U11505 ( .A(n9819), .ZN(n9821) );
  INV_X1 U11506 ( .A(n9819), .ZN(n9822) );
  NAND2_X1 U11507 ( .A1(n12263), .A2(n12262), .ZN(n12268) );
  XNOR2_X1 U11508 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12267) );
  NAND2_X2 U11509 ( .A1(n11279), .A2(n16437), .ZN(n11228) );
  INV_X1 U11510 ( .A(n10863), .ZN(n10887) );
  NAND2_X1 U11511 ( .A1(n13867), .A2(n13866), .ZN(n10042) );
  AND2_X1 U11512 ( .A1(n15882), .A2(n12705), .ZN(n13224) );
  NAND2_X1 U11513 ( .A1(n10059), .A2(n10058), .ZN(n16298) );
  AOI21_X1 U11514 ( .B1(n10060), .B2(n15437), .A(n11199), .ZN(n10058) );
  NAND3_X1 U11515 ( .A1(n10055), .A2(n10053), .A3(n10052), .ZN(n11198) );
  NOR2_X1 U11516 ( .A1(n16358), .A2(n10054), .ZN(n10053) );
  INV_X1 U11517 ( .A(n10057), .ZN(n10054) );
  NOR2_X1 U11518 ( .A1(n18371), .A2(n9849), .ZN(n13000) );
  BUF_X1 U11519 ( .A(n12549), .Z(n12204) );
  BUF_X1 U11520 ( .A(n11673), .Z(n12551) );
  CLKBUF_X2 U11521 ( .A(n11703), .Z(n12548) );
  INV_X1 U11522 ( .A(n11682), .ZN(n12619) );
  AND2_X1 U11523 ( .A1(n11721), .A2(n12671), .ZN(n11729) );
  OR2_X1 U11524 ( .A1(n11780), .A2(n12671), .ZN(n11736) );
  NOR2_X1 U11525 ( .A1(n10423), .A2(n10424), .ZN(n10422) );
  INV_X1 U11526 ( .A(n11680), .ZN(n10423) );
  OR2_X1 U11527 ( .A1(n12258), .A2(n12421), .ZN(n11648) );
  NAND2_X1 U11528 ( .A1(n11792), .A2(n11793), .ZN(n11829) );
  AND2_X2 U11529 ( .A1(n11481), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13380) );
  INV_X1 U11530 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11481) );
  INV_X1 U11531 ( .A(n12303), .ZN(n12295) );
  NAND2_X1 U11532 ( .A1(n10852), .A2(n10855), .ZN(n10853) );
  NAND3_X1 U11533 ( .A1(n9800), .A2(n9947), .A3(n10905), .ZN(n9998) );
  INV_X1 U11534 ( .A(n10786), .ZN(n9947) );
  AND2_X1 U11535 ( .A1(n14337), .A2(n9903), .ZN(n12838) );
  INV_X1 U11536 ( .A(n12254), .ZN(n10442) );
  NOR2_X1 U11537 ( .A1(n12441), .A2(n10445), .ZN(n10444) );
  NAND2_X1 U11538 ( .A1(n10441), .A2(n14411), .ZN(n10440) );
  NOR2_X1 U11539 ( .A1(n14424), .A2(n14439), .ZN(n10441) );
  NAND2_X1 U11540 ( .A1(n10427), .A2(n14453), .ZN(n10426) );
  AND2_X1 U11541 ( .A1(n10429), .A2(n11900), .ZN(n10428) );
  INV_X1 U11542 ( .A(n13864), .ZN(n10429) );
  NAND2_X1 U11543 ( .A1(n14044), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12249) );
  INV_X1 U11544 ( .A(n11991), .ZN(n11951) );
  NOR2_X2 U11545 ( .A1(n11540), .A2(n20189), .ZN(n11991) );
  NAND2_X1 U11546 ( .A1(n10415), .A2(n14646), .ZN(n10028) );
  AND2_X1 U11547 ( .A1(n14635), .A2(n14768), .ZN(n10415) );
  NAND2_X1 U11548 ( .A1(n14683), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U11549 ( .A1(n9960), .A2(n10192), .ZN(n10020) );
  INV_X1 U11550 ( .A(n10027), .ZN(n9960) );
  NAND2_X1 U11551 ( .A1(n16042), .A2(n16041), .ZN(n10033) );
  NAND2_X1 U11552 ( .A1(n12718), .A2(n12404), .ZN(n12403) );
  NAND2_X1 U11553 ( .A1(n10146), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11659) );
  AOI21_X1 U11554 ( .B1(n12268), .B2(n12267), .A(n12264), .ZN(n12299) );
  AND2_X1 U11555 ( .A1(n14204), .A2(n14203), .ZN(n14205) );
  INV_X1 U11556 ( .A(n11041), .ZN(n10143) );
  INV_X1 U11557 ( .A(n15065), .ZN(n10279) );
  AND2_X1 U11558 ( .A1(n9892), .A2(n14884), .ZN(n10263) );
  NAND2_X1 U11559 ( .A1(n9963), .A2(n10372), .ZN(n10041) );
  AND3_X1 U11560 ( .A1(n10368), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n13979), .ZN(n10372) );
  NAND2_X1 U11561 ( .A1(n13289), .A2(n13288), .ZN(n13293) );
  NOR3_X1 U11562 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n19006), .ZN(n12916) );
  NAND2_X1 U11563 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18981), .ZN(
        n12921) );
  OR2_X1 U11564 ( .A1(n15882), .A2(n14306), .ZN(n13322) );
  INV_X1 U11565 ( .A(n11554), .ZN(n14044) );
  NAND2_X1 U11566 ( .A1(n13838), .A2(n12674), .ZN(n12677) );
  AND2_X1 U11567 ( .A1(n10029), .A2(n10028), .ZN(n12814) );
  NAND2_X1 U11568 ( .A1(n12691), .A2(n10154), .ZN(n10029) );
  OR2_X1 U11569 ( .A1(n14317), .A2(n12417), .ZN(n12863) );
  NAND2_X1 U11570 ( .A1(n14319), .A2(n14318), .ZN(n14317) );
  NAND2_X1 U11571 ( .A1(n14646), .A2(n14635), .ZN(n12689) );
  NAND2_X1 U11572 ( .A1(n12711), .A2(n12710), .ZN(n12743) );
  OAI22_X1 U11573 ( .A1(n20000), .A2(n11474), .B1(n19998), .B2(n10923), .ZN(
        n11251) );
  NAND2_X1 U11574 ( .A1(n13532), .A2(n10320), .ZN(n13808) );
  AND2_X1 U11575 ( .A1(n9891), .A2(n13724), .ZN(n10320) );
  OR2_X1 U11576 ( .A1(n10268), .A2(n13476), .ZN(n10267) );
  NAND2_X1 U11577 ( .A1(n10539), .A2(n16411), .ZN(n10546) );
  XNOR2_X1 U11578 ( .A(n11086), .B(n11085), .ZN(n12488) );
  NAND2_X1 U11579 ( .A1(n12485), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11086) );
  OR2_X1 U11580 ( .A1(n10275), .A2(n10274), .ZN(n10270) );
  NAND2_X1 U11581 ( .A1(n15127), .A2(n15125), .ZN(n12454) );
  AND2_X1 U11582 ( .A1(n15154), .A2(n10383), .ZN(n15121) );
  AND2_X1 U11583 ( .A1(n10384), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10383) );
  NOR2_X1 U11584 ( .A1(n15262), .A2(n10385), .ZN(n10384) );
  INV_X1 U11585 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U11586 ( .A1(n15449), .A2(n15454), .ZN(n9996) );
  AND2_X1 U11587 ( .A1(n11475), .A2(n16433), .ZN(n15381) );
  AOI21_X1 U11588 ( .B1(n13222), .B2(n13284), .A(n13221), .ZN(n13271) );
  INV_X1 U11589 ( .A(n13277), .ZN(n13284) );
  NAND2_X1 U11590 ( .A1(n11252), .A2(n11233), .ZN(n16432) );
  INV_X1 U11591 ( .A(n9846), .ZN(n17326) );
  NOR2_X1 U11592 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12912) );
  INV_X1 U11593 ( .A(n13029), .ZN(n12911) );
  NOR2_X1 U11594 ( .A1(n17674), .A2(n18006), .ZN(n18009) );
  INV_X1 U11595 ( .A(n19025), .ZN(n18350) );
  INV_X1 U11596 ( .A(n14602), .ZN(n14618) );
  AND2_X1 U11597 ( .A1(n11198), .A2(n9880), .ZN(n10122) );
  NAND2_X1 U11598 ( .A1(n11842), .A2(n11841), .ZN(n11844) );
  OR2_X1 U11599 ( .A1(n12295), .A2(n11830), .ZN(n11842) );
  OR2_X1 U11600 ( .A1(n11698), .A2(n11697), .ZN(n12606) );
  NAND2_X1 U11601 ( .A1(n11680), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10421) );
  OR2_X1 U11602 ( .A1(n12619), .A2(n11780), .ZN(n11680) );
  NAND2_X1 U11603 ( .A1(n11637), .A2(n14846), .ZN(n11623) );
  NAND2_X1 U11604 ( .A1(n9863), .A2(n9830), .ZN(n9997) );
  INV_X1 U11605 ( .A(n9998), .ZN(n10827) );
  NAND2_X1 U11606 ( .A1(n10808), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n9984) );
  OR2_X1 U11607 ( .A1(n19570), .A2(n9977), .ZN(n9986) );
  INV_X1 U11608 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U11609 ( .A1(n19606), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n9985) );
  NAND2_X1 U11610 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9988) );
  NAND2_X1 U11611 ( .A1(n10800), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9989) );
  NAND2_X1 U11612 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9990) );
  BUF_X1 U11613 ( .A(n11593), .Z(n12199) );
  AND2_X1 U11614 ( .A1(n11866), .A2(n11865), .ZN(n11872) );
  NAND2_X1 U11615 ( .A1(n20204), .A2(n11625), .ZN(n11620) );
  OR2_X1 U11616 ( .A1(n11815), .A2(n11814), .ZN(n12645) );
  NAND2_X1 U11617 ( .A1(n11616), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10196) );
  AND3_X1 U11618 ( .A1(n11624), .A2(n10435), .A3(n10436), .ZN(n12736) );
  OR2_X1 U11619 ( .A1(n12285), .A2(n9812), .ZN(n12301) );
  NOR2_X1 U11620 ( .A1(n10902), .A2(n10901), .ZN(n10904) );
  NAND2_X1 U11621 ( .A1(n10827), .A2(n10826), .ZN(n10852) );
  AND2_X1 U11622 ( .A1(n10660), .A2(n11089), .ZN(n10644) );
  OR2_X1 U11623 ( .A1(n10660), .A2(n11089), .ZN(n10643) );
  AND4_X1 U11624 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10883) );
  NAND2_X1 U11625 ( .A1(n14957), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13215) );
  NAND2_X1 U11626 ( .A1(n10597), .A2(n10591), .ZN(n10533) );
  AOI21_X1 U11627 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19966), .A(
        n10904), .ZN(n10908) );
  INV_X1 U11628 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16412) );
  INV_X1 U11629 ( .A(n15811), .ZN(n15810) );
  AND2_X1 U11630 ( .A1(n15790), .A2(n17510), .ZN(n15788) );
  INV_X1 U11631 ( .A(n17510), .ZN(n15789) );
  AND2_X1 U11632 ( .A1(n10112), .A2(n17514), .ZN(n15790) );
  INV_X1 U11633 ( .A(n12988), .ZN(n10255) );
  INV_X1 U11634 ( .A(n12986), .ZN(n10250) );
  AND2_X1 U11635 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  NAND3_X1 U11636 ( .A1(n10007), .A2(n10006), .A3(n11627), .ZN(n12258) );
  INV_X1 U11637 ( .A(n11876), .ZN(n11877) );
  INV_X1 U11638 ( .A(n12652), .ZN(n12600) );
  INV_X1 U11639 ( .A(n12251), .ZN(n12563) );
  NOR2_X1 U11640 ( .A1(n14465), .A2(n9888), .ZN(n10427) );
  NOR2_X1 U11641 ( .A1(n10090), .A2(n14370), .ZN(n10089) );
  INV_X1 U11642 ( .A(n14385), .ZN(n10090) );
  INV_X1 U11643 ( .A(n10173), .ZN(n10172) );
  NOR2_X1 U11644 ( .A1(n14801), .A2(n14815), .ZN(n10419) );
  AND2_X1 U11645 ( .A1(n16025), .A2(n10187), .ZN(n10027) );
  NOR2_X1 U11646 ( .A1(n10155), .A2(n12679), .ZN(n10187) );
  AND2_X1 U11647 ( .A1(n12687), .A2(n10461), .ZN(n10192) );
  AOI21_X1 U11648 ( .B1(n10155), .B2(n12678), .A(n10154), .ZN(n10153) );
  AND2_X1 U11649 ( .A1(n11729), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12601) );
  INV_X1 U11650 ( .A(n10181), .ZN(n10180) );
  INV_X1 U11651 ( .A(n10179), .ZN(n10178) );
  OR2_X1 U11652 ( .A1(n11720), .A2(n11719), .ZN(n12671) );
  INV_X1 U11653 ( .A(n10175), .ZN(n10174) );
  INV_X1 U11654 ( .A(n10177), .ZN(n10176) );
  INV_X1 U11655 ( .A(n12341), .ZN(n12405) );
  OAI21_X1 U11656 ( .B1(n20180), .B2(n12618), .A(n12604), .ZN(n12630) );
  OR2_X1 U11657 ( .A1(n12404), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U11658 ( .A1(n11616), .A2(n20204), .ZN(n12327) );
  OR2_X1 U11659 ( .A1(n11709), .A2(n11708), .ZN(n12610) );
  INV_X1 U11660 ( .A(n10407), .ZN(n10406) );
  AOI21_X1 U11661 ( .B1(n12605), .B2(n11751), .A(n11741), .ZN(n11743) );
  NAND2_X1 U11662 ( .A1(n10151), .A2(n11791), .ZN(n11792) );
  NAND2_X1 U11663 ( .A1(n20850), .A2(n16196), .ZN(n10151) );
  NAND2_X1 U11664 ( .A1(n10026), .A2(n11829), .ZN(n20180) );
  NAND2_X1 U11665 ( .A1(n20334), .A2(n11794), .ZN(n10026) );
  NOR2_X1 U11666 ( .A1(n20460), .A2(n20459), .ZN(n20554) );
  AOI22_X1 U11667 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U11668 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11563) );
  AND2_X1 U11669 ( .A1(n11681), .A2(n11609), .ZN(n12303) );
  NOR2_X1 U11670 ( .A1(n12696), .A2(n16196), .ZN(n11681) );
  NAND2_X1 U11671 ( .A1(n11721), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11780) );
  OR2_X1 U11672 ( .A1(n10754), .A2(n10753), .ZN(n11302) );
  NOR2_X1 U11673 ( .A1(n10293), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10292) );
  INV_X1 U11674 ( .A(n10294), .ZN(n10293) );
  NOR2_X1 U11675 ( .A1(n10935), .A2(n10297), .ZN(n10296) );
  INV_X1 U11676 ( .A(n11007), .ZN(n10297) );
  NAND2_X1 U11677 ( .A1(n11013), .A2(n11011), .ZN(n11008) );
  OR2_X1 U11678 ( .A1(n11025), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11013) );
  NOR2_X1 U11679 ( .A1(n10968), .A2(n10967), .ZN(n10980) );
  OR2_X1 U11680 ( .A1(n10963), .A2(n10962), .ZN(n10968) );
  NOR2_X1 U11681 ( .A1(n10953), .A2(n10954), .ZN(n10946) );
  NAND2_X1 U11682 ( .A1(n10269), .A2(n13443), .ZN(n10268) );
  INV_X1 U11683 ( .A(n16385), .ZN(n10269) );
  AND2_X2 U11684 ( .A1(n10581), .A2(n10580), .ZN(n10620) );
  AND2_X1 U11685 ( .A1(n14227), .A2(n16437), .ZN(n12484) );
  NOR2_X1 U11686 ( .A1(n9913), .A2(n14932), .ZN(n10360) );
  INV_X1 U11687 ( .A(n14924), .ZN(n10361) );
  NAND2_X1 U11688 ( .A1(n10354), .A2(n10353), .ZN(n10352) );
  INV_X1 U11689 ( .A(n13606), .ZN(n10353) );
  INV_X1 U11690 ( .A(n10355), .ZN(n10354) );
  NOR2_X1 U11691 ( .A1(n11092), .A2(n10341), .ZN(n10340) );
  INV_X1 U11692 ( .A(n13663), .ZN(n10341) );
  AND2_X1 U11693 ( .A1(n10275), .A2(n10274), .ZN(n10272) );
  NAND2_X1 U11694 ( .A1(n16242), .A2(n11078), .ZN(n11059) );
  AND2_X1 U11695 ( .A1(n10460), .A2(n10333), .ZN(n10332) );
  NAND2_X1 U11696 ( .A1(n15437), .A2(n15435), .ZN(n10333) );
  NAND2_X1 U11697 ( .A1(n15243), .A2(n11205), .ZN(n10079) );
  AOI21_X1 U11698 ( .B1(n10076), .B2(n10077), .A(n10075), .ZN(n10074) );
  INV_X1 U11699 ( .A(n11208), .ZN(n10075) );
  INV_X1 U11700 ( .A(n10080), .ZN(n10076) );
  NAND2_X1 U11701 ( .A1(n11203), .A2(n15251), .ZN(n10072) );
  INV_X1 U11702 ( .A(n13922), .ZN(n10264) );
  NOR2_X1 U11703 ( .A1(n13725), .A2(n10349), .ZN(n10348) );
  INV_X1 U11704 ( .A(n13803), .ZN(n10349) );
  NAND2_X1 U11705 ( .A1(n10972), .A2(n9894), .ZN(n10323) );
  NAND2_X1 U11706 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  INV_X1 U11707 ( .A(n13298), .ZN(n10339) );
  NAND2_X1 U11708 ( .A1(n10971), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10972) );
  OR2_X1 U11709 ( .A1(n10838), .A2(n10837), .ZN(n10851) );
  OAI21_X1 U11710 ( .B1(n10961), .B2(n11078), .A(n13795), .ZN(n10965) );
  AND2_X1 U11711 ( .A1(n13570), .A2(n9898), .ZN(n10050) );
  INV_X1 U11712 ( .A(n10050), .ZN(n10047) );
  INV_X1 U11713 ( .A(n10048), .ZN(n10046) );
  INV_X1 U11714 ( .A(n11088), .ZN(n9938) );
  INV_X1 U11715 ( .A(n10643), .ZN(n10614) );
  NAND2_X1 U11716 ( .A1(n10774), .A2(n9992), .ZN(n10775) );
  NAND2_X1 U11717 ( .A1(n10672), .A2(n10671), .ZN(n10674) );
  NOR2_X2 U11718 ( .A1(n10590), .A2(n10589), .ZN(n11260) );
  MUX2_X1 U11719 ( .A(n10588), .B(n10587), .S(n11437), .Z(n10589) );
  NAND2_X1 U11720 ( .A1(n10683), .A2(n10704), .ZN(n10678) );
  AND2_X1 U11721 ( .A1(n14305), .A2(n13579), .ZN(n10705) );
  AND2_X1 U11722 ( .A1(n13222), .A2(n19208), .ZN(n10704) );
  AND2_X1 U11723 ( .A1(n15526), .A2(n13579), .ZN(n10703) );
  NAND2_X1 U11724 ( .A1(n13014), .A2(n18834), .ZN(n14024) );
  NAND2_X1 U11725 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18992), .ZN(
        n12917) );
  OAI21_X1 U11726 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15914) );
  NOR2_X1 U11727 ( .A1(n17656), .A2(n15826), .ZN(n15827) );
  OR2_X1 U11728 ( .A1(n15825), .A2(n15824), .ZN(n15826) );
  NAND2_X1 U11729 ( .A1(n15827), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16532) );
  NOR2_X1 U11730 ( .A1(n15818), .A2(n17793), .ZN(n15816) );
  INV_X1 U11731 ( .A(n15757), .ZN(n15761) );
  AND2_X1 U11732 ( .A1(n9930), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15757) );
  NAND2_X1 U11733 ( .A1(n15810), .A2(n9969), .ZN(n10390) );
  INV_X1 U11734 ( .A(n15807), .ZN(n9969) );
  INV_X1 U11735 ( .A(n17514), .ZN(n15791) );
  NAND2_X1 U11736 ( .A1(n10112), .A2(n15920), .ZN(n15747) );
  NOR2_X1 U11737 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19006), .ZN(
        n14018) );
  NOR2_X1 U11738 ( .A1(n18355), .A2(n18360), .ZN(n18821) );
  NAND3_X1 U11739 ( .A1(n18806), .A2(n19026), .A3(n14024), .ZN(n15917) );
  NAND2_X1 U11740 ( .A1(n18384), .A2(n18360), .ZN(n15764) );
  INV_X1 U11741 ( .A(n13779), .ZN(n12424) );
  OR2_X1 U11742 ( .A1(n20030), .A2(n20189), .ZN(n13779) );
  OR2_X1 U11743 ( .A1(n11616), .A2(n12696), .ZN(n13541) );
  INV_X1 U11744 ( .A(n12249), .ZN(n12569) );
  AND2_X1 U11745 ( .A1(n20189), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12568) );
  NOR2_X1 U11746 ( .A1(n10440), .A2(n10438), .ZN(n10437) );
  INV_X1 U11747 ( .A(n14394), .ZN(n10438) );
  NAND2_X1 U11748 ( .A1(n14730), .A2(n10192), .ZN(n10021) );
  CLKBUF_X1 U11749 ( .A(n14531), .Z(n14532) );
  AND2_X1 U11750 ( .A1(n11901), .A2(n9841), .ZN(n10431) );
  NAND2_X1 U11751 ( .A1(n11867), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11878) );
  NAND2_X1 U11752 ( .A1(n11852), .A2(n11851), .ZN(n13561) );
  INV_X1 U11753 ( .A(n11850), .ZN(n11851) );
  NAND2_X1 U11754 ( .A1(n12643), .A2(n11991), .ZN(n11852) );
  CLKBUF_X1 U11755 ( .A(n13559), .Z(n13560) );
  NAND2_X1 U11756 ( .A1(n11823), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11847) );
  CLKBUF_X1 U11757 ( .A(n13458), .Z(n13459) );
  INV_X1 U11758 ( .A(n13262), .ZN(n11772) );
  NOR2_X2 U11759 ( .A1(n14360), .A2(n12411), .ZN(n14319) );
  NAND2_X1 U11760 ( .A1(n9962), .A2(n10013), .ZN(n9961) );
  NAND2_X1 U11761 ( .A1(n10014), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10013) );
  NAND2_X1 U11762 ( .A1(n12400), .A2(n10182), .ZN(n12401) );
  INV_X1 U11763 ( .A(n14720), .ZN(n10145) );
  NOR2_X1 U11764 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14743) );
  NAND2_X1 U11765 ( .A1(n12677), .A2(n10416), .ZN(n16025) );
  NAND2_X1 U11766 ( .A1(n9957), .A2(n16034), .ZN(n13838) );
  NAND2_X1 U11767 ( .A1(n9959), .A2(n12659), .ZN(n9958) );
  NOR2_X1 U11768 ( .A1(n12355), .A2(n16170), .ZN(n10093) );
  NAND2_X1 U11769 ( .A1(n10033), .A2(n12650), .ZN(n13620) );
  NAND2_X1 U11770 ( .A1(n12642), .A2(n12641), .ZN(n16042) );
  NAND2_X1 U11771 ( .A1(n12629), .A2(n12628), .ZN(n13463) );
  INV_X1 U11772 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10198) );
  XNOR2_X1 U11773 ( .A(n11740), .B(n11738), .ZN(n11751) );
  AND2_X1 U11774 ( .A1(n13333), .A2(n13332), .ZN(n15852) );
  INV_X1 U11775 ( .A(n20586), .ZN(n20660) );
  OR2_X1 U11776 ( .A1(n20456), .A2(n20334), .ZN(n20709) );
  AOI21_X1 U11777 ( .B1(n12299), .B2(n12266), .A(n12298), .ZN(n12319) );
  NAND2_X1 U11778 ( .A1(n11780), .A2(n11779), .ZN(n12274) );
  OAI21_X1 U11779 ( .B1(n11302), .B2(n11228), .A(n10282), .ZN(n10926) );
  NAND2_X1 U11780 ( .A1(n11228), .A2(n11223), .ZN(n10282) );
  INV_X1 U11781 ( .A(n16430), .ZN(n9943) );
  INV_X1 U11782 ( .A(n11228), .ZN(n11259) );
  NOR2_X1 U11783 ( .A1(n11046), .A2(n10283), .ZN(n10940) );
  OR3_X1 U11784 ( .A1(n10938), .A2(P2_EBX_REG_24__SCAN_IN), .A3(
        P2_EBX_REG_25__SCAN_IN), .ZN(n10283) );
  AND2_X1 U11785 ( .A1(n11056), .A2(n11011), .ZN(n11077) );
  AND2_X1 U11786 ( .A1(n12515), .A2(n10212), .ZN(n12495) );
  AND2_X1 U11787 ( .A1(n9840), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10212) );
  INV_X1 U11788 ( .A(n16272), .ZN(n10203) );
  OR2_X1 U11789 ( .A1(n11046), .A2(n10938), .ZN(n11050) );
  INV_X1 U11790 ( .A(n13674), .ZN(n11132) );
  NAND2_X1 U11791 ( .A1(n11011), .A2(n10992), .ZN(n19124) );
  NOR2_X1 U11792 ( .A1(n13633), .A2(n13530), .ZN(n10321) );
  OR2_X1 U11793 ( .A1(n13632), .A2(n13631), .ZN(n13633) );
  NAND2_X1 U11794 ( .A1(n10303), .A2(n9910), .ZN(n10299) );
  NAND2_X1 U11795 ( .A1(n10316), .A2(n14081), .ZN(n10315) );
  INV_X1 U11796 ( .A(n10318), .ZN(n10316) );
  AND3_X1 U11797 ( .A1(n11355), .A2(n11354), .A3(n11353), .ZN(n13476) );
  NOR2_X1 U11798 ( .A1(n12516), .A2(n15219), .ZN(n12515) );
  AND2_X1 U11799 ( .A1(n15006), .A2(n15005), .ZN(n15008) );
  NAND2_X1 U11800 ( .A1(n12513), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12516) );
  NOR2_X1 U11801 ( .A1(n10380), .A2(n15423), .ZN(n10379) );
  AND2_X1 U11802 ( .A1(n11200), .A2(n15435), .ZN(n10060) );
  INV_X1 U11803 ( .A(n13579), .ZN(n13340) );
  NAND2_X1 U11804 ( .A1(n19863), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13277) );
  NOR2_X1 U11805 ( .A1(n11053), .A2(n15153), .ZN(n12769) );
  AND2_X1 U11806 ( .A1(n12766), .A2(n10327), .ZN(n15137) );
  AOI21_X1 U11807 ( .B1(n15153), .B2(n10329), .A(n10328), .ZN(n10327) );
  NAND2_X1 U11808 ( .A1(n15439), .A2(n15435), .ZN(n10331) );
  AOI21_X1 U11809 ( .B1(n10141), .B2(n10143), .A(n9874), .ZN(n10139) );
  INV_X1 U11810 ( .A(n15311), .ZN(n10277) );
  NAND2_X1 U11811 ( .A1(n15177), .A2(n15186), .ZN(n9951) );
  NAND2_X1 U11812 ( .A1(n15084), .A2(n9905), .ZN(n15310) );
  AND2_X1 U11813 ( .A1(n11424), .A2(n11423), .ZN(n15102) );
  NOR2_X2 U11814 ( .A1(n13958), .A2(n13957), .ZN(n15006) );
  INV_X1 U11815 ( .A(n15229), .ZN(n15382) );
  NAND2_X1 U11816 ( .A1(n10069), .A2(n15251), .ZN(n15244) );
  INV_X1 U11817 ( .A(n15452), .ZN(n15424) );
  OR2_X1 U11818 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  INV_X1 U11819 ( .A(n13538), .ZN(n10266) );
  AND2_X1 U11820 ( .A1(n16410), .A2(n13213), .ZN(n15452) );
  NAND2_X1 U11821 ( .A1(n10323), .A2(n10989), .ZN(n10322) );
  OAI21_X1 U11822 ( .B1(n9995), .B2(n10042), .A(n9993), .ZN(n10138) );
  NAND2_X1 U11823 ( .A1(n13963), .A2(n10989), .ZN(n9995) );
  XNOR2_X1 U11824 ( .A(n10886), .B(n10984), .ZN(n16344) );
  NAND2_X1 U11825 ( .A1(n13962), .A2(n9847), .ZN(n9963) );
  INV_X1 U11826 ( .A(n13980), .ZN(n10373) );
  OAI21_X1 U11827 ( .B1(n13657), .B2(n13658), .A(n10960), .ZN(n13867) );
  OAI21_X1 U11828 ( .B1(n10798), .B2(n13873), .A(n9966), .ZN(n10364) );
  NAND2_X1 U11829 ( .A1(n10260), .A2(n9914), .ZN(n13590) );
  INV_X1 U11830 ( .A(n11310), .ZN(n10256) );
  NAND2_X1 U11831 ( .A1(n10948), .A2(n13713), .ZN(n10051) );
  NOR2_X1 U11832 ( .A1(n10049), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10048) );
  INV_X1 U11833 ( .A(n13713), .ZN(n10049) );
  AND2_X1 U11834 ( .A1(n11258), .A2(n19866), .ZN(n11475) );
  NAND2_X1 U11835 ( .A1(n13160), .A2(n19809), .ZN(n13287) );
  NAND2_X1 U11836 ( .A1(n10705), .A2(n10699), .ZN(n19570) );
  INV_X1 U11837 ( .A(n19570), .ZN(n10757) );
  OR2_X1 U11838 ( .A1(n19448), .A2(n19981), .ZN(n19601) );
  OR2_X1 U11839 ( .A1(n19448), .A2(n19447), .ZN(n19669) );
  NAND2_X1 U11840 ( .A1(n19448), .A2(n19447), .ZN(n19726) );
  AND2_X1 U11841 ( .A1(n15913), .A2(n19863), .ZN(n19807) );
  INV_X1 U11842 ( .A(n19807), .ZN(n19546) );
  INV_X1 U11843 ( .A(n15776), .ZN(n18806) );
  OAI21_X1 U11844 ( .B1(n16714), .B2(n10232), .A(n10231), .ZN(n16699) );
  NAND2_X1 U11845 ( .A1(n10233), .A2(n17638), .ZN(n10232) );
  OR2_X1 U11846 ( .A1(n10229), .A2(n16701), .ZN(n10231) );
  INV_X1 U11847 ( .A(n16701), .ZN(n10233) );
  NOR2_X1 U11848 ( .A1(n16723), .A2(n16975), .ZN(n16714) );
  OR2_X1 U11849 ( .A1(n16714), .A2(n16715), .ZN(n10234) );
  AOI21_X1 U11850 ( .B1(n10229), .B2(n17738), .A(n17727), .ZN(n10228) );
  NAND4_X1 U11851 ( .A1(n19020), .A2(n18350), .A3(n18345), .A4(n15914), .ZN(
        n15552) );
  OR2_X2 U11852 ( .A1(n12917), .A2(n13029), .ZN(n17304) );
  NOR3_X1 U11853 ( .A1(n18981), .A2(n18992), .A3(n13029), .ZN(n12913) );
  OR3_X1 U11854 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18828), .ZN(n15688) );
  AOI211_X1 U11855 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15681), .B(n15680), .ZN(n15682) );
  AND2_X1 U11856 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10110) );
  NAND2_X1 U11857 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10401) );
  AND2_X1 U11858 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n9934) );
  INV_X1 U11859 ( .A(n17671), .ZN(n10240) );
  NOR2_X1 U11860 ( .A1(n17737), .A2(n17736), .ZN(n17710) );
  NOR2_X1 U11861 ( .A1(n10237), .A2(n10236), .ZN(n17751) );
  NAND2_X1 U11862 ( .A1(n9828), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10236) );
  NOR3_X1 U11863 ( .A1(n16924), .A2(n17864), .A3(n16909), .ZN(n17831) );
  NOR2_X1 U11864 ( .A1(n16678), .A2(n17929), .ZN(n17894) );
  OR2_X1 U11865 ( .A1(n17945), .A2(n15753), .ZN(n9937) );
  NOR2_X1 U11866 ( .A1(n17748), .A2(n17953), .ZN(n17773) );
  NAND2_X1 U11867 ( .A1(n15899), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16476) );
  INV_X1 U11868 ( .A(n10397), .ZN(n10396) );
  OAI21_X1 U11869 ( .B1(n16532), .B2(n16533), .A(n16531), .ZN(n10397) );
  OR2_X1 U11870 ( .A1(n16535), .A2(n18811), .ZN(n10394) );
  AND2_X1 U11871 ( .A1(n16541), .A2(n16532), .ZN(n17648) );
  NAND2_X1 U11872 ( .A1(n17648), .A2(n17793), .ZN(n17647) );
  AND2_X1 U11873 ( .A1(n15821), .A2(n15822), .ZN(n10446) );
  INV_X1 U11874 ( .A(n18197), .ZN(n18811) );
  OR2_X1 U11875 ( .A1(n15759), .A2(n15758), .ZN(n9930) );
  NOR2_X1 U11876 ( .A1(n17501), .A2(n15745), .ZN(n17925) );
  AND2_X1 U11877 ( .A1(n9937), .A2(n9936), .ZN(n17936) );
  INV_X1 U11878 ( .A(n17937), .ZN(n9936) );
  NOR2_X1 U11879 ( .A1(n17947), .A2(n17946), .ZN(n17945) );
  NAND2_X1 U11880 ( .A1(n18376), .A2(n18371), .ZN(n15778) );
  INV_X1 U11881 ( .A(n15920), .ZN(n15794) );
  OAI21_X1 U11882 ( .B1(n12908), .B2(n12907), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13930) );
  INV_X1 U11883 ( .A(n15963), .ZN(n20070) );
  INV_X1 U11884 ( .A(n14756), .ZN(n14750) );
  AND2_X2 U11885 ( .A1(n12448), .A2(n12705), .ZN(n20092) );
  NAND2_X1 U11886 ( .A1(n13322), .A2(n12447), .ZN(n12448) );
  NAND2_X1 U11887 ( .A1(n12257), .A2(n12256), .ZN(n14505) );
  INV_X1 U11888 ( .A(n14565), .ZN(n14592) );
  OR2_X1 U11889 ( .A1(n12582), .A2(n12581), .ZN(n14602) );
  AOI21_X1 U11890 ( .B1(n13325), .B2(n12574), .A(n20008), .ZN(n12582) );
  AND2_X1 U11891 ( .A1(n13330), .A2(n13224), .ZN(n12581) );
  OR2_X1 U11892 ( .A1(n12565), .A2(n12867), .ZN(n12325) );
  INV_X1 U11893 ( .A(n14505), .ZN(n12812) );
  AND2_X1 U11894 ( .A1(n12444), .A2(n12443), .ZN(n14643) );
  NAND2_X1 U11895 ( .A1(n12440), .A2(n12441), .ZN(n12444) );
  INV_X1 U11896 ( .A(n20141), .ZN(n16043) );
  NAND2_X1 U11897 ( .A1(n20155), .A2(n12816), .ZN(n16047) );
  NAND2_X1 U11898 ( .A1(n16047), .A2(n20151), .ZN(n20141) );
  XNOR2_X1 U11899 ( .A(n10011), .B(n12694), .ZN(n12893) );
  NAND2_X1 U11900 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n12690), .ZN(
        n10148) );
  XNOR2_X1 U11901 ( .A(n9954), .B(n12690), .ZN(n14758) );
  NAND2_X1 U11902 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  NAND2_X1 U11903 ( .A1(n12846), .A2(n16009), .ZN(n9955) );
  OR2_X1 U11904 ( .A1(n12845), .A2(n16009), .ZN(n9956) );
  AND2_X1 U11905 ( .A1(n12743), .A2(n12716), .ZN(n16182) );
  INV_X1 U11906 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20856) );
  NAND2_X1 U11907 ( .A1(n19216), .A2(n19199), .ZN(n10207) );
  OR2_X1 U11908 ( .A1(n19179), .A2(n11194), .ZN(n10206) );
  NAND2_X1 U11909 ( .A1(n12524), .A2(n12525), .ZN(n16208) );
  AOI21_X1 U11910 ( .B1(n19152), .B2(n15173), .A(n10203), .ZN(n10202) );
  NAND2_X1 U11911 ( .A1(n16279), .A2(n19152), .ZN(n16271) );
  NAND2_X1 U11912 ( .A1(n16280), .A2(n16281), .ZN(n16279) );
  NAND2_X1 U11913 ( .A1(n10199), .A2(n15844), .ZN(n15843) );
  INV_X1 U11914 ( .A(n19197), .ZN(n19179) );
  OR2_X1 U11915 ( .A1(n11277), .A2(n11276), .ZN(n13482) );
  NOR2_X1 U11916 ( .A1(n13360), .A2(n13359), .ZN(n13361) );
  INV_X1 U11917 ( .A(n15012), .ZN(n14961) );
  AND2_X1 U11918 ( .A1(n15501), .A2(n13167), .ZN(n19316) );
  INV_X1 U11919 ( .A(n11197), .ZN(n10133) );
  NOR2_X1 U11920 ( .A1(n10129), .A2(n11080), .ZN(n10128) );
  OR2_X1 U11921 ( .A1(n12454), .A2(n10131), .ZN(n10130) );
  NAND2_X1 U11922 ( .A1(n11080), .A2(n10132), .ZN(n10131) );
  AND2_X1 U11923 ( .A1(n16365), .A2(n19975), .ZN(n19290) );
  OR2_X1 U11924 ( .A1(n15121), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10055) );
  NOR2_X1 U11925 ( .A1(n10891), .A2(n12851), .ZN(n10056) );
  NAND2_X1 U11926 ( .A1(n15013), .A2(n15014), .ZN(n12482) );
  XNOR2_X1 U11927 ( .A(n9999), .B(n12456), .ZN(n12858) );
  NAND2_X1 U11928 ( .A1(n12454), .A2(n15124), .ZN(n9999) );
  OR2_X1 U11929 ( .A1(n15405), .A2(n9964), .ZN(n15387) );
  NOR2_X1 U11930 ( .A1(n16410), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9964) );
  AND2_X1 U11931 ( .A1(n11475), .A2(n19997), .ZN(n16391) );
  NAND2_X1 U11932 ( .A1(n11475), .A2(n19999), .ZN(n19311) );
  INV_X1 U11933 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19994) );
  NOR2_X1 U11934 ( .A1(n18805), .A2(n17560), .ZN(n19040) );
  INV_X1 U11935 ( .A(n19040), .ZN(n19036) );
  INV_X1 U11936 ( .A(n17030), .ZN(n17003) );
  INV_X1 U11937 ( .A(n17007), .ZN(n17036) );
  INV_X1 U11938 ( .A(n16498), .ZN(n9971) );
  NOR2_X1 U11939 ( .A1(n17783), .A2(n9920), .ZN(n17665) );
  AOI21_X1 U11940 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17773), .A(
        n18752), .ZN(n17833) );
  NOR2_X2 U11941 ( .A1(n17999), .A2(n17494), .ZN(n17859) );
  INV_X1 U11942 ( .A(n17861), .ZN(n17905) );
  XNOR2_X1 U11943 ( .A(n9972), .B(n16517), .ZN(n16499) );
  NAND2_X1 U11944 ( .A1(n9973), .A2(n16476), .ZN(n9972) );
  INV_X1 U11945 ( .A(n16474), .ZN(n9973) );
  CLKBUF_X1 U11946 ( .A(n18325), .Z(n18315) );
  AOI21_X1 U11947 ( .B1(n18011), .B2(n18197), .A(n9896), .ZN(n18024) );
  NAND2_X1 U11948 ( .A1(n16531), .A2(n18315), .ZN(n18229) );
  INV_X1 U11949 ( .A(n18229), .ZN(n18241) );
  INV_X1 U11950 ( .A(n18334), .ZN(n18322) );
  INV_X1 U11951 ( .A(n17019), .ZN(n18878) );
  AND4_X1 U11952 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10882) );
  NAND2_X1 U11953 ( .A1(n10895), .A2(n10894), .ZN(n10900) );
  OR2_X1 U11954 ( .A1(n11216), .A2(n10911), .ZN(n10895) );
  OAI21_X1 U11955 ( .B1(n18992), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n13016), .ZN(n13017) );
  AOI21_X1 U11956 ( .B1(n17281), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n10254), .ZN(n10253) );
  NOR2_X1 U11957 ( .A1(n17287), .A2(n18709), .ZN(n10254) );
  NAND2_X1 U11958 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10252) );
  AND2_X1 U11959 ( .A1(n11817), .A2(n11816), .ZN(n11828) );
  OR2_X1 U11960 ( .A1(n12295), .A2(n11805), .ZN(n11817) );
  OR2_X1 U11961 ( .A1(n11840), .A2(n11839), .ZN(n12653) );
  NAND2_X1 U11962 ( .A1(n10450), .A2(n11621), .ZN(n11637) );
  OAI21_X1 U11963 ( .B1(n11667), .B2(n10408), .A(n10412), .ZN(n10407) );
  INV_X1 U11964 ( .A(n10420), .ZN(n10412) );
  AOI22_X1 U11965 ( .A1(n11684), .A2(n10421), .B1(n11680), .B2(n10424), .ZN(
        n10420) );
  NOR2_X1 U11966 ( .A1(n13400), .A2(n16196), .ZN(n10009) );
  OR2_X1 U11967 ( .A1(n11790), .A2(n11789), .ZN(n12633) );
  AOI22_X1 U11968 ( .A1(n11534), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U11969 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U11970 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11528) );
  AND2_X1 U11971 ( .A1(n11598), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11495) );
  AND2_X2 U11972 ( .A1(n13380), .A2(n13397), .ZN(n11668) );
  OAI21_X1 U11973 ( .B1(n10900), .B2(n10899), .A(n10898), .ZN(n10902) );
  AND2_X1 U11974 ( .A1(n15529), .A2(n19973), .ZN(n10899) );
  XNOR2_X1 U11975 ( .A(n16411), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10901) );
  INV_X1 U11976 ( .A(n14959), .ZN(n10312) );
  INV_X1 U11977 ( .A(n10616), .ZN(n10617) );
  AOI22_X1 U11978 ( .A1(n16416), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16452), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10622) );
  INV_X1 U11979 ( .A(n16344), .ZN(n10368) );
  NOR2_X1 U11980 ( .A1(n9987), .A2(n9982), .ZN(n9981) );
  NAND4_X1 U11981 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9982)
         );
  AOI21_X1 U11982 ( .B1(n10683), .B2(n9834), .A(n9992), .ZN(n9991) );
  INV_X1 U11983 ( .A(n10620), .ZN(n11234) );
  NAND2_X1 U11984 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19994), .ZN(
        n10911) );
  NAND2_X1 U11985 ( .A1(n13042), .A2(n10620), .ZN(n11236) );
  NAND2_X1 U11986 ( .A1(n15788), .A2(n15787), .ZN(n15805) );
  NAND2_X1 U11987 ( .A1(n18384), .A2(n15915), .ZN(n12999) );
  INV_X1 U11988 ( .A(n12999), .ZN(n13003) );
  INV_X1 U11989 ( .A(n13376), .ZN(n12727) );
  AND2_X1 U11990 ( .A1(n14316), .A2(n10444), .ZN(n10443) );
  OR2_X1 U11991 ( .A1(n11895), .A2(n13739), .ZN(n11902) );
  NAND2_X1 U11992 ( .A1(n11901), .A2(n10428), .ZN(n10432) );
  INV_X1 U11993 ( .A(n14623), .ZN(n10014) );
  INV_X1 U11994 ( .A(n10183), .ZN(n10182) );
  NOR2_X1 U11995 ( .A1(n10087), .A2(n14514), .ZN(n10086) );
  INV_X1 U11996 ( .A(n15934), .ZN(n10087) );
  INV_X1 U11997 ( .A(n11872), .ZN(n10024) );
  INV_X1 U11998 ( .A(n11873), .ZN(n10025) );
  AND2_X1 U11999 ( .A1(n16016), .A2(n16017), .ZN(n14833) );
  INV_X1 U12000 ( .A(n12676), .ZN(n10417) );
  NOR2_X1 U12001 ( .A1(n10189), .A2(n10032), .ZN(n10031) );
  INV_X1 U12002 ( .A(n12650), .ZN(n10032) );
  INV_X1 U12003 ( .A(n13619), .ZN(n9959) );
  NAND2_X1 U12004 ( .A1(n10185), .A2(n12638), .ZN(n12640) );
  NAND2_X1 U12005 ( .A1(n10193), .A2(n10194), .ZN(n12615) );
  AND2_X1 U12006 ( .A1(n10195), .A2(n12609), .ZN(n10194) );
  OR2_X1 U12007 ( .A1(n9856), .A2(n10196), .ZN(n10195) );
  AOI211_X1 U12008 ( .C1(n11725), .C2(n12601), .A(n11724), .B(n11723), .ZN(
        n11768) );
  INV_X1 U12009 ( .A(n12610), .ZN(n11725) );
  AND2_X1 U12010 ( .A1(n11731), .A2(n11730), .ZN(n11767) );
  OR2_X1 U12011 ( .A1(n12295), .A2(n11726), .ZN(n11731) );
  OR2_X1 U12012 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  AND3_X1 U12013 ( .A1(n11737), .A2(n11736), .A3(n11735), .ZN(n11738) );
  NAND2_X1 U12014 ( .A1(n11769), .A2(n11732), .ZN(n11740) );
  INV_X1 U12015 ( .A(n12601), .ZN(n11732) );
  NAND2_X1 U12016 ( .A1(n11645), .A2(n11651), .ZN(n11652) );
  NOR2_X1 U12017 ( .A1(n11650), .A2(n11649), .ZN(n11651) );
  INV_X1 U12018 ( .A(n11648), .ZN(n11649) );
  AOI22_X1 U12019 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U12020 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U12021 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11511) );
  AND2_X1 U12022 ( .A1(n11776), .A2(n20700), .ZN(n20461) );
  INV_X1 U12023 ( .A(n11792), .ZN(n20334) );
  NOR2_X1 U12024 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12265), .ZN(
        n12298) );
  OR3_X1 U12025 ( .A1(n12292), .A2(n12316), .A3(n12291), .ZN(n12293) );
  NOR2_X1 U12026 ( .A1(n10295), .A2(n10936), .ZN(n10294) );
  INV_X1 U12027 ( .A(n10296), .ZN(n10295) );
  NAND2_X1 U12028 ( .A1(n11008), .A2(n11007), .ZN(n11010) );
  NOR2_X1 U12029 ( .A1(n10287), .A2(n10286), .ZN(n10285) );
  INV_X1 U12030 ( .A(n11022), .ZN(n10286) );
  INV_X1 U12031 ( .A(n10288), .ZN(n10287) );
  NOR2_X1 U12032 ( .A1(n10291), .A2(n11018), .ZN(n10290) );
  INV_X1 U12033 ( .A(n10934), .ZN(n10291) );
  NOR2_X1 U12034 ( .A1(n10289), .A2(n11016), .ZN(n10288) );
  INV_X1 U12035 ( .A(n10290), .ZN(n10289) );
  AND2_X1 U12036 ( .A1(n13926), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11018) );
  AND2_X1 U12037 ( .A1(n9860), .A2(n11114), .ZN(n10284) );
  NAND2_X1 U12038 ( .A1(n10926), .A2(n11267), .ZN(n10928) );
  NAND2_X1 U12039 ( .A1(n14946), .A2(n14182), .ZN(n14204) );
  INV_X1 U12040 ( .A(n14178), .ZN(n14181) );
  INV_X1 U12041 ( .A(n14929), .ZN(n10309) );
  NAND2_X1 U12042 ( .A1(n14060), .A2(n10319), .ZN(n10318) );
  INV_X1 U12043 ( .A(n14998), .ZN(n10319) );
  NAND2_X1 U12044 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U12045 ( .A1(n11084), .A2(n10214), .ZN(n10213) );
  INV_X1 U12046 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12047 ( .A1(n19126), .A2(n10210), .ZN(n10209) );
  INV_X1 U12048 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U12049 ( .A1(n10356), .A2(n13601), .ZN(n10355) );
  INV_X1 U12050 ( .A(n13533), .ZN(n10356) );
  NOR2_X1 U12051 ( .A1(n16364), .A2(n10220), .ZN(n10223) );
  INV_X1 U12052 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10220) );
  INV_X1 U12053 ( .A(n11302), .ZN(n10897) );
  NOR2_X1 U12054 ( .A1(n9869), .A2(n10135), .ZN(n10134) );
  INV_X1 U12055 ( .A(n15124), .ZN(n10135) );
  INV_X1 U12056 ( .A(n12828), .ZN(n10274) );
  INV_X1 U12057 ( .A(n15054), .ZN(n10278) );
  NAND2_X1 U12058 ( .A1(n9926), .A2(n10066), .ZN(n10065) );
  INV_X1 U12059 ( .A(n10067), .ZN(n10066) );
  INV_X1 U12060 ( .A(n10375), .ZN(n10374) );
  NAND2_X1 U12061 ( .A1(n10378), .A2(n15349), .ZN(n10377) );
  INV_X1 U12062 ( .A(n11455), .ZN(n10378) );
  NOR2_X1 U12063 ( .A1(n15236), .A2(n10081), .ZN(n10080) );
  INV_X1 U12064 ( .A(n11205), .ZN(n10081) );
  INV_X1 U12065 ( .A(n10607), .ZN(n11147) );
  OR2_X1 U12066 ( .A1(n10382), .A2(n15443), .ZN(n10380) );
  NAND2_X1 U12067 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10382) );
  NOR2_X1 U12068 ( .A1(n10966), .A2(n10324), .ZN(n9994) );
  NAND2_X1 U12069 ( .A1(n13964), .A2(n13963), .ZN(n10973) );
  XNOR2_X1 U12070 ( .A(n10863), .B(n11078), .ZN(n10884) );
  INV_X1 U12071 ( .A(n10854), .ZN(n10144) );
  NAND2_X1 U12072 ( .A1(n10863), .A2(n10853), .ZN(n10854) );
  NOR2_X1 U12073 ( .A1(n10849), .A2(n10848), .ZN(n11323) );
  NAND2_X1 U12074 ( .A1(n10970), .A2(n13683), .ZN(n10971) );
  NAND2_X1 U12075 ( .A1(n9998), .A2(n9946), .ZN(n10334) );
  OAI211_X1 U12076 ( .C1(n10642), .C2(n19863), .A(n10641), .B(n10640), .ZN(
        n10671) );
  AOI21_X1 U12077 ( .B1(n10634), .B2(n11442), .A(n10633), .ZN(n10642) );
  NAND2_X1 U12078 ( .A1(n10493), .A2(n10492), .ZN(n11237) );
  AND2_X1 U12079 ( .A1(n13164), .A2(n10669), .ZN(n10702) );
  AND2_X1 U12080 ( .A1(n19304), .A2(n19208), .ZN(n10699) );
  NAND2_X1 U12081 ( .A1(n10563), .A2(n16411), .ZN(n10570) );
  NAND2_X1 U12082 ( .A1(n10568), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10569) );
  NAND2_X1 U12083 ( .A1(n10530), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10531) );
  AOI22_X1 U12084 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U12085 ( .A1(n19974), .A2(n19807), .ZN(n19314) );
  AOI221_X1 U12086 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10908), 
        .C1(n13099), .C2(n10908), .A(n10907), .ZN(n11232) );
  NAND3_X1 U12087 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18999), .ZN(n12918) );
  NAND2_X1 U12088 ( .A1(n16650), .A2(n10241), .ZN(n17524) );
  AOI211_X1 U12089 ( .C1(n18365), .C2(n15919), .A(n15764), .B(n14013), .ZN(
        n15784) );
  NOR3_X1 U12090 ( .A1(n15764), .A2(n18819), .A3(n15772), .ZN(n15767) );
  NAND2_X1 U12091 ( .A1(n17524), .A2(n10095), .ZN(n13013) );
  AOI21_X1 U12092 ( .B1(n13001), .B2(n13003), .A(n10096), .ZN(n10095) );
  NOR2_X1 U12093 ( .A1(n18350), .A2(n15550), .ZN(n13001) );
  INV_X1 U12094 ( .A(n13014), .ZN(n10096) );
  NAND2_X1 U12095 ( .A1(n10255), .A2(n9865), .ZN(n10249) );
  INV_X1 U12096 ( .A(n17524), .ZN(n14025) );
  NAND2_X1 U12097 ( .A1(n18819), .A2(n14012), .ZN(n13010) );
  CLKBUF_X1 U12098 ( .A(n12312), .Z(n12313) );
  NAND2_X1 U12099 ( .A1(n12445), .A2(n12579), .ZN(n14306) );
  AND2_X1 U12100 ( .A1(n12718), .A2(n11613), .ZN(n12445) );
  CLKBUF_X1 U12101 ( .A(n12258), .Z(n12259) );
  OR2_X1 U12102 ( .A1(n14332), .A2(n12426), .ZN(n12868) );
  AND2_X1 U12103 ( .A1(n12373), .A2(n12372), .ZN(n14526) );
  NAND2_X1 U12104 ( .A1(n10166), .A2(n10165), .ZN(n12366) );
  NAND2_X1 U12105 ( .A1(n12404), .A2(n10167), .ZN(n10166) );
  MUX2_X1 U12106 ( .A(n12253), .B(n12821), .S(n12566), .Z(n12254) );
  INV_X1 U12107 ( .A(n14313), .ZN(n13777) );
  MUX2_X1 U12108 ( .A(n12214), .B(n14639), .S(n12566), .Z(n12441) );
  NAND2_X1 U12109 ( .A1(n12195), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12229) );
  AND2_X1 U12110 ( .A1(n12141), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12142) );
  INV_X1 U12111 ( .A(n12140), .ZN(n12141) );
  AOI21_X1 U12112 ( .B1(n12566), .B2(n14671), .A(n12160), .ZN(n14365) );
  CLKBUF_X1 U12113 ( .A(n14350), .Z(n14351) );
  NOR2_X1 U12114 ( .A1(n12096), .A2(n14695), .ZN(n12097) );
  NAND2_X1 U12115 ( .A1(n12097), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12140) );
  AND2_X1 U12116 ( .A1(n10418), .A2(n14815), .ZN(n10038) );
  AND2_X1 U12117 ( .A1(n12095), .A2(n12094), .ZN(n14411) );
  AND2_X1 U12118 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n12061), .ZN(
        n12062) );
  NAND2_X1 U12119 ( .A1(n12062), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12096) );
  INV_X1 U12120 ( .A(n10441), .ZN(n10439) );
  CLKBUF_X1 U12121 ( .A(n14436), .Z(n14437) );
  NAND2_X1 U12122 ( .A1(n12030), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12060) );
  INV_X1 U12123 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14736) );
  INV_X1 U12124 ( .A(n10427), .ZN(n10425) );
  NOR2_X1 U12125 ( .A1(n11998), .A2(n15938), .ZN(n11999) );
  NAND2_X1 U12126 ( .A1(n11982), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11998) );
  CLKBUF_X1 U12127 ( .A(n14523), .Z(n14524) );
  NOR2_X1 U12128 ( .A1(n11968), .A2(n15953), .ZN(n11982) );
  OR2_X1 U12129 ( .A1(n11962), .A2(n15964), .ZN(n11968) );
  CLKBUF_X1 U12130 ( .A(n14521), .Z(n14522) );
  AND2_X1 U12131 ( .A1(n11918), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11919) );
  NOR2_X1 U12132 ( .A1(n11902), .A2(n11903), .ZN(n11918) );
  AOI21_X1 U12133 ( .B1(n13891), .B2(n12566), .A(n11917), .ZN(n13864) );
  INV_X1 U12134 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13739) );
  CLKBUF_X1 U12135 ( .A(n13613), .Z(n13614) );
  OR2_X1 U12136 ( .A1(n11878), .A2(n11881), .ZN(n11895) );
  AOI21_X1 U12137 ( .B1(n12651), .B2(n11991), .A(n11871), .ZN(n13645) );
  CLKBUF_X1 U12138 ( .A(n13611), .Z(n13612) );
  AND2_X1 U12139 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11506), .ZN(
        n11823) );
  NAND2_X1 U12140 ( .A1(n12845), .A2(n10154), .ZN(n12692) );
  NAND2_X1 U12141 ( .A1(n14647), .A2(n12690), .ZN(n12693) );
  INV_X1 U12142 ( .A(n10028), .ZN(n12844) );
  NAND2_X1 U12143 ( .A1(n10171), .A2(n10170), .ZN(n12410) );
  NAND2_X1 U12144 ( .A1(n12404), .A2(n21212), .ZN(n10171) );
  NAND2_X1 U12145 ( .A1(n14396), .A2(n9909), .ZN(n14360) );
  INV_X1 U12146 ( .A(n14358), .ZN(n10088) );
  NAND2_X1 U12147 ( .A1(n14396), .A2(n10089), .ZN(n14371) );
  NAND2_X1 U12148 ( .A1(n12395), .A2(n10172), .ZN(n12396) );
  NAND2_X1 U12149 ( .A1(n14396), .A2(n14385), .ZN(n14387) );
  NAND2_X1 U12150 ( .A1(n10169), .A2(n10168), .ZN(n12394) );
  NAND2_X1 U12151 ( .A1(n12404), .A2(n21168), .ZN(n10169) );
  AND2_X1 U12152 ( .A1(n14416), .A2(n14395), .ZN(n14396) );
  NAND2_X1 U12153 ( .A1(n10018), .A2(n10154), .ZN(n14683) );
  NOR2_X1 U12154 ( .A1(n10191), .A2(n15889), .ZN(n10019) );
  NOR2_X1 U12155 ( .A1(n14427), .A2(n14414), .ZN(n14416) );
  OR2_X1 U12156 ( .A1(n14442), .A2(n14426), .ZN(n14427) );
  NOR2_X1 U12157 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10418) );
  AND2_X1 U12158 ( .A1(n14469), .A2(n14455), .ZN(n14457) );
  AND2_X1 U12159 ( .A1(n12389), .A2(n12388), .ZN(n14440) );
  NAND2_X1 U12160 ( .A1(n14457), .A2(n14440), .ZN(n14442) );
  AND2_X1 U12161 ( .A1(n15935), .A2(n10084), .ZN(n14469) );
  NOR2_X1 U12162 ( .A1(n10085), .A2(n14467), .ZN(n10084) );
  INV_X1 U12163 ( .A(n10086), .ZN(n10085) );
  NAND2_X1 U12164 ( .A1(n15935), .A2(n10086), .ZN(n14515) );
  NAND2_X1 U12165 ( .A1(n15935), .A2(n15934), .ZN(n15937) );
  AND2_X1 U12166 ( .A1(n16188), .A2(n16196), .ZN(n12815) );
  NAND2_X1 U12167 ( .A1(n12363), .A2(n10180), .ZN(n12364) );
  NOR2_X1 U12168 ( .A1(n15972), .A2(n15971), .ZN(n15974) );
  OR2_X1 U12169 ( .A1(n13918), .A2(n13917), .ZN(n15972) );
  NAND2_X1 U12170 ( .A1(n12357), .A2(n10178), .ZN(n12358) );
  OR2_X1 U12171 ( .A1(n13883), .A2(n13882), .ZN(n13918) );
  NAND2_X1 U12172 ( .A1(n10163), .A2(n10162), .ZN(n12356) );
  NAND2_X1 U12173 ( .A1(n12404), .A2(n10164), .ZN(n10163) );
  NAND2_X1 U12174 ( .A1(n12350), .A2(n10174), .ZN(n12351) );
  NAND2_X1 U12175 ( .A1(n10160), .A2(n10159), .ZN(n12354) );
  NAND2_X1 U12176 ( .A1(n12404), .A2(n10161), .ZN(n10160) );
  NAND2_X1 U12177 ( .A1(n12347), .A2(n10176), .ZN(n12348) );
  OR2_X1 U12178 ( .A1(n10094), .A2(n13512), .ZN(n16173) );
  NAND2_X1 U12179 ( .A1(n12346), .A2(n10092), .ZN(n10094) );
  INV_X1 U12180 ( .A(n16170), .ZN(n10092) );
  INV_X1 U12181 ( .A(n12723), .ZN(n11650) );
  OR2_X1 U12182 ( .A1(n13512), .A2(n13511), .ZN(n16171) );
  NAND2_X1 U12183 ( .A1(n10186), .A2(n12631), .ZN(n13510) );
  XNOR2_X1 U12184 ( .A(n12640), .B(n12639), .ZN(n13509) );
  NAND2_X1 U12185 ( .A1(n13471), .A2(n13470), .ZN(n13512) );
  XNOR2_X1 U12186 ( .A(n12630), .B(n13469), .ZN(n13464) );
  AOI21_X1 U12187 ( .B1(n13780), .B2(n12718), .A(n12337), .ZN(n13347) );
  NAND2_X1 U12188 ( .A1(n10157), .A2(n10156), .ZN(n12339) );
  NAND2_X1 U12189 ( .A1(n12404), .A2(n10158), .ZN(n10157) );
  INV_X1 U12190 ( .A(n16140), .ZN(n16117) );
  OR2_X1 U12191 ( .A1(n12744), .A2(n20171), .ZN(n13352) );
  NAND2_X1 U12192 ( .A1(n12626), .A2(n12625), .ZN(n13344) );
  AND2_X1 U12193 ( .A1(n14810), .A2(n20161), .ZN(n16140) );
  OR2_X1 U12194 ( .A1(n13316), .A2(n11647), .ZN(n12723) );
  NAND2_X1 U12195 ( .A1(n11742), .A2(n9952), .ZN(n11744) );
  INV_X1 U12196 ( .A(n10015), .ZN(n9952) );
  OR2_X1 U12197 ( .A1(n20456), .A2(n11792), .ZN(n20432) );
  BUF_X1 U12198 ( .A(n11570), .Z(n20213) );
  CLKBUF_X1 U12199 ( .A(n11617), .Z(n11618) );
  AOI22_X1 U12200 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11562) );
  INV_X1 U12201 ( .A(n20557), .ZN(n20847) );
  AND2_X1 U12202 ( .A1(n13427), .A2(n20859), .ZN(n20560) );
  INV_X1 U12203 ( .A(n20560), .ZN(n20426) );
  INV_X1 U12204 ( .A(n20513), .ZN(n20659) );
  INV_X1 U12205 ( .A(n20342), .ZN(n20236) );
  NOR2_X1 U12206 ( .A1(n20189), .A2(n16195), .ZN(n15874) );
  NOR2_X1 U12207 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16452) );
  NAND2_X1 U12208 ( .A1(n10556), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U12209 ( .A1(n10551), .A2(n16411), .ZN(n10558) );
  XNOR2_X1 U12210 ( .A(n11075), .B(n11072), .ZN(n12535) );
  NOR2_X1 U12211 ( .A1(n11066), .A2(n11065), .ZN(n11070) );
  NOR2_X1 U12212 ( .A1(n12521), .A2(n10217), .ZN(n12523) );
  NAND2_X1 U12213 ( .A1(n11008), .A2(n10296), .ZN(n11004) );
  NOR2_X1 U12214 ( .A1(n12509), .A2(n15257), .ZN(n12512) );
  NAND2_X1 U12215 ( .A1(n19124), .A2(n10290), .ZN(n10467) );
  AND2_X1 U12216 ( .A1(n19124), .A2(n10288), .ZN(n11023) );
  NAND2_X1 U12217 ( .A1(n19124), .A2(n10934), .ZN(n11019) );
  NAND2_X1 U12218 ( .A1(n10980), .A2(n9860), .ZN(n10987) );
  NAND2_X1 U12219 ( .A1(n10360), .A2(n10362), .ZN(n10359) );
  INV_X1 U12220 ( .A(n12457), .ZN(n10362) );
  OR2_X1 U12221 ( .A1(n11366), .A2(n11365), .ZN(n13630) );
  NAND2_X1 U12222 ( .A1(n10303), .A2(n9911), .ZN(n10304) );
  NOR2_X1 U12223 ( .A1(n14922), .A2(n10309), .ZN(n10305) );
  NAND2_X1 U12224 ( .A1(n10310), .A2(n10308), .ZN(n10307) );
  NOR2_X1 U12225 ( .A1(n10309), .A2(n14934), .ZN(n10308) );
  INV_X1 U12226 ( .A(n14922), .ZN(n10310) );
  INV_X1 U12227 ( .A(n14934), .ZN(n10301) );
  INV_X1 U12228 ( .A(n14229), .ZN(n10302) );
  NAND2_X1 U12229 ( .A1(n14138), .A2(n10314), .ZN(n10313) );
  NAND2_X1 U12230 ( .A1(n14968), .A2(n14970), .ZN(n14969) );
  NAND2_X1 U12231 ( .A1(n15084), .A2(n11430), .ZN(n15064) );
  NOR2_X2 U12232 ( .A1(n14974), .A2(n14975), .ZN(n14138) );
  NAND2_X1 U12233 ( .A1(n10317), .A2(n14060), .ZN(n14997) );
  INV_X1 U12234 ( .A(n14049), .ZN(n10317) );
  OR2_X1 U12235 ( .A1(n13954), .A2(n13953), .ZN(n13956) );
  OR2_X1 U12236 ( .A1(n16384), .A2(n10268), .ZN(n13475) );
  NOR2_X1 U12237 ( .A1(n14222), .A2(n13296), .ZN(n13593) );
  NAND2_X1 U12238 ( .A1(n11288), .A2(n11287), .ZN(n13186) );
  AND2_X1 U12239 ( .A1(n13186), .A2(n13185), .ZN(n13188) );
  INV_X1 U12240 ( .A(n11213), .ZN(n13150) );
  NOR2_X1 U12241 ( .A1(n16430), .A2(n13144), .ZN(n13038) );
  INV_X1 U12242 ( .A(n13930), .ZN(n19315) );
  INV_X1 U12243 ( .A(n10134), .ZN(n10129) );
  INV_X1 U12244 ( .A(n12455), .ZN(n10132) );
  NOR3_X1 U12245 ( .A1(n12521), .A2(n10219), .A3(n10216), .ZN(n12485) );
  OR2_X1 U12246 ( .A1(n10217), .A2(n10218), .ZN(n10216) );
  NOR3_X1 U12247 ( .A1(n12521), .A2(n10219), .A3(n10217), .ZN(n12490) );
  INV_X1 U12248 ( .A(n10360), .ZN(n10358) );
  AND2_X1 U12249 ( .A1(n12785), .A2(n12784), .ZN(n12783) );
  OR2_X1 U12250 ( .A1(n12493), .A2(n15156), .ZN(n12521) );
  NAND2_X1 U12251 ( .A1(n12515), .A2(n9840), .ZN(n12519) );
  NAND2_X1 U12252 ( .A1(n12515), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12517) );
  NAND2_X1 U12253 ( .A1(n9810), .A2(n10335), .ZN(n14995) );
  INV_X1 U12254 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15219) );
  NAND2_X1 U12255 ( .A1(n12512), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12511) );
  INV_X1 U12256 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12496) );
  NOR2_X1 U12257 ( .A1(n12511), .A2(n12496), .ZN(n12513) );
  NAND2_X1 U12258 ( .A1(n10890), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10067) );
  NOR2_X1 U12259 ( .A1(n13726), .A2(n13725), .ZN(n13804) );
  NAND2_X1 U12260 ( .A1(n12510), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12509) );
  AND2_X1 U12261 ( .A1(n12507), .A2(n10208), .ZN(n12510) );
  AND2_X1 U12262 ( .A1(n9837), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10208) );
  NAND2_X1 U12263 ( .A1(n12507), .A2(n9837), .ZN(n12508) );
  INV_X1 U12264 ( .A(n10352), .ZN(n10351) );
  OR2_X1 U12265 ( .A1(n13483), .A2(n10355), .ZN(n13605) );
  NAND2_X1 U12266 ( .A1(n12507), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12506) );
  NOR2_X1 U12267 ( .A1(n12504), .A2(n16335), .ZN(n12507) );
  NOR2_X1 U12268 ( .A1(n13483), .A2(n13533), .ZN(n13600) );
  NAND2_X1 U12269 ( .A1(n10221), .A2(n10222), .ZN(n12504) );
  AND2_X1 U12270 ( .A1(n9833), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10221) );
  AND2_X1 U12271 ( .A1(n10222), .A2(n9833), .ZN(n12505) );
  NAND2_X1 U12272 ( .A1(n10222), .A2(n10223), .ZN(n12502) );
  NOR2_X1 U12273 ( .A1(n12500), .A2(n16364), .ZN(n12503) );
  INV_X1 U12274 ( .A(n10338), .ZN(n10336) );
  NAND2_X1 U12275 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12499) );
  NOR2_X1 U12276 ( .A1(n12499), .A2(n14033), .ZN(n12501) );
  INV_X1 U12277 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14033) );
  OAI22_X1 U12278 ( .A1(n10126), .A2(n10129), .B1(n11080), .B2(n10134), .ZN(
        n10125) );
  NOR2_X1 U12279 ( .A1(n11080), .A2(n10132), .ZN(n10126) );
  AND2_X1 U12280 ( .A1(n9921), .A2(n12777), .ZN(n10275) );
  INV_X1 U12281 ( .A(n12481), .ZN(n10276) );
  NOR2_X1 U12282 ( .A1(n12775), .A2(n12794), .ZN(n15123) );
  AND2_X1 U12283 ( .A1(n12474), .A2(n12473), .ZN(n15029) );
  NAND2_X1 U12284 ( .A1(n14949), .A2(n14950), .ZN(n14952) );
  AOI21_X1 U12285 ( .B1(n10003), .B2(n10142), .A(n10001), .ZN(n10000) );
  INV_X1 U12286 ( .A(n10003), .ZN(n10002) );
  INV_X1 U12287 ( .A(n15165), .ZN(n10001) );
  OR3_X1 U12288 ( .A1(n16253), .A2(n11326), .A3(n15155), .ZN(n15150) );
  AND2_X1 U12289 ( .A1(n12469), .A2(n12468), .ZN(n15311) );
  NAND2_X1 U12290 ( .A1(n15084), .A2(n9904), .ZN(n15062) );
  INV_X1 U12291 ( .A(n10065), .ZN(n10064) );
  NAND2_X1 U12292 ( .A1(n10140), .A2(n11041), .ZN(n15176) );
  NAND2_X1 U12293 ( .A1(n10331), .A2(n10332), .ZN(n10140) );
  NAND2_X1 U12294 ( .A1(n10376), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10375) );
  INV_X1 U12295 ( .A(n10377), .ZN(n10376) );
  AND2_X1 U12296 ( .A1(n15214), .A2(n15226), .ZN(n15202) );
  INV_X1 U12297 ( .A(n10071), .ZN(n10070) );
  OAI21_X1 U12298 ( .B1(n10078), .B2(n10072), .A(n10074), .ZN(n10071) );
  AND2_X1 U12299 ( .A1(n11427), .A2(n11426), .ZN(n14872) );
  AND2_X1 U12300 ( .A1(n10263), .A2(n10262), .ZN(n10261) );
  INV_X1 U12301 ( .A(n15102), .ZN(n10262) );
  NAND2_X1 U12302 ( .A1(n16366), .A2(n10263), .ZN(n15101) );
  NAND2_X1 U12303 ( .A1(n10073), .A2(n10077), .ZN(n15228) );
  NAND2_X1 U12304 ( .A1(n15244), .A2(n10080), .ZN(n10073) );
  AND2_X1 U12305 ( .A1(n16366), .A2(n9892), .ZN(n14885) );
  AND2_X1 U12306 ( .A1(n10348), .A2(n10346), .ZN(n10345) );
  INV_X1 U12307 ( .A(n13909), .ZN(n10346) );
  NAND2_X1 U12308 ( .A1(n10347), .A2(n10348), .ZN(n13910) );
  NAND2_X1 U12309 ( .A1(n16366), .A2(n13832), .ZN(n13923) );
  AND2_X1 U12310 ( .A1(n15464), .A2(n15463), .ZN(n15486) );
  NAND2_X1 U12311 ( .A1(n10973), .A2(n10325), .ZN(n15464) );
  INV_X1 U12312 ( .A(n10323), .ZN(n10325) );
  NOR2_X1 U12313 ( .A1(n16384), .A2(n16385), .ZN(n16383) );
  NOR2_X1 U12314 ( .A1(n10338), .A2(n10343), .ZN(n10337) );
  INV_X1 U12315 ( .A(n13364), .ZN(n10343) );
  NAND2_X1 U12316 ( .A1(n10042), .A2(n10966), .ZN(n13964) );
  INV_X1 U12317 ( .A(n10860), .ZN(n13870) );
  NOR2_X1 U12318 ( .A1(n11310), .A2(n10257), .ZN(n10259) );
  NAND2_X1 U12319 ( .A1(n13493), .A2(n10258), .ZN(n10257) );
  INV_X1 U12320 ( .A(n13591), .ZN(n10258) );
  NAND2_X1 U12321 ( .A1(n9800), .A2(n9947), .ZN(n10040) );
  NAND2_X1 U12322 ( .A1(n10050), .A2(n13577), .ZN(n10044) );
  NAND2_X1 U12323 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  OAI21_X1 U12324 ( .B1(n10614), .B2(n11090), .A(n10120), .ZN(n10119) );
  NAND2_X1 U12325 ( .A1(n9938), .A2(n10645), .ZN(n10646) );
  OR2_X1 U12326 ( .A1(n15381), .A2(n15386), .ZN(n19302) );
  XNOR2_X1 U12327 ( .A(n13293), .B(n13290), .ZN(n13338) );
  AND2_X2 U12328 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15521) );
  NOR2_X2 U12329 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15511) );
  CLKBUF_X1 U12330 ( .A(n14270), .Z(n15518) );
  OR2_X1 U12331 ( .A1(n19963), .A2(n19316), .ZN(n19449) );
  OR2_X1 U12332 ( .A1(n19963), .A2(n19988), .ZN(n19480) );
  INV_X1 U12333 ( .A(n19449), .ZN(n19508) );
  INV_X1 U12334 ( .A(n19480), .ZN(n19539) );
  INV_X1 U12335 ( .A(n10800), .ZN(n19697) );
  INV_X1 U12336 ( .A(n10803), .ZN(n19758) );
  INV_X2 U12337 ( .A(n16437), .ZN(n19317) );
  AND2_X1 U12338 ( .A1(n19963), .A2(n19988), .ZN(n19752) );
  NOR2_X2 U12339 ( .A1(n19315), .A2(n19314), .ZN(n19349) );
  NOR2_X2 U12340 ( .A1(n19313), .A2(n19314), .ZN(n19350) );
  NAND2_X1 U12341 ( .A1(n19963), .A2(n19316), .ZN(n19727) );
  AOI21_X1 U12342 ( .B1(n15770), .B2(n14023), .A(n15769), .ZN(n18812) );
  NOR2_X1 U12343 ( .A1(n14025), .A2(n14024), .ZN(n18805) );
  OR2_X1 U12344 ( .A1(n16800), .A2(n17738), .ZN(n10230) );
  NOR2_X1 U12345 ( .A1(n19036), .A2(n15915), .ZN(n13030) );
  AND2_X1 U12346 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17152), .ZN(n17125) );
  NOR2_X1 U12347 ( .A1(n17583), .A2(n10098), .ZN(n10097) );
  AOI21_X1 U12348 ( .B1(n15917), .B2(n15916), .A(n18874), .ZN(n17513) );
  INV_X1 U12349 ( .A(n17513), .ZN(n17372) );
  NOR3_X1 U12350 ( .A1(n17524), .A2(n19023), .A3(n17560), .ZN(n17542) );
  NOR2_X1 U12351 ( .A1(n17561), .A2(n17560), .ZN(n17562) );
  NOR2_X1 U12352 ( .A1(n18006), .A2(n17667), .ZN(n17641) );
  NAND2_X1 U12353 ( .A1(n17710), .A2(n9826), .ZN(n17634) );
  OR2_X1 U12354 ( .A1(n18150), .A2(n18029), .ZN(n17667) );
  INV_X1 U12355 ( .A(n18150), .ZN(n18068) );
  NAND2_X1 U12356 ( .A1(n17710), .A2(n9887), .ZN(n17670) );
  NAND2_X1 U12357 ( .A1(n17894), .A2(n9895), .ZN(n10237) );
  NOR2_X1 U12358 ( .A1(n17834), .A2(n17815), .ZN(n10238) );
  INV_X1 U12359 ( .A(n17954), .ZN(n16987) );
  INV_X1 U12360 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17956) );
  NAND2_X1 U12361 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17954) );
  INV_X1 U12362 ( .A(n17995), .ZN(n17953) );
  INV_X1 U12363 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17016) );
  NOR2_X1 U12364 ( .A1(n15900), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16474) );
  NOR2_X1 U12365 ( .A1(n16532), .A2(n10457), .ZN(n15899) );
  NAND2_X1 U12366 ( .A1(n17792), .A2(n17686), .ZN(n10108) );
  NAND2_X1 U12367 ( .A1(n17729), .A2(n9919), .ZN(n17698) );
  NAND2_X1 U12368 ( .A1(n17860), .A2(n18115), .ZN(n18150) );
  INV_X1 U12369 ( .A(n18224), .ZN(n18841) );
  NOR2_X1 U12370 ( .A1(n15816), .A2(n18237), .ZN(n17862) );
  NAND2_X1 U12371 ( .A1(n10115), .A2(n17857), .ZN(n10113) );
  NAND2_X1 U12372 ( .A1(n18831), .A2(n18821), .ZN(n10245) );
  NAND2_X1 U12373 ( .A1(n15760), .A2(n9928), .ZN(n17900) );
  NAND2_X1 U12374 ( .A1(n15757), .A2(n9929), .ZN(n9928) );
  INV_X1 U12375 ( .A(n15762), .ZN(n9929) );
  INV_X1 U12376 ( .A(n17793), .ZN(n17902) );
  AND2_X1 U12377 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  NAND2_X1 U12378 ( .A1(n17921), .A2(n9873), .ZN(n10391) );
  NAND2_X1 U12379 ( .A1(n17910), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17909) );
  NOR2_X1 U12380 ( .A1(n17936), .A2(n15755), .ZN(n17924) );
  XNOR2_X1 U12381 ( .A(n15797), .B(n18291), .ZN(n17966) );
  NOR2_X1 U12382 ( .A1(n17973), .A2(n15749), .ZN(n17963) );
  NOR2_X1 U12383 ( .A1(n17962), .A2(n17963), .ZN(n17961) );
  XNOR2_X1 U12384 ( .A(n15748), .B(n18304), .ZN(n17974) );
  NOR2_X1 U12385 ( .A1(n17975), .A2(n17974), .ZN(n17973) );
  OAI21_X1 U12386 ( .B1(n14021), .B2(n13026), .A(n14022), .ZN(n15776) );
  AOI211_X1 U12387 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n12980), .B(n12979), .ZN(n15779) );
  INV_X1 U12388 ( .A(n13013), .ZN(n18831) );
  AND2_X1 U12389 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18817) );
  INV_X1 U12390 ( .A(n18817), .ZN(n18832) );
  NAND2_X1 U12391 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15645) );
  NOR2_X1 U12392 ( .A1(n13013), .A2(n15768), .ZN(n14010) );
  AOI22_X1 U12393 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12939) );
  AOI211_X1 U12394 ( .C1(n15554), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12937), .B(n12936), .ZN(n12938) );
  OAI211_X1 U12395 ( .C1(n15688), .C2(n17285), .A(n12998), .B(n12997), .ZN(
        n18355) );
  AOI211_X1 U12396 ( .C1(n15554), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12996), .B(n12995), .ZN(n12997) );
  OAI211_X1 U12397 ( .C1(n17287), .C2(n18696), .A(n12959), .B(n12958), .ZN(
        n18360) );
  NOR2_X1 U12398 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18343), .ZN(n18511) );
  INV_X1 U12399 ( .A(n15779), .ZN(n18365) );
  OAI211_X1 U12400 ( .C1(n17283), .C2(n18374), .A(n12969), .B(n12968), .ZN(
        n18371) );
  AOI211_X1 U12401 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n12967), .B(n12966), .ZN(n12968) );
  INV_X1 U12402 ( .A(n18511), .ZN(n18653) );
  OAI22_X1 U12403 ( .A1(n16473), .A2(n18807), .B1(n18811), .B2(n16472), .ZN(
        n18862) );
  NOR2_X1 U12404 ( .A1(n13010), .A2(n10102), .ZN(n18867) );
  NAND2_X1 U12405 ( .A1(n18345), .A2(n10103), .ZN(n10102) );
  NOR2_X1 U12406 ( .A1(n15764), .A2(n18371), .ZN(n10103) );
  NOR2_X1 U12407 ( .A1(n18869), .A2(n17994), .ZN(n19020) );
  NOR3_X1 U12408 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18903), .A3(n18885), 
        .ZN(n15775) );
  OR3_X1 U12409 ( .A1(n12313), .A2(n20008), .A3(n14311), .ZN(n13108) );
  AND2_X1 U12410 ( .A1(n13543), .A2(n13108), .ZN(n20875) );
  OR2_X1 U12411 ( .A1(n20030), .A2(n20466), .ZN(n20057) );
  INV_X1 U12412 ( .A(n20059), .ZN(n20073) );
  OR2_X1 U12413 ( .A1(n20030), .A2(n13738), .ZN(n20055) );
  INV_X1 U12414 ( .A(n15978), .ZN(n20047) );
  INV_X1 U12415 ( .A(n20057), .ZN(n20069) );
  INV_X1 U12416 ( .A(n20032), .ZN(n20077) );
  NAND2_X1 U12417 ( .A1(n20032), .A2(n13814), .ZN(n20029) );
  NAND2_X1 U12418 ( .A1(n12424), .A2(n12420), .ZN(n15963) );
  INV_X1 U12419 ( .A(n14546), .ZN(n20088) );
  CLKBUF_X1 U12420 ( .A(n14543), .Z(n14544) );
  INV_X1 U12421 ( .A(n14604), .ZN(n14620) );
  CLKBUF_X1 U12422 ( .A(n13455), .Z(n13456) );
  AND3_X1 U12423 ( .A1(n13226), .A2(n13225), .A3(n13224), .ZN(n20095) );
  INV_X1 U12424 ( .A(n13748), .ZN(n20135) );
  INV_X1 U12425 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14695) );
  NAND2_X1 U12426 ( .A1(n10021), .A2(n9835), .ZN(n14692) );
  NAND2_X1 U12427 ( .A1(n10145), .A2(n10038), .ZN(n14693) );
  CLKBUF_X1 U12428 ( .A(n14613), .Z(n14616) );
  NAND2_X1 U12429 ( .A1(n12677), .A2(n12676), .ZN(n13889) );
  INV_X1 U12430 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20056) );
  CLKBUF_X1 U12431 ( .A(n13518), .Z(n13519) );
  INV_X1 U12432 ( .A(n16047), .ZN(n20152) );
  XNOR2_X1 U12433 ( .A(n10082), .B(n12865), .ZN(n14756) );
  AOI21_X1 U12434 ( .B1(n12863), .B2(n13172), .A(n10083), .ZN(n10082) );
  INV_X1 U12435 ( .A(n12689), .ZN(n14636) );
  NAND2_X1 U12436 ( .A1(n10145), .A2(n10418), .ZN(n14704) );
  NAND2_X1 U12437 ( .A1(n10023), .A2(n16016), .ZN(n16020) );
  INV_X1 U12438 ( .A(n14743), .ZN(n10023) );
  INV_X1 U12439 ( .A(n20149), .ZN(n20140) );
  NAND2_X1 U12440 ( .A1(n10188), .A2(n12659), .ZN(n16037) );
  NOR2_X1 U12441 ( .A1(n12328), .A2(n14788), .ZN(n13467) );
  NAND2_X1 U12442 ( .A1(n16140), .A2(n20162), .ZN(n20157) );
  CLKBUF_X1 U12443 ( .A(n11758), .Z(n11759) );
  INV_X1 U12444 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20866) );
  INV_X1 U12445 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20514) );
  NOR2_X2 U12446 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20858) );
  INV_X1 U12447 ( .A(n20858), .ZN(n20852) );
  AND2_X1 U12448 ( .A1(n10037), .A2(n11666), .ZN(n10035) );
  OR2_X1 U12449 ( .A1(n20466), .A2(n14307), .ZN(n20841) );
  NOR2_X1 U12450 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16188) );
  INV_X1 U12451 ( .A(n20291), .ZN(n20262) );
  INV_X1 U12452 ( .A(n20425), .ZN(n20390) );
  OR2_X1 U12453 ( .A1(n20432), .A2(n20426), .ZN(n20455) );
  INV_X1 U12454 ( .A(n20455), .ZN(n20483) );
  INV_X1 U12455 ( .A(n20547), .ZN(n20508) );
  INV_X1 U12456 ( .A(n20626), .ZN(n20577) );
  OAI211_X1 U12457 ( .C1(n20693), .C2(n20667), .A(n20666), .B(n20665), .ZN(
        n20696) );
  INV_X1 U12458 ( .A(n20583), .ZN(n20706) );
  INV_X1 U12459 ( .A(n20595), .ZN(n20718) );
  INV_X1 U12460 ( .A(n20599), .ZN(n20724) );
  OR2_X1 U12461 ( .A1(n20709), .A2(n20426), .ZN(n20735) );
  INV_X1 U12462 ( .A(n20603), .ZN(n20730) );
  INV_X1 U12463 ( .A(n20607), .ZN(n20738) );
  INV_X1 U12464 ( .A(n20539), .ZN(n20744) );
  INV_X1 U12465 ( .A(n20615), .ZN(n20750) );
  OR2_X1 U12466 ( .A1(n20709), .A2(n20659), .ZN(n20764) );
  INV_X1 U12467 ( .A(n20735), .ZN(n20760) );
  NAND2_X1 U12468 ( .A1(n12311), .A2(n12310), .ZN(n15882) );
  NAND2_X1 U12469 ( .A1(n12297), .A2(n12319), .ZN(n12311) );
  OR2_X1 U12470 ( .A1(n20766), .A2(n16196), .ZN(n20008) );
  NAND2_X1 U12471 ( .A1(n16195), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20766) );
  AOI21_X1 U12472 ( .B1(n16432), .B2(n16431), .A(n9940), .ZN(n16436) );
  NAND2_X1 U12473 ( .A1(n16246), .A2(n19152), .ZN(n16236) );
  NAND2_X1 U12474 ( .A1(n16236), .A2(n16237), .ZN(n16235) );
  AND2_X1 U12475 ( .A1(n10941), .A2(n11077), .ZN(n16242) );
  NOR2_X1 U12476 ( .A1(n10203), .A2(n15173), .ZN(n10201) );
  NAND2_X1 U12477 ( .A1(n16259), .A2(n16260), .ZN(n16258) );
  INV_X1 U12478 ( .A(n19141), .ZN(n19205) );
  NAND2_X1 U12479 ( .A1(n14867), .A2(n19152), .ZN(n10199) );
  NAND2_X1 U12480 ( .A1(n14868), .A2(n15195), .ZN(n14867) );
  NAND2_X1 U12481 ( .A1(n19152), .A2(n10464), .ZN(n19074) );
  INV_X1 U12482 ( .A(n19210), .ZN(n19167) );
  INV_X1 U12483 ( .A(n19207), .ZN(n19185) );
  AND2_X1 U12484 ( .A1(n19043), .A2(n12532), .ZN(n19197) );
  NAND2_X1 U12485 ( .A1(n16200), .A2(n12531), .ZN(n19183) );
  XNOR2_X1 U12486 ( .A(n13496), .B(n13498), .ZN(n19448) );
  NOR2_X1 U12487 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  OR2_X1 U12488 ( .A1(n11403), .A2(n11402), .ZN(n13724) );
  CLKBUF_X1 U12489 ( .A(n13808), .Z(n13806) );
  OR2_X1 U12490 ( .A1(n11390), .A2(n11389), .ZN(n13676) );
  AND2_X1 U12491 ( .A1(n13532), .A2(n10321), .ZN(n13677) );
  AND2_X1 U12492 ( .A1(n10342), .A2(n11091), .ZN(n13664) );
  OR2_X1 U12493 ( .A1(n13301), .A2(n19352), .ZN(n15012) );
  OAI21_X1 U12494 ( .B1(n14935), .B2(n10300), .A(n10299), .ZN(n10298) );
  NAND2_X1 U12495 ( .A1(n10301), .A2(n14929), .ZN(n10300) );
  AND2_X1 U12496 ( .A1(n19249), .A2(n13931), .ZN(n19217) );
  AND2_X1 U12497 ( .A1(n19249), .A2(n13927), .ZN(n16286) );
  NOR2_X1 U12498 ( .A1(n16384), .A2(n10267), .ZN(n13539) );
  AND2_X1 U12499 ( .A1(n13181), .A2(n19866), .ZN(n19249) );
  INV_X1 U12500 ( .A(n15120), .ZN(n19246) );
  INV_X1 U12501 ( .A(n15023), .ZN(n19245) );
  INV_X1 U12502 ( .A(n19249), .ZN(n19231) );
  OR2_X1 U12503 ( .A1(n13046), .A2(n14227), .ZN(n13143) );
  XNOR2_X1 U12504 ( .A(n15229), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15241) );
  NAND2_X1 U12505 ( .A1(n10061), .A2(n15435), .ZN(n15429) );
  NAND2_X1 U12506 ( .A1(n10062), .A2(n10995), .ZN(n10061) );
  INV_X1 U12507 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16335) );
  INV_X1 U12508 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16364) );
  INV_X1 U12509 ( .A(n16355), .ZN(n19296) );
  NAND2_X1 U12510 ( .A1(n13045), .A2(n11082), .ZN(n16365) );
  AND2_X1 U12511 ( .A1(n16365), .A2(n13105), .ZN(n16355) );
  INV_X1 U12512 ( .A(n19290), .ZN(n15258) );
  INV_X1 U12513 ( .A(n16365), .ZN(n19287) );
  AOI211_X1 U12514 ( .C1(n16390), .C2(n16205), .A(n12830), .B(n12829), .ZN(
        n12833) );
  NAND2_X1 U12515 ( .A1(n10891), .A2(n12851), .ZN(n10057) );
  OR2_X1 U12516 ( .A1(n15013), .A2(n12778), .ZN(n16222) );
  NAND2_X1 U12517 ( .A1(n10004), .A2(n10139), .ZN(n15167) );
  NAND2_X1 U12518 ( .A1(n10331), .A2(n10141), .ZN(n10004) );
  INV_X1 U12519 ( .A(n9949), .ZN(n15179) );
  NOR2_X1 U12520 ( .A1(n9949), .A2(n15181), .ZN(n15329) );
  OAI22_X1 U12521 ( .A1(n15229), .A2(n19311), .B1(n15388), .B2(n15415), .ZN(
        n15395) );
  OAI21_X1 U12522 ( .B1(n15244), .B2(n15243), .A(n11205), .ZN(n15235) );
  OR2_X1 U12523 ( .A1(n15384), .A2(n9899), .ZN(n15405) );
  AND2_X1 U12524 ( .A1(n15386), .A2(n15385), .ZN(n9965) );
  OR2_X1 U12525 ( .A1(n10138), .A2(n10136), .ZN(n15451) );
  INV_X1 U12526 ( .A(n10322), .ZN(n10136) );
  NAND2_X1 U12527 ( .A1(n10369), .A2(n10888), .ZN(n15481) );
  NOR2_X1 U12528 ( .A1(n10371), .A2(n16344), .ZN(n10370) );
  AND2_X1 U12529 ( .A1(n11475), .A2(n11461), .ZN(n16390) );
  NOR2_X1 U12530 ( .A1(n13195), .A2(n11310), .ZN(n13494) );
  NAND2_X1 U12531 ( .A1(n10948), .A2(n10048), .ZN(n13569) );
  AND2_X1 U12532 ( .A1(n11452), .A2(n19297), .ZN(n13213) );
  INV_X1 U12533 ( .A(n16390), .ZN(n19305) );
  INV_X1 U12534 ( .A(n19316), .ZN(n19988) );
  INV_X1 U12535 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19984) );
  NOR2_X1 U12536 ( .A1(n19756), .A2(n19633), .ZN(n19974) );
  XNOR2_X1 U12537 ( .A(n13272), .B(n13271), .ZN(n19981) );
  INV_X1 U12538 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19973) );
  INV_X1 U12539 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19966) );
  XNOR2_X1 U12540 ( .A(n13337), .B(n13339), .ZN(n19963) );
  INV_X1 U12541 ( .A(n13338), .ZN(n13339) );
  INV_X1 U12542 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16426) );
  INV_X1 U12543 ( .A(n13162), .ZN(n13163) );
  NAND2_X2 U12544 ( .A1(n9941), .A2(n10595), .ZN(n16416) );
  INV_X1 U12545 ( .A(n19981), .ZN(n19447) );
  INV_X1 U12546 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13099) );
  INV_X1 U12547 ( .A(n19381), .ZN(n19384) );
  OR2_X1 U12548 ( .A1(n19396), .A2(n19546), .ZN(n19414) );
  OR2_X1 U12549 ( .A1(n19449), .A2(n19669), .ZN(n19446) );
  OR2_X1 U12550 ( .A1(n19480), .A2(n19726), .ZN(n19507) );
  INV_X1 U12551 ( .A(n19538), .ZN(n19565) );
  AOI22_X1 U12552 ( .A1(n19579), .A2(n19578), .B1(n19577), .B2(n19798), .ZN(
        n19595) );
  INV_X1 U12553 ( .A(n19624), .ZN(n19625) );
  INV_X1 U12554 ( .A(n19825), .ZN(n19732) );
  INV_X1 U12555 ( .A(n19831), .ZN(n19736) );
  INV_X1 U12556 ( .A(n19813), .ZN(n19753) );
  INV_X1 U12557 ( .A(n19819), .ZN(n19767) );
  INV_X1 U12558 ( .A(n19849), .ZN(n19785) );
  OAI21_X1 U12559 ( .B1(n19763), .B2(n19762), .A(n19761), .ZN(n19792) );
  INV_X1 U12560 ( .A(n19776), .ZN(n19790) );
  INV_X1 U12561 ( .A(n19860), .ZN(n19791) );
  AND2_X1 U12562 ( .A1(n13285), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19851) );
  NOR2_X2 U12563 ( .A1(n19543), .A2(n19727), .ZN(n19855) );
  AND3_X1 U12564 ( .A1(n15506), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19866) );
  INV_X1 U12565 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19633) );
  INV_X1 U12566 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19809) );
  INV_X2 U12567 ( .A(n20006), .ZN(n20005) );
  NAND2_X1 U12568 ( .A1(n19020), .A2(n18862), .ZN(n16651) );
  AND2_X1 U12569 ( .A1(n10234), .A2(n10229), .ZN(n16700) );
  INV_X1 U12570 ( .A(n10234), .ZN(n16713) );
  NOR2_X1 U12571 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16789), .ZN(n16782) );
  OAI21_X1 U12572 ( .B1(n16800), .B2(n10227), .A(n10229), .ZN(n10226) );
  AND2_X1 U12573 ( .A1(n10230), .A2(n10229), .ZN(n16788) );
  NOR2_X1 U12574 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16906), .ZN(n16889) );
  NOR2_X1 U12575 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16932), .ZN(n16910) );
  NOR2_X1 U12576 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16956), .ZN(n16938) );
  NOR2_X1 U12577 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16982), .ZN(n16965) );
  INV_X1 U12578 ( .A(n17026), .ZN(n16998) );
  NOR2_X2 U12579 ( .A1(n18975), .A2(n17035), .ZN(n17030) );
  OAI211_X1 U12580 ( .C1(n18877), .C2(n18870), .A(n13027), .B(n19036), .ZN(
        n17017) );
  INV_X1 U12581 ( .A(n18384), .ZN(n17371) );
  NOR2_X1 U12582 ( .A1(n16750), .A2(n17092), .ZN(n17097) );
  INV_X1 U12583 ( .A(n17168), .ZN(n17152) );
  NOR2_X1 U12584 ( .A1(n17211), .A2(n17225), .ZN(n17197) );
  NAND2_X1 U12585 ( .A1(n10106), .A2(n10104), .ZN(n18384) );
  NOR2_X1 U12586 ( .A1(n12949), .A2(n10105), .ZN(n10104) );
  INV_X1 U12587 ( .A(n12948), .ZN(n10106) );
  AND2_X1 U12588 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10105) );
  NOR3_X1 U12589 ( .A1(n17248), .A2(n15643), .A3(n17243), .ZN(n17226) );
  NAND2_X1 U12590 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17226), .ZN(n17225) );
  INV_X1 U12591 ( .A(n15552), .ZN(n17368) );
  INV_X1 U12592 ( .A(n17381), .ZN(n17376) );
  AND2_X1 U12593 ( .A1(n17399), .A2(n9843), .ZN(n17384) );
  NAND2_X1 U12594 ( .A1(n17399), .A2(n9842), .ZN(n17390) );
  INV_X1 U12595 ( .A(n17403), .ZN(n17399) );
  NAND2_X1 U12596 ( .A1(n17399), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17398) );
  NOR2_X1 U12597 ( .A1(n18384), .A2(n17408), .ZN(n17404) );
  NOR2_X1 U12598 ( .A1(n17446), .A2(n10100), .ZN(n17409) );
  INV_X1 U12599 ( .A(n17419), .ZN(n10101) );
  NAND2_X1 U12600 ( .A1(n17409), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17408) );
  NOR3_X1 U12601 ( .A1(n18384), .A2(n17566), .A3(n17446), .ZN(n17438) );
  NAND2_X1 U12602 ( .A1(n17450), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17446) );
  INV_X1 U12603 ( .A(n17402), .ZN(n17444) );
  NOR2_X1 U12604 ( .A1(n17458), .A2(n17627), .ZN(n17450) );
  NOR2_X1 U12605 ( .A1(n17372), .A2(n17371), .ZN(n17485) );
  NOR2_X1 U12606 ( .A1(n15673), .A2(n9974), .ZN(n17501) );
  OR2_X1 U12607 ( .A1(n15674), .A2(n9975), .ZN(n9974) );
  AND2_X1 U12608 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9975) );
  NAND2_X1 U12609 ( .A1(n10111), .A2(n10109), .ZN(n17510) );
  INV_X1 U12610 ( .A(n15684), .ZN(n10111) );
  NOR2_X1 U12611 ( .A1(n15685), .A2(n10110), .ZN(n10109) );
  NOR2_X1 U12612 ( .A1(n10399), .A2(n15720), .ZN(n15721) );
  INV_X1 U12613 ( .A(n17485), .ZN(n17520) );
  NOR2_X1 U12614 ( .A1(n15711), .A2(n9934), .ZN(n9933) );
  INV_X1 U12615 ( .A(n15710), .ZN(n9935) );
  NOR2_X2 U12616 ( .A1(n15919), .A2(n17372), .ZN(n17517) );
  INV_X1 U12617 ( .A(n17509), .ZN(n17518) );
  NOR2_X1 U12618 ( .A1(n19025), .A2(n17615), .ZN(n17616) );
  OAI21_X1 U12619 ( .B1(n19025), .B2(n19026), .A(n17562), .ZN(n17623) );
  CLKBUF_X1 U12620 ( .A(n17616), .Z(n17624) );
  AND2_X1 U12621 ( .A1(n17710), .A2(n9902), .ZN(n16510) );
  INV_X1 U12622 ( .A(n17635), .ZN(n10239) );
  NAND2_X1 U12623 ( .A1(n17891), .A2(n18115), .ZN(n17783) );
  NAND2_X1 U12624 ( .A1(n10235), .A2(n9828), .ZN(n17776) );
  INV_X1 U12625 ( .A(n10237), .ZN(n10235) );
  INV_X1 U12626 ( .A(n17783), .ZN(n17795) );
  NAND2_X1 U12627 ( .A1(n17894), .A2(n17831), .ZN(n17832) );
  OAI21_X1 U12628 ( .B1(n17861), .B2(n18198), .A(n10248), .ZN(n17891) );
  NAND2_X1 U12629 ( .A1(n17986), .A2(n17860), .ZN(n10248) );
  INV_X1 U12630 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17912) );
  INV_X1 U12631 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17929) );
  INV_X1 U12632 ( .A(n9937), .ZN(n17938) );
  INV_X1 U12633 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17971) );
  INV_X1 U12634 ( .A(n18680), .ZN(n18752) );
  NOR2_X1 U12635 ( .A1(n19025), .A2(n16651), .ZN(n17978) );
  NAND2_X1 U12636 ( .A1(n17995), .A2(n17830), .ZN(n17989) );
  INV_X1 U12637 ( .A(n17986), .ZN(n18000) );
  NAND2_X1 U12638 ( .A1(n10247), .A2(n10246), .ZN(n18249) );
  INV_X1 U12639 ( .A(n18316), .ZN(n10246) );
  NAND2_X1 U12640 ( .A1(n10395), .A2(n10393), .ZN(n16536) );
  AND2_X1 U12641 ( .A1(n10394), .A2(n16534), .ZN(n10393) );
  NAND2_X1 U12642 ( .A1(n17628), .A2(n10396), .ZN(n10395) );
  NAND2_X1 U12643 ( .A1(n10245), .A2(n10243), .ZN(n18316) );
  NOR2_X1 U12644 ( .A1(n18820), .A2(n10244), .ZN(n10243) );
  INV_X1 U12645 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18129) );
  INV_X1 U12646 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18142) );
  AND2_X1 U12647 ( .A1(n18112), .A2(n18288), .ZN(n18166) );
  NAND2_X1 U12648 ( .A1(n10116), .A2(n10115), .ZN(n10114) );
  AND2_X1 U12649 ( .A1(n10245), .A2(n10242), .ZN(n18224) );
  INV_X1 U12650 ( .A(n18820), .ZN(n10242) );
  INV_X1 U12651 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18237) );
  INV_X1 U12652 ( .A(n9930), .ZN(n17914) );
  NAND2_X1 U12653 ( .A1(n18293), .A2(n18294), .ZN(n18292) );
  INV_X2 U12654 ( .A(n18216), .ZN(n18330) );
  AND2_X1 U12655 ( .A1(n18979), .A2(n16647), .ZN(n19019) );
  INV_X1 U12656 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18847) );
  INV_X1 U12657 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18852) );
  INV_X1 U12658 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18856) );
  INV_X1 U12659 ( .A(n19004), .ZN(n19007) );
  INV_X1 U12660 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18368) );
  INV_X1 U12661 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18374) );
  INV_X1 U12662 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18975) );
  CLKBUF_X1 U12663 ( .A(n16631), .Z(n16637) );
  NAND2_X1 U12664 ( .A1(n14643), .A2(n20089), .ZN(n12453) );
  INV_X1 U12665 ( .A(n14643), .ZN(n14553) );
  OAI21_X1 U12666 ( .B1(n12893), .B2(n20155), .A(n9875), .ZN(P1_U2968) );
  OAI21_X1 U12667 ( .B1(n14758), .B2(n20155), .A(n9877), .ZN(P1_U2969) );
  NOR2_X1 U12668 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  INV_X1 U12669 ( .A(n12823), .ZN(n12824) );
  AND2_X1 U12670 ( .A1(n12764), .A2(n10448), .ZN(n10010) );
  NAND2_X1 U12671 ( .A1(n12725), .A2(n20169), .ZN(n12764) );
  OAI21_X1 U12672 ( .B1(n16208), .B2(n16207), .A(n10204), .ZN(P2_U2824) );
  INV_X1 U12673 ( .A(n10205), .ZN(n10204) );
  OAI21_X1 U12674 ( .B1(n16206), .B2(n19207), .A(n9876), .ZN(n10205) );
  OAI21_X1 U12675 ( .B1(n16280), .B2(n19165), .A(n10202), .ZN(n16270) );
  CLKBUF_X1 U12676 ( .A(n13529), .Z(n13481) );
  NAND2_X1 U12677 ( .A1(n11198), .A2(n9831), .ZN(n10123) );
  OR2_X1 U12678 ( .A1(n12859), .A2(n16358), .ZN(n12461) );
  OR2_X1 U12679 ( .A1(n12859), .A2(n19311), .ZN(n12860) );
  INV_X1 U12680 ( .A(n16650), .ZN(n16645) );
  OR2_X1 U12681 ( .A1(n16706), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10224) );
  AOI21_X1 U12682 ( .B1(n16499), .B2(n17859), .A(n9970), .ZN(n16500) );
  NAND2_X1 U12683 ( .A1(n9878), .A2(n9971), .ZN(n9970) );
  AOI21_X1 U12684 ( .B1(n16499), .B2(n18241), .A(n10117), .ZN(n15903) );
  OR2_X1 U12685 ( .A1(n15902), .A2(n16494), .ZN(n10117) );
  AOI21_X1 U12686 ( .B1(n18013), .B2(n18241), .A(n9931), .ZN(n18015) );
  AOI21_X1 U12687 ( .B1(n18024), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9932), .ZN(n9931) );
  OAI21_X1 U12688 ( .B1(n18012), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18315), .ZN(n9932) );
  INV_X1 U12689 ( .A(n12338), .ZN(n12717) );
  INV_X1 U12690 ( .A(n12913), .ZN(n17317) );
  INV_X1 U12691 ( .A(n16008), .ZN(n14647) );
  AND4_X1 U12692 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n9825) );
  AND2_X1 U12693 ( .A1(n9838), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9826) );
  NAND2_X2 U12694 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18824), .ZN(
        n15691) );
  INV_X2 U12695 ( .A(n9848), .ZN(n15716) );
  NOR2_X2 U12696 ( .A1(n18981), .A2(n12918), .ZN(n15607) );
  AND2_X1 U12697 ( .A1(n17831), .A2(n10238), .ZN(n9828) );
  NOR2_X1 U12698 ( .A1(n14437), .A2(n10440), .ZN(n14393) );
  NOR2_X1 U12699 ( .A1(n10381), .A2(n10380), .ZN(n15421) );
  INV_X1 U12700 ( .A(n11570), .ZN(n11646) );
  NOR2_X1 U12701 ( .A1(n14437), .A2(n10439), .ZN(n14409) );
  AND2_X1 U12702 ( .A1(n10889), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9829) );
  NAND2_X1 U12703 ( .A1(n14719), .A2(n10419), .ZN(n10191) );
  OR2_X1 U12704 ( .A1(n14523), .A2(n9888), .ZN(n14464) );
  AND4_X1 U12705 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n9830) );
  AND2_X1 U12706 ( .A1(n10133), .A2(n16356), .ZN(n9831) );
  NAND2_X1 U12708 ( .A1(n10022), .A2(n10192), .ZN(n14720) );
  AND2_X1 U12709 ( .A1(n10223), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9833) );
  AND2_X1 U12710 ( .A1(n10693), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U12711 ( .A1(n10851), .A2(n10850), .ZN(n10855) );
  AND2_X1 U12712 ( .A1(n10020), .A2(n10190), .ZN(n9835) );
  NAND2_X1 U12713 ( .A1(n10063), .A2(n9925), .ZN(n15162) );
  INV_X1 U12714 ( .A(n12696), .ZN(n10434) );
  INV_X1 U12715 ( .A(n13195), .ZN(n10260) );
  NAND2_X1 U12716 ( .A1(n13532), .A2(n13531), .ZN(n13634) );
  OR2_X1 U12717 ( .A1(n14049), .A2(n10318), .ZN(n9836) );
  AND2_X1 U12718 ( .A1(n10209), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9837) );
  AND2_X1 U12719 ( .A1(n9887), .A2(n10240), .ZN(n9838) );
  AND2_X1 U12720 ( .A1(n13593), .A2(n13361), .ZN(n9839) );
  AND2_X1 U12721 ( .A1(n10213), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9840) );
  AND2_X1 U12722 ( .A1(n10428), .A2(n13915), .ZN(n9841) );
  AND2_X1 U12723 ( .A1(n10097), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9842) );
  AND2_X1 U12724 ( .A1(n9842), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9843) );
  OR2_X1 U12725 ( .A1(n15039), .A2(n15038), .ZN(n9845) );
  AND2_X1 U12726 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10721) );
  INV_X1 U12727 ( .A(n12915), .ZN(n17158) );
  INV_X2 U12728 ( .A(n17158), .ZN(n17280) );
  NOR2_X1 U12729 ( .A1(n15229), .A2(n11455), .ZN(n15208) );
  NAND2_X1 U12730 ( .A1(n14720), .A2(n14719), .ZN(n14701) );
  OR2_X1 U12731 ( .A1(n12921), .A2(n13029), .ZN(n9846) );
  AND2_X1 U12732 ( .A1(n10862), .A2(n10373), .ZN(n9847) );
  OR2_X1 U12733 ( .A1(n12920), .A2(n15645), .ZN(n9848) );
  NOR2_X1 U12734 ( .A1(n15229), .A2(n10375), .ZN(n11473) );
  AND3_X2 U12735 ( .A1(n10892), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10716) );
  CLKBUF_X3 U12736 ( .A(n10716), .Z(n14276) );
  NOR2_X1 U12737 ( .A1(n12985), .A2(n10249), .ZN(n9849) );
  OR2_X1 U12738 ( .A1(n12921), .A2(n12920), .ZN(n9850) );
  NAND2_X1 U12739 ( .A1(n10973), .A2(n10972), .ZN(n13982) );
  OR2_X1 U12740 ( .A1(n14943), .A2(n10359), .ZN(n9851) );
  OR2_X1 U12741 ( .A1(n15422), .A2(n16292), .ZN(n9852) );
  OR3_X1 U12742 ( .A1(n11046), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n10938), .ZN(
        n9853) );
  NAND2_X1 U12743 ( .A1(n12059), .A2(n12058), .ZN(n14423) );
  OR2_X1 U12744 ( .A1(n14523), .A2(n14600), .ZN(n14518) );
  NOR2_X1 U12745 ( .A1(n15422), .A2(n10065), .ZN(n15172) );
  NAND2_X1 U12746 ( .A1(n15142), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12775) );
  NAND2_X1 U12747 ( .A1(n16025), .A2(n13886), .ZN(n16026) );
  NOR2_X1 U12748 ( .A1(n15229), .A2(n10377), .ZN(n9854) );
  OR2_X1 U12749 ( .A1(n10381), .A2(n10382), .ZN(n9855) );
  NOR2_X1 U12750 ( .A1(n11780), .A2(n11734), .ZN(n9856) );
  AND2_X1 U12751 ( .A1(n17399), .A2(n10097), .ZN(n9857) );
  AND2_X1 U12752 ( .A1(n11611), .A2(n11554), .ZN(n11621) );
  NOR2_X1 U12753 ( .A1(n14523), .A2(n10425), .ZN(n9858) );
  AND2_X1 U12754 ( .A1(n15747), .A2(n15791), .ZN(n9859) );
  AND2_X1 U12755 ( .A1(n10978), .A2(n10975), .ZN(n9860) );
  INV_X2 U12756 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16411) );
  XNOR2_X1 U12757 ( .A(n14204), .B(n14202), .ZN(n14939) );
  NAND2_X1 U12758 ( .A1(n14969), .A2(n10313), .ZN(n14955) );
  INV_X1 U12759 ( .A(n17922), .ZN(n15806) );
  INV_X1 U12760 ( .A(n13511), .ZN(n12346) );
  OR2_X1 U12761 ( .A1(n14289), .A2(n19158), .ZN(n9861) );
  INV_X1 U12762 ( .A(n11610), .ZN(n11634) );
  AND2_X1 U12763 ( .A1(n11008), .A2(n10294), .ZN(n9862) );
  AND2_X2 U12764 ( .A1(n10005), .A2(n11486), .ZN(n11559) );
  AND4_X1 U12765 ( .A1(n10814), .A2(n10812), .A3(n10811), .A4(n10813), .ZN(
        n9863) );
  NAND2_X1 U12766 ( .A1(n18831), .A2(n15768), .ZN(n18826) );
  INV_X1 U12767 ( .A(n18826), .ZN(n10247) );
  AND4_X1 U12768 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9864) );
  AND3_X1 U12769 ( .A1(n12987), .A2(n10251), .A3(n10250), .ZN(n9865) );
  AND4_X1 U12770 ( .A1(n11632), .A2(n12728), .A3(n13778), .A4(n11623), .ZN(
        n9866) );
  OR2_X1 U12771 ( .A1(n17317), .A2(n10402), .ZN(n9867) );
  AND2_X1 U12772 ( .A1(n16209), .A2(n10206), .ZN(n9868) );
  NOR3_X1 U12773 ( .A1(n11073), .A2(n11326), .A3(n12851), .ZN(n9869) );
  NOR2_X1 U12774 ( .A1(n13176), .A2(n10594), .ZN(n10621) );
  INV_X1 U12775 ( .A(n10142), .ZN(n10141) );
  OAI21_X1 U12776 ( .B1(n10332), .B2(n10143), .A(n11047), .ZN(n10142) );
  AND2_X1 U12777 ( .A1(n10492), .A2(n19339), .ZN(n9870) );
  AND2_X1 U12778 ( .A1(n10061), .A2(n10060), .ZN(n9871) );
  INV_X1 U12779 ( .A(n17860), .ZN(n18196) );
  NAND2_X1 U12780 ( .A1(n17899), .A2(n15763), .ZN(n17860) );
  OR2_X1 U12781 ( .A1(n10888), .A2(n11453), .ZN(n9872) );
  NAND2_X1 U12782 ( .A1(n13283), .A2(n13282), .ZN(n13337) );
  AND2_X1 U12783 ( .A1(n15810), .A2(n17922), .ZN(n9873) );
  INV_X1 U12784 ( .A(n11684), .ZN(n10424) );
  AOI22_X1 U12785 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11683), .B2(n11682), .ZN(n11684) );
  NAND2_X1 U12786 ( .A1(n11634), .A2(n11570), .ZN(n11608) );
  AND2_X2 U12787 ( .A1(n13397), .A2(n11486), .ZN(n11598) );
  INV_X1 U12788 ( .A(n18345), .ZN(n15915) );
  OAI211_X1 U12789 ( .C1(n17287), .C2(n18685), .A(n12939), .B(n12938), .ZN(
        n18345) );
  NOR2_X1 U12790 ( .A1(n15178), .A2(n15324), .ZN(n9874) );
  AND2_X1 U12791 ( .A1(n12895), .A2(n12894), .ZN(n9875) );
  INV_X1 U12792 ( .A(n10191), .ZN(n10190) );
  AND2_X1 U12793 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13887) );
  AND2_X1 U12794 ( .A1(n10207), .A2(n9868), .ZN(n9876) );
  AND2_X1 U12795 ( .A1(n12850), .A2(n12849), .ZN(n9877) );
  NAND3_X1 U12796 ( .A1(n16517), .A2(n16493), .A3(n17652), .ZN(n9878) );
  INV_X1 U12797 ( .A(n10298), .ZN(n14921) );
  OR2_X1 U12798 ( .A1(n10961), .A2(n13874), .ZN(n10860) );
  AND3_X1 U12799 ( .A1(n11528), .A2(n11521), .A3(n11523), .ZN(n9879) );
  AND2_X1 U12800 ( .A1(n10133), .A2(n10125), .ZN(n9880) );
  AND2_X1 U12801 ( .A1(n15701), .A2(n15700), .ZN(n15793) );
  INV_X1 U12802 ( .A(n15793), .ZN(n10112) );
  AND2_X1 U12803 ( .A1(n10702), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9881) );
  AND2_X1 U12804 ( .A1(n10424), .A2(n16196), .ZN(n9882) );
  AND2_X1 U12805 ( .A1(n11088), .A2(n10660), .ZN(n9883) );
  AND2_X1 U12806 ( .A1(n10860), .A2(n10144), .ZN(n9884) );
  AND2_X1 U12807 ( .A1(n9997), .A2(n10825), .ZN(n10826) );
  INV_X1 U12808 ( .A(n10826), .ZN(n9946) );
  AND2_X1 U12809 ( .A1(n10351), .A2(n13641), .ZN(n9885) );
  INV_X1 U12810 ( .A(n12767), .ZN(n10329) );
  AND2_X1 U12811 ( .A1(n16232), .A2(n11078), .ZN(n12767) );
  NAND2_X1 U12812 ( .A1(n10041), .A2(n9872), .ZN(n10889) );
  INV_X1 U12813 ( .A(n10889), .ZN(n10381) );
  BUF_X1 U12814 ( .A(n11535), .Z(n12235) );
  INV_X1 U12815 ( .A(n11291), .ZN(n11329) );
  AND3_X1 U12816 ( .A1(n11295), .A2(n14227), .A3(n11265), .ZN(n11327) );
  INV_X1 U12817 ( .A(n12500), .ZN(n10222) );
  NAND2_X1 U12818 ( .A1(n11901), .A2(n11900), .ZN(n13730) );
  AND2_X1 U12819 ( .A1(n12507), .A2(n10209), .ZN(n9886) );
  AND3_X1 U12820 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9887) );
  OAI21_X1 U12821 ( .B1(n15236), .B2(n10079), .A(n11207), .ZN(n10078) );
  OR2_X1 U12822 ( .A1(n14520), .A2(n14600), .ZN(n9888) );
  NAND2_X1 U12823 ( .A1(n13962), .A2(n10862), .ZN(n13978) );
  OR3_X1 U12824 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17717), .ZN(n9889) );
  OR2_X1 U12825 ( .A1(n11052), .A2(n12790), .ZN(n9890) );
  AND2_X1 U12826 ( .A1(n13269), .A2(n13219), .ZN(n13272) );
  INV_X1 U12827 ( .A(n13979), .ZN(n10371) );
  INV_X1 U12828 ( .A(n13726), .ZN(n10347) );
  NAND2_X1 U12829 ( .A1(n13095), .A2(n11228), .ZN(n11439) );
  OR2_X1 U12830 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13886) );
  INV_X1 U12831 ( .A(n13886), .ZN(n10155) );
  AND2_X1 U12832 ( .A1(n10321), .A2(n13676), .ZN(n9891) );
  AND2_X1 U12833 ( .A1(n10264), .A2(n13832), .ZN(n9892) );
  OR2_X1 U12834 ( .A1(n18204), .A2(n17884), .ZN(n9893) );
  AND2_X1 U12835 ( .A1(n16337), .A2(n16338), .ZN(n9894) );
  INV_X1 U12836 ( .A(n10989), .ZN(n10324) );
  AND2_X1 U12837 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9895) );
  OR2_X1 U12838 ( .A1(n18010), .A2(n18027), .ZN(n9896) );
  AND2_X1 U12839 ( .A1(n16366), .A2(n10261), .ZN(n11425) );
  INV_X1 U12840 ( .A(n14439), .ZN(n12058) );
  INV_X1 U12841 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13984) );
  OR2_X1 U12842 ( .A1(n15466), .A2(n15482), .ZN(n9897) );
  INV_X1 U12843 ( .A(n10905), .ZN(n11317) );
  OR2_X1 U12844 ( .A1(n10796), .A2(n10795), .ZN(n10905) );
  OR2_X1 U12845 ( .A1(n13713), .A2(n13577), .ZN(n9898) );
  OR2_X1 U12846 ( .A1(n15409), .A2(n9965), .ZN(n9899) );
  NOR2_X1 U12847 ( .A1(n9856), .A2(n9812), .ZN(n9900) );
  OR2_X1 U12848 ( .A1(n15449), .A2(n15454), .ZN(n9901) );
  AND2_X1 U12849 ( .A1(n9826), .A2(n10239), .ZN(n9902) );
  AND2_X1 U12850 ( .A1(n10442), .A2(n10443), .ZN(n9903) );
  INV_X1 U12851 ( .A(n10078), .ZN(n10077) );
  INV_X1 U12852 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16311) );
  NAND2_X1 U12853 ( .A1(n15767), .A2(n19034), .ZN(n18835) );
  INV_X1 U12854 ( .A(n18835), .ZN(n10244) );
  NAND2_X2 U12855 ( .A1(n12526), .A2(n13145), .ZN(n9942) );
  NAND2_X1 U12856 ( .A1(n13594), .A2(n13593), .ZN(n13358) );
  NAND2_X1 U12857 ( .A1(n10342), .A2(n10340), .ZN(n13297) );
  INV_X1 U12858 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16196) );
  AND2_X1 U12859 ( .A1(n11081), .A2(n14957), .ZN(n19291) );
  AND2_X1 U12860 ( .A1(n10279), .A2(n11430), .ZN(n9904) );
  AND2_X1 U12861 ( .A1(n9904), .A2(n10278), .ZN(n9905) );
  AND2_X1 U12862 ( .A1(n10342), .A2(n10337), .ZN(n13363) );
  AND2_X1 U12863 ( .A1(n13363), .A2(n13447), .ZN(n13446) );
  AND2_X1 U12864 ( .A1(n14959), .A2(n14970), .ZN(n9906) );
  NAND2_X1 U12865 ( .A1(n11778), .A2(n11777), .ZN(n20336) );
  INV_X1 U12866 ( .A(n20336), .ZN(n10037) );
  INV_X1 U12867 ( .A(n14994), .ZN(n10335) );
  OR3_X1 U12868 ( .A1(n10465), .A2(n14956), .A3(n14157), .ZN(n9907) );
  AND2_X1 U12869 ( .A1(n13532), .A2(n9891), .ZN(n13723) );
  AND2_X1 U12870 ( .A1(n10698), .A2(n10702), .ZN(n10828) );
  OR2_X1 U12871 ( .A1(n12521), .A2(n12491), .ZN(n9908) );
  AND2_X1 U12872 ( .A1(n10089), .A2(n10088), .ZN(n9909) );
  AND2_X1 U12873 ( .A1(n10302), .A2(n14929), .ZN(n9910) );
  OAI211_X1 U12874 ( .C1(n11520), .C2(n11951), .A(n11519), .B(n11518), .ZN(
        n13915) );
  AND2_X1 U12875 ( .A1(n10305), .A2(n10302), .ZN(n9911) );
  INV_X1 U12876 ( .A(n12258), .ZN(n11614) );
  NOR2_X1 U12877 ( .A1(n14542), .A2(n14536), .ZN(n12370) );
  AND2_X1 U12878 ( .A1(n10225), .A2(n10228), .ZN(n9912) );
  OR2_X1 U12879 ( .A1(n10363), .A2(n10361), .ZN(n9913) );
  AND2_X1 U12880 ( .A1(n10256), .A2(n13493), .ZN(n9914) );
  INV_X1 U12881 ( .A(n19152), .ZN(n19165) );
  NAND2_X1 U12882 ( .A1(n12515), .A2(n10213), .ZN(n10215) );
  NAND2_X1 U12883 ( .A1(n11721), .A2(n11570), .ZN(n12712) );
  NAND2_X1 U12884 ( .A1(n10342), .A2(n10336), .ZN(n10344) );
  AND3_X1 U12885 ( .A1(n10436), .A2(n10435), .A3(n12730), .ZN(n9915) );
  AND2_X1 U12886 ( .A1(n10260), .A2(n10259), .ZN(n9916) );
  OR2_X1 U12887 ( .A1(n13483), .A2(n10352), .ZN(n10357) );
  OR2_X1 U12888 ( .A1(n10603), .A2(n10602), .ZN(n11091) );
  AND2_X1 U12889 ( .A1(n9905), .A2(n10277), .ZN(n9917) );
  INV_X1 U12890 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15175) );
  XNOR2_X1 U12891 ( .A(n19025), .B(n15915), .ZN(n19034) );
  INV_X1 U12892 ( .A(n19034), .ZN(n10241) );
  AND2_X1 U12893 ( .A1(n17710), .A2(n9838), .ZN(n9918) );
  AND3_X1 U12894 ( .A1(n15831), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n9919) );
  OR2_X1 U12895 ( .A1(n18029), .A2(n18034), .ZN(n9920) );
  AND2_X1 U12896 ( .A1(n10276), .A2(n15014), .ZN(n9921) );
  NAND2_X1 U12897 ( .A1(n10459), .A2(n10398), .ZN(n9922) );
  INV_X1 U12898 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n10158) );
  INV_X1 U12899 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n10164) );
  INV_X1 U12900 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n10167) );
  INV_X1 U12901 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n10161) );
  INV_X1 U12902 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10398) );
  AND2_X1 U12903 ( .A1(n9828), .A2(n17894), .ZN(n9923) );
  AND2_X1 U12904 ( .A1(n10038), .A2(n15889), .ZN(n9924) );
  AND2_X1 U12905 ( .A1(n10064), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9925) );
  AND2_X1 U12906 ( .A1(n10374), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9926) );
  INV_X1 U12907 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10098) );
  INV_X1 U12908 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n10099) );
  INV_X1 U12909 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10211) );
  INV_X1 U12910 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10218) );
  INV_X1 U12911 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10402) );
  INV_X1 U12912 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10219) );
  AOI22_X2 U12913 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20224), .B1(DATAI_26_), 
        .B2(n20225), .ZN(n20642) );
  NOR3_X2 U12914 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18745), .A3(
        n18416), .ZN(n18411) );
  NOR3_X2 U12915 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18745), .A3(
        n18652), .ZN(n18594) );
  NOR3_X2 U12916 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18745), .A3(
        n18508), .ZN(n18502) );
  AOI22_X2 U12917 ( .A1(DATAI_31_), .A2(n20225), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20224), .ZN(n20765) );
  NOR2_X1 U12918 ( .A1(n19339), .A2(n19351), .ZN(n9927) );
  NAND2_X1 U12919 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19807), .ZN(n19351) );
  INV_X2 U12920 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18992) );
  INV_X2 U12921 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18999) );
  AND2_X2 U12922 ( .A1(n9939), .A2(n10662), .ZN(n11088) );
  NAND2_X1 U12923 ( .A1(n10669), .A2(n10674), .ZN(n9939) );
  NAND2_X1 U12924 ( .A1(n9942), .A2(n14957), .ZN(n11263) );
  NAND2_X1 U12925 ( .A1(n13083), .A2(n9942), .ZN(n13084) );
  NAND3_X1 U12926 ( .A1(n13081), .A2(n13043), .A3(n9942), .ZN(n13044) );
  NAND2_X1 U12927 ( .A1(n13038), .A2(n9942), .ZN(n19043) );
  NOR2_X1 U12928 ( .A1(n9943), .A2(n9941), .ZN(n9940) );
  NAND2_X1 U12929 ( .A1(n10853), .A2(n9944), .ZN(n10970) );
  NOR2_X1 U12930 ( .A1(n10855), .A2(n9946), .ZN(n9945) );
  NAND4_X1 U12931 ( .A1(n10713), .A2(n10711), .A3(n10714), .A4(n10712), .ZN(
        n9948) );
  OAI21_X2 U12933 ( .B1(n10137), .B2(n10138), .A(n9996), .ZN(n15439) );
  NAND2_X1 U12934 ( .A1(n10683), .A2(n10702), .ZN(n19419) );
  NAND2_X2 U12935 ( .A1(n9953), .A2(n11658), .ZN(n11667) );
  NAND2_X1 U12936 ( .A1(n20364), .A2(n9953), .ZN(n13426) );
  NAND2_X1 U12937 ( .A1(n11686), .A2(n11685), .ZN(n9953) );
  INV_X1 U12938 ( .A(n11608), .ZN(n11558) );
  NAND2_X2 U12939 ( .A1(n9832), .A2(n9825), .ZN(n11570) );
  NAND3_X1 U12940 ( .A1(n10030), .A2(n16035), .A3(n9958), .ZN(n9957) );
  AND2_X2 U12941 ( .A1(n10005), .A2(n13382), .ZN(n11542) );
  AND2_X2 U12942 ( .A1(n11479), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13382) );
  NAND3_X1 U12943 ( .A1(n10021), .A2(n10019), .A3(n10020), .ZN(n10018) );
  NAND3_X1 U12944 ( .A1(n12688), .A2(n14684), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U12945 ( .A1(n9963), .A2(n13979), .ZN(n16343) );
  NAND2_X1 U12946 ( .A1(n9963), .A2(n10370), .ZN(n10369) );
  OAI21_X1 U12947 ( .B1(n10797), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n9968), .ZN(n9966) );
  NAND2_X1 U12948 ( .A1(n10785), .A2(n10784), .ZN(n9968) );
  NAND2_X1 U12949 ( .A1(n9968), .A2(n10797), .ZN(n13659) );
  NAND2_X1 U12950 ( .A1(n9967), .A2(n10798), .ZN(n13660) );
  INV_X1 U12951 ( .A(n9968), .ZN(n9967) );
  NAND3_X1 U12952 ( .A1(n15247), .A2(n15229), .A3(n10925), .ZN(n15248) );
  INV_X2 U12953 ( .A(n10678), .ZN(n10802) );
  XNOR2_X2 U12954 ( .A(n9800), .B(n10786), .ZN(n13574) );
  XNOR2_X2 U12955 ( .A(n15818), .B(n18237), .ZN(n18243) );
  NAND3_X1 U12956 ( .A1(n10388), .A2(n10387), .A3(n10391), .ZN(n17910) );
  NOR2_X4 U12957 ( .A1(n16533), .A2(n17494), .ZN(n17793) );
  NAND4_X2 U12958 ( .A1(n18992), .A2(n18999), .A3(n18981), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17306) );
  INV_X2 U12959 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18981) );
  NAND2_X1 U12960 ( .A1(n10587), .A2(n11441), .ZN(n11245) );
  NAND2_X1 U12961 ( .A1(n19323), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9978) );
  NAND2_X1 U12962 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n9979) );
  NAND2_X1 U12963 ( .A1(n10683), .A2(n9881), .ZN(n9983) );
  NAND4_X1 U12964 ( .A1(n9981), .A2(n9980), .A3(n10759), .A4(n10756), .ZN(
        n10367) );
  NAND4_X1 U12965 ( .A1(n9991), .A2(n9990), .A3(n9989), .A4(n9988), .ZN(n9987)
         );
  INV_X1 U12966 ( .A(n14957), .ZN(n9992) );
  NAND3_X1 U12967 ( .A1(n10281), .A2(n11064), .A3(n12766), .ZN(n15127) );
  OAI21_X2 U12968 ( .B1(n10331), .B2(n10002), .A(n10000), .ZN(n15153) );
  INV_X1 U12969 ( .A(n15153), .ZN(n10330) );
  AND2_X2 U12970 ( .A1(n10139), .A2(n9890), .ZN(n10003) );
  AND2_X2 U12971 ( .A1(n10005), .A2(n11488), .ZN(n11703) );
  NOR2_X1 U12972 ( .A1(n12575), .A2(n10404), .ZN(n13315) );
  INV_X1 U12973 ( .A(n10404), .ZN(n10006) );
  INV_X1 U12974 ( .A(n12575), .ZN(n10007) );
  NAND2_X1 U12975 ( .A1(n10008), .A2(n11644), .ZN(n11653) );
  NAND2_X1 U12976 ( .A1(n10146), .A2(n10009), .ZN(n10008) );
  OAI21_X1 U12977 ( .B1(n11659), .B2(n10198), .A(n11629), .ZN(n11758) );
  OAI21_X1 U12978 ( .B1(n12893), .B2(n20176), .A(n10010), .ZN(P1_U3000) );
  NAND2_X1 U12979 ( .A1(n10012), .A2(n10148), .ZN(n10011) );
  NAND2_X1 U12980 ( .A1(n10405), .A2(n10422), .ZN(n10017) );
  NAND3_X1 U12981 ( .A1(n10409), .A2(n13416), .A3(n9882), .ZN(n10016) );
  NAND2_X1 U12982 ( .A1(n12684), .A2(n10027), .ZN(n10022) );
  AND2_X2 U12983 ( .A1(n13382), .A2(n13397), .ZN(n11592) );
  AND2_X2 U12984 ( .A1(n11487), .A2(n13382), .ZN(n11529) );
  NAND2_X1 U12985 ( .A1(n10033), .A2(n10031), .ZN(n10030) );
  NAND2_X1 U12986 ( .A1(n11667), .A2(n11666), .ZN(n13416) );
  NAND2_X1 U12987 ( .A1(n11667), .A2(n10035), .ZN(n10034) );
  NAND2_X1 U12988 ( .A1(n10410), .A2(n20336), .ZN(n10036) );
  XNOR2_X1 U12989 ( .A(n10040), .B(n10905), .ZN(n10797) );
  NAND2_X1 U12990 ( .A1(n10948), .A2(n10045), .ZN(n10043) );
  NAND2_X1 U12991 ( .A1(n10043), .A2(n10044), .ZN(n13657) );
  NAND2_X1 U12992 ( .A1(n10051), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13568) );
  NAND2_X1 U12993 ( .A1(n15121), .A2(n10056), .ZN(n10052) );
  NAND3_X1 U12994 ( .A1(n10055), .A2(n10057), .A3(n10052), .ZN(n12837) );
  NAND2_X1 U12995 ( .A1(n15439), .A2(n10060), .ZN(n10059) );
  INV_X1 U12996 ( .A(n15439), .ZN(n10062) );
  INV_X1 U12997 ( .A(n15422), .ZN(n10063) );
  OR2_X1 U12998 ( .A1(n15253), .A2(n11203), .ZN(n10069) );
  NAND2_X1 U12999 ( .A1(n10068), .A2(n10070), .ZN(n15203) );
  NAND3_X1 U13000 ( .A1(n15253), .A2(n10077), .A3(n15251), .ZN(n10068) );
  NOR2_X1 U13001 ( .A1(n14317), .A2(n12864), .ZN(n10083) );
  INV_X1 U13002 ( .A(n13512), .ZN(n10091) );
  AND3_X2 U13003 ( .A1(n10091), .A2(n12346), .A3(n10093), .ZN(n16162) );
  NAND3_X1 U13004 ( .A1(n10101), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_17__SCAN_IN), .ZN(n10100) );
  NOR3_X2 U13005 ( .A1(n17688), .A2(n18002), .A3(n17698), .ZN(n17676) );
  NAND2_X1 U13006 ( .A1(n17744), .A2(n17728), .ZN(n17729) );
  NAND2_X1 U13007 ( .A1(n17792), .A2(n18120), .ZN(n17728) );
  NAND2_X1 U13008 ( .A1(n10108), .A2(n9889), .ZN(n10107) );
  NAND2_X1 U13009 ( .A1(n15822), .A2(n15820), .ZN(n17792) );
  NAND2_X2 U13010 ( .A1(n17779), .A2(n17902), .ZN(n17744) );
  AND2_X1 U13011 ( .A1(n10114), .A2(n9893), .ZN(n17858) );
  NOR2_X1 U13012 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10115) );
  INV_X1 U13013 ( .A(n17883), .ZN(n10116) );
  INV_X1 U13014 ( .A(n10386), .ZN(n10392) );
  NAND2_X1 U13015 ( .A1(n15811), .A2(n15807), .ZN(n10386) );
  INV_X2 U13016 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19006) );
  NAND3_X2 U13017 ( .A1(n10646), .A2(n10119), .A3(n10118), .ZN(n13579) );
  NAND2_X1 U13018 ( .A1(n10468), .A2(n11088), .ZN(n10118) );
  NAND2_X1 U13019 ( .A1(n10613), .A2(n11090), .ZN(n10120) );
  NAND2_X1 U13020 ( .A1(n12454), .A2(n10128), .ZN(n10127) );
  NAND2_X1 U13021 ( .A1(n10130), .A2(n10121), .ZN(n12826) );
  NAND3_X1 U13022 ( .A1(n10130), .A2(n10127), .A3(n10122), .ZN(n10124) );
  AND2_X1 U13023 ( .A1(n10124), .A2(n10123), .ZN(P2_U2983) );
  NAND2_X1 U13024 ( .A1(n10322), .A2(n9901), .ZN(n10137) );
  NAND2_X1 U13025 ( .A1(n10861), .A2(n10144), .ZN(n10862) );
  NAND4_X1 U13026 ( .A1(n9866), .A2(n11645), .A3(n10147), .A4(n11648), .ZN(
        n10146) );
  INV_X1 U13027 ( .A(n11628), .ZN(n10147) );
  AND2_X2 U13028 ( .A1(n11615), .A2(n12572), .ZN(n11645) );
  NAND2_X1 U13029 ( .A1(n11843), .A2(n11844), .ZN(n11873) );
  NAND2_X1 U13030 ( .A1(n10149), .A2(n12648), .ZN(n12649) );
  NAND3_X1 U13031 ( .A1(n10150), .A2(n12695), .A3(n11873), .ZN(n10149) );
  NAND2_X1 U13032 ( .A1(n11846), .A2(n11845), .ZN(n10150) );
  NAND3_X1 U13033 ( .A1(n12677), .A2(n10416), .A3(n12678), .ZN(n10152) );
  NAND2_X1 U13034 ( .A1(n10152), .A2(n10153), .ZN(n12687) );
  NAND2_X2 U13035 ( .A1(n12327), .A2(n10184), .ZN(n12341) );
  OR2_X1 U13036 ( .A1(n9816), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12329) );
  OR2_X1 U13037 ( .A1(n12413), .A2(n20995), .ZN(n12334) );
  OR2_X1 U13038 ( .A1(n12413), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12383) );
  OR2_X1 U13039 ( .A1(n12413), .A2(n10158), .ZN(n10156) );
  OR2_X1 U13040 ( .A1(n12413), .A2(n10161), .ZN(n10159) );
  OR2_X1 U13041 ( .A1(n12413), .A2(n10164), .ZN(n10162) );
  OR2_X1 U13042 ( .A1(n9816), .A2(n10167), .ZN(n10165) );
  OR2_X1 U13043 ( .A1(n9816), .A2(n21168), .ZN(n10168) );
  OR2_X1 U13044 ( .A1(n9816), .A2(n21212), .ZN(n10170) );
  OAI21_X1 U13045 ( .B1(n13172), .B2(n14673), .A(n10184), .ZN(n10173) );
  OAI21_X1 U13046 ( .B1(n13172), .B2(n16168), .A(n10184), .ZN(n10175) );
  OAI21_X1 U13047 ( .B1(n13172), .B2(n16179), .A(n10184), .ZN(n10177) );
  OAI21_X1 U13048 ( .B1(n13172), .B2(n16157), .A(n10184), .ZN(n10179) );
  OAI21_X1 U13049 ( .B1(n13172), .B2(n12742), .A(n10184), .ZN(n10181) );
  OAI21_X1 U13050 ( .B1(n13172), .B2(n16049), .A(n10184), .ZN(n10183) );
  NAND2_X1 U13051 ( .A1(n13510), .A2(n13509), .ZN(n12642) );
  NAND2_X1 U13052 ( .A1(n12632), .A2(n12695), .ZN(n10185) );
  NAND2_X1 U13053 ( .A1(n13463), .A2(n13464), .ZN(n10186) );
  NAND2_X1 U13054 ( .A1(n13620), .A2(n13619), .ZN(n10188) );
  INV_X1 U13055 ( .A(n12659), .ZN(n10189) );
  INV_X1 U13056 ( .A(n13426), .ZN(n10197) );
  NAND2_X1 U13057 ( .A1(n13426), .A2(n9900), .ZN(n10193) );
  AOI21_X2 U13058 ( .B1(n10197), .B2(n16196), .A(n9856), .ZN(n12605) );
  OAI211_X1 U13059 ( .C1(n10199), .C2(n15844), .A(n15843), .B(n19108), .ZN(
        n15845) );
  AOI21_X4 U13060 ( .B1(n12488), .B2(n19863), .A(n12487), .ZN(n19152) );
  NAND2_X1 U13061 ( .A1(n16280), .A2(n10201), .ZN(n10200) );
  NAND2_X1 U13062 ( .A1(n10200), .A2(n19152), .ZN(n16259) );
  INV_X1 U13063 ( .A(n10215), .ZN(n12520) );
  NAND3_X1 U13064 ( .A1(n16698), .A2(n16697), .A3(n10224), .ZN(P3_U2641) );
  NAND2_X1 U13065 ( .A1(n16800), .A2(n17001), .ZN(n10225) );
  INV_X1 U13066 ( .A(n10226), .ZN(n16781) );
  INV_X1 U13067 ( .A(n10228), .ZN(n10227) );
  INV_X1 U13068 ( .A(n10230), .ZN(n16799) );
  INV_X1 U13069 ( .A(n16975), .ZN(n10229) );
  INV_X1 U13070 ( .A(n18249), .ZN(n18144) );
  NAND3_X1 U13071 ( .A1(n10260), .A2(n10259), .A3(n13794), .ZN(n13793) );
  AND2_X1 U13072 ( .A1(n15031), .A2(n10275), .ZN(n12827) );
  NAND3_X1 U13073 ( .A1(n10273), .A2(n10271), .A3(n10270), .ZN(n16204) );
  NAND2_X1 U13074 ( .A1(n15031), .A2(n10272), .ZN(n10271) );
  OR2_X1 U13075 ( .A1(n15031), .A2(n10274), .ZN(n10273) );
  AND2_X2 U13076 ( .A1(n15031), .A2(n12777), .ZN(n15013) );
  AND2_X2 U13077 ( .A1(n15084), .A2(n9917), .ZN(n15309) );
  NAND2_X1 U13078 ( .A1(n15144), .A2(n15151), .ZN(n11053) );
  INV_X1 U13079 ( .A(n11053), .ZN(n10280) );
  NAND3_X1 U13080 ( .A1(n10330), .A2(n10280), .A3(n12767), .ZN(n12766) );
  NAND2_X1 U13081 ( .A1(n12769), .A2(n15264), .ZN(n10281) );
  NAND2_X1 U13082 ( .A1(n10980), .A2(n10284), .ZN(n10981) );
  NAND2_X1 U13083 ( .A1(n19124), .A2(n10285), .ZN(n11025) );
  NAND2_X1 U13084 ( .A1(n11008), .A2(n10292), .ZN(n10996) );
  INV_X1 U13085 ( .A(n14228), .ZN(n10303) );
  OAI211_X1 U13086 ( .C1(n14935), .C2(n10307), .A(n10304), .B(n10463), .ZN(
        n14286) );
  XNOR2_X2 U13087 ( .A(n14228), .B(n14229), .ZN(n14935) );
  AOI21_X2 U13088 ( .B1(n14968), .B2(n9906), .A(n10311), .ZN(n14178) );
  OAI21_X2 U13089 ( .B1(n10313), .B2(n10312), .A(n9907), .ZN(n10311) );
  INV_X1 U13090 ( .A(n14138), .ZN(n14976) );
  INV_X1 U13091 ( .A(n10465), .ZN(n10314) );
  NOR2_X2 U13092 ( .A1(n14049), .A2(n10315), .ZN(n14986) );
  NAND2_X2 U13093 ( .A1(n13295), .A2(n13294), .ZN(n13594) );
  NOR2_X4 U13094 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U13095 ( .A1(n11053), .A2(n10329), .ZN(n10326) );
  NAND2_X1 U13096 ( .A1(n10326), .A2(n12765), .ZN(n10328) );
  OR2_X2 U13097 ( .A1(n14995), .A2(n11459), .ZN(n14980) );
  INV_X1 U13098 ( .A(n10344), .ZN(n13299) );
  INV_X1 U13099 ( .A(n13483), .ZN(n10350) );
  NAND2_X1 U13100 ( .A1(n10350), .A2(n9885), .ZN(n13673) );
  INV_X1 U13101 ( .A(n10357), .ZN(n13640) );
  NOR2_X1 U13102 ( .A1(n14943), .A2(n14932), .ZN(n12785) );
  INV_X1 U13103 ( .A(n12784), .ZN(n10363) );
  OAI22_X1 U13104 ( .A1(n13869), .A2(n10364), .B1(n13871), .B2(n13870), .ZN(
        n16359) );
  AND2_X4 U13105 ( .A1(n10365), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10509) );
  NOR2_X1 U13106 ( .A1(n10721), .A2(n10365), .ZN(n15517) );
  INV_X1 U13107 ( .A(n10366), .ZN(n10593) );
  NOR2_X1 U13108 ( .A1(n10366), .A2(n13930), .ZN(n13931) );
  NOR2_X1 U13109 ( .A1(n13926), .A2(n10366), .ZN(n10579) );
  NOR2_X1 U13110 ( .A1(n19315), .A2(n10366), .ZN(n13929) );
  NOR2_X2 U13111 ( .A1(n10572), .A2(n10366), .ZN(n13097) );
  NAND2_X1 U13112 ( .A1(n13574), .A2(n13572), .ZN(n10785) );
  NAND2_X1 U13113 ( .A1(n10889), .A2(n10379), .ZN(n15422) );
  AND2_X2 U13114 ( .A1(n15154), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15142) );
  OR2_X1 U13115 ( .A1(n17921), .A2(n10386), .ZN(n10387) );
  NAND2_X1 U13116 ( .A1(n17921), .A2(n17922), .ZN(n17920) );
  NAND2_X1 U13117 ( .A1(n10392), .A2(n15806), .ZN(n10389) );
  NAND2_X1 U13118 ( .A1(n17920), .A2(n15807), .ZN(n17790) );
  NAND2_X1 U13119 ( .A1(n17647), .A2(n16541), .ZN(n17629) );
  OAI21_X1 U13120 ( .B1(n17850), .B2(n9922), .A(n17902), .ZN(n15822) );
  NOR2_X1 U13121 ( .A1(n17850), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17812) );
  XNOR2_X1 U13122 ( .A(n15792), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18294) );
  XNOR2_X1 U13123 ( .A(n15791), .B(n15793), .ZN(n15792) );
  NAND4_X1 U13124 ( .A1(n10401), .A2(n15718), .A3(n10403), .A4(n10400), .ZN(
        n10399) );
  AND3_X1 U13125 ( .A1(n15719), .A2(n15717), .A3(n9867), .ZN(n10400) );
  NAND2_X1 U13126 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13127 ( .A1(n11613), .A2(n11612), .ZN(n10404) );
  NAND2_X1 U13128 ( .A1(n10409), .A2(n13416), .ZN(n13398) );
  INV_X1 U13129 ( .A(n13416), .ZN(n10405) );
  NAND2_X1 U13130 ( .A1(n10410), .A2(n10422), .ZN(n10408) );
  INV_X1 U13131 ( .A(n11666), .ZN(n10410) );
  INV_X1 U13132 ( .A(n11667), .ZN(n10411) );
  NAND3_X1 U13133 ( .A1(n10414), .A2(n10413), .A3(n9879), .ZN(n11617) );
  OR2_X2 U13134 ( .A1(n14523), .A2(n10426), .ZN(n14436) );
  INV_X1 U13135 ( .A(n10432), .ZN(n13916) );
  OAI21_X1 U13136 ( .B1(n10431), .B2(n11922), .A(n11936), .ZN(n14613) );
  OR2_X1 U13137 ( .A1(n10432), .A2(n10430), .ZN(n11936) );
  NAND2_X1 U13138 ( .A1(n11922), .A2(n13915), .ZN(n10430) );
  NAND2_X1 U13139 ( .A1(n11622), .A2(n20204), .ZN(n10436) );
  NOR2_X1 U13140 ( .A1(n12712), .A2(n10434), .ZN(n10433) );
  NAND3_X1 U13141 ( .A1(n10436), .A2(n10435), .A3(n10433), .ZN(n12312) );
  NAND2_X1 U13142 ( .A1(n14337), .A2(n10443), .ZN(n12255) );
  AND2_X1 U13143 ( .A1(n14337), .A2(n10444), .ZN(n12442) );
  NAND2_X1 U13144 ( .A1(n14337), .A2(n14339), .ZN(n12440) );
  INV_X1 U13145 ( .A(n14339), .ZN(n10445) );
  CLKBUF_X1 U13146 ( .A(n15422), .Z(n16293) );
  INV_X1 U13147 ( .A(n12442), .ZN(n12443) );
  OAI22_X1 U13148 ( .A1(n10628), .A2(n10627), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10607), .ZN(n10631) );
  NAND2_X1 U13149 ( .A1(n11133), .A2(n11132), .ZN(n13726) );
  INV_X1 U13150 ( .A(n13673), .ZN(n11133) );
  NAND2_X1 U13151 ( .A1(n12812), .A2(n20047), .ZN(n12439) );
  NAND2_X1 U13152 ( .A1(n12255), .A2(n12254), .ZN(n12257) );
  INV_X2 U13153 ( .A(n13925), .ZN(n19352) );
  OAI21_X1 U13154 ( .B1(n10653), .B2(n11087), .A(n10647), .ZN(n10656) );
  NAND2_X1 U13155 ( .A1(n10653), .A2(n10660), .ZN(n10648) );
  NOR2_X1 U13156 ( .A1(n19339), .A2(n19351), .ZN(n19832) );
  AND3_X1 U13157 ( .A1(n19339), .A2(n19332), .A3(n11437), .ZN(n10581) );
  AND2_X1 U13158 ( .A1(n10586), .A2(n13925), .ZN(n10580) );
  INV_X1 U13159 ( .A(n10669), .ZN(n10675) );
  NAND2_X1 U13160 ( .A1(n11609), .A2(n11554), .ZN(n11556) );
  AOI22_X1 U13161 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11551) );
  NAND4_X1 U13162 ( .A1(n19339), .A2(n11265), .A3(n19352), .A4(n13291), .ZN(
        n10597) );
  OAI21_X1 U13163 ( .B1(n11608), .B2(n11609), .A(n11621), .ZN(n12575) );
  CLKBUF_X1 U13164 ( .A(n13579), .Z(n15545) );
  NAND2_X1 U13165 ( .A1(n13579), .A2(n13284), .ZN(n13289) );
  NAND2_X1 U13166 ( .A1(n12838), .A2(n12839), .ZN(n12841) );
  AOI22_X1 U13167 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11543) );
  AND2_X1 U13168 ( .A1(n9915), .A2(n12726), .ZN(n13403) );
  INV_X1 U13169 ( .A(n11278), .ZN(n11328) );
  INV_X1 U13170 ( .A(n11301), .ZN(n11406) );
  INV_X2 U13171 ( .A(n17365), .ZN(n17360) );
  NOR2_X1 U13172 ( .A1(n12763), .A2(n12762), .ZN(n10448) );
  AND2_X1 U13173 ( .A1(n14602), .A2(n14044), .ZN(n10449) );
  NAND2_X2 U13174 ( .A1(n14602), .A2(n13259), .ZN(n14622) );
  OR2_X1 U13175 ( .A1(n13779), .A2(n12429), .ZN(n14471) );
  INV_X1 U13176 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20703) );
  AND2_X1 U13177 ( .A1(n11608), .A2(n11721), .ZN(n10450) );
  AND2_X1 U13178 ( .A1(n10618), .A2(n10617), .ZN(n10451) );
  AND4_X1 U13179 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n10452) );
  AND3_X1 U13180 ( .A1(n10475), .A2(n10474), .A3(n16411), .ZN(n10453) );
  OR2_X1 U13181 ( .A1(n11406), .A2(n11326), .ZN(n10454) );
  NOR2_X1 U13182 ( .A1(n20553), .A2(n20856), .ZN(n10455) );
  OR2_X1 U13183 ( .A1(n17287), .A2(n17316), .ZN(n10456) );
  OR2_X1 U13184 ( .A1(n17902), .A2(n16538), .ZN(n10457) );
  AND2_X1 U13185 ( .A1(n11211), .A2(n11210), .ZN(n10458) );
  AND3_X1 U13186 ( .A1(n18170), .A2(n18195), .A3(n15817), .ZN(n10459) );
  AND4_X1 U13187 ( .A1(n11211), .A2(n15205), .A3(n15202), .A4(n11028), .ZN(
        n10460) );
  INV_X1 U13188 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n12265) );
  INV_X1 U13189 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11795) );
  INV_X1 U13190 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15817) );
  INV_X2 U13191 ( .A(n19033), .ZN(n18966) );
  AND2_X1 U13192 ( .A1(n14731), .A2(n14833), .ZN(n10461) );
  NAND2_X1 U13193 ( .A1(n20776), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20814) );
  INV_X1 U13194 ( .A(n20814), .ZN(n20887) );
  INV_X1 U13195 ( .A(n15388), .ZN(n10890) );
  INV_X1 U13196 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12694) );
  INV_X1 U13197 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12690) );
  INV_X1 U13198 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11084) );
  INV_X1 U13199 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11881) );
  NOR2_X1 U13200 ( .A1(n16163), .A2(n16162), .ZN(n10462) );
  INV_X1 U13201 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15856) );
  OR2_X1 U13202 ( .A1(n14263), .A2(n14262), .ZN(n10463) );
  INV_X1 U13203 ( .A(n11267), .ZN(n11071) );
  OR2_X1 U13204 ( .A1(n14877), .A2(n15221), .ZN(n10464) );
  INV_X1 U13205 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19798) );
  INV_X1 U13206 ( .A(n13530), .ZN(n13531) );
  NAND2_X1 U13207 ( .A1(n14136), .A2(n14135), .ZN(n10465) );
  OR2_X2 U13208 ( .A1(n10996), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10466) );
  INV_X1 U13209 ( .A(n10933), .ZN(n11326) );
  AND2_X2 U13210 ( .A1(n11487), .A2(n11486), .ZN(n11535) );
  NAND2_X1 U13211 ( .A1(n20092), .A2(n14044), .ZN(n14546) );
  NAND2_X1 U13212 ( .A1(n11554), .A2(n20092), .ZN(n14539) );
  INV_X1 U13213 ( .A(n14539), .ZN(n20089) );
  OR2_X2 U13214 ( .A1(n13543), .A2(n13542), .ZN(n20134) );
  INV_X1 U13215 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15506) );
  AND2_X2 U13216 ( .A1(n10674), .A2(n10673), .ZN(n13164) );
  AND2_X1 U13217 ( .A1(n11090), .A2(n10643), .ZN(n10468) );
  INV_X1 U13218 ( .A(n11507), .ZN(n12178) );
  INV_X1 U13219 ( .A(n12178), .ZN(n12566) );
  NOR2_X1 U13220 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11507) );
  NOR2_X1 U13221 ( .A1(n9812), .A2(n12696), .ZN(n12338) );
  NAND2_X1 U13222 ( .A1(n12341), .A2(n11620), .ZN(n12728) );
  INV_X1 U13223 ( .A(n12696), .ZN(n11627) );
  NAND2_X1 U13224 ( .A1(n11556), .A2(n11647), .ZN(n12576) );
  AOI22_X1 U13225 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11531) );
  OR2_X1 U13226 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15856), .ZN(
        n12261) );
  INV_X1 U13227 ( .A(n12606), .ZN(n11734) );
  OR2_X1 U13228 ( .A1(n12295), .A2(n11733), .ZN(n11737) );
  AOI22_X1 U13229 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11503) );
  INV_X1 U13230 ( .A(n12301), .ZN(n12302) );
  INV_X1 U13231 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13400) );
  OR2_X1 U13232 ( .A1(n11679), .A2(n11678), .ZN(n11682) );
  OR2_X1 U13233 ( .A1(n14115), .A2(n14114), .ZN(n14133) );
  AND4_X1 U13234 ( .A1(n10876), .A2(n10875), .A3(n10874), .A4(n10873), .ZN(
        n10881) );
  AOI22_X1 U13235 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10522) );
  OR2_X1 U13236 ( .A1(n13021), .A2(n13020), .ZN(n13016) );
  INV_X1 U13237 ( .A(n18006), .ZN(n15823) );
  INV_X1 U13238 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U13239 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11510) );
  OR2_X1 U13240 ( .A1(n12295), .A2(n11854), .ZN(n11866) );
  OR2_X1 U13241 ( .A1(n11864), .A2(n11863), .ZN(n12661) );
  INV_X1 U13242 ( .A(n14179), .ZN(n14180) );
  INV_X1 U13243 ( .A(n11285), .ZN(n11286) );
  AND2_X1 U13244 ( .A1(n10914), .A2(n10913), .ZN(n11226) );
  NAND2_X1 U13245 ( .A1(n13926), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U13246 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n15696) );
  AND2_X1 U13247 ( .A1(n12299), .A2(n12298), .ZN(n12317) );
  INV_X1 U13248 ( .A(n11659), .ZN(n11775) );
  OR2_X1 U13249 ( .A1(n12154), .A2(n12153), .ZN(n12161) );
  NOR2_X1 U13250 ( .A1(n12698), .A2(n12577), .ZN(n13327) );
  OR2_X1 U13251 ( .A1(n12229), .A2(n14641), .ZN(n12230) );
  INV_X1 U13252 ( .A(n12060), .ZN(n12061) );
  INV_X1 U13253 ( .A(n13731), .ZN(n11900) );
  AND2_X1 U13254 ( .A1(n20213), .A2(n11616), .ZN(n12695) );
  INV_X1 U13255 ( .A(n11751), .ZN(n11752) );
  AND2_X1 U13256 ( .A1(n12303), .A2(n12695), .ZN(n12297) );
  NAND2_X1 U13257 ( .A1(n14181), .A2(n14180), .ZN(n14182) );
  OR2_X1 U13258 ( .A1(n14199), .A2(n14201), .ZN(n14223) );
  INV_X1 U13259 ( .A(n14991), .ZN(n14081) );
  NAND2_X1 U13260 ( .A1(n11301), .A2(n11286), .ZN(n11287) );
  NOR2_X1 U13261 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16426), .ZN(
        n10907) );
  AND2_X1 U13262 ( .A1(n11421), .A2(n11420), .ZN(n13922) );
  NAND2_X1 U13263 ( .A1(n10579), .A2(n10581), .ZN(n10910) );
  AND2_X2 U13264 ( .A1(n10591), .A2(n19332), .ZN(n11444) );
  AND2_X1 U13265 ( .A1(n13164), .A2(n10675), .ZN(n10693) );
  NAND2_X1 U13266 ( .A1(n10525), .A2(n16411), .ZN(n10532) );
  AOI21_X1 U13267 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18847), .A(
        n13015), .ZN(n13021) );
  INV_X1 U13268 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15602) );
  INV_X1 U13269 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U13270 ( .A1(n15820), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n18142), .B2(n17793), .ZN(n15821) );
  INV_X1 U13271 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17235) );
  OAI211_X1 U13272 ( .C1(n11659), .C2(n11660), .A(n11665), .B(n11664), .ZN(
        n11666) );
  AND2_X1 U13273 ( .A1(n12376), .A2(n12375), .ZN(n15934) );
  NOR2_X1 U13274 ( .A1(n14846), .A2(n16196), .ZN(n12251) );
  NAND2_X1 U13275 ( .A1(n14614), .A2(n11936), .ZN(n14543) );
  OR2_X1 U13276 ( .A1(n12230), .A2(n14320), .ZN(n12323) );
  AND2_X1 U13277 ( .A1(n12194), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12195) );
  NOR2_X1 U13278 ( .A1(n12029), .A2(n14736), .ZN(n12030) );
  INV_X1 U13279 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11903) );
  NOR2_X1 U13280 ( .A1(n11847), .A2(n20056), .ZN(n11867) );
  INV_X1 U13281 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20189) );
  AND2_X1 U13282 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20342), .ZN(n20226) );
  NAND2_X2 U13283 ( .A1(n10976), .A2(n11267), .ZN(n11011) );
  OR2_X1 U13284 ( .A1(n11378), .A2(n11377), .ZN(n13629) );
  NOR2_X1 U13285 ( .A1(n13215), .A2(n13291), .ZN(n14174) );
  INV_X1 U13286 ( .A(n14277), .ZN(n14268) );
  AND2_X1 U13289 ( .A1(n13703), .A2(n10991), .ZN(n15482) );
  INV_X1 U13290 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13577) );
  INV_X1 U13291 ( .A(n10910), .ZN(n16438) );
  NOR2_X1 U13292 ( .A1(n11434), .A2(n11433), .ZN(n16433) );
  AND2_X1 U13293 ( .A1(n11248), .A2(n11247), .ZN(n13087) );
  AND2_X2 U13294 ( .A1(n10683), .A2(n10699), .ZN(n19323) );
  AOI22_X1 U13295 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18856), .B1(
        n13025), .B2(n13024), .ZN(n14022) );
  INV_X1 U13296 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17051) );
  NOR2_X1 U13297 ( .A1(n15699), .A2(n15698), .ZN(n15700) );
  NAND2_X1 U13298 ( .A1(n15806), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15807) );
  INV_X1 U13299 ( .A(n18296), .ZN(n18231) );
  OR2_X1 U13300 ( .A1(n14369), .A2(n14321), .ZN(n14332) );
  INV_X1 U13301 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15953) );
  OR2_X1 U13302 ( .A1(n20030), .A2(n12430), .ZN(n20059) );
  AND2_X1 U13303 ( .A1(n12397), .A2(n12396), .ZN(n14385) );
  AND3_X1 U13304 ( .A1(n11967), .A2(n11966), .A3(n11965), .ZN(n14533) );
  AND2_X1 U13305 ( .A1(n13541), .A2(n20876), .ZN(n13542) );
  INV_X1 U13306 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14641) );
  NAND2_X1 U13307 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12193) );
  INV_X1 U13308 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15938) );
  INV_X1 U13309 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15964) );
  AND4_X1 U13310 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n13731) );
  INV_X1 U13311 ( .A(n20169), .ZN(n16151) );
  NAND2_X1 U13312 ( .A1(n12743), .A2(n12741), .ZN(n20162) );
  OAI22_X1 U13313 ( .A1(n15874), .A2(n20884), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n20841), .ZN(n20342) );
  INV_X1 U13314 ( .A(n15882), .ZN(n14307) );
  OR2_X1 U13315 ( .A1(n20180), .A2(n20457), .ZN(n20557) );
  AOI21_X1 U13316 ( .B1(n20866), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20236), 
        .ZN(n20710) );
  OR2_X1 U13317 ( .A1(n16201), .A2(n14920), .ZN(n19141) );
  NAND2_X1 U13318 ( .A1(n19179), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19210) );
  OR2_X1 U13319 ( .A1(n11232), .A2(n10915), .ZN(n16430) );
  INV_X1 U13320 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15257) );
  INV_X1 U13321 ( .A(n10674), .ZN(n10670) );
  INV_X1 U13322 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U13323 ( .A1(n11475), .A2(n11264), .ZN(n16400) );
  AND2_X1 U13324 ( .A1(n11475), .A2(n11451), .ZN(n15386) );
  NAND2_X1 U13325 ( .A1(n16457), .A2(n15912), .ZN(n15913) );
  NAND2_X1 U13326 ( .A1(n19798), .A2(n19809), .ZN(n19756) );
  AND2_X1 U13327 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19797), .ZN(
        n13285) );
  NOR2_X1 U13328 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16815), .ZN(n16796) );
  INV_X1 U13329 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16885) );
  INV_X1 U13330 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17121) );
  INV_X1 U13331 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17185) );
  INV_X1 U13332 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17273) );
  INV_X1 U13333 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17736) );
  INV_X1 U13334 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17775) );
  INV_X1 U13335 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17815) );
  INV_X1 U13336 ( .A(n17862), .ZN(n18198) );
  NOR2_X1 U13337 ( .A1(n18067), .A2(n17685), .ZN(n18044) );
  NOR2_X1 U13338 ( .A1(n18841), .A2(n18826), .ZN(n18296) );
  INV_X1 U13339 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18170) );
  INV_X1 U13340 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17857) );
  INV_X1 U13341 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15813) );
  NAND2_X1 U13342 ( .A1(n17965), .A2(n17966), .ZN(n17964) );
  INV_X1 U13343 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17285) );
  AOI221_X1 U13344 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18869), .C1(n18985), 
        .C2(P3_STATE2_REG_2__SCAN_IN), .A(n19000), .ZN(n18343) );
  OAI21_X1 U13345 ( .B1(n14504), .B2(n15963), .A(n12884), .ZN(n12885) );
  OR2_X1 U13346 ( .A1(n14762), .A2(n15963), .ZN(n12437) );
  NOR2_X1 U13347 ( .A1(n13839), .A2(n13939), .ZN(n14479) );
  AND2_X1 U13348 ( .A1(n20875), .A2(n12322), .ZN(n20030) );
  NAND2_X1 U13349 ( .A1(n12424), .A2(n12423), .ZN(n20032) );
  INV_X1 U13350 ( .A(n20008), .ZN(n12705) );
  INV_X1 U13351 ( .A(n13588), .ZN(n13766) );
  NAND2_X1 U13352 ( .A1(n11999), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12029) );
  NAND2_X1 U13353 ( .A1(n11919), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11962) );
  AND2_X1 U13354 ( .A1(n12713), .A2(n12730), .ZN(n15862) );
  OAI21_X1 U13355 ( .B1(n13468), .B2(n20162), .A(n16116), .ZN(n13625) );
  AND2_X1 U13356 ( .A1(n12743), .A2(n12724), .ZN(n20169) );
  INV_X1 U13357 ( .A(n20260), .ZN(n20859) );
  OAI22_X1 U13358 ( .A1(n20192), .A2(n20191), .B1(n20522), .B2(n20337), .ZN(
        n20231) );
  INV_X1 U13359 ( .A(n20298), .ZN(n20181) );
  OAI22_X1 U13360 ( .A1(n20269), .A2(n20268), .B1(n20522), .B2(n20396), .ZN(
        n20293) );
  NAND2_X1 U13361 ( .A1(n20180), .A2(n20456), .ZN(n20298) );
  INV_X1 U13362 ( .A(n20338), .ZN(n20360) );
  OAI22_X1 U13363 ( .A1(n20398), .A2(n20397), .B1(n20396), .B2(n20661), .ZN(
        n20421) );
  INV_X1 U13364 ( .A(n20448), .ZN(n20451) );
  OAI211_X1 U13365 ( .C1(n20481), .C2(n20466), .A(n20518), .B(n20465), .ZN(
        n20484) );
  INV_X1 U13366 ( .A(n20582), .ZN(n20458) );
  OAI22_X1 U13367 ( .A1(n20524), .A2(n20523), .B1(n20522), .B2(n20662), .ZN(
        n20549) );
  AND2_X1 U13368 ( .A1(n13427), .A2(n20260), .ZN(n20513) );
  OAI22_X1 U13369 ( .A1(n20592), .A2(n20591), .B1(n20590), .B2(n20661), .ZN(
        n20622) );
  OR2_X1 U13370 ( .A1(n13427), .A2(n20859), .ZN(n20582) );
  NOR2_X2 U13371 ( .A1(n20709), .A2(n20634), .ZN(n20695) );
  INV_X1 U13372 ( .A(n20620), .ZN(n20758) );
  INV_X1 U13373 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20776) );
  NOR2_X1 U13374 ( .A1(n20888), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20812) );
  INV_X1 U13375 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U13376 ( .B1(n14292), .B2(n19207), .A(n12536), .ZN(n12537) );
  INV_X1 U13377 ( .A(n19158), .ZN(n19199) );
  INV_X1 U13378 ( .A(n19869), .ZN(n19108) );
  INV_X1 U13379 ( .A(n19112), .ZN(n16371) );
  AND2_X1 U13380 ( .A1(n19249), .A2(n13929), .ZN(n19215) );
  INV_X1 U13381 ( .A(n13834), .ZN(n19243) );
  AOI21_X1 U13382 ( .B1(n13149), .B2(n13148), .A(n19877), .ZN(n19250) );
  INV_X1 U13383 ( .A(n13143), .ZN(n13077) );
  AND2_X1 U13384 ( .A1(n13607), .A2(n10357), .ZN(n16319) );
  NOR2_X1 U13385 ( .A1(n11467), .A2(n15470), .ZN(n16377) );
  INV_X1 U13386 ( .A(n19311), .ZN(n16388) );
  INV_X1 U13387 ( .A(n16400), .ZN(n19308) );
  INV_X1 U13388 ( .A(n19756), .ZN(n19961) );
  AND2_X1 U13389 ( .A1(n10922), .A2(n10921), .ZN(n19998) );
  NAND2_X1 U13390 ( .A1(n16432), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16457) );
  OAI21_X1 U13391 ( .B1(n19326), .B2(n19325), .A(n19324), .ZN(n19355) );
  INV_X1 U13392 ( .A(n19391), .ZN(n19413) );
  OAI21_X1 U13393 ( .B1(n19425), .B2(n19424), .A(n19423), .ZN(n19442) );
  INV_X1 U13394 ( .A(n19454), .ZN(n19476) );
  OAI21_X1 U13395 ( .B1(n19486), .B2(n19485), .A(n19484), .ZN(n19503) );
  INV_X1 U13396 ( .A(n19507), .ZN(n19534) );
  NOR2_X1 U13397 ( .A1(n19545), .A2(n19542), .ZN(n19564) );
  INV_X1 U13398 ( .A(n19601), .ZN(n19569) );
  INV_X1 U13399 ( .A(n19634), .ZN(n19656) );
  INV_X1 U13400 ( .A(n19669), .ZN(n19957) );
  NOR2_X1 U13401 ( .A1(n19726), .A2(n19690), .ZN(n19744) );
  INV_X1 U13402 ( .A(n19843), .ZN(n19781) );
  AND2_X1 U13403 ( .A1(n19448), .A2(n19981), .ZN(n19802) );
  INV_X1 U13404 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19889) );
  NAND2_X1 U13405 ( .A1(n19020), .A2(n18806), .ZN(n17560) );
  NOR2_X1 U13406 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16770), .ZN(n16756) );
  NOR2_X1 U13407 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16838), .ZN(n16823) );
  NOR2_X1 U13408 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16859), .ZN(n16845) );
  NOR2_X1 U13409 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16881), .ZN(n16865) );
  INV_X1 U13410 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17277) );
  INV_X1 U13411 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16933) );
  INV_X1 U13412 ( .A(n17017), .ZN(n17035) );
  NAND2_X1 U13413 ( .A1(n13030), .A2(n18866), .ZN(n17026) );
  NOR2_X1 U13414 ( .A1(n16791), .A2(n17139), .ZN(n17105) );
  NAND2_X1 U13415 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17197), .ZN(n17196) );
  AND3_X1 U13416 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17349), .A3(n17323), .ZN(
        n17321) );
  NAND3_X1 U13417 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17368), .A3(n17353), .ZN(
        n15643) );
  INV_X1 U13418 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17848) );
  NOR2_X1 U13419 ( .A1(n18979), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19037) );
  INV_X1 U13420 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17987) );
  INV_X1 U13421 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18088) );
  NOR2_X1 U13422 ( .A1(n18057), .A2(n18305), .ZN(n18064) );
  INV_X1 U13423 ( .A(n17791), .ZN(n18115) );
  INV_X1 U13424 ( .A(n18114), .ZN(n18221) );
  AOI21_X1 U13425 ( .B1(n15783), .B2(n15782), .A(n18874), .ZN(n18325) );
  INV_X1 U13426 ( .A(n18325), .ZN(n18305) );
  NOR2_X1 U13427 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18975), .ZN(
        n19000) );
  CLKBUF_X1 U13428 ( .A(n18421), .Z(n18455) );
  CLKBUF_X1 U13429 ( .A(n18462), .Z(n18478) );
  INV_X1 U13430 ( .A(n18501), .ZN(n18572) );
  CLKBUF_X1 U13431 ( .A(n18711), .Z(n18697) );
  OR2_X1 U13432 ( .A1(n18653), .A2(n18720), .ZN(n18680) );
  AND2_X1 U13433 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18752), .ZN(n18764) );
  AND2_X1 U13434 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18752), .ZN(n18796) );
  INV_X1 U13435 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18985) );
  AND2_X1 U13436 ( .A1(n18966), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18903) );
  NOR2_X1 U13437 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12909), .ZN(n16631)
         );
  NAND2_X1 U13438 ( .A1(n11614), .A2(n13224), .ZN(n13543) );
  INV_X1 U13439 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21003) );
  INV_X1 U13440 ( .A(n12885), .ZN(n12886) );
  AND2_X1 U13441 ( .A1(n12437), .A2(n12436), .ZN(n12438) );
  OR2_X1 U13442 ( .A1(n20030), .A2(n12326), .ZN(n15978) );
  INV_X1 U13443 ( .A(n12451), .ZN(n12452) );
  OR2_X1 U13444 ( .A1(n14618), .A2(n13259), .ZN(n14604) );
  NAND2_X1 U13445 ( .A1(n20095), .A2(n11627), .ZN(n13375) );
  INV_X1 U13446 ( .A(n20095), .ZN(n20122) );
  INV_X1 U13447 ( .A(n20134), .ZN(n13587) );
  OR2_X1 U13448 ( .A1(n20134), .A2(n11616), .ZN(n13748) );
  NAND2_X1 U13449 ( .A1(n12811), .A2(n20858), .ZN(n20142) );
  NAND2_X2 U13450 ( .A1(n15862), .A2(n13224), .ZN(n20155) );
  NAND2_X1 U13451 ( .A1(n13626), .A2(n13625), .ZN(n16138) );
  INV_X1 U13452 ( .A(n16182), .ZN(n20176) );
  NAND2_X1 U13453 ( .A1(n20181), .A2(n20458), .ZN(n20259) );
  OR2_X1 U13454 ( .A1(n20298), .A2(n20634), .ZN(n20291) );
  OR2_X1 U13455 ( .A1(n20298), .A2(n20659), .ZN(n20328) );
  OR2_X1 U13456 ( .A1(n20298), .A2(n20426), .ZN(n20338) );
  NAND2_X1 U13457 ( .A1(n20335), .A2(n20458), .ZN(n20388) );
  OR2_X1 U13458 ( .A1(n20432), .A2(n20634), .ZN(n20425) );
  OR2_X1 U13459 ( .A1(n20432), .A2(n20659), .ZN(n20448) );
  NAND2_X1 U13460 ( .A1(n20847), .A2(n20458), .ZN(n20512) );
  NAND2_X1 U13461 ( .A1(n20847), .A2(n20491), .ZN(n20547) );
  NAND2_X1 U13462 ( .A1(n20847), .A2(n20513), .ZN(n20581) );
  NAND2_X1 U13463 ( .A1(n20847), .A2(n20560), .ZN(n20626) );
  OR2_X1 U13464 ( .A1(n20709), .A2(n20582), .ZN(n20658) );
  INV_X1 U13465 ( .A(n20739), .ZN(n20683) );
  INV_X1 U13466 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16195) );
  INV_X1 U13467 ( .A(n20829), .ZN(n20769) );
  NAND2_X1 U13468 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20880) );
  INV_X1 U13469 ( .A(n11439), .ZN(n14043) );
  NAND2_X1 U13470 ( .A1(n11251), .A2(n10924), .ZN(n13045) );
  OR3_X1 U13471 ( .A1(n19043), .A2(n14854), .A3(n16450), .ZN(n19158) );
  OR2_X1 U13472 ( .A1(n13143), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19207) );
  INV_X1 U13473 ( .A(n14983), .ZN(n15010) );
  INV_X1 U13474 ( .A(n13301), .ZN(n14983) );
  INV_X1 U13475 ( .A(n13301), .ZN(n15000) );
  NAND2_X1 U13476 ( .A1(n19249), .A2(n13184), .ZN(n15120) );
  AND2_X1 U13477 ( .A1(n15120), .A2(n15023), .ZN(n19239) );
  NAND2_X1 U13478 ( .A1(n19249), .A2(n13183), .ZN(n13834) );
  INV_X1 U13479 ( .A(n19250), .ZN(n19284) );
  NAND2_X1 U13480 ( .A1(n13038), .A2(n12528), .ZN(n13148) );
  INV_X1 U13481 ( .A(n19291), .ZN(n16356) );
  INV_X1 U13482 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19126) );
  OR2_X1 U13483 ( .A1(n13045), .A2(n14957), .ZN(n16358) );
  OR2_X1 U13484 ( .A1(n12802), .A2(n19300), .ZN(n12801) );
  XNOR2_X1 U13485 ( .A(n11212), .B(n10458), .ZN(n15201) );
  INV_X1 U13486 ( .A(n16391), .ZN(n19300) );
  INV_X1 U13487 ( .A(n19302), .ZN(n16410) );
  NAND2_X1 U13488 ( .A1(n19569), .A2(n19508), .ZN(n19381) );
  NAND2_X1 U13489 ( .A1(n19569), .A2(n19539), .ZN(n19391) );
  OR2_X1 U13490 ( .A1(n19480), .A2(n19669), .ZN(n19454) );
  OR2_X1 U13491 ( .A1(n19449), .A2(n19726), .ZN(n19497) );
  NAND2_X1 U13492 ( .A1(n19508), .A2(n19802), .ZN(n19538) );
  NAND2_X1 U13493 ( .A1(n19802), .A2(n19539), .ZN(n19599) );
  OR2_X1 U13494 ( .A1(n19727), .A2(n19601), .ZN(n19634) );
  NAND2_X1 U13495 ( .A1(n19752), .A2(n19957), .ZN(n19689) );
  INV_X1 U13496 ( .A(n19744), .ZN(n19751) );
  OR2_X1 U13497 ( .A1(n19727), .A2(n19726), .ZN(n19776) );
  NAND2_X1 U13498 ( .A1(n19752), .A2(n19802), .ZN(n19859) );
  NOR2_X1 U13499 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15910) );
  INV_X1 U13500 ( .A(n19956), .ZN(n19870) );
  NAND2_X1 U13501 ( .A1(n19878), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20006) );
  NAND2_X1 U13502 ( .A1(n18985), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17994) );
  INV_X1 U13503 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16909) );
  NAND2_X1 U13504 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18882), .ZN(n17019) );
  INV_X1 U13505 ( .A(n17014), .ZN(n17037) );
  NOR2_X1 U13506 ( .A1(n16729), .A2(n17082), .ZN(n17087) );
  NOR2_X1 U13507 ( .A1(n17170), .A2(n17196), .ZN(n17183) );
  NOR2_X2 U13508 ( .A1(n15552), .A2(n17371), .ZN(n17365) );
  NOR2_X1 U13509 ( .A1(n17456), .A2(n17475), .ZN(n17479) );
  INV_X1 U13510 ( .A(n17517), .ZN(n17506) );
  NAND2_X1 U13511 ( .A1(n17542), .A2(n18345), .ZN(n17541) );
  INV_X1 U13512 ( .A(n17542), .ZN(n17559) );
  INV_X1 U13513 ( .A(n17808), .ZN(n17845) );
  INV_X1 U13514 ( .A(n17859), .ZN(n17903) );
  INV_X1 U13515 ( .A(n17978), .ZN(n17999) );
  NAND2_X1 U13516 ( .A1(n18216), .A2(n18305), .ZN(n18317) );
  NAND2_X1 U13517 ( .A1(n18809), .A2(n18315), .ZN(n18332) );
  INV_X1 U13518 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18354) );
  INV_X1 U13519 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18379) );
  INV_X1 U13520 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18415) );
  INV_X1 U13521 ( .A(n18527), .ZN(n18459) );
  INV_X1 U13522 ( .A(n18550), .ZN(n18482) );
  INV_X1 U13523 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18507) );
  INV_X1 U13524 ( .A(n18673), .ZN(n18602) );
  INV_X1 U13525 ( .A(n18739), .ZN(n18651) );
  INV_X1 U13526 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18685) );
  INV_X1 U13527 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18709) );
  INV_X1 U13528 ( .A(n19020), .ZN(n18874) );
  INV_X1 U13529 ( .A(n18971), .ZN(n18883) );
  INV_X1 U13530 ( .A(n15775), .ZN(n19023) );
  AND2_X2 U13531 ( .A1(n12592), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20177)
         );
  INV_X1 U13532 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U13533 ( .A1(n12439), .A2(n12438), .ZN(P1_U2811) );
  NAND2_X1 U13534 ( .A1(n12453), .A2(n12452), .ZN(P1_U2845) );
  NAND2_X1 U13535 ( .A1(n12861), .A2(n12860), .ZN(P2_U3016) );
  OAI21_X1 U13536 ( .B1(n15201), .B2(n19300), .A(n11478), .ZN(P2_U3025) );
  OR4_X1 U13537 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        P3_U2670) );
  NOR2_X2 U13538 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10469) );
  AND2_X4 U13539 ( .A1(n10469), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14254) );
  AOI22_X1 U13540 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10472) );
  AND2_X4 U13541 ( .A1(n15521), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14270) );
  AOI22_X1 U13542 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10471) );
  BUF_X4 U13543 ( .A(n10520), .Z(n14247) );
  AND2_X4 U13544 ( .A1(n15521), .A2(n16412), .ZN(n10715) );
  AOI22_X1 U13545 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10470) );
  INV_X1 U13546 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13547 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U13548 ( .A1(n9864), .A2(n10473), .ZN(n10479) );
  AOI22_X1 U13549 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13550 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13551 ( .A1(n9809), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13552 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10476) );
  NAND3_X1 U13553 ( .A1(n10453), .A2(n10477), .A3(n10476), .ZN(n10478) );
  AND2_X4 U13554 ( .A1(n10479), .A2(n10478), .ZN(n11267) );
  AOI22_X1 U13555 ( .A1(n9804), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U13556 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U13557 ( .A1(n10509), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13558 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10480) );
  NAND4_X1 U13559 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10484) );
  NAND2_X1 U13560 ( .A1(n10484), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10491) );
  AOI22_X1 U13561 ( .A1(n9809), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13562 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13563 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13564 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13565 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10489) );
  NAND2_X1 U13566 ( .A1(n10489), .A2(n16411), .ZN(n10490) );
  NAND2_X2 U13567 ( .A1(n10491), .A2(n10490), .ZN(n13291) );
  NOR2_X2 U13568 ( .A1(n11267), .A2(n13291), .ZN(n10586) );
  INV_X1 U13569 ( .A(n10586), .ZN(n10493) );
  NAND2_X1 U13570 ( .A1(n13291), .A2(n11267), .ZN(n10492) );
  AOI22_X1 U13571 ( .A1(n10509), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10494) );
  INV_X1 U13572 ( .A(n10494), .ZN(n10499) );
  AOI22_X1 U13573 ( .A1(n9809), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13574 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13575 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10495) );
  NAND3_X1 U13576 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(n10498) );
  NOR2_X1 U13577 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  NAND2_X1 U13578 ( .A1(n10500), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10508) );
  BUF_X4 U13579 ( .A(n10520), .Z(n14273) );
  AOI22_X1 U13580 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13581 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13582 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10502) );
  AND4_X1 U13583 ( .A1(n10505), .A2(n10504), .A3(n10503), .A4(n10502), .ZN(
        n10506) );
  NAND2_X1 U13584 ( .A1(n10506), .A2(n16411), .ZN(n10507) );
  INV_X1 U13585 ( .A(n13291), .ZN(n13165) );
  BUF_X8 U13586 ( .A(n10509), .Z(n14271) );
  AOI22_X1 U13587 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13588 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13589 ( .A1(n9806), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13590 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10510) );
  NAND4_X1 U13591 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10519) );
  AOI22_X1 U13592 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13593 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13594 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13595 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10514) );
  NAND4_X1 U13596 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10518) );
  MUX2_X2 U13597 ( .A(n10519), .B(n10518), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13925) );
  AOI22_X1 U13598 ( .A1(n9804), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13599 ( .A1(n10520), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13600 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10521) );
  NAND4_X1 U13601 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10525) );
  AOI22_X1 U13602 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13603 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13604 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13605 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10526) );
  NAND4_X1 U13606 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10530) );
  NAND2_X2 U13607 ( .A1(n10532), .A2(n10531), .ZN(n11437) );
  NAND2_X1 U13608 ( .A1(n11435), .A2(n11437), .ZN(n10534) );
  INV_X2 U13609 ( .A(n11267), .ZN(n11265) );
  NAND2_X1 U13610 ( .A1(n10534), .A2(n10533), .ZN(n10634) );
  AOI22_X1 U13611 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13612 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13613 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13614 ( .A1(n9820), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13615 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  AOI22_X1 U13616 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13617 ( .A1(n9809), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13618 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13619 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13620 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  NAND2_X1 U13621 ( .A1(n10544), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10545) );
  AOI22_X1 U13622 ( .A1(n9806), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13623 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13624 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13625 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10547) );
  NAND4_X1 U13626 ( .A1(n10550), .A2(n10549), .A3(n10548), .A4(n10547), .ZN(
        n10551) );
  AOI22_X1 U13627 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13628 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13629 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13630 ( .A1(n9804), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10552) );
  NAND4_X1 U13631 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10556) );
  NAND2_X1 U13632 ( .A1(n10634), .A2(n11259), .ZN(n10577) );
  NAND2_X1 U13633 ( .A1(n13182), .A2(n11437), .ZN(n10571) );
  AOI22_X1 U13634 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13635 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13636 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13637 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10559) );
  NAND4_X1 U13638 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10563) );
  AOI22_X1 U13639 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13640 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10715), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13641 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13642 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10564) );
  NAND4_X1 U13643 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10568) );
  AND2_X1 U13644 ( .A1(n19332), .A2(n13925), .ZN(n11240) );
  NAND2_X1 U13645 ( .A1(n10571), .A2(n11240), .ZN(n10575) );
  MUX2_X1 U13646 ( .A(n19339), .B(n11267), .S(n13291), .Z(n10574) );
  NAND4_X1 U13647 ( .A1(n10591), .A2(n19339), .A3(n11440), .A4(n11267), .ZN(
        n10572) );
  INV_X1 U13648 ( .A(n13097), .ZN(n10573) );
  OAI211_X2 U13649 ( .C1(n10575), .C2(n10574), .A(n10573), .B(n19317), .ZN(
        n11448) );
  NAND2_X1 U13650 ( .A1(n13182), .A2(n14227), .ZN(n11442) );
  NAND2_X1 U13651 ( .A1(n11442), .A2(n19317), .ZN(n10576) );
  AND2_X2 U13652 ( .A1(n11448), .A2(n10576), .ZN(n10632) );
  NAND2_X1 U13653 ( .A1(n10577), .A2(n10632), .ZN(n10578) );
  NAND2_X1 U13654 ( .A1(n10578), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10583) );
  NAND3_X1 U13655 ( .A1(n10910), .A2(n19332), .A3(n14957), .ZN(n10582) );
  NAND2_X1 U13656 ( .A1(n16437), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11213) );
  NAND2_X2 U13657 ( .A1(n10583), .A2(n10638), .ZN(n10628) );
  NAND2_X1 U13658 ( .A1(n10628), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10585) );
  NAND2_X1 U13659 ( .A1(n16452), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10584) );
  NAND2_X1 U13660 ( .A1(n10585), .A2(n10584), .ZN(n10603) );
  NAND2_X2 U13661 ( .A1(n14227), .A2(n19317), .ZN(n13095) );
  NAND3_X1 U13662 ( .A1(n11439), .A2(n11441), .A3(n13925), .ZN(n10590) );
  NAND2_X1 U13663 ( .A1(n10586), .A2(n14227), .ZN(n10588) );
  NAND2_X2 U13664 ( .A1(n11260), .A2(n11444), .ZN(n15520) );
  NAND2_X2 U13665 ( .A1(n13097), .A2(n19317), .ZN(n13145) );
  INV_X1 U13666 ( .A(n13095), .ZN(n10592) );
  NAND2_X1 U13667 ( .A1(n10592), .A2(n11444), .ZN(n13176) );
  NAND2_X1 U13668 ( .A1(n10593), .A2(n13926), .ZN(n10594) );
  INV_X1 U13669 ( .A(n10621), .ZN(n10595) );
  AND3_X2 U13670 ( .A1(n16451), .A2(n13145), .A3(n10595), .ZN(n10596) );
  AOI21_X4 U13671 ( .B1(n15520), .B2(n10596), .A(n19863), .ZN(n11096) );
  INV_X1 U13672 ( .A(n11096), .ZN(n10601) );
  AND2_X4 U13673 ( .A1(n10620), .A2(n10624), .ZN(n11188) );
  AOI22_X1 U13674 ( .A1(n11188), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10600) );
  INV_X1 U13675 ( .A(n10597), .ZN(n13177) );
  INV_X1 U13676 ( .A(n11444), .ZN(n10625) );
  NOR2_X1 U13677 ( .A1(n10625), .A2(n11228), .ZN(n10598) );
  AND2_X2 U13678 ( .A1(n13177), .A2(n10598), .ZN(n13168) );
  NAND2_X1 U13679 ( .A1(n10607), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13680 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  NAND2_X1 U13681 ( .A1(n10628), .A2(n15529), .ZN(n10606) );
  AOI21_X1 U13682 ( .B1(n19863), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10605) );
  NAND2_X2 U13683 ( .A1(n10606), .A2(n10605), .ZN(n10660) );
  NAND2_X1 U13684 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10612) );
  INV_X2 U13685 ( .A(n11095), .ZN(n10607) );
  INV_X1 U13686 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U13687 ( .A1(n11188), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13688 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10608) );
  OAI211_X1 U13689 ( .C1(n11095), .C2(n14907), .A(n10609), .B(n10608), .ZN(
        n10610) );
  INV_X1 U13690 ( .A(n10610), .ZN(n10611) );
  NAND2_X2 U13691 ( .A1(n10612), .A2(n10611), .ZN(n11089) );
  INV_X1 U13692 ( .A(n10644), .ZN(n10613) );
  NAND2_X1 U13693 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10619) );
  NAND2_X1 U13694 ( .A1(n11188), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10618) );
  INV_X1 U13695 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10929) );
  NAND2_X1 U13696 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10615) );
  AND2_X2 U13697 ( .A1(n10619), .A2(n10451), .ZN(n10647) );
  NAND2_X1 U13698 ( .A1(n10628), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10623) );
  NAND2_X2 U13699 ( .A1(n10620), .A2(n16437), .ZN(n12526) );
  NAND2_X2 U13700 ( .A1(n10623), .A2(n10622), .ZN(n10653) );
  INV_X1 U13701 ( .A(n10624), .ZN(n10626) );
  NOR2_X1 U13702 ( .A1(n10626), .A2(n10625), .ZN(n10627) );
  INV_X1 U13703 ( .A(n15520), .ZN(n10629) );
  AOI22_X1 U13704 ( .A1(n10629), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16452), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10630) );
  NAND2_X1 U13705 ( .A1(n10631), .A2(n10630), .ZN(n10672) );
  INV_X1 U13706 ( .A(n10632), .ZN(n10633) );
  NAND2_X1 U13707 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13708 ( .A1(n10607), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10639) );
  NAND2_X1 U13709 ( .A1(n11188), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10637) );
  AND2_X1 U13710 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10635) );
  NOR2_X1 U13711 ( .A1(n16452), .A2(n10635), .ZN(n10636) );
  NOR2_X1 U13712 ( .A1(n11090), .A2(n10644), .ZN(n10645) );
  OAI21_X1 U13713 ( .B1(n10660), .B2(n10653), .A(n10647), .ZN(n10650) );
  NAND2_X1 U13714 ( .A1(n10648), .A2(n10654), .ZN(n10649) );
  NAND2_X1 U13715 ( .A1(n10650), .A2(n10649), .ZN(n10652) );
  INV_X1 U13716 ( .A(n11089), .ZN(n10651) );
  NAND2_X1 U13717 ( .A1(n10652), .A2(n10651), .ZN(n10659) );
  INV_X1 U13718 ( .A(n10660), .ZN(n11087) );
  INV_X1 U13719 ( .A(n10653), .ZN(n10665) );
  OAI21_X1 U13720 ( .B1(n10665), .B2(n10660), .A(n10654), .ZN(n10655) );
  NAND2_X1 U13721 ( .A1(n10656), .A2(n10655), .ZN(n10657) );
  NAND2_X1 U13722 ( .A1(n10657), .A2(n11089), .ZN(n10658) );
  NAND2_X1 U13723 ( .A1(n10659), .A2(n10658), .ZN(n10668) );
  XNOR2_X1 U13724 ( .A(n10660), .B(n11089), .ZN(n10663) );
  INV_X1 U13725 ( .A(n10663), .ZN(n10661) );
  NAND3_X1 U13726 ( .A1(n10662), .A2(n10661), .A3(n10670), .ZN(n10667) );
  OAI211_X1 U13727 ( .C1(n10665), .C2(n10647), .A(n10663), .B(n10674), .ZN(
        n10666) );
  XNOR2_X2 U13728 ( .A(n10675), .B(n10670), .ZN(n13222) );
  OR2_X2 U13729 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  INV_X1 U13730 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10677) );
  INV_X1 U13731 ( .A(n19606), .ZN(n19603) );
  INV_X1 U13732 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10676) );
  OAI22_X1 U13733 ( .A1(n10678), .A2(n10677), .B1(n19603), .B2(n10676), .ZN(
        n10682) );
  INV_X1 U13734 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10680) );
  INV_X1 U13735 ( .A(n13278), .ZN(n15526) );
  INV_X1 U13736 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10679) );
  OAI22_X1 U13737 ( .A1(n19419), .A2(n10680), .B1(n19758), .B2(n10679), .ZN(
        n10681) );
  NOR2_X1 U13738 ( .A1(n10682), .A2(n10681), .ZN(n10714) );
  INV_X1 U13739 ( .A(n13222), .ZN(n19304) );
  INV_X1 U13740 ( .A(n19323), .ZN(n19320) );
  INV_X1 U13741 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U13742 ( .A1(n19362), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10684) );
  OAI211_X1 U13743 ( .C1(n19320), .C2(n10685), .A(n10684), .B(n14957), .ZN(
        n10690) );
  INV_X1 U13744 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10688) );
  INV_X1 U13745 ( .A(n19663), .ZN(n10687) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10686) );
  OAI22_X1 U13747 ( .A1(n10688), .A2(n19697), .B1(n10687), .B2(n10686), .ZN(
        n10689) );
  NOR2_X1 U13748 ( .A1(n10690), .A2(n10689), .ZN(n10713) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10692) );
  INV_X1 U13750 ( .A(n10809), .ZN(n19456) );
  INV_X1 U13751 ( .A(n10808), .ZN(n19481) );
  INV_X1 U13752 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10691) );
  INV_X1 U13753 ( .A(n10828), .ZN(n19540) );
  INV_X1 U13754 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10695) );
  INV_X1 U13755 ( .A(n10799), .ZN(n19721) );
  INV_X1 U13756 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10694) );
  OAI22_X1 U13757 ( .A1(n19540), .A2(n10695), .B1(n19721), .B2(n10694), .ZN(
        n10696) );
  NOR2_X1 U13758 ( .A1(n10697), .A2(n10696), .ZN(n10712) );
  INV_X1 U13759 ( .A(n19511), .ZN(n19516) );
  INV_X1 U13760 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10701) );
  INV_X1 U13761 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10700) );
  OAI22_X1 U13762 ( .A1(n19516), .A2(n10701), .B1(n19570), .B2(n10700), .ZN(
        n10710) );
  INV_X1 U13763 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10708) );
  INV_X1 U13764 ( .A(n10801), .ZN(n10707) );
  INV_X1 U13765 ( .A(n10810), .ZN(n19638) );
  INV_X1 U13766 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10706) );
  OAI22_X1 U13767 ( .A1(n10708), .A2(n10707), .B1(n19638), .B2(n10706), .ZN(
        n10709) );
  NOR2_X1 U13768 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  AND2_X2 U13769 ( .A1(n14272), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10762) );
  AOI22_X1 U13770 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10720) );
  AND2_X2 U13771 ( .A1(n14270), .A2(n16411), .ZN(n15540) );
  AND2_X2 U13772 ( .A1(n14254), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14109) );
  AOI22_X1 U13773 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14109), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10719) );
  AND2_X2 U13774 ( .A1(n14273), .A2(n16411), .ZN(n10761) );
  AOI22_X1 U13775 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10718) );
  AND2_X2 U13776 ( .A1(n9820), .A2(n16411), .ZN(n10747) );
  AOI22_X1 U13777 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10717) );
  NAND4_X1 U13778 ( .A1(n10720), .A2(n10719), .A3(n10718), .A4(n10717), .ZN(
        n10728) );
  AND2_X2 U13779 ( .A1(n14271), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10733) );
  AND2_X2 U13780 ( .A1(n14272), .A2(n16411), .ZN(n10742) );
  AOI22_X1 U13781 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10726) );
  INV_X1 U13782 ( .A(n10721), .ZN(n10722) );
  NOR2_X1 U13783 ( .A1(n10722), .A2(n16411), .ZN(n10920) );
  AND2_X2 U13784 ( .A1(n10920), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14096) );
  NOR4_X2 U13785 ( .A1(n15529), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U13786 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10725) );
  AND2_X2 U13787 ( .A1(n14264), .A2(n16411), .ZN(n10760) );
  AND2_X2 U13788 ( .A1(n14276), .A2(n16411), .ZN(n10748) );
  AOI22_X1 U13789 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10724) );
  AND2_X2 U13790 ( .A1(n9808), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10839) );
  AND2_X2 U13791 ( .A1(n14273), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10864) );
  AOI22_X1 U13792 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10723) );
  NAND4_X1 U13793 ( .A1(n10726), .A2(n10725), .A3(n10724), .A4(n10723), .ZN(
        n10727) );
  NOR2_X1 U13794 ( .A1(n10728), .A2(n10727), .ZN(n11285) );
  OR2_X1 U13795 ( .A1(n11285), .A2(n14957), .ZN(n13102) );
  INV_X1 U13796 ( .A(n13102), .ZN(n10741) );
  AOI22_X1 U13797 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13798 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10864), .B1(
        n14109), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13799 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13800 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10729) );
  NAND4_X1 U13801 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10740) );
  AOI22_X1 U13802 ( .A1(n10742), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14108), .ZN(n10738) );
  AOI22_X1 U13803 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10762), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13804 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13805 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10735) );
  NAND4_X1 U13806 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10739) );
  NOR2_X1 U13807 ( .A1(n10740), .A2(n10739), .ZN(n11294) );
  INV_X1 U13808 ( .A(n11294), .ZN(n10776) );
  NAND2_X1 U13809 ( .A1(n10741), .A2(n10776), .ZN(n10780) );
  AOI22_X1 U13810 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13811 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13812 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10762), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13813 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10761), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13814 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10754) );
  AOI22_X1 U13815 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13816 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14109), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13817 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10748), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13818 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n11360), .ZN(n10749) );
  NAND4_X1 U13819 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n10753) );
  NAND2_X1 U13820 ( .A1(n10780), .A2(n10897), .ZN(n10755) );
  AOI22_X1 U13821 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10828), .B1(
        n19511), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13822 ( .A1(n10809), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n19663), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13823 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10799), .B1(
        n10810), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13824 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13825 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13826 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10742), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10761), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10763) );
  NAND4_X1 U13828 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10773) );
  AOI22_X1 U13829 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14108), .ZN(n10771) );
  AOI22_X1 U13830 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n9823), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13831 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14109), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13832 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10748), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10768) );
  NAND4_X1 U13833 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n10772) );
  INV_X1 U13834 ( .A(n11311), .ZN(n10774) );
  INV_X1 U13835 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13214) );
  INV_X1 U13836 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12498) );
  NAND2_X1 U13837 ( .A1(n13102), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13101) );
  INV_X1 U13838 ( .A(n13101), .ZN(n10777) );
  XNOR2_X1 U13839 ( .A(n11285), .B(n10776), .ZN(n10778) );
  NAND2_X1 U13840 ( .A1(n10777), .A2(n10778), .ZN(n10779) );
  XOR2_X1 U13841 ( .A(n10778), .B(n10777), .Z(n13111) );
  NAND2_X1 U13842 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13111), .ZN(
        n13110) );
  NAND2_X1 U13843 ( .A1(n10779), .A2(n13110), .ZN(n10781) );
  XNOR2_X1 U13844 ( .A(n13214), .B(n10781), .ZN(n13199) );
  XNOR2_X1 U13845 ( .A(n10897), .B(n10780), .ZN(n13198) );
  NAND2_X1 U13846 ( .A1(n13199), .A2(n13198), .ZN(n13197) );
  NAND2_X1 U13847 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10781), .ZN(
        n10782) );
  NAND2_X1 U13848 ( .A1(n13197), .A2(n10782), .ZN(n10783) );
  XNOR2_X1 U13849 ( .A(n10783), .B(n13577), .ZN(n13572) );
  NAND2_X1 U13850 ( .A1(n10783), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10784) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13852 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13853 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13854 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10761), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10787) );
  NAND4_X1 U13855 ( .A1(n10790), .A2(n10789), .A3(n10788), .A4(n10787), .ZN(
        n10796) );
  AOI22_X1 U13856 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13858 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13859 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n11360), .ZN(n10791) );
  NAND4_X1 U13860 ( .A1(n10794), .A2(n10793), .A3(n10792), .A4(n10791), .ZN(
        n10795) );
  INV_X1 U13861 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13873) );
  INV_X1 U13862 ( .A(n10797), .ZN(n10798) );
  AOI22_X1 U13863 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10828), .B1(
        n19511), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10799), .B1(
        n19663), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13865 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10800), .B1(
        n10801), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13866 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13867 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19422), .B1(
        n10808), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13868 ( .A1(n19362), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13869 ( .A1(n10809), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10810), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13870 ( .A1(n19323), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n19606), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13871 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13872 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13873 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13874 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10815) );
  NAND4_X1 U13875 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10824) );
  AOI22_X1 U13876 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13877 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13878 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13879 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13880 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10823) );
  NOR2_X1 U13881 ( .A1(n10824), .A2(n10823), .ZN(n11319) );
  NAND2_X1 U13882 ( .A1(n11319), .A2(n14227), .ZN(n10825) );
  INV_X1 U13883 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13874) );
  NAND2_X1 U13884 ( .A1(n10961), .A2(n13874), .ZN(n13868) );
  AOI22_X1 U13885 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19422), .B1(
        n19362), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13886 ( .A1(n10828), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10810), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13887 ( .A1(n19323), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10800), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13888 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10829) );
  NAND4_X1 U13889 ( .A1(n10832), .A2(n10831), .A3(n10830), .A4(n10829), .ZN(
        n10838) );
  AOI22_X1 U13890 ( .A1(n10808), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13891 ( .A1(n10809), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10799), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13892 ( .A1(n19511), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n19663), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13893 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10801), .B1(
        n19606), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10833) );
  NAND4_X1 U13894 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10837) );
  AOI22_X1 U13895 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13896 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13897 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13898 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10840) );
  NAND4_X1 U13899 ( .A1(n10843), .A2(n10842), .A3(n10841), .A4(n10840), .ZN(
        n10849) );
  AOI22_X1 U13900 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13901 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13902 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13903 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10844) );
  NAND4_X1 U13904 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10848) );
  NAND2_X1 U13905 ( .A1(n11323), .A2(n9992), .ZN(n10850) );
  NAND2_X1 U13906 ( .A1(n13871), .A2(n9884), .ZN(n10858) );
  NAND2_X1 U13907 ( .A1(n10859), .A2(n10854), .ZN(n10857) );
  NAND2_X1 U13908 ( .A1(n13870), .A2(n10855), .ZN(n10856) );
  NAND3_X1 U13909 ( .A1(n10858), .A2(n10857), .A3(n10856), .ZN(n13961) );
  NAND2_X1 U13910 ( .A1(n13961), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13962) );
  INV_X1 U13911 ( .A(n10859), .ZN(n13871) );
  NAND2_X1 U13912 ( .A1(n13871), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U13913 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10868) );
  NAND2_X1 U13914 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10867) );
  NAND2_X1 U13915 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10866) );
  NAND2_X1 U13916 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10865) );
  NAND2_X1 U13917 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10872) );
  NAND2_X1 U13918 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10871) );
  NAND2_X1 U13919 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10870) );
  NAND2_X1 U13920 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10869) );
  NAND2_X1 U13921 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10876) );
  NAND2_X1 U13922 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10875) );
  NAND2_X1 U13923 ( .A1(n10734), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10874) );
  NAND2_X1 U13924 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14108), .ZN(
        n10873) );
  NAND2_X1 U13925 ( .A1(n10742), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10880) );
  NAND2_X1 U13926 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10879) );
  NAND2_X1 U13927 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10878) );
  NAND2_X1 U13928 ( .A1(n10762), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10877) );
  NAND4_X1 U13929 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10452), .ZN(
        n10933) );
  AND2_X1 U13930 ( .A1(n10884), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13980) );
  INV_X1 U13931 ( .A(n10884), .ZN(n10885) );
  INV_X1 U13932 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U13933 ( .A1(n10885), .A2(n13992), .ZN(n13979) );
  NAND2_X1 U13934 ( .A1(n10887), .A2(n11078), .ZN(n10886) );
  INV_X1 U13935 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10984) );
  INV_X2 U13936 ( .A(n11326), .ZN(n11078) );
  NAND3_X1 U13937 ( .A1(n10887), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11078), .ZN(n10888) );
  INV_X1 U13938 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15462) );
  INV_X1 U13939 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15454) );
  INV_X1 U13940 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16292) );
  NAND2_X1 U13941 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15388) );
  NAND2_X1 U13942 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11455) );
  AND2_X1 U13943 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15349) );
  INV_X1 U13944 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15328) );
  INV_X1 U13945 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12790) );
  NOR2_X2 U13946 ( .A1(n15162), .A2(n12790), .ZN(n15154) );
  AND2_X1 U13947 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15264) );
  NAND2_X1 U13948 ( .A1(n15264), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15262) );
  INV_X1 U13949 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10891) );
  OAI21_X1 U13950 ( .B1(n19994), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10911), .ZN(n10916) );
  MUX2_X1 U13951 ( .A(n11285), .B(n10916), .S(n11228), .Z(n10949) );
  NAND2_X1 U13952 ( .A1(n19984), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10894) );
  NAND2_X1 U13953 ( .A1(n10892), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10893) );
  NAND2_X1 U13954 ( .A1(n10894), .A2(n10893), .ZN(n11216) );
  NAND2_X1 U13955 ( .A1(n16412), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10898) );
  OAI21_X1 U13956 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16412), .A(
        n10898), .ZN(n10896) );
  XNOR2_X1 U13957 ( .A(n10900), .B(n10896), .ZN(n11214) );
  INV_X1 U13958 ( .A(n11214), .ZN(n11223) );
  OAI21_X1 U13959 ( .B1(n10949), .B2(n11216), .A(n10926), .ZN(n10906) );
  AND2_X1 U13960 ( .A1(n10902), .A2(n10901), .ZN(n10903) );
  NOR2_X1 U13961 ( .A1(n10904), .A2(n10903), .ZN(n10913) );
  MUX2_X1 U13962 ( .A(n11311), .B(n10913), .S(n11228), .Z(n10931) );
  NAND3_X1 U13963 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10908), .A3(
        n13099), .ZN(n10914) );
  MUX2_X1 U13964 ( .A(n10914), .B(n10905), .S(n11259), .Z(n10932) );
  NAND3_X1 U13965 ( .A1(n10906), .A2(n10931), .A3(n10932), .ZN(n10909) );
  INV_X1 U13966 ( .A(n11232), .ZN(n11230) );
  NAND2_X1 U13967 ( .A1(n10909), .A2(n11230), .ZN(n20000) );
  NAND2_X1 U13968 ( .A1(n16438), .A2(n12484), .ZN(n11474) );
  INV_X1 U13969 ( .A(n10911), .ZN(n10912) );
  XNOR2_X1 U13970 ( .A(n11216), .B(n10912), .ZN(n11219) );
  AND2_X1 U13971 ( .A1(n11214), .A2(n11226), .ZN(n10917) );
  AND2_X1 U13972 ( .A1(n11219), .A2(n10917), .ZN(n10915) );
  INV_X1 U13973 ( .A(n10916), .ZN(n11220) );
  AOI21_X1 U13974 ( .B1(n11220), .B2(n10917), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n10918) );
  INV_X1 U13975 ( .A(n10918), .ZN(n10919) );
  OR2_X1 U13976 ( .A1(n16430), .A2(n10919), .ZN(n10922) );
  OR2_X1 U13977 ( .A1(n10920), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13093) );
  INV_X1 U13978 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13089) );
  OAI21_X1 U13979 ( .B1(n9824), .B2(n13093), .A(n13089), .ZN(n19990) );
  NAND2_X1 U13980 ( .A1(n19990), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U13981 ( .A1(n16438), .A2(n14957), .ZN(n10923) );
  AND2_X1 U13982 ( .A1(n16437), .A2(n19866), .ZN(n10924) );
  INV_X1 U13983 ( .A(n16358), .ZN(n10925) );
  INV_X1 U13984 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n19201) );
  NAND2_X1 U13985 ( .A1(n10929), .A2(n19201), .ZN(n10930) );
  MUX2_X1 U13986 ( .A(n11294), .B(n10930), .S(n13926), .Z(n10954) );
  INV_X1 U13987 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13714) );
  MUX2_X1 U13988 ( .A(n10931), .B(n13714), .S(n13926), .Z(n10945) );
  INV_X1 U13989 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14040) );
  MUX2_X1 U13990 ( .A(n10932), .B(n14040), .S(n13926), .Z(n10957) );
  NAND2_X1 U13991 ( .A1(n10958), .A2(n10957), .ZN(n10963) );
  MUX2_X1 U13992 ( .A(n11319), .B(P2_EBX_REG_5__SCAN_IN), .S(n13926), .Z(
        n10962) );
  MUX2_X1 U13993 ( .A(n11323), .B(P2_EBX_REG_6__SCAN_IN), .S(n13926), .Z(
        n10967) );
  INV_X1 U13994 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13449) );
  MUX2_X1 U13995 ( .A(n10933), .B(n13449), .S(n13926), .Z(n10978) );
  NAND2_X1 U13996 ( .A1(n11071), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10975) );
  NOR2_X2 U13997 ( .A1(n10981), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n19123) );
  INV_X1 U13998 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U13999 ( .A1(n19123), .A2(n13608), .ZN(n10992) );
  NAND2_X1 U14000 ( .A1(n11071), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10934) );
  AND2_X1 U14001 ( .A1(n11265), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U14002 ( .A1(n13926), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11022) );
  NAND2_X1 U14003 ( .A1(n11071), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U14004 ( .A1(n11071), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11005) );
  INV_X1 U14005 ( .A(n11005), .ZN(n10935) );
  NAND2_X1 U14006 ( .A1(n11071), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11003) );
  INV_X1 U14007 ( .A(n11003), .ZN(n10936) );
  INV_X1 U14008 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U14009 ( .A1(n11011), .A2(n10466), .ZN(n10937) );
  NAND2_X1 U14010 ( .A1(n11071), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14011 ( .A1(n10937), .A2(n11043), .ZN(n11046) );
  NAND2_X1 U14012 ( .A1(n11071), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11042) );
  INV_X1 U14013 ( .A(n11042), .ZN(n10938) );
  NAND2_X1 U14014 ( .A1(n11071), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10939) );
  OR2_X1 U14015 ( .A1(n10940), .A2(n10939), .ZN(n10941) );
  INV_X1 U14016 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14017 ( .A1(n10940), .A2(n11174), .ZN(n11056) );
  XNOR2_X1 U14018 ( .A(n11059), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15144) );
  NAND2_X1 U14019 ( .A1(n11071), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10942) );
  MUX2_X1 U14020 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n10942), .S(n9853), .Z(
        n10943) );
  NAND2_X1 U14021 ( .A1(n10943), .A2(n11011), .ZN(n16253) );
  OR2_X1 U14022 ( .A1(n16253), .A2(n11326), .ZN(n10944) );
  INV_X1 U14023 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15155) );
  NAND2_X1 U14024 ( .A1(n10944), .A2(n15155), .ZN(n15151) );
  NAND2_X1 U14025 ( .A1(n13574), .A2(n11326), .ZN(n10948) );
  NOR2_X1 U14026 ( .A1(n10946), .A2(n10945), .ZN(n10947) );
  OR2_X1 U14027 ( .A1(n10958), .A2(n10947), .ZN(n13713) );
  INV_X1 U14028 ( .A(n10949), .ZN(n10950) );
  MUX2_X1 U14029 ( .A(n10950), .B(P2_EBX_REG_0__SCAN_IN), .S(n13926), .Z(
        n19204) );
  NAND2_X1 U14030 ( .A1(n19204), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13113) );
  NAND3_X1 U14031 ( .A1(n11265), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U14032 ( .A1(n10954), .A2(n10951), .ZN(n19182) );
  NOR2_X1 U14033 ( .A1(n13113), .A2(n19182), .ZN(n10952) );
  NAND2_X1 U14034 ( .A1(n13113), .A2(n19182), .ZN(n13112) );
  OAI21_X1 U14035 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10952), .A(
        n13112), .ZN(n13201) );
  XNOR2_X1 U14036 ( .A(n10954), .B(n10953), .ZN(n14906) );
  XNOR2_X1 U14037 ( .A(n14906), .B(n13214), .ZN(n13200) );
  OR2_X1 U14038 ( .A1(n13201), .A2(n13200), .ZN(n14302) );
  INV_X1 U14039 ( .A(n14906), .ZN(n10955) );
  NAND2_X1 U14040 ( .A1(n10955), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10956) );
  AND2_X1 U14041 ( .A1(n14302), .A2(n10956), .ZN(n13570) );
  XNOR2_X1 U14042 ( .A(n10958), .B(n10957), .ZN(n10959) );
  XNOR2_X1 U14043 ( .A(n10959), .B(n13873), .ZN(n13658) );
  INV_X1 U14044 ( .A(n10959), .ZN(n19169) );
  NAND2_X1 U14045 ( .A1(n19169), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10960) );
  NAND2_X1 U14046 ( .A1(n10963), .A2(n10962), .ZN(n10964) );
  NAND2_X1 U14047 ( .A1(n10968), .A2(n10964), .ZN(n13795) );
  XNOR2_X1 U14048 ( .A(n10965), .B(n13874), .ZN(n13866) );
  NAND2_X1 U14049 ( .A1(n10965), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10966) );
  AND2_X1 U14050 ( .A1(n10968), .A2(n10967), .ZN(n10969) );
  OR2_X1 U14051 ( .A1(n10969), .A2(n10980), .ZN(n13683) );
  INV_X1 U14052 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13973) );
  INV_X1 U14053 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U14054 ( .A1(n10976), .A2(n11111), .ZN(n10974) );
  OAI211_X1 U14055 ( .C1(n10976), .C2(n10975), .A(n10974), .B(n11011), .ZN(
        n19142) );
  OR2_X1 U14056 ( .A1(n19142), .A2(n11326), .ZN(n10985) );
  INV_X1 U14057 ( .A(n10985), .ZN(n10977) );
  NAND2_X1 U14058 ( .A1(n10977), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16337) );
  INV_X1 U14059 ( .A(n10978), .ZN(n10979) );
  XNOR2_X1 U14060 ( .A(n10980), .B(n10979), .ZN(n19155) );
  NAND2_X1 U14061 ( .A1(n19155), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16338) );
  NAND3_X1 U14062 ( .A1(n10981), .A2(n11265), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n10982) );
  NAND2_X1 U14063 ( .A1(n10982), .A2(n11011), .ZN(n10983) );
  OR2_X1 U14064 ( .A1(n10983), .A2(n19123), .ZN(n13693) );
  OAI21_X1 U14065 ( .B1(n13693), .B2(n11326), .A(n15462), .ZN(n15465) );
  NAND2_X1 U14066 ( .A1(n10985), .A2(n10984), .ZN(n16336) );
  OR2_X1 U14067 ( .A1(n19155), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16340) );
  AND2_X1 U14068 ( .A1(n16336), .A2(n16340), .ZN(n15463) );
  NAND2_X1 U14069 ( .A1(n11071), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10986) );
  XNOR2_X1 U14070 ( .A(n10987), .B(n10986), .ZN(n13703) );
  NAND2_X1 U14071 ( .A1(n13703), .A2(n11078), .ZN(n10988) );
  INV_X1 U14072 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14073 ( .A1(n10988), .A2(n11453), .ZN(n15483) );
  AND3_X1 U14074 ( .A1(n15465), .A2(n15463), .A3(n15483), .ZN(n10989) );
  NAND2_X1 U14075 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10990) );
  NOR2_X1 U14076 ( .A1(n13693), .A2(n10990), .ZN(n15466) );
  AND2_X1 U14077 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10991) );
  OR2_X1 U14078 ( .A1(n19124), .A2(n11326), .ZN(n15449) );
  NAND3_X1 U14079 ( .A1(n11265), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n10992), 
        .ZN(n10993) );
  NAND2_X1 U14080 ( .A1(n11019), .A2(n10993), .ZN(n19113) );
  OR2_X1 U14081 ( .A1(n19113), .A2(n11326), .ZN(n10994) );
  INV_X1 U14082 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15443) );
  AND2_X1 U14083 ( .A1(n10994), .A2(n15443), .ZN(n15437) );
  INV_X1 U14084 ( .A(n15437), .ZN(n10995) );
  OR3_X1 U14085 ( .A1(n19113), .A2(n11326), .A3(n15443), .ZN(n15435) );
  NAND3_X1 U14086 ( .A1(n10996), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11265), 
        .ZN(n10997) );
  NAND3_X1 U14087 ( .A1(n10466), .A2(n10997), .A3(n11011), .ZN(n14864) );
  OR2_X1 U14088 ( .A1(n14864), .A2(n11326), .ZN(n10998) );
  INV_X1 U14089 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14090 ( .A1(n10998), .A2(n11472), .ZN(n11211) );
  NAND2_X1 U14091 ( .A1(n11071), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10999) );
  MUX2_X1 U14092 ( .A(n10999), .B(n11265), .S(n9862), .Z(n11000) );
  NAND2_X1 U14093 ( .A1(n11000), .A2(n10996), .ZN(n19068) );
  OR2_X1 U14094 ( .A1(n19068), .A2(n11326), .ZN(n11002) );
  INV_X1 U14095 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11001) );
  NAND2_X1 U14096 ( .A1(n11002), .A2(n11001), .ZN(n15205) );
  XNOR2_X1 U14097 ( .A(n11004), .B(n11003), .ZN(n14874) );
  NAND2_X1 U14098 ( .A1(n14874), .A2(n11078), .ZN(n11030) );
  INV_X1 U14099 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U14100 ( .A1(n11030), .A2(n15363), .ZN(n15214) );
  XNOR2_X1 U14101 ( .A(n11010), .B(n11005), .ZN(n19081) );
  NAND2_X1 U14102 ( .A1(n19081), .A2(n11078), .ZN(n11006) );
  INV_X1 U14103 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U14104 ( .A1(n11006), .A2(n11151), .ZN(n15226) );
  OR2_X1 U14105 ( .A1(n11008), .A2(n11007), .ZN(n11009) );
  NAND2_X1 U14106 ( .A1(n11010), .A2(n11009), .ZN(n14889) );
  INV_X1 U14107 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15394) );
  OAI21_X1 U14108 ( .B1(n14889), .B2(n11326), .A(n15394), .ZN(n11207) );
  AND2_X1 U14109 ( .A1(n11265), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11012) );
  INV_X1 U14110 ( .A(n11011), .ZN(n11048) );
  AOI21_X1 U14111 ( .B1(n11025), .B2(n11012), .A(n11048), .ZN(n11014) );
  NAND2_X1 U14112 ( .A1(n11014), .A2(n11013), .ZN(n19094) );
  OR2_X1 U14113 ( .A1(n19094), .A2(n11326), .ZN(n11015) );
  XNOR2_X1 U14114 ( .A(n11015), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11204) );
  AND2_X1 U14115 ( .A1(n10467), .A2(n11016), .ZN(n11017) );
  OR2_X1 U14116 ( .A1(n11017), .A2(n11023), .ZN(n19103) );
  OAI21_X1 U14117 ( .B1(n19103), .B2(n11326), .A(n16292), .ZN(n16296) );
  NAND2_X1 U14118 ( .A1(n11019), .A2(n11018), .ZN(n11020) );
  NAND2_X1 U14119 ( .A1(n10467), .A2(n11020), .ZN(n13852) );
  OR2_X1 U14120 ( .A1(n13852), .A2(n11326), .ZN(n11021) );
  INV_X1 U14121 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15423) );
  NAND2_X1 U14122 ( .A1(n11021), .A2(n15423), .ZN(n11201) );
  AND2_X1 U14123 ( .A1(n16296), .A2(n11201), .ZN(n11027) );
  OR2_X1 U14124 ( .A1(n11023), .A2(n11022), .ZN(n11024) );
  NAND2_X1 U14125 ( .A1(n11025), .A2(n11024), .ZN(n14899) );
  OR2_X1 U14126 ( .A1(n14899), .A2(n11326), .ZN(n11026) );
  INV_X1 U14127 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U14128 ( .A1(n11026), .A2(n15385), .ZN(n15251) );
  AND4_X1 U14129 ( .A1(n11207), .A2(n11204), .A3(n11027), .A4(n15251), .ZN(
        n11028) );
  NAND2_X1 U14130 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11029) );
  OR2_X1 U14131 ( .A1(n14864), .A2(n11029), .ZN(n11210) );
  OR2_X1 U14132 ( .A1(n11030), .A2(n15363), .ZN(n15215) );
  AND2_X1 U14133 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U14134 ( .A1(n19081), .A2(n11031), .ZN(n15225) );
  AND2_X1 U14135 ( .A1(n15215), .A2(n15225), .ZN(n11208) );
  NAND2_X1 U14136 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11032) );
  OR2_X1 U14137 ( .A1(n14889), .A2(n11032), .ZN(n11206) );
  NAND2_X1 U14138 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11033) );
  OR2_X1 U14139 ( .A1(n14899), .A2(n11033), .ZN(n15250) );
  INV_X1 U14140 ( .A(n19103), .ZN(n11035) );
  AND2_X1 U14141 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14142 ( .A1(n11035), .A2(n11034), .ZN(n16295) );
  NAND2_X1 U14143 ( .A1(n15250), .A2(n16295), .ZN(n11203) );
  NAND2_X1 U14144 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11036) );
  NOR2_X1 U14145 ( .A1(n13852), .A2(n11036), .ZN(n15430) );
  NOR2_X1 U14146 ( .A1(n11203), .A2(n15430), .ZN(n11038) );
  NAND2_X1 U14147 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11037) );
  OR2_X1 U14148 ( .A1(n19094), .A2(n11037), .ZN(n11205) );
  AND3_X1 U14149 ( .A1(n11206), .A2(n11038), .A3(n11205), .ZN(n11040) );
  NAND2_X1 U14150 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11039) );
  AND4_X1 U14151 ( .A1(n11210), .A2(n11208), .A3(n11040), .A4(n15204), .ZN(
        n11041) );
  XNOR2_X1 U14152 ( .A(n11046), .B(n11042), .ZN(n16276) );
  NAND2_X1 U14153 ( .A1(n16276), .A2(n11078), .ZN(n15178) );
  INV_X1 U14154 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15340) );
  INV_X1 U14155 ( .A(n11043), .ZN(n11044) );
  NAND2_X1 U14156 ( .A1(n11044), .A2(n10466), .ZN(n11045) );
  AND2_X1 U14157 ( .A1(n11046), .A2(n11045), .ZN(n15840) );
  NAND2_X1 U14158 ( .A1(n15840), .A2(n11078), .ZN(n15186) );
  AOI22_X1 U14159 ( .A1(n15178), .A2(n15328), .B1(n15340), .B2(n15186), .ZN(
        n11047) );
  NOR2_X1 U14160 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15324) );
  AND2_X1 U14161 ( .A1(n11265), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11049) );
  AOI21_X1 U14162 ( .B1(n11050), .B2(n11049), .A(n11048), .ZN(n11051) );
  NAND2_X1 U14163 ( .A1(n9853), .A2(n11051), .ZN(n16265) );
  NAND2_X1 U14164 ( .A1(n11052), .A2(n12790), .ZN(n15165) );
  INV_X1 U14165 ( .A(n15264), .ZN(n12794) );
  INV_X1 U14166 ( .A(n11077), .ZN(n11054) );
  NAND2_X1 U14167 ( .A1(n11071), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U14168 ( .A1(n11054), .A2(n11055), .ZN(n11066) );
  INV_X1 U14169 ( .A(n11055), .ZN(n11057) );
  NAND2_X1 U14170 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  AND2_X1 U14171 ( .A1(n11066), .A2(n11058), .ZN(n16232) );
  INV_X1 U14172 ( .A(n11059), .ZN(n11060) );
  NAND2_X1 U14173 ( .A1(n11060), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11061) );
  NAND2_X1 U14174 ( .A1(n11061), .A2(n15150), .ZN(n12768) );
  AND2_X1 U14175 ( .A1(n13926), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11065) );
  INV_X1 U14176 ( .A(n11065), .ZN(n11062) );
  XNOR2_X1 U14177 ( .A(n11066), .B(n11062), .ZN(n16225) );
  NAND2_X1 U14178 ( .A1(n16225), .A2(n11078), .ZN(n12771) );
  NOR2_X1 U14179 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12793) );
  NOR2_X1 U14180 ( .A1(n12771), .A2(n12793), .ZN(n11063) );
  NOR2_X1 U14181 ( .A1(n12768), .A2(n11063), .ZN(n11064) );
  INV_X1 U14182 ( .A(n11070), .ZN(n11067) );
  NAND2_X1 U14183 ( .A1(n11071), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11069) );
  XNOR2_X1 U14184 ( .A(n11067), .B(n11069), .ZN(n16210) );
  NAND2_X1 U14185 ( .A1(n16210), .A2(n11078), .ZN(n11068) );
  INV_X1 U14186 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U14187 ( .A1(n11068), .A2(n15269), .ZN(n15125) );
  NAND2_X1 U14188 ( .A1(n11070), .A2(n11069), .ZN(n11075) );
  NAND2_X1 U14189 ( .A1(n11071), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11072) );
  AOI21_X1 U14190 ( .B1(n12535), .B2(n11078), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12455) );
  INV_X1 U14191 ( .A(n12535), .ZN(n11073) );
  INV_X1 U14192 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12851) );
  AND2_X1 U14193 ( .A1(n11078), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U14194 ( .A1(n16210), .A2(n11074), .ZN(n15124) );
  NOR2_X1 U14195 ( .A1(n11075), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11076) );
  MUX2_X1 U14196 ( .A(n11077), .B(n11076), .S(n13926), .Z(n16199) );
  NAND2_X1 U14197 ( .A1(n16199), .A2(n11078), .ZN(n11079) );
  XOR2_X1 U14198 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11079), .Z(
        n11080) );
  INV_X1 U14199 ( .A(n13045), .ZN(n11081) );
  NAND2_X1 U14200 ( .A1(n15506), .A2(n19809), .ZN(n19958) );
  NAND2_X1 U14201 ( .A1(n19958), .A2(n19756), .ZN(n19985) );
  NAND2_X1 U14202 ( .A1(n19985), .A2(n19863), .ZN(n11082) );
  NAND2_X1 U14203 ( .A1(n19633), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14204 ( .A1(n13277), .A2(n11083), .ZN(n13105) );
  NAND2_X1 U14205 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12501), .ZN(
        n12500) );
  NAND2_X1 U14206 ( .A1(n12495), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12493) );
  INV_X1 U14207 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15156) );
  INV_X1 U14208 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12491) );
  INV_X1 U14209 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15135) );
  INV_X1 U14210 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U14211 ( .A1(n9883), .A2(n11089), .B1(n11088), .B2(n10660), .ZN(
        n11094) );
  INV_X1 U14212 ( .A(n11090), .ZN(n11093) );
  INV_X1 U14213 ( .A(n11091), .ZN(n11092) );
  NAND2_X1 U14214 ( .A1(n11138), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11098) );
  AOI22_X1 U14215 ( .A1(n11188), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11097) );
  OAI211_X1 U14216 ( .C1(n14040), .C2(n11147), .A(n11098), .B(n11097), .ZN(
        n13663) );
  INV_X1 U14217 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13302) );
  NAND2_X1 U14218 ( .A1(n11188), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U14219 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11099) );
  OAI211_X1 U14220 ( .C1(n11147), .C2(n13302), .A(n11100), .B(n11099), .ZN(
        n11101) );
  AOI21_X1 U14221 ( .B1(n11138), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11101), .ZN(n13298) );
  NAND2_X1 U14222 ( .A1(n11138), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11106) );
  INV_X1 U14223 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13368) );
  NAND2_X1 U14224 ( .A1(n11188), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U14225 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11102) );
  OAI211_X1 U14226 ( .C1(n11147), .C2(n13368), .A(n11103), .B(n11102), .ZN(
        n11104) );
  INV_X1 U14227 ( .A(n11104), .ZN(n11105) );
  NAND2_X1 U14228 ( .A1(n11106), .A2(n11105), .ZN(n13364) );
  NAND2_X1 U14229 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11108) );
  AOI22_X1 U14230 ( .A1(n11188), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11107) );
  OAI211_X1 U14231 ( .C1(n11147), .C2(n13449), .A(n11108), .B(n11107), .ZN(
        n13447) );
  NAND2_X1 U14232 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11110) );
  AOI22_X1 U14233 ( .A1(n11188), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11109) );
  OAI211_X1 U14234 ( .C1(n11111), .C2(n11147), .A(n11110), .B(n11109), .ZN(
        n13484) );
  INV_X1 U14235 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11114) );
  NAND2_X1 U14236 ( .A1(n11188), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U14237 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11112) );
  OAI211_X1 U14238 ( .C1(n11147), .C2(n11114), .A(n11113), .B(n11112), .ZN(
        n11115) );
  AOI21_X1 U14239 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11115), .ZN(n13533) );
  INV_X1 U14240 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U14241 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11117) );
  AOI22_X1 U14242 ( .A1(n11188), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11116) );
  OAI211_X1 U14243 ( .C1(n11118), .C2(n11147), .A(n11117), .B(n11116), .ZN(
        n13601) );
  NAND2_X1 U14244 ( .A1(n11188), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14245 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11119) );
  OAI211_X1 U14246 ( .C1(n11147), .C2(n13608), .A(n11120), .B(n11119), .ZN(
        n11121) );
  AOI21_X1 U14247 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11121), .ZN(n13606) );
  NAND2_X1 U14248 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11127) );
  INV_X1 U14249 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U14250 ( .A1(n11188), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14251 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11122) );
  OAI211_X1 U14252 ( .C1(n11147), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        n11125) );
  INV_X1 U14253 ( .A(n11125), .ZN(n11126) );
  NAND2_X1 U14254 ( .A1(n11127), .A2(n11126), .ZN(n13641) );
  INV_X1 U14255 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U14256 ( .A1(n11188), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U14257 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11128) );
  OAI211_X1 U14258 ( .C1(n11147), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        n11131) );
  AOI21_X1 U14259 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11131), .ZN(n13674) );
  INV_X1 U14260 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14261 ( .A1(n11188), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14262 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11134) );
  OAI211_X1 U14263 ( .C1(n11147), .C2(n11136), .A(n11135), .B(n11134), .ZN(
        n11137) );
  AOI21_X1 U14264 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11137), .ZN(n13725) );
  AOI22_X1 U14265 ( .A1(n11188), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11140) );
  NAND2_X1 U14266 ( .A1(n10607), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11139) );
  OAI211_X1 U14267 ( .C1(n9814), .C2(n15385), .A(n11140), .B(n11139), .ZN(
        n13803) );
  INV_X1 U14268 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13912) );
  NAND2_X1 U14269 ( .A1(n11188), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11142) );
  NAND2_X1 U14270 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11141) );
  OAI211_X1 U14271 ( .C1(n11147), .C2(n13912), .A(n11142), .B(n11141), .ZN(
        n11143) );
  AOI21_X1 U14272 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11143), .ZN(n13909) );
  INV_X1 U14273 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U14274 ( .A1(n11188), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U14275 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11144) );
  OAI211_X1 U14276 ( .C1(n11147), .C2(n11146), .A(n11145), .B(n11144), .ZN(
        n11148) );
  AOI21_X1 U14277 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11148), .ZN(n13957) );
  AOI22_X1 U14278 ( .A1(n11188), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11150) );
  NAND2_X1 U14279 ( .A1(n10607), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11149) );
  OAI211_X1 U14280 ( .C1(n9814), .C2(n11151), .A(n11150), .B(n11149), .ZN(
        n15005) );
  AOI22_X1 U14281 ( .A1(n11188), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11153) );
  NAND2_X1 U14282 ( .A1(n10607), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11152) );
  OAI211_X1 U14283 ( .C1(n9814), .C2(n15363), .A(n11153), .B(n11152), .ZN(
        n14879) );
  NAND2_X1 U14284 ( .A1(n11188), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U14285 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11154) );
  OAI211_X1 U14286 ( .C1(n11147), .C2(n11156), .A(n11155), .B(n11154), .ZN(
        n11157) );
  AOI21_X1 U14287 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11157), .ZN(n14994) );
  INV_X1 U14288 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11160) );
  NAND2_X1 U14289 ( .A1(n11188), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14290 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11158) );
  OAI211_X1 U14291 ( .C1(n11147), .C2(n11160), .A(n11159), .B(n11158), .ZN(
        n11161) );
  AOI21_X1 U14292 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11161), .ZN(n11459) );
  INV_X1 U14293 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U14294 ( .A1(n11188), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U14295 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11162) );
  OAI211_X1 U14296 ( .C1(n11147), .C2(n11164), .A(n11163), .B(n11162), .ZN(
        n11165) );
  AOI21_X1 U14297 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11165), .ZN(n14979) );
  NOR2_X4 U14298 ( .A1(n14980), .A2(n14979), .ZN(n14982) );
  AOI22_X1 U14299 ( .A1(n11188), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11167) );
  NAND2_X1 U14300 ( .A1(n10607), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11166) );
  OAI211_X1 U14301 ( .C1(n9814), .C2(n15328), .A(n11167), .B(n11166), .ZN(
        n14971) );
  AND2_X2 U14302 ( .A1(n14982), .A2(n14971), .ZN(n14963) );
  AOI22_X1 U14303 ( .A1(n11188), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11169) );
  NAND2_X1 U14304 ( .A1(n10607), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11168) );
  OAI211_X1 U14305 ( .C1(n9814), .C2(n12790), .A(n11169), .B(n11168), .ZN(
        n14962) );
  AND2_X2 U14306 ( .A1(n14963), .A2(n14962), .ZN(n14949) );
  AOI22_X1 U14307 ( .A1(n11188), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11171) );
  NAND2_X1 U14308 ( .A1(n10607), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11170) );
  OAI211_X1 U14309 ( .C1(n9814), .C2(n15155), .A(n11171), .B(n11170), .ZN(
        n14950) );
  NAND2_X1 U14310 ( .A1(n11188), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U14311 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11172) );
  OAI211_X1 U14312 ( .C1(n11147), .C2(n11174), .A(n11173), .B(n11172), .ZN(
        n11175) );
  AOI21_X1 U14313 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11175), .ZN(n14941) );
  OR2_X2 U14314 ( .A1(n14952), .A2(n14941), .ZN(n14943) );
  INV_X1 U14315 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U14316 ( .A1(n11188), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14317 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11176) );
  OAI211_X1 U14318 ( .C1(n11147), .C2(n11178), .A(n11177), .B(n11176), .ZN(
        n11179) );
  AOI21_X1 U14319 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11179), .ZN(n14932) );
  INV_X1 U14320 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U14321 ( .A1(n11188), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11181) );
  NAND2_X1 U14322 ( .A1(n10607), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11180) );
  OAI211_X1 U14323 ( .C1(n9814), .C2(n12776), .A(n11181), .B(n11180), .ZN(
        n12784) );
  AOI22_X1 U14324 ( .A1(n11188), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11183) );
  NAND2_X1 U14325 ( .A1(n10607), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11182) );
  OAI211_X1 U14326 ( .C1(n9814), .C2(n15269), .A(n11183), .B(n11182), .ZN(
        n14924) );
  INV_X1 U14327 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U14328 ( .A1(n11188), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14329 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11184) );
  OAI211_X1 U14330 ( .C1(n11147), .C2(n11186), .A(n11185), .B(n11184), .ZN(
        n11187) );
  AOI21_X1 U14331 ( .B1(n9815), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11187), .ZN(n12457) );
  AOI22_X1 U14332 ( .A1(n11188), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11190) );
  NAND2_X1 U14333 ( .A1(n10607), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11189) );
  OAI211_X1 U14334 ( .C1(n9814), .C2(n10891), .A(n11190), .B(n11189), .ZN(
        n11192) );
  XNOR2_X2 U14335 ( .A(n9851), .B(n11192), .ZN(n16205) );
  AND2_X1 U14336 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19975) );
  NAND2_X1 U14337 ( .A1(n16205), .A2(n19290), .ZN(n11196) );
  NOR2_X1 U14338 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15909) );
  INV_X1 U14339 ( .A(n15909), .ZN(n11193) );
  OR2_X2 U14340 ( .A1(n19958), .A2(n11193), .ZN(n19170) );
  INV_X1 U14341 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11194) );
  NOR2_X1 U14342 ( .A1(n19170), .A2(n11194), .ZN(n12830) );
  AOI21_X1 U14343 ( .B1(n19287), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12830), .ZN(n11195) );
  OAI211_X1 U14344 ( .C1(n19296), .C2(n12488), .A(n11196), .B(n11195), .ZN(
        n11197) );
  INV_X1 U14345 ( .A(n11201), .ZN(n11199) );
  NOR2_X1 U14346 ( .A1(n11199), .A2(n15430), .ZN(n11200) );
  INV_X1 U14347 ( .A(n16296), .ZN(n11202) );
  NOR2_X1 U14348 ( .A1(n16298), .A2(n11202), .ZN(n15253) );
  INV_X1 U14349 ( .A(n11204), .ZN(n15243) );
  NAND2_X1 U14350 ( .A1(n11207), .A2(n11206), .ZN(n15236) );
  NAND3_X1 U14351 ( .A1(n15203), .A2(n15202), .A3(n15205), .ZN(n11209) );
  NAND2_X1 U14352 ( .A1(n11209), .A2(n15204), .ZN(n11212) );
  NAND2_X1 U14353 ( .A1(n11213), .A2(n14957), .ZN(n11215) );
  MUX2_X1 U14354 ( .A(n11215), .B(n11228), .S(n11214), .Z(n11225) );
  INV_X1 U14355 ( .A(n11216), .ZN(n11217) );
  NAND2_X1 U14356 ( .A1(n11217), .A2(n11220), .ZN(n11218) );
  NAND2_X1 U14357 ( .A1(n11259), .A2(n11218), .ZN(n11222) );
  OAI211_X1 U14358 ( .C1(n14957), .C2(n11220), .A(n19317), .B(n11219), .ZN(
        n11221) );
  OAI211_X1 U14359 ( .C1(n13095), .C2(n11223), .A(n11222), .B(n11221), .ZN(
        n11224) );
  NAND2_X1 U14360 ( .A1(n11225), .A2(n11224), .ZN(n11227) );
  MUX2_X1 U14361 ( .A(n11228), .B(n11227), .S(n11226), .Z(n11229) );
  NAND2_X1 U14362 ( .A1(n11230), .A2(n11229), .ZN(n11231) );
  MUX2_X1 U14363 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11231), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11252) );
  NAND2_X1 U14364 ( .A1(n11232), .A2(n13150), .ZN(n11233) );
  AND2_X1 U14365 ( .A1(n16432), .A2(n14957), .ZN(n13147) );
  NAND2_X1 U14366 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16455) );
  INV_X1 U14367 ( .A(n16455), .ZN(n19872) );
  INV_X1 U14368 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19878) );
  NAND2_X2 U14369 ( .A1(n20005), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19946) );
  NOR2_X1 U14370 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19873) );
  INV_X1 U14371 ( .A(n19873), .ZN(n19883) );
  NAND3_X1 U14372 ( .A1(n19878), .A2(n19946), .A3(n19883), .ZN(n19877) );
  NOR2_X1 U14373 ( .A1(n19872), .A2(n19877), .ZN(n13042) );
  NAND3_X1 U14374 ( .A1(n13147), .A2(n13042), .A3(n11440), .ZN(n11257) );
  MUX2_X1 U14375 ( .A(n11234), .B(n19332), .S(n9992), .Z(n11235) );
  OR2_X1 U14376 ( .A1(n11235), .A2(n19872), .ZN(n11249) );
  OR2_X1 U14377 ( .A1(n16430), .A2(n11236), .ZN(n11248) );
  NAND2_X1 U14378 ( .A1(n11237), .A2(n13925), .ZN(n11238) );
  NAND2_X1 U14379 ( .A1(n11238), .A2(n12484), .ZN(n11436) );
  AND2_X1 U14380 ( .A1(n11239), .A2(n11436), .ZN(n11244) );
  NAND2_X1 U14381 ( .A1(n9992), .A2(n11441), .ZN(n11431) );
  NAND2_X1 U14382 ( .A1(n11431), .A2(n19317), .ZN(n11241) );
  NAND3_X1 U14383 ( .A1(n11241), .A2(n11240), .A3(n11437), .ZN(n11242) );
  NAND2_X1 U14384 ( .A1(n13145), .A2(n11242), .ZN(n11243) );
  NAND2_X1 U14385 ( .A1(n11244), .A2(n11243), .ZN(n11434) );
  INV_X1 U14386 ( .A(n11245), .ZN(n11246) );
  NOR2_X1 U14387 ( .A1(n11434), .A2(n11246), .ZN(n11247) );
  OAI21_X1 U14388 ( .B1(n16430), .B2(n11249), .A(n13087), .ZN(n11250) );
  NOR2_X1 U14389 ( .A1(n11251), .A2(n11250), .ZN(n11256) );
  INV_X1 U14390 ( .A(n13147), .ZN(n11254) );
  AOI21_X1 U14391 ( .B1(n11252), .B2(n19317), .A(n19339), .ZN(n11253) );
  NAND2_X1 U14392 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  NAND3_X1 U14393 ( .A1(n11257), .A2(n11256), .A3(n11255), .ZN(n11258) );
  AND2_X1 U14394 ( .A1(n16438), .A2(n11259), .ZN(n19997) );
  INV_X1 U14395 ( .A(n11261), .ZN(n11262) );
  NAND2_X1 U14396 ( .A1(n11260), .A2(n11262), .ZN(n13086) );
  NAND2_X1 U14397 ( .A1(n13086), .A2(n11263), .ZN(n11264) );
  AND2_X1 U14398 ( .A1(n13925), .A2(n19809), .ZN(n11295) );
  INV_X1 U14399 ( .A(n11305), .ZN(n12477) );
  NOR2_X1 U14400 ( .A1(n14957), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11266) );
  AND2_X1 U14401 ( .A1(n11267), .A2(n11266), .ZN(n11301) );
  AOI22_X1 U14402 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14403 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14404 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14405 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11268) );
  NAND4_X1 U14406 ( .A1(n11271), .A2(n11270), .A3(n11269), .A4(n11268), .ZN(
        n11277) );
  AOI22_X1 U14407 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14408 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14409 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14410 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11272) );
  NAND4_X1 U14411 ( .A1(n11275), .A2(n11274), .A3(n11273), .A4(n11272), .ZN(
        n11276) );
  INV_X1 U14412 ( .A(n13482), .ZN(n11281) );
  NOR2_X1 U14413 ( .A1(n13925), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11278) );
  INV_X2 U14414 ( .A(n11328), .ZN(n12478) );
  AND2_X2 U14415 ( .A1(n11279), .A2(n19809), .ZN(n11291) );
  AOI22_X1 U14416 ( .A1(n12478), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11280) );
  OAI21_X1 U14417 ( .B1(n11406), .B2(n11281), .A(n11280), .ZN(n11282) );
  AOI21_X1 U14418 ( .B1(n12477), .B2(P2_REIP_REG_8__SCAN_IN), .A(n11282), .ZN(
        n16385) );
  INV_X1 U14419 ( .A(n13182), .ZN(n13184) );
  NAND2_X1 U14420 ( .A1(n13184), .A2(n11291), .ZN(n11303) );
  INV_X1 U14421 ( .A(n11295), .ZN(n11283) );
  NAND2_X1 U14422 ( .A1(n19994), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19986) );
  NAND2_X1 U14423 ( .A1(n11283), .A2(n19986), .ZN(n11284) );
  AND2_X1 U14424 ( .A1(n11303), .A2(n11284), .ZN(n11288) );
  INV_X1 U14425 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19060) );
  NAND2_X1 U14426 ( .A1(n11327), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11290) );
  AOI21_X1 U14427 ( .B1(n19352), .B2(P2_EAX_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11289) );
  OAI211_X1 U14428 ( .C1(n14227), .C2(n12498), .A(n11290), .B(n11289), .ZN(
        n13185) );
  NAND2_X1 U14429 ( .A1(n12477), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11293) );
  INV_X1 U14430 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19298) );
  AOI22_X1 U14431 ( .A1(n11278), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11292) );
  NAND2_X1 U14432 ( .A1(n11293), .A2(n11292), .ZN(n11298) );
  XNOR2_X1 U14433 ( .A(n13188), .B(n11298), .ZN(n13307) );
  OR2_X1 U14434 ( .A1(n11294), .A2(n11406), .ZN(n11297) );
  AOI22_X1 U14435 ( .A1(n13182), .A2(n11295), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U14436 ( .A1(n11297), .A2(n11296), .ZN(n13306) );
  NOR2_X1 U14437 ( .A1(n13307), .A2(n13306), .ZN(n11300) );
  NOR2_X1 U14438 ( .A1(n13188), .A2(n11298), .ZN(n11299) );
  NAND2_X1 U14439 ( .A1(n11301), .A2(n11302), .ZN(n11304) );
  OAI211_X1 U14440 ( .C1(n19809), .C2(n19973), .A(n11304), .B(n11303), .ZN(
        n11308) );
  XNOR2_X1 U14441 ( .A(n11309), .B(n11308), .ZN(n13194) );
  NAND2_X1 U14442 ( .A1(n11327), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14443 ( .A1(n12478), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U14444 ( .A1(n11307), .A2(n11306), .ZN(n13193) );
  NOR2_X1 U14445 ( .A1(n13194), .A2(n13193), .ZN(n13195) );
  NOR2_X1 U14446 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  NAND2_X1 U14447 ( .A1(n11327), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11315) );
  NAND2_X1 U14448 ( .A1(n11301), .A2(n11311), .ZN(n11314) );
  AOI22_X1 U14449 ( .A1(n11291), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11313) );
  NAND2_X1 U14450 ( .A1(n12478), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11312) );
  NAND4_X1 U14451 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n13493) );
  AOI22_X1 U14452 ( .A1(n12478), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11316) );
  OAI21_X1 U14453 ( .B1(n11406), .B2(n11317), .A(n11316), .ZN(n11318) );
  AOI21_X1 U14454 ( .B1(n12477), .B2(P2_REIP_REG_4__SCAN_IN), .A(n11318), .ZN(
        n13591) );
  AOI22_X1 U14455 ( .A1(n11327), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11322) );
  INV_X1 U14456 ( .A(n11319), .ZN(n11320) );
  AOI22_X1 U14457 ( .A1(n11301), .A2(n11320), .B1(n12478), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U14458 ( .A1(n11322), .A2(n11321), .ZN(n13794) );
  INV_X1 U14459 ( .A(n13793), .ZN(n13239) );
  NOR2_X1 U14460 ( .A1(n11406), .A2(n11323), .ZN(n13238) );
  NAND2_X1 U14461 ( .A1(n11327), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14462 ( .A1(n12478), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14463 ( .A1(n11325), .A2(n11324), .ZN(n13237) );
  OAI21_X1 U14464 ( .B1(n13239), .B2(n13238), .A(n13237), .ZN(n13241) );
  INV_X1 U14465 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19269) );
  INV_X1 U14466 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19902) );
  OAI222_X1 U14467 ( .A1(n13992), .A2(n11329), .B1(n11328), .B2(n19269), .C1(
        n11305), .C2(n19902), .ZN(n13267) );
  NAND2_X1 U14468 ( .A1(n11327), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14469 ( .A1(n12478), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14470 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10760), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14471 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14472 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10742), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14473 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10864), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11330) );
  NAND4_X1 U14474 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11339) );
  AOI22_X1 U14475 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14476 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14477 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14478 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14108), .ZN(n11334) );
  NAND4_X1 U14479 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  NOR2_X1 U14480 ( .A1(n11339), .A2(n11338), .ZN(n13530) );
  NAND2_X1 U14481 ( .A1(n11301), .A2(n13531), .ZN(n11340) );
  NAND3_X1 U14482 ( .A1(n11342), .A2(n11341), .A3(n11340), .ZN(n13443) );
  NAND2_X1 U14483 ( .A1(n11327), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14484 ( .A1(n12478), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14486 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14487 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14488 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10761), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11343) );
  NAND4_X1 U14489 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n11352) );
  AOI22_X1 U14490 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14491 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14492 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14493 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n11360), .ZN(n11347) );
  NAND4_X1 U14494 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11351) );
  NOR2_X1 U14495 ( .A1(n11352), .A2(n11351), .ZN(n13631) );
  INV_X1 U14496 ( .A(n13631), .ZN(n13598) );
  NAND2_X1 U14497 ( .A1(n11301), .A2(n13598), .ZN(n11353) );
  AOI22_X1 U14498 ( .A1(n11327), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n12478), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14499 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10839), .B1(
        n10760), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14500 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14501 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14502 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10761), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14503 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11366) );
  AOI22_X1 U14504 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14505 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14506 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14507 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n11360), .ZN(n11361) );
  NAND4_X1 U14508 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  AOI22_X1 U14509 ( .A1(n11301), .A2(n13630), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n11291), .ZN(n11367) );
  NAND2_X1 U14510 ( .A1(n11368), .A2(n11367), .ZN(n13538) );
  AOI22_X1 U14511 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14512 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14513 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10761), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11369) );
  NAND4_X1 U14515 ( .A1(n11372), .A2(n11371), .A3(n11370), .A4(n11369), .ZN(
        n11378) );
  AOI22_X1 U14516 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14517 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14518 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14519 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14108), .ZN(n11373) );
  NAND4_X1 U14520 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  INV_X1 U14521 ( .A(n13629), .ZN(n13635) );
  AOI22_X1 U14522 ( .A1(n12478), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11379) );
  OAI21_X1 U14523 ( .B1(n11406), .B2(n13635), .A(n11379), .ZN(n11380) );
  AOI21_X1 U14524 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n11327), .A(n11380), 
        .ZN(n15440) );
  INV_X1 U14525 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14526 ( .A1(n12478), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14527 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14528 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14529 ( .A1(n10742), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14530 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11381) );
  NAND4_X1 U14531 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11390) );
  AOI22_X1 U14532 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14533 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14109), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14534 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14535 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11385) );
  NAND4_X1 U14536 ( .A1(n11388), .A2(n11387), .A3(n11386), .A4(n11385), .ZN(
        n11389) );
  NAND2_X1 U14537 ( .A1(n11301), .A2(n13676), .ZN(n11391) );
  OAI211_X1 U14538 ( .C1(n11305), .C2(n11393), .A(n11392), .B(n11391), .ZN(
        n13648) );
  AOI22_X1 U14539 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14540 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14541 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14542 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14543 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11403) );
  AOI22_X1 U14544 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14545 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14546 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14547 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14548 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11402) );
  INV_X1 U14549 ( .A(n13724), .ZN(n11405) );
  AOI22_X1 U14550 ( .A1(n12478), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11404) );
  OAI21_X1 U14551 ( .B1(n11406), .B2(n11405), .A(n11404), .ZN(n11407) );
  AOI21_X1 U14552 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n11327), .A(n11407), 
        .ZN(n16368) );
  NOR2_X4 U14553 ( .A1(n16367), .A2(n16368), .ZN(n16366) );
  AOI22_X1 U14554 ( .A1(n11327), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n12478), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14555 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14556 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14558 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10762), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11408) );
  NAND4_X1 U14559 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11417) );
  AOI22_X1 U14560 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14561 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14562 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14563 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14564 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11416) );
  NOR2_X1 U14565 ( .A1(n11417), .A2(n11416), .ZN(n13807) );
  INV_X1 U14566 ( .A(n13807), .ZN(n13809) );
  AOI22_X1 U14567 ( .A1(n11301), .A2(n13809), .B1(n11291), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14568 ( .A1(n11419), .A2(n11418), .ZN(n13832) );
  NAND2_X1 U14569 ( .A1(n11327), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14570 ( .A1(n12478), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11420) );
  INV_X1 U14571 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19921) );
  AOI22_X1 U14572 ( .A1(n12478), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11422) );
  OAI21_X1 U14573 ( .B1(n11305), .B2(n19921), .A(n11422), .ZN(n14884) );
  NAND2_X1 U14574 ( .A1(n11327), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14575 ( .A1(n12478), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11423) );
  INV_X1 U14576 ( .A(n11425), .ZN(n15100) );
  NAND2_X1 U14577 ( .A1(n11327), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14578 ( .A1(n12478), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11426) );
  NOR2_X2 U14579 ( .A1(n15100), .A2(n14872), .ZN(n15082) );
  INV_X1 U14580 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U14581 ( .A1(n12478), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11428) );
  OAI21_X1 U14582 ( .B1(n11305), .B2(n19927), .A(n11428), .ZN(n15081) );
  AND2_X2 U14583 ( .A1(n15082), .A2(n15081), .ZN(n15084) );
  INV_X1 U14584 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U14585 ( .A1(n12478), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11429) );
  OAI21_X1 U14586 ( .B1(n11305), .B2(n19929), .A(n11429), .ZN(n11430) );
  OAI21_X1 U14587 ( .B1(n15084), .B2(n11430), .A(n15064), .ZN(n14871) );
  INV_X1 U14588 ( .A(n14871), .ZN(n15078) );
  INV_X1 U14589 ( .A(n11431), .ZN(n11432) );
  NAND2_X1 U14590 ( .A1(n11432), .A2(n13184), .ZN(n11433) );
  NAND2_X1 U14591 ( .A1(n11435), .A2(n14957), .ZN(n15497) );
  NAND2_X1 U14592 ( .A1(n15497), .A2(n11436), .ZN(n11438) );
  NAND2_X1 U14593 ( .A1(n11438), .A2(n11437), .ZN(n11450) );
  AOI22_X1 U14594 ( .A1(n14043), .A2(n11441), .B1(n16437), .B2(n11440), .ZN(
        n11447) );
  NAND2_X1 U14595 ( .A1(n11442), .A2(n10597), .ZN(n11443) );
  NAND2_X1 U14596 ( .A1(n11443), .A2(n11439), .ZN(n11445) );
  NAND2_X1 U14597 ( .A1(n11445), .A2(n11444), .ZN(n11446) );
  AND3_X1 U14598 ( .A1(n11448), .A2(n11447), .A3(n11446), .ZN(n11449) );
  NAND2_X1 U14599 ( .A1(n11450), .A2(n11449), .ZN(n15544) );
  OR2_X1 U14600 ( .A1(n15544), .A2(n13168), .ZN(n11451) );
  NOR2_X1 U14601 ( .A1(n13874), .A2(n13873), .ZN(n13872) );
  INV_X1 U14602 ( .A(n13872), .ZN(n13968) );
  NOR3_X1 U14603 ( .A1(n13973), .A2(n13577), .A3(n13968), .ZN(n13990) );
  NOR2_X1 U14604 ( .A1(n12498), .A2(n19298), .ZN(n11463) );
  NOR2_X1 U14605 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11463), .ZN(
        n13576) );
  INV_X1 U14606 ( .A(n13576), .ZN(n13204) );
  NAND4_X1 U14607 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n13990), .A4(n13204), .ZN(
        n11454) );
  INV_X1 U14608 ( .A(n11463), .ZN(n19301) );
  NAND2_X1 U14609 ( .A1(n15386), .A2(n19301), .ZN(n11452) );
  INV_X2 U14610 ( .A(n19170), .ZN(n19286) );
  OR2_X1 U14611 ( .A1(n11475), .A2(n19286), .ZN(n19297) );
  NAND2_X1 U14612 ( .A1(n15386), .A2(n13214), .ZN(n13209) );
  NAND2_X1 U14613 ( .A1(n13213), .A2(n13209), .ZN(n13575) );
  AOI211_X1 U14614 ( .C1(n19302), .C2(n11454), .A(n11453), .B(n13575), .ZN(
        n15487) );
  NAND2_X1 U14615 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11467) );
  INV_X1 U14616 ( .A(n11467), .ZN(n15453) );
  NAND2_X1 U14617 ( .A1(n15487), .A2(n15453), .ZN(n15425) );
  AND2_X1 U14618 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16378) );
  NAND2_X1 U14619 ( .A1(n16378), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16376) );
  NOR2_X1 U14620 ( .A1(n15425), .A2(n16376), .ZN(n15380) );
  OR2_X1 U14621 ( .A1(n15388), .A2(n11455), .ZN(n11469) );
  INV_X1 U14622 ( .A(n11469), .ZN(n11456) );
  NAND2_X1 U14623 ( .A1(n15380), .A2(n11456), .ZN(n15358) );
  NAND2_X1 U14624 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15349), .ZN(
        n11457) );
  NOR2_X1 U14625 ( .A1(n15358), .A2(n11457), .ZN(n12780) );
  OR2_X1 U14626 ( .A1(n12780), .A2(n15452), .ZN(n15341) );
  INV_X1 U14627 ( .A(n14980), .ZN(n11458) );
  AOI21_X1 U14628 ( .B1(n11459), .B2(n14995), .A(n11458), .ZN(n15199) );
  NAND2_X1 U14629 ( .A1(n16416), .A2(n9992), .ZN(n11460) );
  NAND2_X1 U14630 ( .A1(n11460), .A2(n15520), .ZN(n11461) );
  NAND2_X1 U14631 ( .A1(n19286), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15194) );
  INV_X1 U14632 ( .A(n15194), .ZN(n11462) );
  AOI21_X1 U14633 ( .B1(n15199), .B2(n16390), .A(n11462), .ZN(n11471) );
  NAND2_X1 U14634 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16393) );
  NAND2_X1 U14635 ( .A1(n15381), .A2(n13204), .ZN(n11466) );
  NAND2_X1 U14636 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11463), .ZN(
        n13205) );
  INV_X1 U14637 ( .A(n13205), .ZN(n11464) );
  NAND2_X1 U14638 ( .A1(n15386), .A2(n11464), .ZN(n11465) );
  NAND2_X1 U14639 ( .A1(n11466), .A2(n11465), .ZN(n13662) );
  NAND2_X1 U14640 ( .A1(n13990), .A2(n13662), .ZN(n13991) );
  NOR2_X1 U14641 ( .A1(n16393), .A2(n13991), .ZN(n15489) );
  NAND2_X1 U14642 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15489), .ZN(
        n15470) );
  INV_X1 U14643 ( .A(n16376), .ZN(n11468) );
  NAND2_X1 U14644 ( .A1(n16377), .A2(n11468), .ZN(n15415) );
  NOR2_X1 U14645 ( .A1(n15415), .A2(n11469), .ZN(n15364) );
  NAND3_X1 U14646 ( .A1(n15364), .A2(n15349), .A3(n11472), .ZN(n11470) );
  OAI211_X1 U14647 ( .C1(n15341), .C2(n11472), .A(n11471), .B(n11470), .ZN(
        n11477) );
  NOR2_X1 U14648 ( .A1(n9854), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15196) );
  INV_X1 U14649 ( .A(n11474), .ZN(n19999) );
  NOR3_X1 U14650 ( .A1(n15196), .A2(n11473), .A3(n19311), .ZN(n11476) );
  AOI211_X1 U14651 ( .C1(n19308), .C2(n15078), .A(n11477), .B(n11476), .ZN(
        n11478) );
  INV_X1 U14652 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11479) );
  INV_X1 U14653 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14654 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11485) );
  AND2_X2 U14655 ( .A1(n11487), .A2(n11488), .ZN(n11547) );
  BUF_X4 U14656 ( .A(n11547), .Z(n11593) );
  AOI22_X1 U14657 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11484) );
  NOR2_X4 U14658 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U14659 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11483) );
  BUF_X4 U14660 ( .A(n11529), .Z(n12549) );
  AOI22_X1 U14661 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14662 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11494) );
  AOI22_X1 U14664 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11492) );
  AND2_X2 U14665 ( .A1(n13377), .A2(n13380), .ZN(n11714) );
  AOI22_X1 U14666 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11491) );
  AND2_X2 U14667 ( .A1(n11486), .A2(n13377), .ZN(n11534) );
  AOI22_X1 U14668 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11490) );
  AND2_X2 U14669 ( .A1(n11487), .A2(n13380), .ZN(n11583) );
  AOI22_X1 U14670 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11489) );
  NAND4_X1 U14671 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11493) );
  NOR2_X1 U14672 ( .A1(n11494), .A2(n11493), .ZN(n11520) );
  AOI21_X1 U14673 ( .B1(n11559), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n11495), .ZN(n11499) );
  AOI22_X1 U14674 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14675 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14676 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14677 ( .A1(n11592), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14678 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14679 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14680 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11796) );
  INV_X1 U14681 ( .A(n11796), .ZN(n11506) );
  XNOR2_X1 U14682 ( .A(n11918), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14004) );
  NAND2_X1 U14683 ( .A1(n14004), .A2(n12566), .ZN(n11519) );
  AOI22_X1 U14684 ( .A1(n11714), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14685 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11592), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14686 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14687 ( .A1(n11668), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11547), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14688 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14689 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11512) );
  NAND2_X2 U14690 ( .A1(n11517), .A2(n11516), .ZN(n11554) );
  AOI22_X1 U14691 ( .A1(n12569), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12568), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14692 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14693 ( .A1(n11592), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14694 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14695 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14696 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14697 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14698 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14699 ( .A1(n11592), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14700 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14701 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14702 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14703 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11598), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11536) );
  NAND3_X1 U14704 ( .A1(n11625), .A2(n11540), .A3(n11570), .ZN(n11555) );
  AOI22_X1 U14705 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14706 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14707 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14708 ( .A1(n11592), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14709 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11600), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11548) );
  NAND2_X2 U14710 ( .A1(n11553), .A2(n11552), .ZN(n11609) );
  INV_X1 U14711 ( .A(n11556), .ZN(n11557) );
  NAND2_X1 U14712 ( .A1(n11558), .A2(n11557), .ZN(n11622) );
  AOI22_X1 U14713 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14714 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U14715 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11569) );
  AOI22_X1 U14716 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14717 ( .A1(n11592), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14718 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11565) );
  NAND4_X1 U14719 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(
        n11568) );
  OR2_X4 U14720 ( .A1(n11569), .A2(n11568), .ZN(n20204) );
  NAND2_X1 U14721 ( .A1(n11541), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U14722 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14723 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11572) );
  NAND2_X1 U14724 ( .A1(n11534), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14725 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U14726 ( .A1(n11668), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11577) );
  NAND2_X1 U14727 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11576) );
  NAND2_X1 U14728 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U14729 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U14730 ( .A1(n11592), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11581) );
  NAND2_X1 U14731 ( .A1(n11703), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U14732 ( .A1(n11673), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11579) );
  NAND2_X1 U14733 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11587) );
  NAND2_X1 U14734 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11586) );
  NAND2_X1 U14735 ( .A1(n11714), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11585) );
  NAND2_X1 U14736 ( .A1(n11600), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11584) );
  AND4_X4 U14737 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n12696) );
  INV_X1 U14738 ( .A(n12312), .ZN(n11607) );
  AOI22_X1 U14739 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11592), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14740 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14741 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14742 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U14743 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11606) );
  AOI22_X1 U14744 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11541), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14745 ( .A1(n11714), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14746 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14747 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n11605) );
  NAND2_X1 U14748 ( .A1(n11607), .A2(n9812), .ZN(n12572) );
  NAND2_X1 U14749 ( .A1(n11646), .A2(n11610), .ZN(n11611) );
  INV_X1 U14750 ( .A(n11620), .ZN(n11613) );
  INV_X1 U14751 ( .A(n12576), .ZN(n11612) );
  NAND2_X1 U14752 ( .A1(n11614), .A2(n11616), .ZN(n11615) );
  NAND2_X1 U14753 ( .A1(n10434), .A2(n11618), .ZN(n12729) );
  OAI211_X1 U14754 ( .C1(n13541), .C2(n11721), .A(n12737), .B(n12729), .ZN(
        n11619) );
  INV_X1 U14755 ( .A(n11619), .ZN(n11632) );
  NAND2_X1 U14756 ( .A1(n12696), .A2(n11616), .ZN(n13778) );
  INV_X1 U14757 ( .A(n11621), .ZN(n11633) );
  NAND2_X1 U14758 ( .A1(n12712), .A2(n11618), .ZN(n11624) );
  INV_X1 U14759 ( .A(n20204), .ZN(n11626) );
  NAND2_X1 U14760 ( .A1(n11625), .A2(n11626), .ZN(n13376) );
  XNOR2_X1 U14761 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12421) );
  MUX2_X1 U14762 ( .A(n20766), .B(n12815), .S(n20866), .Z(n11722) );
  INV_X1 U14763 ( .A(n11722), .ZN(n11629) );
  INV_X1 U14764 ( .A(n12736), .ZN(n11631) );
  AND2_X2 U14765 ( .A1(n12696), .A2(n9812), .ZN(n14313) );
  NAND3_X1 U14766 ( .A1(n13777), .A2(n11608), .A3(n20204), .ZN(n11630) );
  NAND2_X1 U14767 ( .A1(n11631), .A2(n11630), .ZN(n11641) );
  INV_X1 U14768 ( .A(n13541), .ZN(n12666) );
  NAND2_X1 U14769 ( .A1(n12666), .A2(n11633), .ZN(n11636) );
  NAND2_X1 U14770 ( .A1(n16188), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20011) );
  INV_X1 U14771 ( .A(n20011), .ZN(n11635) );
  NAND2_X1 U14772 ( .A1(n12727), .A2(n11634), .ZN(n12738) );
  AND4_X1 U14773 ( .A1(n11636), .A2(n11635), .A3(n12738), .A4(n13778), .ZN(
        n11639) );
  NAND3_X1 U14774 ( .A1(n11637), .A2(n11616), .A3(n14846), .ZN(n11638) );
  AND3_X1 U14775 ( .A1(n11632), .A2(n11639), .A3(n11638), .ZN(n11640) );
  NAND2_X1 U14776 ( .A1(n11641), .A2(n11640), .ZN(n11760) );
  INV_X1 U14777 ( .A(n12815), .ZN(n11642) );
  NAND2_X1 U14778 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11662) );
  OAI21_X1 U14779 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11662), .ZN(n20520) );
  NAND2_X1 U14780 ( .A1(n20766), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11655) );
  OAI21_X1 U14781 ( .B1(n11642), .B2(n20520), .A(n11655), .ZN(n11643) );
  INV_X1 U14782 ( .A(n11643), .ZN(n11644) );
  NAND3_X1 U14783 ( .A1(n14313), .A2(n12727), .A3(n11646), .ZN(n13316) );
  XNOR2_X2 U14784 ( .A(n11653), .B(n11654), .ZN(n11685) );
  INV_X1 U14785 ( .A(n11654), .ZN(n11657) );
  NAND2_X1 U14786 ( .A1(n11655), .A2(n13400), .ZN(n11656) );
  NAND2_X1 U14787 ( .A1(n11657), .A2(n11656), .ZN(n11658) );
  INV_X1 U14788 ( .A(n11662), .ZN(n11661) );
  NAND2_X1 U14789 ( .A1(n11661), .A2(n15856), .ZN(n20553) );
  NAND2_X1 U14790 ( .A1(n11662), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11663) );
  NAND2_X1 U14791 ( .A1(n20553), .A2(n11663), .ZN(n20190) );
  NAND2_X1 U14792 ( .A1(n20190), .A2(n12815), .ZN(n11665) );
  NAND2_X1 U14793 ( .A1(n20766), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11664) );
  AOI22_X1 U14794 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14795 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14796 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14797 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14798 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11679) );
  AOI22_X1 U14799 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14800 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14801 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14802 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11674) );
  NAND4_X1 U14803 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11678) );
  NAND2_X1 U14804 ( .A1(n12696), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11779) );
  INV_X1 U14805 ( .A(n11779), .ZN(n11683) );
  INV_X1 U14806 ( .A(n11685), .ZN(n11688) );
  INV_X1 U14807 ( .A(n11686), .ZN(n11687) );
  AOI22_X1 U14808 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14809 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11593), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14810 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14811 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14812 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11698) );
  AOI22_X1 U14813 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14814 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14815 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14816 ( .A1(n12084), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14817 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11697) );
  AOI22_X1 U14818 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14819 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14820 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14821 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11699) );
  NAND4_X1 U14822 ( .A1(n11702), .A2(n11701), .A3(n11700), .A4(n11699), .ZN(
        n11709) );
  AOI22_X1 U14823 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14824 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11593), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14825 ( .A1(n12084), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11534), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14826 ( .A1(n11703), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11704) );
  NAND4_X1 U14827 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11708) );
  AOI22_X1 U14828 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14829 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14830 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14831 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U14832 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11720) );
  AOI22_X1 U14833 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14834 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14835 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14836 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11715) );
  NAND4_X1 U14837 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n11719) );
  NOR2_X1 U14838 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11722), .ZN(n11724) );
  NOR2_X1 U14839 ( .A1(n11736), .A2(n11725), .ZN(n11723) );
  INV_X1 U14840 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U14841 ( .A1(n12696), .A2(n12610), .ZN(n11727) );
  NAND2_X1 U14842 ( .A1(n11727), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11728) );
  NOR2_X1 U14843 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  INV_X1 U14844 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11733) );
  OR2_X1 U14845 ( .A1(n11734), .A2(n11779), .ZN(n11735) );
  INV_X1 U14846 ( .A(n11738), .ZN(n11739) );
  NOR2_X1 U14847 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  INV_X1 U14848 ( .A(n11743), .ZN(n11742) );
  NAND2_X1 U14849 ( .A1(n11744), .A2(n11794), .ZN(n12617) );
  INV_X1 U14850 ( .A(n11647), .ZN(n11745) );
  NAND2_X1 U14851 ( .A1(n11745), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11822) );
  XNOR2_X1 U14852 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13816) );
  AOI21_X1 U14853 ( .B1(n11507), .B2(n13816), .A(n12568), .ZN(n11747) );
  NAND2_X1 U14854 ( .A1(n12569), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11746) );
  OAI211_X1 U14855 ( .C1(n11822), .C2(n11660), .A(n11747), .B(n11746), .ZN(
        n11748) );
  INV_X1 U14856 ( .A(n11748), .ZN(n11749) );
  OAI21_X1 U14857 ( .B1(n12617), .B2(n11951), .A(n11749), .ZN(n11750) );
  NAND2_X1 U14858 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14859 ( .A1(n11750), .A2(n11774), .ZN(n13435) );
  INV_X1 U14860 ( .A(n13435), .ZN(n11773) );
  INV_X1 U14861 ( .A(n12605), .ZN(n11753) );
  XNOR2_X2 U14862 ( .A(n11753), .B(n11752), .ZN(n13427) );
  NAND2_X1 U14863 ( .A1(n13427), .A2(n11991), .ZN(n11757) );
  AOI22_X1 U14864 ( .A1(n12569), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20703), .ZN(n11755) );
  INV_X1 U14865 ( .A(n11822), .ZN(n11762) );
  NAND2_X1 U14866 ( .A1(n11762), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11754) );
  AND2_X1 U14867 ( .A1(n11755), .A2(n11754), .ZN(n11756) );
  NAND2_X1 U14868 ( .A1(n11757), .A2(n11756), .ZN(n13264) );
  INV_X1 U14869 ( .A(n11760), .ZN(n11761) );
  XNOR2_X1 U14870 ( .A(n11759), .B(n11761), .ZN(n20861) );
  NAND2_X1 U14871 ( .A1(n20861), .A2(n11991), .ZN(n11766) );
  AOI22_X1 U14872 ( .A1(n12569), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20703), .ZN(n11764) );
  NAND2_X1 U14873 ( .A1(n11762), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11763) );
  AND2_X1 U14874 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  NAND2_X1 U14875 ( .A1(n11766), .A2(n11765), .ZN(n13258) );
  NAND2_X1 U14876 ( .A1(n11768), .A2(n11767), .ZN(n11770) );
  NAND2_X1 U14877 ( .A1(n11770), .A2(n11769), .ZN(n20260) );
  AOI21_X1 U14878 ( .B1(n20260), .B2(n11634), .A(n20703), .ZN(n13257) );
  NAND2_X1 U14879 ( .A1(n13258), .A2(n13257), .ZN(n13256) );
  OR2_X1 U14880 ( .A1(n13258), .A2(n12178), .ZN(n11771) );
  NAND2_X1 U14881 ( .A1(n13256), .A2(n11771), .ZN(n13263) );
  NAND2_X1 U14882 ( .A1(n13264), .A2(n13263), .ZN(n13262) );
  NAND2_X1 U14883 ( .A1(n11773), .A2(n11772), .ZN(n13436) );
  NAND2_X1 U14884 ( .A1(n13436), .A2(n11774), .ZN(n13455) );
  INV_X1 U14885 ( .A(n11794), .ZN(n11793) );
  NAND2_X1 U14886 ( .A1(n11775), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11778) );
  NAND3_X1 U14887 ( .A1(n20856), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20429) );
  INV_X1 U14888 ( .A(n20429), .ZN(n20433) );
  NAND2_X1 U14889 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20433), .ZN(
        n20430) );
  NAND2_X1 U14890 ( .A1(n20856), .A2(n20430), .ZN(n11776) );
  NOR3_X1 U14891 ( .A1(n20856), .A2(n15856), .A3(n20514), .ZN(n20712) );
  NAND2_X1 U14892 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20712), .ZN(
        n20700) );
  AOI22_X1 U14893 ( .A1(n12815), .A2(n20461), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20766), .ZN(n11777) );
  AOI22_X1 U14894 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14895 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14896 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14897 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11781) );
  NAND4_X1 U14898 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11790) );
  AOI22_X1 U14899 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14900 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14901 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14902 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11785) );
  NAND4_X1 U14903 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11789) );
  AOI22_X1 U14904 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12274), .B2(n12633), .ZN(n11791) );
  INV_X1 U14905 ( .A(n20180), .ZN(n20846) );
  NAND2_X1 U14906 ( .A1(n20846), .A2(n11991), .ZN(n11804) );
  INV_X1 U14907 ( .A(n11823), .ZN(n11799) );
  INV_X1 U14908 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11797) );
  NAND2_X1 U14909 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  NAND2_X1 U14910 ( .A1(n11799), .A2(n11798), .ZN(n20072) );
  AOI22_X1 U14911 ( .A1(n20072), .A2(n12566), .B1(n12568), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U14912 ( .A1(n12569), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11800) );
  OAI211_X1 U14913 ( .C1(n11822), .C2(n11795), .A(n11801), .B(n11800), .ZN(
        n11802) );
  INV_X1 U14914 ( .A(n11802), .ZN(n11803) );
  NAND2_X1 U14915 ( .A1(n11804), .A2(n11803), .ZN(n13457) );
  NAND2_X1 U14916 ( .A1(n13455), .A2(n13457), .ZN(n13458) );
  INV_X1 U14917 ( .A(n13458), .ZN(n11827) );
  INV_X1 U14918 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U14919 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14920 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14921 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14922 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12241), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11806) );
  NAND4_X1 U14923 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11815) );
  AOI22_X1 U14924 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12204), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14925 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12100), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14926 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14927 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11810) );
  NAND4_X1 U14928 ( .A1(n11813), .A2(n11812), .A3(n11811), .A4(n11810), .ZN(
        n11814) );
  NAND2_X1 U14929 ( .A1(n12274), .A2(n12645), .ZN(n11816) );
  INV_X1 U14930 ( .A(n11828), .ZN(n11818) );
  XNOR2_X1 U14931 ( .A(n11829), .B(n11818), .ZN(n12632) );
  INV_X1 U14932 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U14933 ( .A1(n20703), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U14934 ( .A1(n12569), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11819) );
  OAI211_X1 U14935 ( .C1(n11822), .C2(n11821), .A(n11820), .B(n11819), .ZN(
        n11824) );
  OAI21_X1 U14936 ( .B1(n11823), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11847), .ZN(n14493) );
  MUX2_X1 U14937 ( .A(n11824), .B(n14493), .S(n11507), .Z(n11825) );
  AOI21_X1 U14938 ( .B1(n12632), .B2(n11991), .A(n11825), .ZN(n13520) );
  INV_X1 U14939 ( .A(n13520), .ZN(n11826) );
  NAND2_X1 U14940 ( .A1(n11827), .A2(n11826), .ZN(n13518) );
  INV_X1 U14941 ( .A(n13518), .ZN(n11853) );
  NOR2_X2 U14942 ( .A1(n11829), .A2(n11828), .ZN(n11843) );
  INV_X1 U14943 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14944 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14945 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14946 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14947 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11831) );
  NAND4_X1 U14948 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11840) );
  AOI22_X1 U14949 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14950 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14951 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14952 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U14953 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11839) );
  NAND2_X1 U14954 ( .A1(n12274), .A2(n12653), .ZN(n11841) );
  INV_X1 U14955 ( .A(n11843), .ZN(n11846) );
  INV_X1 U14956 ( .A(n11844), .ZN(n11845) );
  INV_X1 U14957 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13566) );
  AND2_X1 U14958 ( .A1(n11847), .A2(n20056), .ZN(n11848) );
  OR2_X1 U14959 ( .A1(n11848), .A2(n11867), .ZN(n20058) );
  AOI22_X1 U14960 ( .A1(n20058), .A2(n12566), .B1(n12568), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11849) );
  OAI21_X1 U14961 ( .B1(n12249), .B2(n13566), .A(n11849), .ZN(n11850) );
  NAND2_X1 U14962 ( .A1(n11853), .A2(n13561), .ZN(n13559) );
  INV_X1 U14963 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14964 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14965 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14966 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14967 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11855) );
  NAND4_X1 U14968 ( .A1(n11858), .A2(n11857), .A3(n11856), .A4(n11855), .ZN(
        n11864) );
  AOI22_X1 U14969 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14970 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14971 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14972 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11859) );
  NAND4_X1 U14973 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11863) );
  NAND2_X1 U14974 ( .A1(n12274), .A2(n12661), .ZN(n11865) );
  NAND2_X1 U14975 ( .A1(n11873), .A2(n11872), .ZN(n12651) );
  INV_X1 U14976 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11870) );
  OR2_X1 U14977 ( .A1(n11867), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11868) );
  NAND2_X1 U14978 ( .A1(n11878), .A2(n11868), .ZN(n20041) );
  AOI22_X1 U14979 ( .A1(n20041), .A2(n12566), .B1(n12568), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11869) );
  OAI21_X1 U14980 ( .B1(n12249), .B2(n11870), .A(n11869), .ZN(n11871) );
  NOR2_X1 U14981 ( .A1(n13559), .A2(n13645), .ZN(n13611) );
  INV_X1 U14982 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U14983 ( .A1(n12274), .A2(n12671), .ZN(n11874) );
  OAI21_X1 U14984 ( .B1(n12295), .B2(n11875), .A(n11874), .ZN(n11876) );
  XNOR2_X1 U14985 ( .A(n12600), .B(n11877), .ZN(n12660) );
  NAND2_X1 U14986 ( .A1(n12660), .A2(n11991), .ZN(n11884) );
  INV_X1 U14987 ( .A(n12568), .ZN(n11963) );
  NAND2_X1 U14988 ( .A1(n11878), .A2(n11881), .ZN(n11879) );
  NAND2_X1 U14989 ( .A1(n11895), .A2(n11879), .ZN(n20033) );
  NAND2_X1 U14990 ( .A1(n20033), .A2(n12566), .ZN(n11880) );
  OAI21_X1 U14991 ( .B1(n11881), .B2(n11963), .A(n11880), .ZN(n11882) );
  AOI21_X1 U14992 ( .B1(n12569), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11882), .ZN(
        n11883) );
  NAND2_X1 U14993 ( .A1(n11884), .A2(n11883), .ZN(n13615) );
  NAND2_X1 U14994 ( .A1(n13611), .A2(n13615), .ZN(n13613) );
  INV_X1 U14995 ( .A(n13613), .ZN(n11901) );
  AOI22_X1 U14996 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14997 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U14998 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14999 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U15000 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11894) );
  AOI22_X1 U15001 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U15002 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15003 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U15004 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11889) );
  NAND4_X1 U15005 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11893) );
  OAI21_X1 U15006 ( .B1(n11894), .B2(n11893), .A(n11991), .ZN(n11899) );
  NAND2_X1 U15007 ( .A1(n12569), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11898) );
  XNOR2_X1 U15008 ( .A(n11895), .B(n13739), .ZN(n13858) );
  NAND2_X1 U15009 ( .A1(n13858), .A2(n12566), .ZN(n11897) );
  NAND2_X1 U15010 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11896) );
  XOR2_X1 U15011 ( .A(n11903), .B(n11902), .Z(n14480) );
  INV_X1 U15012 ( .A(n14480), .ZN(n13891) );
  AOI22_X1 U15013 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U15014 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15015 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15016 ( .A1(n12084), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U15017 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11913) );
  AOI22_X1 U15018 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15019 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15020 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15021 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U15022 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11912) );
  OAI21_X1 U15023 ( .B1(n11913), .B2(n11912), .A(n11991), .ZN(n11916) );
  NAND2_X1 U15024 ( .A1(n12569), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U15025 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11914) );
  NAND3_X1 U15026 ( .A1(n11916), .A2(n11915), .A3(n11914), .ZN(n11917) );
  NAND2_X1 U15027 ( .A1(n12569), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11921) );
  OAI21_X1 U15028 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11919), .A(
        n11962), .ZN(n16033) );
  AOI22_X1 U15029 ( .A1(n11507), .A2(n16033), .B1(n12568), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U15030 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  INV_X1 U15031 ( .A(n14613), .ZN(n11935) );
  AOI22_X1 U15032 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15033 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15034 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15035 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U15036 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11932) );
  AOI22_X1 U15037 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11593), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15038 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15039 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15040 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U15041 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  OR2_X1 U15042 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  NAND2_X1 U15043 ( .A1(n11991), .A2(n11933), .ZN(n14617) );
  INV_X1 U15044 ( .A(n14617), .ZN(n11934) );
  NAND2_X1 U15045 ( .A1(n11935), .A2(n11934), .ZN(n14614) );
  AOI22_X1 U15046 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12199), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15047 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12204), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15048 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15049 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11937) );
  NAND4_X1 U15050 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n11946) );
  AOI22_X1 U15051 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15052 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13379), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15053 ( .A1(n12542), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15054 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11941) );
  NAND4_X1 U15055 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n11941), .ZN(
        n11945) );
  NOR2_X1 U15056 ( .A1(n11946), .A2(n11945), .ZN(n11950) );
  XOR2_X1 U15057 ( .A(n15964), .B(n11962), .Z(n16021) );
  INV_X1 U15058 ( .A(n16021), .ZN(n11947) );
  AOI22_X1 U15059 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12566), .B2(n11947), .ZN(n11949) );
  NAND2_X1 U15060 ( .A1(n12569), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11948) );
  OAI211_X1 U15061 ( .C1(n11951), .C2(n11950), .A(n11949), .B(n11948), .ZN(
        n14545) );
  NAND2_X1 U15062 ( .A1(n14543), .A2(n14545), .ZN(n14531) );
  AOI22_X1 U15063 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15064 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15065 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15066 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11952) );
  NAND4_X1 U15067 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11961) );
  AOI22_X1 U15068 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15069 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15070 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15071 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U15072 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  OAI21_X1 U15073 ( .B1(n11961), .B2(n11960), .A(n11991), .ZN(n11967) );
  NAND2_X1 U15074 ( .A1(n12569), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11966) );
  XNOR2_X1 U15075 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11968), .ZN(
        n15958) );
  OAI22_X1 U15076 ( .A1(n15958), .A2(n12178), .B1(n11963), .B2(n15953), .ZN(
        n11964) );
  INV_X1 U15077 ( .A(n11964), .ZN(n11965) );
  NOR2_X2 U15078 ( .A1(n14531), .A2(n14533), .ZN(n14521) );
  XOR2_X1 U15079 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11982), .Z(
        n16012) );
  AOI22_X1 U15080 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15081 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15082 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15083 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U15084 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11978) );
  AOI22_X1 U15085 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15086 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15087 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15088 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15089 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11977) );
  OR2_X1 U15090 ( .A1(n11978), .A2(n11977), .ZN(n11979) );
  AOI22_X1 U15091 ( .A1(n11991), .A2(n11979), .B1(n12568), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U15092 ( .A1(n12569), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11980) );
  OAI211_X1 U15093 ( .C1(n16012), .C2(n12178), .A(n11981), .B(n11980), .ZN(
        n14525) );
  NAND2_X1 U15094 ( .A1(n14521), .A2(n14525), .ZN(n14523) );
  XNOR2_X1 U15095 ( .A(n11998), .B(n15938), .ZN(n15999) );
  AOI22_X1 U15096 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15097 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15098 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15099 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11983) );
  NAND4_X1 U15100 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n11993) );
  AOI22_X1 U15101 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15102 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15103 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15104 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U15105 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11992) );
  OAI21_X1 U15106 ( .B1(n11993), .B2(n11992), .A(n11991), .ZN(n11996) );
  NAND2_X1 U15107 ( .A1(n12569), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U15108 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11994) );
  NAND3_X1 U15109 ( .A1(n11996), .A2(n11995), .A3(n11994), .ZN(n11997) );
  AOI21_X1 U15110 ( .B1(n15999), .B2(n12566), .A(n11997), .ZN(n14600) );
  OAI21_X1 U15111 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11999), .A(
        n12029), .ZN(n15993) );
  INV_X1 U15112 ( .A(n15993), .ZN(n15923) );
  AOI22_X1 U15113 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15114 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15115 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15116 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U15117 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12009) );
  AOI22_X1 U15118 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15119 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15120 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15121 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12004) );
  NAND4_X1 U15122 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(
        n12008) );
  OR2_X1 U15123 ( .A1(n12009), .A2(n12008), .ZN(n12012) );
  INV_X1 U15124 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12010) );
  INV_X1 U15125 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15925) );
  OAI22_X1 U15126 ( .A1(n12249), .A2(n12010), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15925), .ZN(n12011) );
  AOI21_X1 U15127 ( .B1(n12251), .B2(n12012), .A(n12011), .ZN(n12013) );
  MUX2_X1 U15128 ( .A(n15923), .B(n12013), .S(n12178), .Z(n14520) );
  AOI22_X1 U15129 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15130 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15131 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15132 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U15133 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12023) );
  AOI22_X1 U15134 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15135 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15136 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15137 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U15138 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  OR2_X1 U15139 ( .A1(n12023), .A2(n12022), .ZN(n12028) );
  INV_X1 U15140 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12026) );
  INV_X1 U15141 ( .A(n12029), .ZN(n12024) );
  XNOR2_X1 U15142 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12024), .ZN(
        n14470) );
  AOI22_X1 U15143 ( .A1(n12566), .A2(n14470), .B1(n12568), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12025) );
  OAI21_X1 U15144 ( .B1(n12249), .B2(n12026), .A(n12025), .ZN(n12027) );
  AOI21_X1 U15145 ( .B1(n12251), .B2(n12028), .A(n12027), .ZN(n14465) );
  OAI21_X1 U15146 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12030), .A(
        n12060), .ZN(n14722) );
  AOI22_X1 U15147 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15148 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15149 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15150 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U15151 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n12040) );
  AOI22_X1 U15152 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15153 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15154 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15155 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U15156 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12039) );
  NOR2_X1 U15157 ( .A1(n12040), .A2(n12039), .ZN(n12042) );
  AOI22_X1 U15158 ( .A1(n12569), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20703), .ZN(n12041) );
  OAI21_X1 U15159 ( .B1(n12563), .B2(n12042), .A(n12041), .ZN(n12043) );
  MUX2_X1 U15160 ( .A(n14722), .B(n12043), .S(n12178), .Z(n14453) );
  XNOR2_X1 U15161 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12060), .ZN(
        n14716) );
  AOI22_X1 U15162 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15163 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15164 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15165 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U15166 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12053) );
  AOI22_X1 U15167 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15168 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15169 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15170 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12048) );
  NAND4_X1 U15171 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12052) );
  OR2_X1 U15172 ( .A1(n12053), .A2(n12052), .ZN(n12056) );
  INV_X1 U15173 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12054) );
  INV_X1 U15174 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14714) );
  OAI22_X1 U15175 ( .A1(n12249), .A2(n12054), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14714), .ZN(n12055) );
  AOI21_X1 U15176 ( .B1(n12251), .B2(n12056), .A(n12055), .ZN(n12057) );
  MUX2_X1 U15177 ( .A(n14716), .B(n12057), .S(n12178), .Z(n14439) );
  OAI21_X1 U15178 ( .B1(n12062), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12096), .ZN(n14707) );
  INV_X1 U15179 ( .A(n14707), .ZN(n12078) );
  AOI22_X1 U15180 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15181 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12199), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15182 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12204), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15183 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12064) );
  NAND4_X1 U15184 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12073) );
  AOI22_X1 U15185 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15186 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15187 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12084), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15188 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U15189 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12072) );
  OR2_X1 U15190 ( .A1(n12073), .A2(n12072), .ZN(n12076) );
  INV_X1 U15191 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12074) );
  INV_X1 U15192 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14425) );
  OAI22_X1 U15193 ( .A1(n12249), .A2(n12074), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14425), .ZN(n12075) );
  AOI21_X1 U15194 ( .B1(n12251), .B2(n12076), .A(n12075), .ZN(n12077) );
  MUX2_X1 U15195 ( .A(n12078), .B(n12077), .S(n12178), .Z(n14424) );
  AOI22_X1 U15196 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15197 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15198 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15199 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12079) );
  NAND4_X1 U15200 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n12090) );
  AOI22_X1 U15201 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15202 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15203 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15204 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U15205 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12089) );
  NOR2_X1 U15206 ( .A1(n12090), .A2(n12089), .ZN(n12093) );
  AOI21_X1 U15207 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14695), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12091) );
  AOI21_X1 U15208 ( .B1(n12569), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12091), .ZN(
        n12092) );
  OAI21_X1 U15209 ( .B1(n12563), .B2(n12093), .A(n12092), .ZN(n12095) );
  XNOR2_X1 U15210 ( .A(n12096), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14699) );
  NAND2_X1 U15211 ( .A1(n14699), .A2(n12566), .ZN(n12094) );
  INV_X1 U15212 ( .A(n12097), .ZN(n12098) );
  INV_X1 U15213 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U15214 ( .A1(n12098), .A2(n14401), .ZN(n12099) );
  NAND2_X1 U15215 ( .A1(n12140), .A2(n12099), .ZN(n14688) );
  AOI22_X1 U15216 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15217 ( .A1(n12199), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15218 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15219 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15220 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12111) );
  AOI22_X1 U15221 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15222 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15223 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15224 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12106) );
  NAND4_X1 U15225 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  NOR2_X1 U15226 ( .A1(n12111), .A2(n12110), .ZN(n12113) );
  AOI22_X1 U15227 ( .A1(n12569), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20703), .ZN(n12112) );
  OAI21_X1 U15228 ( .B1(n12563), .B2(n12113), .A(n12112), .ZN(n12114) );
  MUX2_X1 U15229 ( .A(n14688), .B(n12114), .S(n12178), .Z(n14394) );
  AOI22_X1 U15230 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15231 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15232 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15233 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12115) );
  NAND4_X1 U15234 ( .A1(n12118), .A2(n12117), .A3(n12116), .A4(n12115), .ZN(
        n12124) );
  AOI22_X1 U15235 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15236 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15237 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15238 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12119) );
  NAND4_X1 U15239 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12123) );
  NOR2_X1 U15240 ( .A1(n12124), .A2(n12123), .ZN(n12155) );
  AOI22_X1 U15241 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15242 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15243 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15244 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12125) );
  NAND4_X1 U15245 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(
        n12135) );
  AOI22_X1 U15246 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15247 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15248 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15249 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12130) );
  NAND4_X1 U15250 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12134) );
  NOR2_X1 U15251 ( .A1(n12135), .A2(n12134), .ZN(n12156) );
  XOR2_X1 U15252 ( .A(n12155), .B(n12156), .Z(n12138) );
  INV_X1 U15253 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12136) );
  INV_X1 U15254 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14677) );
  OAI22_X1 U15255 ( .A1(n12249), .A2(n12136), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14677), .ZN(n12137) );
  AOI21_X1 U15256 ( .B1(n12138), .B2(n12251), .A(n12137), .ZN(n12139) );
  XNOR2_X1 U15257 ( .A(n12140), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14681) );
  MUX2_X1 U15258 ( .A(n12139), .B(n14681), .S(n12566), .Z(n14379) );
  NOR2_X2 U15259 ( .A1(n14377), .A2(n14379), .ZN(n14364) );
  INV_X1 U15260 ( .A(n12142), .ZN(n12143) );
  INV_X1 U15261 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U15262 ( .A1(n12143), .A2(n14667), .ZN(n12144) );
  AND2_X1 U15263 ( .A1(n12193), .A2(n12144), .ZN(n14671) );
  AOI22_X1 U15264 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15265 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15266 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15267 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U15268 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12154) );
  AOI22_X1 U15269 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15270 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15271 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15272 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12149) );
  NAND4_X1 U15273 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12153) );
  NOR2_X1 U15274 ( .A1(n12156), .A2(n12155), .ZN(n12162) );
  XOR2_X1 U15275 ( .A(n12161), .B(n12162), .Z(n12159) );
  INV_X1 U15276 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21019) );
  NOR2_X1 U15277 ( .A1(n21003), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12157) );
  OAI22_X1 U15278 ( .A1(n12249), .A2(n21019), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12157), .ZN(n12158) );
  AOI21_X1 U15279 ( .B1(n12159), .B2(n12251), .A(n12158), .ZN(n12160) );
  NAND2_X1 U15280 ( .A1(n14364), .A2(n14365), .ZN(n14350) );
  INV_X1 U15281 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14354) );
  XNOR2_X1 U15282 ( .A(n12193), .B(n14354), .ZN(n14660) );
  INV_X1 U15283 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U15284 ( .A1(n12162), .A2(n12161), .ZN(n12179) );
  AOI22_X1 U15285 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15286 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15287 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15288 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U15289 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12172) );
  AOI22_X1 U15290 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15291 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15292 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15293 ( .A1(n12204), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U15294 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  NOR2_X1 U15295 ( .A1(n12172), .A2(n12171), .ZN(n12180) );
  XOR2_X1 U15296 ( .A(n12179), .B(n12180), .Z(n12173) );
  NAND2_X1 U15297 ( .A1(n12173), .A2(n12251), .ZN(n12175) );
  OAI21_X1 U15298 ( .B1(n21003), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20703), .ZN(n12174) );
  OAI211_X1 U15299 ( .C1(n12249), .C2(n12176), .A(n12175), .B(n12174), .ZN(
        n12177) );
  OAI21_X1 U15300 ( .B1(n12178), .B2(n14660), .A(n12177), .ZN(n14352) );
  NOR2_X2 U15301 ( .A1(n14350), .A2(n14352), .ZN(n14337) );
  NOR2_X1 U15302 ( .A1(n12180), .A2(n12179), .ZN(n12198) );
  AOI22_X1 U15303 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15304 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15305 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15306 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12181) );
  NAND4_X1 U15307 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12190) );
  AOI22_X1 U15308 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13379), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15309 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15310 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15311 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U15312 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12189) );
  OR2_X1 U15313 ( .A1(n12190), .A2(n12189), .ZN(n12197) );
  XNOR2_X1 U15314 ( .A(n12198), .B(n12197), .ZN(n12192) );
  AOI22_X1 U15315 ( .A1(n12569), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20703), .ZN(n12191) );
  OAI21_X1 U15316 ( .B1(n12192), .B2(n12563), .A(n12191), .ZN(n12196) );
  INV_X1 U15317 ( .A(n12193), .ZN(n12194) );
  OAI21_X1 U15318 ( .B1(n12195), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12229), .ZN(n14651) );
  MUX2_X1 U15319 ( .A(n12196), .B(n14651), .S(n12566), .Z(n14339) );
  NAND2_X1 U15320 ( .A1(n12198), .A2(n12197), .ZN(n12215) );
  AOI22_X1 U15321 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12199), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15322 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15323 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15324 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U15325 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12210) );
  AOI22_X1 U15326 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15327 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15328 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12204), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15329 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15330 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12209) );
  NOR2_X1 U15331 ( .A1(n12210), .A2(n12209), .ZN(n12216) );
  XOR2_X1 U15332 ( .A(n12215), .B(n12216), .Z(n12213) );
  INV_X1 U15333 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12211) );
  OAI22_X1 U15334 ( .A1(n12249), .A2(n12211), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14641), .ZN(n12212) );
  AOI21_X1 U15335 ( .B1(n12213), .B2(n12251), .A(n12212), .ZN(n12214) );
  XNOR2_X1 U15336 ( .A(n12229), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14639) );
  NOR2_X1 U15337 ( .A1(n12216), .A2(n12215), .ZN(n12234) );
  AOI22_X1 U15338 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15339 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15340 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15341 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15342 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12226) );
  AOI22_X1 U15343 ( .A1(n11535), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15344 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15345 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15346 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11598), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12221) );
  NAND4_X1 U15347 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12225) );
  OR2_X1 U15348 ( .A1(n12226), .A2(n12225), .ZN(n12233) );
  XNOR2_X1 U15349 ( .A(n12234), .B(n12233), .ZN(n12228) );
  AOI22_X1 U15350 ( .A1(n12569), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20703), .ZN(n12227) );
  OAI21_X1 U15351 ( .B1(n12228), .B2(n12563), .A(n12227), .ZN(n12232) );
  INV_X1 U15352 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U15353 ( .A1(n12230), .A2(n14320), .ZN(n12231) );
  NAND2_X1 U15354 ( .A1(n12323), .A2(n12231), .ZN(n14631) );
  MUX2_X1 U15355 ( .A(n12232), .B(n14631), .S(n12566), .Z(n14316) );
  NAND2_X1 U15356 ( .A1(n12234), .A2(n12233), .ZN(n12558) );
  AOI22_X1 U15357 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12550), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15358 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12541), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15359 ( .A1(n13379), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15360 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12237) );
  NAND4_X1 U15361 ( .A1(n12240), .A2(n12239), .A3(n12238), .A4(n12237), .ZN(
        n12247) );
  AOI22_X1 U15362 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15363 ( .A1(n12540), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15364 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11598), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15365 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12242) );
  NAND4_X1 U15366 ( .A1(n12245), .A2(n12244), .A3(n12243), .A4(n12242), .ZN(
        n12246) );
  NOR2_X1 U15367 ( .A1(n12247), .A2(n12246), .ZN(n12559) );
  XOR2_X1 U15368 ( .A(n12558), .B(n12559), .Z(n12252) );
  INV_X1 U15369 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12248) );
  INV_X1 U15370 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12819) );
  OAI22_X1 U15371 ( .A1(n12249), .A2(n12248), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12819), .ZN(n12250) );
  AOI21_X1 U15372 ( .B1(n12252), .B2(n12251), .A(n12250), .ZN(n12253) );
  XNOR2_X1 U15373 ( .A(n12323), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12821) );
  INV_X1 U15374 ( .A(n12838), .ZN(n12256) );
  MUX2_X1 U15375 ( .A(n20514), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12271) );
  NAND2_X1 U15376 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20866), .ZN(
        n12275) );
  INV_X1 U15377 ( .A(n12275), .ZN(n12270) );
  NAND2_X1 U15378 ( .A1(n12271), .A2(n12270), .ZN(n12269) );
  NAND2_X1 U15379 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20514), .ZN(
        n12260) );
  NAND2_X1 U15380 ( .A1(n12269), .A2(n12260), .ZN(n12283) );
  NAND2_X1 U15381 ( .A1(n12283), .A2(n12261), .ZN(n12263) );
  NAND2_X1 U15382 ( .A1(n15856), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12262) );
  NOR2_X1 U15383 ( .A1(n11795), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12264) );
  NAND2_X1 U15384 ( .A1(n12265), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12266) );
  NAND2_X1 U15385 ( .A1(n12319), .A2(n12274), .ZN(n12309) );
  XNOR2_X1 U15386 ( .A(n12268), .B(n12267), .ZN(n12315) );
  OAI21_X1 U15387 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12314) );
  NAND2_X1 U15388 ( .A1(n12274), .A2(n11616), .ZN(n12273) );
  NAND2_X1 U15389 ( .A1(n11646), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12272) );
  NAND2_X1 U15390 ( .A1(n12273), .A2(n12272), .ZN(n12285) );
  NOR2_X1 U15391 ( .A1(n12314), .A2(n12285), .ZN(n12281) );
  INV_X1 U15392 ( .A(n12274), .ZN(n12292) );
  OAI21_X1 U15393 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20866), .A(
        n12275), .ZN(n12276) );
  NOR2_X1 U15394 ( .A1(n12292), .A2(n12276), .ZN(n12280) );
  INV_X1 U15395 ( .A(n12276), .ZN(n12278) );
  OR2_X1 U15396 ( .A1(n20213), .A2(n12696), .ZN(n12277) );
  NAND2_X1 U15397 ( .A1(n12277), .A2(n9812), .ZN(n12291) );
  OAI211_X1 U15398 ( .C1(n12696), .C2(n12712), .A(n12278), .B(n12291), .ZN(
        n12279) );
  OAI21_X1 U15399 ( .B1(n12297), .B2(n12280), .A(n12279), .ZN(n12286) );
  NAND2_X1 U15400 ( .A1(n12281), .A2(n12286), .ZN(n12290) );
  MUX2_X1 U15401 ( .A(n15856), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12282) );
  XNOR2_X1 U15402 ( .A(n12283), .B(n12282), .ZN(n12316) );
  NAND2_X1 U15403 ( .A1(n12303), .A2(n12316), .ZN(n12284) );
  OAI211_X1 U15404 ( .C1(n12292), .C2(n12316), .A(n12291), .B(n12284), .ZN(
        n12289) );
  INV_X1 U15405 ( .A(n12285), .ZN(n12287) );
  OAI211_X1 U15406 ( .C1(n12287), .C2(n12286), .A(n12314), .B(n12301), .ZN(
        n12288) );
  NAND3_X1 U15407 ( .A1(n12290), .A2(n12289), .A3(n12288), .ZN(n12294) );
  AOI22_X1 U15408 ( .A1(n12295), .A2(n12315), .B1(n12294), .B2(n12293), .ZN(
        n12296) );
  AOI21_X1 U15409 ( .B1(n12297), .B2(n12315), .A(n12296), .ZN(n12306) );
  INV_X1 U15410 ( .A(n12317), .ZN(n12300) );
  NOR2_X1 U15411 ( .A1(n12303), .A2(n12300), .ZN(n12305) );
  NAND3_X1 U15412 ( .A1(n12303), .A2(n12302), .A3(n12317), .ZN(n12304) );
  OAI21_X1 U15413 ( .B1(n12306), .B2(n12305), .A(n12304), .ZN(n12307) );
  AOI21_X1 U15414 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16196), .A(
        n12307), .ZN(n12308) );
  NAND2_X1 U15415 ( .A1(n12309), .A2(n12308), .ZN(n12310) );
  NOR4_X1 U15416 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12318) );
  OR2_X1 U15417 ( .A1(n12319), .A2(n12318), .ZN(n14311) );
  OR2_X1 U15418 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n16195), .ZN(n12817) );
  NOR2_X1 U15419 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n12817), .ZN(n12320) );
  INV_X1 U15420 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20466) );
  NOR3_X1 U15421 ( .A1(n20466), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15883) );
  MUX2_X1 U15422 ( .A(n12320), .B(n15883), .S(P1_STATE2_REG_0__SCAN_IN), .Z(
        n12321) );
  NOR2_X1 U15423 ( .A1(n20149), .A2(n12321), .ZN(n12322) );
  INV_X1 U15424 ( .A(n12323), .ZN(n12324) );
  NAND2_X1 U15425 ( .A1(n12324), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12565) );
  INV_X1 U15426 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12867) );
  NAND2_X1 U15427 ( .A1(n12892), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12326) );
  INV_X1 U15428 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21235) );
  NAND2_X1 U15429 ( .A1(n12338), .A2(n21235), .ZN(n12330) );
  INV_X1 U15430 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12328) );
  NAND3_X1 U15431 ( .A1(n12330), .A2(n12404), .A3(n12329), .ZN(n12332) );
  NAND2_X1 U15432 ( .A1(n12332), .A2(n12331), .ZN(n12336) );
  INV_X1 U15433 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n20995) );
  NAND2_X1 U15434 ( .A1(n12404), .A2(n20995), .ZN(n12333) );
  NAND2_X1 U15435 ( .A1(n12334), .A2(n12333), .ZN(n13343) );
  XNOR2_X1 U15436 ( .A(n12336), .B(n13343), .ZN(n13780) );
  INV_X1 U15437 ( .A(n13343), .ZN(n12335) );
  NOR2_X1 U15438 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  INV_X1 U15439 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U15440 ( .B1(n12718), .B2(n13356), .A(n12339), .ZN(n13346) );
  AND2_X1 U15441 ( .A1(n13347), .A2(n13346), .ZN(n13471) );
  INV_X1 U15442 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12340) );
  MUX2_X1 U15443 ( .A(n12404), .B(n12403), .S(n12340), .Z(n12343) );
  INV_X1 U15444 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U15445 ( .A1(n12405), .A2(n13469), .ZN(n12342) );
  AND2_X1 U15446 ( .A1(n12343), .A2(n12342), .ZN(n13470) );
  MUX2_X1 U15447 ( .A(n13172), .B(n12413), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12345) );
  INV_X1 U15448 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12639) );
  NOR2_X1 U15449 ( .A1(n12718), .A2(n12639), .ZN(n12344) );
  NOR2_X1 U15450 ( .A1(n12345), .A2(n12344), .ZN(n13511) );
  OR2_X1 U15451 ( .A1(n12403), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12349) );
  INV_X1 U15452 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16179) );
  INV_X1 U15453 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21242) );
  NAND2_X1 U15454 ( .A1(n12718), .A2(n21242), .ZN(n12347) );
  NAND2_X1 U15455 ( .A1(n12349), .A2(n12348), .ZN(n16170) );
  OR2_X1 U15456 ( .A1(n12403), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12352) );
  INV_X1 U15457 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16168) );
  INV_X1 U15458 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21021) );
  NAND2_X1 U15459 ( .A1(n12718), .A2(n21021), .ZN(n12350) );
  AND2_X1 U15460 ( .A1(n12352), .A2(n12351), .ZN(n16159) );
  INV_X1 U15461 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13841) );
  OR2_X1 U15462 ( .A1(n12718), .A2(n13841), .ZN(n12353) );
  NAND2_X1 U15463 ( .A1(n12354), .A2(n12353), .ZN(n16160) );
  NAND2_X1 U15464 ( .A1(n16159), .A2(n16160), .ZN(n12355) );
  INV_X1 U15465 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13835) );
  OAI21_X1 U15466 ( .B1(n12718), .B2(n13835), .A(n12356), .ZN(n13736) );
  NAND2_X1 U15467 ( .A1(n16162), .A2(n13736), .ZN(n13883) );
  OR2_X1 U15468 ( .A1(n12403), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n12359) );
  INV_X1 U15469 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16157) );
  INV_X1 U15470 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21227) );
  NAND2_X1 U15471 ( .A1(n12718), .A2(n21227), .ZN(n12357) );
  NAND2_X1 U15472 ( .A1(n12359), .A2(n12358), .ZN(n13882) );
  INV_X1 U15473 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n20979) );
  NAND2_X1 U15474 ( .A1(n12718), .A2(n20979), .ZN(n12360) );
  OAI211_X1 U15475 ( .C1(n12413), .C2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12360), .B(n12404), .ZN(n12362) );
  NAND2_X1 U15476 ( .A1(n13172), .A2(n20979), .ZN(n12361) );
  AND2_X1 U15477 ( .A1(n12362), .A2(n12361), .ZN(n13917) );
  OR2_X1 U15478 ( .A1(n12403), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n12365) );
  INV_X1 U15479 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12742) );
  INV_X1 U15480 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21230) );
  NAND2_X1 U15481 ( .A1(n12718), .A2(n21230), .ZN(n12363) );
  NAND2_X1 U15482 ( .A1(n12365), .A2(n12364), .ZN(n15971) );
  OAI21_X1 U15483 ( .B1(n12718), .B2(n16126), .A(n12366), .ZN(n14540) );
  NAND2_X1 U15484 ( .A1(n15974), .A2(n14540), .ZN(n14542) );
  INV_X1 U15485 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n12367) );
  MUX2_X1 U15486 ( .A(n12404), .B(n12403), .S(n12367), .Z(n12369) );
  INV_X1 U15487 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14821) );
  NAND2_X1 U15488 ( .A1(n12405), .A2(n14821), .ZN(n12368) );
  NAND2_X1 U15489 ( .A1(n12369), .A2(n12368), .ZN(n14536) );
  INV_X1 U15490 ( .A(n12370), .ZN(n14535) );
  INV_X1 U15491 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U15492 ( .A1(n12718), .A2(n14530), .ZN(n12371) );
  OAI211_X1 U15493 ( .C1(n9816), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12371), .B(n12404), .ZN(n12373) );
  NAND2_X1 U15494 ( .A1(n13172), .A2(n14530), .ZN(n12372) );
  NOR2_X2 U15495 ( .A1(n14535), .A2(n14526), .ZN(n15935) );
  INV_X1 U15496 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n12374) );
  MUX2_X1 U15497 ( .A(n12404), .B(n12403), .S(n12374), .Z(n12376) );
  INV_X1 U15498 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U15499 ( .A1(n12405), .A2(n16098), .ZN(n12375) );
  MUX2_X1 U15500 ( .A(n13172), .B(n9816), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12379) );
  INV_X1 U15501 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12377) );
  NOR2_X1 U15502 ( .A1(n12718), .A2(n12377), .ZN(n12378) );
  NOR2_X1 U15503 ( .A1(n12379), .A2(n12378), .ZN(n14514) );
  INV_X1 U15504 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n12380) );
  MUX2_X1 U15505 ( .A(n12404), .B(n12403), .S(n12380), .Z(n12382) );
  NAND2_X1 U15506 ( .A1(n12405), .A2(n12679), .ZN(n12381) );
  NAND2_X1 U15507 ( .A1(n12382), .A2(n12381), .ZN(n14467) );
  INV_X1 U15508 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21043) );
  NAND2_X1 U15509 ( .A1(n12718), .A2(n21043), .ZN(n12384) );
  INV_X1 U15510 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14825) );
  NAND3_X1 U15511 ( .A1(n12384), .A2(n12404), .A3(n12383), .ZN(n12386) );
  NAND2_X1 U15512 ( .A1(n13172), .A2(n21043), .ZN(n12385) );
  NAND2_X1 U15513 ( .A1(n12386), .A2(n12385), .ZN(n14455) );
  INV_X1 U15514 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n12387) );
  MUX2_X1 U15515 ( .A(n12404), .B(n12403), .S(n12387), .Z(n12389) );
  INV_X1 U15516 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U15517 ( .A1(n12405), .A2(n14801), .ZN(n12388) );
  MUX2_X1 U15518 ( .A(n13172), .B(n9816), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12391) );
  INV_X1 U15519 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14815) );
  NOR2_X1 U15520 ( .A1(n12718), .A2(n14815), .ZN(n12390) );
  NOR2_X1 U15521 ( .A1(n12391), .A2(n12390), .ZN(n14426) );
  MUX2_X1 U15522 ( .A(n12403), .B(n12404), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12393) );
  INV_X1 U15523 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15889) );
  NAND2_X1 U15524 ( .A1(n12405), .A2(n15889), .ZN(n12392) );
  NAND2_X1 U15525 ( .A1(n12393), .A2(n12392), .ZN(n14414) );
  INV_X1 U15526 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14804) );
  OAI21_X1 U15527 ( .B1(n12718), .B2(n14804), .A(n12394), .ZN(n14395) );
  OR2_X1 U15528 ( .A1(n12403), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12397) );
  INV_X1 U15529 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14673) );
  INV_X1 U15530 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21214) );
  NAND2_X1 U15531 ( .A1(n12718), .A2(n21214), .ZN(n12395) );
  MUX2_X1 U15532 ( .A(n13172), .B(n12413), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12399) );
  INV_X1 U15533 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14794) );
  NOR2_X1 U15534 ( .A1(n12718), .A2(n14794), .ZN(n12398) );
  NOR2_X1 U15535 ( .A1(n12399), .A2(n12398), .ZN(n14370) );
  OR2_X1 U15536 ( .A1(n12403), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n12402) );
  INV_X1 U15537 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16049) );
  INV_X1 U15538 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21211) );
  NAND2_X1 U15539 ( .A1(n12718), .A2(n21211), .ZN(n12400) );
  NAND2_X1 U15540 ( .A1(n12402), .A2(n12401), .ZN(n14358) );
  INV_X1 U15541 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14331) );
  MUX2_X1 U15542 ( .A(n12404), .B(n12403), .S(n14331), .Z(n12407) );
  INV_X1 U15543 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14783) );
  NAND2_X1 U15544 ( .A1(n12405), .A2(n14783), .ZN(n12406) );
  AND2_X1 U15545 ( .A1(n12407), .A2(n12406), .ZN(n12449) );
  INV_X1 U15546 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12408) );
  OR2_X1 U15547 ( .A1(n12718), .A2(n12408), .ZN(n12409) );
  NAND2_X1 U15548 ( .A1(n12410), .A2(n12409), .ZN(n14344) );
  NAND2_X1 U15549 ( .A1(n12449), .A2(n14344), .ZN(n12411) );
  INV_X1 U15550 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U15551 ( .A1(n12718), .A2(n14506), .ZN(n12412) );
  OAI211_X1 U15552 ( .C1(n12413), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12412), .B(n12404), .ZN(n12415) );
  NAND2_X1 U15553 ( .A1(n13172), .A2(n14506), .ZN(n12414) );
  NAND2_X1 U15554 ( .A1(n12415), .A2(n12414), .ZN(n14318) );
  INV_X1 U15555 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n21165) );
  NAND2_X1 U15556 ( .A1(n12718), .A2(n21165), .ZN(n12416) );
  OAI21_X1 U15557 ( .B1(n12341), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12416), .ZN(n12864) );
  MUX2_X1 U15558 ( .A(n12864), .B(P1_EBX_REG_29__SCAN_IN), .S(n13172), .Z(
        n12417) );
  NAND2_X1 U15559 ( .A1(n14317), .A2(n12417), .ZN(n12418) );
  NAND2_X1 U15560 ( .A1(n12863), .A2(n12418), .ZN(n14762) );
  AND2_X1 U15561 ( .A1(n20880), .A2(n21003), .ZN(n15878) );
  INV_X1 U15562 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n21167) );
  NOR2_X1 U15563 ( .A1(n15878), .A2(n21167), .ZN(n12419) );
  AND2_X1 U15564 ( .A1(n12718), .A2(n12419), .ZN(n12420) );
  INV_X1 U15565 ( .A(n12421), .ZN(n12422) );
  NAND2_X1 U15566 ( .A1(n12422), .A2(n20776), .ZN(n20879) );
  NAND2_X1 U15567 ( .A1(n9812), .A2(n20879), .ZN(n12707) );
  NAND2_X1 U15568 ( .A1(n12707), .A2(n15878), .ZN(n12428) );
  NOR2_X1 U15569 ( .A1(n12428), .A2(n12696), .ZN(n12423) );
  INV_X1 U15570 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21181) );
  INV_X1 U15571 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20951) );
  NAND4_X1 U15572 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20053)
         );
  NOR2_X1 U15573 ( .A1(n20951), .A2(n20053), .ZN(n20049) );
  NAND2_X1 U15574 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20049), .ZN(n20031) );
  NOR2_X1 U15575 ( .A1(n21181), .A2(n20031), .ZN(n13735) );
  NAND2_X1 U15576 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13735), .ZN(n13734) );
  INV_X1 U15577 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15960) );
  INV_X1 U15578 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21232) );
  INV_X1 U15579 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n16122) );
  INV_X1 U15580 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15984) );
  NOR4_X1 U15581 ( .A1(n15960), .A2(n21232), .A3(n16122), .A4(n15984), .ZN(
        n15929) );
  NAND4_X1 U15582 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15929), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n14444) );
  INV_X1 U15583 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21007) );
  INV_X1 U15584 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21251) );
  NOR2_X1 U15585 ( .A1(n21007), .A2(n21251), .ZN(n14421) );
  NAND4_X1 U15586 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .A4(n14421), .ZN(n12425) );
  NOR3_X1 U15587 ( .A1(n13734), .A2(n14444), .A3(n12425), .ZN(n14413) );
  INV_X1 U15588 ( .A(n14413), .ZN(n14403) );
  NOR2_X1 U15589 ( .A1(n20032), .A2(n14403), .ZN(n14381) );
  NAND2_X1 U15590 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14382) );
  INV_X1 U15591 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14676) );
  NOR2_X1 U15592 ( .A1(n14382), .A2(n14676), .ZN(n12427) );
  NAND2_X1 U15593 ( .A1(n14381), .A2(n12427), .ZN(n14369) );
  NAND3_X1 U15594 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .ZN(n14321) );
  NAND2_X1 U15595 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12426) );
  INV_X1 U15596 ( .A(n12868), .ZN(n12435) );
  INV_X1 U15597 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21187) );
  INV_X1 U15598 ( .A(n20030), .ZN(n13814) );
  NOR2_X1 U15599 ( .A1(n20030), .A2(n14403), .ZN(n14399) );
  NAND2_X1 U15600 ( .A1(n14399), .A2(n12427), .ZN(n14353) );
  NOR2_X1 U15601 ( .A1(n14353), .A2(n14321), .ZN(n14329) );
  NAND3_X1 U15602 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n14329), .ZN(n12869) );
  NAND2_X1 U15603 ( .A1(n20029), .A2(n12869), .ZN(n14325) );
  OAI211_X1 U15604 ( .C1(n9812), .C2(n21167), .A(n12428), .B(n11627), .ZN(
        n12429) );
  INV_X2 U15605 ( .A(n14471), .ZN(n20043) );
  OR2_X1 U15606 ( .A1(n12892), .A2(n16195), .ZN(n12430) );
  INV_X1 U15607 ( .A(n12821), .ZN(n12431) );
  OAI22_X1 U15608 ( .A1(n12819), .A2(n20057), .B1(n20059), .B2(n12431), .ZN(
        n12432) );
  AOI21_X1 U15609 ( .B1(n20043), .B2(P1_EBX_REG_29__SCAN_IN), .A(n12432), .ZN(
        n12433) );
  OAI21_X1 U15610 ( .B1(n14325), .B2(n21187), .A(n12433), .ZN(n12434) );
  AOI21_X1 U15611 ( .B1(n12435), .B2(n21187), .A(n12434), .ZN(n12436) );
  INV_X1 U15612 ( .A(n14846), .ZN(n12579) );
  NOR2_X1 U15613 ( .A1(n11609), .A2(n20213), .ZN(n12446) );
  NAND4_X1 U15614 ( .A1(n12727), .A2(n14044), .A3(n12446), .A4(n11540), .ZN(
        n12573) );
  OR2_X1 U15615 ( .A1(n12717), .A2(n12573), .ZN(n12447) );
  INV_X1 U15616 ( .A(n14360), .ZN(n14345) );
  AOI21_X1 U15617 ( .B1(n14345), .B2(n14344), .A(n12449), .ZN(n12450) );
  OR2_X1 U15618 ( .A1(n12450), .A2(n14319), .ZN(n14780) );
  OAI22_X1 U15619 ( .A1(n14780), .A2(n14546), .B1(n14331), .B2(n20092), .ZN(
        n12451) );
  OR2_X1 U15620 ( .A1(n12455), .A2(n9869), .ZN(n12456) );
  NAND2_X1 U15621 ( .A1(n12858), .A2(n19291), .ZN(n12463) );
  XNOR2_X2 U15622 ( .A(n14923), .B(n12457), .ZN(n14292) );
  NOR2_X1 U15623 ( .A1(n14292), .A2(n15258), .ZN(n12460) );
  XNOR2_X1 U15624 ( .A(n12485), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12525) );
  NAND2_X1 U15625 ( .A1(n19286), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12852) );
  NAND2_X1 U15626 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12458) );
  OAI211_X1 U15627 ( .C1(n19296), .C2(n12525), .A(n12852), .B(n12458), .ZN(
        n12459) );
  NOR2_X1 U15628 ( .A1(n12460), .A2(n12459), .ZN(n12462) );
  XNOR2_X1 U15629 ( .A(n15121), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12859) );
  NAND3_X1 U15630 ( .A1(n12463), .A2(n12462), .A3(n12461), .ZN(P2_U2984) );
  NAND2_X1 U15631 ( .A1(n11327), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15632 ( .A1(n12478), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12464) );
  AND2_X1 U15633 ( .A1(n12465), .A2(n12464), .ZN(n15065) );
  NAND2_X1 U15634 ( .A1(n11327), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15635 ( .A1(n12478), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12466) );
  AND2_X1 U15636 ( .A1(n12467), .A2(n12466), .ZN(n15054) );
  NAND2_X1 U15637 ( .A1(n11327), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15638 ( .A1(n12478), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12468) );
  INV_X1 U15639 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19936) );
  AOI22_X1 U15640 ( .A1(n12478), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12470) );
  OAI21_X1 U15641 ( .B1(n11305), .B2(n19936), .A(n12470), .ZN(n15047) );
  NAND2_X1 U15642 ( .A1(n15309), .A2(n15047), .ZN(n15039) );
  NAND2_X1 U15643 ( .A1(n12477), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15644 ( .A1(n12478), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12471) );
  AND2_X1 U15645 ( .A1(n12472), .A2(n12471), .ZN(n15038) );
  NAND2_X1 U15646 ( .A1(n11327), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15647 ( .A1(n12478), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12473) );
  NOR2_X4 U15648 ( .A1(n9845), .A2(n15029), .ZN(n15031) );
  INV_X1 U15649 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19942) );
  AOI22_X1 U15650 ( .A1(n12478), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12475) );
  OAI21_X1 U15651 ( .B1(n11305), .B2(n19942), .A(n12475), .ZN(n12777) );
  INV_X1 U15652 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19944) );
  AOI22_X1 U15653 ( .A1(n12478), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12476) );
  OAI21_X1 U15654 ( .B1(n11305), .B2(n19944), .A(n12476), .ZN(n15014) );
  NAND2_X1 U15655 ( .A1(n12477), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15656 ( .A1(n12478), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11291), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12479) );
  AND2_X1 U15657 ( .A1(n12480), .A2(n12479), .ZN(n12481) );
  AND2_X1 U15658 ( .A1(n12482), .A2(n12481), .ZN(n12483) );
  OR2_X2 U15659 ( .A1(n12827), .A2(n12483), .ZN(n14289) );
  INV_X1 U15660 ( .A(n19866), .ZN(n13144) );
  INV_X1 U15661 ( .A(n12484), .ZN(n14854) );
  NAND2_X1 U15662 ( .A1(n19633), .A2(n13042), .ZN(n16450) );
  INV_X1 U15663 ( .A(n12490), .ZN(n12486) );
  AOI21_X1 U15664 ( .B1(n10218), .B2(n12486), .A(n12485), .ZN(n15128) );
  INV_X1 U15665 ( .A(n15128), .ZN(n16215) );
  AND2_X1 U15666 ( .A1(n10891), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12487) );
  NOR2_X1 U15667 ( .A1(n12523), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12489) );
  OR2_X1 U15668 ( .A1(n12490), .A2(n12489), .ZN(n16228) );
  NAND2_X1 U15669 ( .A1(n12521), .A2(n12491), .ZN(n12492) );
  NAND2_X1 U15670 ( .A1(n9908), .A2(n12492), .ZN(n16248) );
  OR2_X1 U15671 ( .A1(n12495), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12494) );
  NAND2_X1 U15672 ( .A1(n12493), .A2(n12494), .ZN(n16272) );
  AOI21_X1 U15673 ( .B1(n15175), .B2(n12519), .A(n12495), .ZN(n15173) );
  INV_X1 U15674 ( .A(n15173), .ZN(n16281) );
  OAI21_X1 U15675 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12515), .A(
        n12517), .ZN(n19075) );
  AND2_X1 U15676 ( .A1(n12511), .A2(n12496), .ZN(n12497) );
  OR2_X1 U15677 ( .A1(n12497), .A2(n12513), .ZN(n15238) );
  AOI21_X1 U15678 ( .B1(n15257), .B2(n12509), .A(n12512), .ZN(n14896) );
  AOI21_X1 U15679 ( .B1(n16311), .B2(n12508), .A(n12510), .ZN(n16304) );
  AOI21_X1 U15680 ( .B1(n19126), .B2(n12506), .A(n9886), .ZN(n19136) );
  AOI21_X1 U15681 ( .B1(n16335), .B2(n12504), .A(n12507), .ZN(n16328) );
  AOI21_X1 U15682 ( .B1(n13984), .B2(n12502), .A(n12505), .ZN(n19153) );
  AOI21_X1 U15683 ( .B1(n16364), .B2(n12500), .A(n12503), .ZN(n16354) );
  AOI21_X1 U15684 ( .B1(n14033), .B2(n12499), .A(n12501), .ZN(n14035) );
  INV_X1 U15685 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19209) );
  AOI22_X1 U15686 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12498), .B1(n19209), 
        .B2(n19863), .ZN(n19196) );
  INV_X1 U15687 ( .A(n19196), .ZN(n15510) );
  INV_X1 U15688 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19180) );
  OAI22_X1 U15689 ( .A1(n19863), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19180), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15509) );
  AND2_X1 U15690 ( .A1(n15510), .A2(n15509), .ZN(n14912) );
  OAI21_X1 U15691 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12499), .ZN(n14914) );
  NAND2_X1 U15692 ( .A1(n14912), .A2(n14914), .ZN(n13711) );
  NOR2_X1 U15693 ( .A1(n14035), .A2(n13711), .ZN(n19164) );
  OAI21_X1 U15694 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12501), .A(
        n12500), .ZN(n19295) );
  NAND2_X1 U15695 ( .A1(n19164), .A2(n19295), .ZN(n13791) );
  NOR2_X1 U15696 ( .A1(n16354), .A2(n13791), .ZN(n13681) );
  OAI21_X1 U15697 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12503), .A(
        n12502), .ZN(n16353) );
  NAND2_X1 U15698 ( .A1(n13681), .A2(n16353), .ZN(n19151) );
  NOR2_X1 U15699 ( .A1(n19153), .A2(n19151), .ZN(n19144) );
  OAI21_X1 U15700 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12505), .A(
        n12504), .ZN(n19145) );
  NAND2_X1 U15701 ( .A1(n19144), .A2(n19145), .ZN(n13701) );
  NOR2_X1 U15702 ( .A1(n16328), .A2(n13701), .ZN(n13691) );
  OAI21_X1 U15703 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12507), .A(
        n12506), .ZN(n16327) );
  NAND2_X1 U15704 ( .A1(n13691), .A2(n16327), .ZN(n19132) );
  NOR2_X1 U15705 ( .A1(n19136), .A2(n19132), .ZN(n19115) );
  OAI21_X1 U15706 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9886), .A(
        n12508), .ZN(n19116) );
  NAND2_X1 U15707 ( .A1(n19115), .A2(n19116), .ZN(n13847) );
  NOR2_X1 U15708 ( .A1(n16304), .A2(n13847), .ZN(n19105) );
  OAI21_X1 U15709 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12510), .A(
        n12509), .ZN(n19106) );
  NAND2_X1 U15710 ( .A1(n19105), .A2(n19106), .ZN(n14897) );
  NOR2_X1 U15711 ( .A1(n14896), .A2(n14897), .ZN(n19090) );
  OAI21_X1 U15712 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12512), .A(
        n12511), .ZN(n19091) );
  AND2_X1 U15713 ( .A1(n19090), .A2(n19091), .ZN(n14888) );
  AND2_X1 U15714 ( .A1(n15238), .A2(n14888), .ZN(n14887) );
  OR2_X1 U15715 ( .A1(n12513), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12514) );
  NAND2_X1 U15716 ( .A1(n12516), .A2(n12514), .ZN(n19079) );
  NAND2_X1 U15717 ( .A1(n14887), .A2(n19079), .ZN(n14877) );
  AOI21_X1 U15718 ( .B1(n15219), .B2(n12516), .A(n12515), .ZN(n15221) );
  NAND2_X1 U15719 ( .A1(n19075), .A2(n19074), .ZN(n19073) );
  NAND2_X1 U15720 ( .A1(n19152), .A2(n19073), .ZN(n14868) );
  NAND2_X1 U15721 ( .A1(n11084), .A2(n12517), .ZN(n12518) );
  NAND2_X1 U15722 ( .A1(n10215), .A2(n12518), .ZN(n15195) );
  OAI21_X1 U15723 ( .B1(n12520), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12519), .ZN(n15844) );
  NAND2_X1 U15724 ( .A1(n19152), .A2(n15843), .ZN(n16280) );
  INV_X1 U15725 ( .A(n12521), .ZN(n12522) );
  AOI21_X1 U15726 ( .B1(n15156), .B2(n12493), .A(n12522), .ZN(n15159) );
  INV_X1 U15727 ( .A(n15159), .ZN(n16260) );
  NAND2_X1 U15728 ( .A1(n19152), .A2(n16258), .ZN(n16247) );
  NAND2_X1 U15729 ( .A1(n16248), .A2(n16247), .ZN(n16246) );
  AOI21_X1 U15730 ( .B1(n15135), .B2(n9908), .A(n12523), .ZN(n15133) );
  INV_X1 U15731 ( .A(n15133), .ZN(n16237) );
  NAND2_X1 U15732 ( .A1(n19152), .A2(n16235), .ZN(n16227) );
  NAND2_X1 U15733 ( .A1(n16228), .A2(n16227), .ZN(n16226) );
  NAND2_X1 U15734 ( .A1(n19152), .A2(n16226), .ZN(n16214) );
  NAND2_X1 U15735 ( .A1(n16215), .A2(n16214), .ZN(n16213) );
  NAND2_X1 U15736 ( .A1(n16213), .A2(n19152), .ZN(n12524) );
  NAND3_X1 U15737 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15909), .A3(n19633), 
        .ZN(n19869) );
  OAI211_X1 U15738 ( .C1(n12525), .C2(n12524), .A(n19108), .B(n16208), .ZN(
        n12539) );
  INV_X1 U15739 ( .A(n12526), .ZN(n12527) );
  NAND2_X1 U15740 ( .A1(n13038), .A2(n12527), .ZN(n13040) );
  OR2_X1 U15741 ( .A1(n13040), .A2(n19872), .ZN(n13046) );
  NOR2_X1 U15742 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19872), .ZN(n12530) );
  OR3_X1 U15743 ( .A1(n13040), .A2(n14227), .A3(n12530), .ZN(n16201) );
  INV_X1 U15744 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14920) );
  INV_X1 U15745 ( .A(n16451), .ZN(n12528) );
  INV_X1 U15746 ( .A(n16450), .ZN(n12529) );
  OR2_X1 U15747 ( .A1(n13148), .A2(n12529), .ZN(n16200) );
  OR3_X1 U15748 ( .A1(n13040), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12530), .ZN(
        n12531) );
  INV_X1 U15749 ( .A(n19183), .ZN(n19202) );
  NOR2_X1 U15750 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19863), .ZN(n19862) );
  NAND3_X1 U15751 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19862), .A3(n15506), 
        .ZN(n16466) );
  AND3_X1 U15752 ( .A1(n16466), .A2(n19869), .A3(n19170), .ZN(n12532) );
  AOI22_X1 U15753 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19197), .ZN(n12533) );
  OAI21_X1 U15754 ( .B1(n11186), .B2(n19202), .A(n12533), .ZN(n12534) );
  AOI21_X1 U15755 ( .B1(n12535), .B2(n19205), .A(n12534), .ZN(n12536) );
  INV_X1 U15756 ( .A(n12537), .ZN(n12538) );
  NAND3_X1 U15757 ( .A1(n9861), .A2(n12539), .A3(n12538), .ZN(P2_U2825) );
  AOI22_X1 U15758 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12540), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15759 ( .A1(n12541), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15760 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15761 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12544) );
  NAND4_X1 U15762 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n12557) );
  AOI22_X1 U15763 ( .A1(n12083), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12199), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15764 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15765 ( .A1(n12550), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12084), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15766 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12551), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12552) );
  NAND4_X1 U15767 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12556) );
  NOR2_X1 U15768 ( .A1(n12557), .A2(n12556), .ZN(n12561) );
  NOR2_X1 U15769 ( .A1(n12559), .A2(n12558), .ZN(n12560) );
  XOR2_X1 U15770 ( .A(n12561), .B(n12560), .Z(n12564) );
  AOI22_X1 U15771 ( .A1(n12569), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20703), .ZN(n12562) );
  OAI21_X1 U15772 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n12567) );
  XNOR2_X1 U15773 ( .A(n12565), .B(n12867), .ZN(n12866) );
  MUX2_X1 U15774 ( .A(n12567), .B(n12866), .S(n12566), .Z(n12839) );
  AOI22_X1 U15775 ( .A1(n12569), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12568), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12570) );
  INV_X1 U15776 ( .A(n12570), .ZN(n12571) );
  XNOR2_X2 U15777 ( .A(n12841), .B(n12571), .ZN(n12888) );
  INV_X1 U15778 ( .A(n12572), .ZN(n16187) );
  INV_X1 U15779 ( .A(n20880), .ZN(n20876) );
  NOR2_X1 U15780 ( .A1(n20876), .A2(n14311), .ZN(n12701) );
  NAND2_X1 U15781 ( .A1(n16187), .A2(n12701), .ZN(n13325) );
  OR2_X1 U15782 ( .A1(n12573), .A2(n13777), .ZN(n12574) );
  OR2_X1 U15783 ( .A1(n12575), .A2(n11620), .ZN(n12698) );
  NAND2_X1 U15784 ( .A1(n11612), .A2(n20880), .ZN(n12577) );
  NAND2_X1 U15785 ( .A1(n13327), .A2(n12718), .ZN(n12580) );
  NOR2_X1 U15786 ( .A1(n13777), .A2(n11620), .ZN(n12578) );
  NAND2_X1 U15787 ( .A1(n12579), .A2(n12578), .ZN(n13386) );
  NAND2_X1 U15788 ( .A1(n12580), .A2(n13386), .ZN(n13330) );
  NAND2_X1 U15789 ( .A1(n12888), .A2(n10449), .ZN(n12599) );
  NOR4_X1 U15790 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12586) );
  NOR4_X1 U15791 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12585) );
  NOR4_X1 U15792 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12584) );
  NOR4_X1 U15793 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12583) );
  AND4_X1 U15794 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        n12591) );
  NOR4_X1 U15795 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12589) );
  NOR4_X1 U15796 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12588) );
  NOR4_X1 U15797 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12587) );
  INV_X1 U15798 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20785) );
  AND4_X1 U15799 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n20785), .ZN(
        n12590) );
  NAND2_X1 U15800 ( .A1(n12591), .A2(n12590), .ZN(n12592) );
  NOR3_X1 U15801 ( .A1(n14618), .A2(n20177), .A3(n11647), .ZN(n12593) );
  AOI22_X1 U15802 ( .A1(n14593), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14618), .ZN(n12594) );
  INV_X1 U15803 ( .A(n12594), .ZN(n12597) );
  INV_X1 U15804 ( .A(n20177), .ZN(n20179) );
  NOR2_X1 U15805 ( .A1(n11647), .A2(n20179), .ZN(n12595) );
  NAND2_X1 U15806 ( .A1(n14602), .A2(n12595), .ZN(n14565) );
  INV_X1 U15807 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16548) );
  NOR2_X1 U15808 ( .A1(n14565), .A2(n16548), .ZN(n12596) );
  NOR2_X1 U15809 ( .A1(n12597), .A2(n12596), .ZN(n12598) );
  NAND2_X1 U15810 ( .A1(n12599), .A2(n12598), .ZN(P1_U2873) );
  INV_X1 U15811 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12843) );
  AND2_X1 U15812 ( .A1(n12601), .A2(n12695), .ZN(n12602) );
  NOR2_X1 U15813 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12678) );
  INV_X1 U15814 ( .A(n12695), .ZN(n12618) );
  NAND2_X1 U15815 ( .A1(n12610), .A2(n12606), .ZN(n12620) );
  AND2_X1 U15816 ( .A1(n12620), .A2(n12619), .ZN(n12634) );
  XNOR2_X1 U15817 ( .A(n12634), .B(n12633), .ZN(n12603) );
  NAND2_X1 U15818 ( .A1(n12603), .A2(n12666), .ZN(n12604) );
  XNOR2_X1 U15819 ( .A(n12610), .B(n12606), .ZN(n12607) );
  OAI211_X1 U15820 ( .C1(n12607), .C2(n13541), .A(n11613), .B(n20213), .ZN(
        n12608) );
  INV_X1 U15821 ( .A(n12608), .ZN(n12609) );
  OR2_X1 U15822 ( .A1(n20260), .A2(n12618), .ZN(n12613) );
  NAND2_X1 U15823 ( .A1(n12696), .A2(n20204), .ZN(n12622) );
  OAI21_X1 U15824 ( .B1(n13541), .B2(n12610), .A(n12622), .ZN(n12611) );
  INV_X1 U15825 ( .A(n12611), .ZN(n12612) );
  NAND2_X1 U15826 ( .A1(n12613), .A2(n12612), .ZN(n20147) );
  NAND2_X1 U15827 ( .A1(n20147), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20146) );
  XNOR2_X1 U15828 ( .A(n12615), .B(n20146), .ZN(n20139) );
  NAND2_X1 U15829 ( .A1(n20139), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20138) );
  INV_X1 U15830 ( .A(n20146), .ZN(n12614) );
  NAND2_X1 U15831 ( .A1(n12615), .A2(n12614), .ZN(n12616) );
  NAND2_X1 U15832 ( .A1(n20138), .A2(n12616), .ZN(n12627) );
  XNOR2_X1 U15833 ( .A(n12627), .B(n13356), .ZN(n13345) );
  OR2_X1 U15834 ( .A1(n20456), .A2(n12618), .ZN(n12626) );
  NOR2_X1 U15835 ( .A1(n12620), .A2(n12619), .ZN(n12621) );
  OR2_X1 U15836 ( .A1(n12634), .A2(n12621), .ZN(n12624) );
  INV_X1 U15837 ( .A(n12622), .ZN(n12623) );
  AOI21_X1 U15838 ( .B1(n12624), .B2(n12666), .A(n12623), .ZN(n12625) );
  NAND2_X1 U15839 ( .A1(n13345), .A2(n13344), .ZN(n12629) );
  NAND2_X1 U15840 ( .A1(n12627), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12628) );
  NAND2_X1 U15841 ( .A1(n12630), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12631) );
  INV_X1 U15842 ( .A(n12633), .ZN(n12635) );
  NOR2_X1 U15843 ( .A1(n12635), .A2(n12634), .ZN(n12644) );
  INV_X1 U15844 ( .A(n12644), .ZN(n12636) );
  XNOR2_X1 U15845 ( .A(n12645), .B(n12636), .ZN(n12637) );
  NAND2_X1 U15846 ( .A1(n12666), .A2(n12637), .ZN(n12638) );
  NAND2_X1 U15847 ( .A1(n12640), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12641) );
  AND2_X1 U15848 ( .A1(n12645), .A2(n12644), .ZN(n12654) );
  INV_X1 U15849 ( .A(n12654), .ZN(n12646) );
  XNOR2_X1 U15850 ( .A(n12653), .B(n12646), .ZN(n12647) );
  NAND2_X1 U15851 ( .A1(n12666), .A2(n12647), .ZN(n12648) );
  XNOR2_X1 U15852 ( .A(n12649), .B(n16179), .ZN(n16041) );
  NAND2_X1 U15853 ( .A1(n12649), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12650) );
  NAND3_X1 U15854 ( .A1(n12652), .A2(n12651), .A3(n12695), .ZN(n12657) );
  NAND2_X1 U15855 ( .A1(n12654), .A2(n12653), .ZN(n12662) );
  XNOR2_X1 U15856 ( .A(n12661), .B(n12662), .ZN(n12655) );
  NAND2_X1 U15857 ( .A1(n12666), .A2(n12655), .ZN(n12656) );
  NAND2_X1 U15858 ( .A1(n12657), .A2(n12656), .ZN(n12658) );
  XNOR2_X1 U15859 ( .A(n12658), .B(n13841), .ZN(n13619) );
  NAND2_X1 U15860 ( .A1(n12658), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12659) );
  NAND2_X1 U15861 ( .A1(n12660), .A2(n12695), .ZN(n12668) );
  INV_X1 U15862 ( .A(n12661), .ZN(n12663) );
  NOR2_X1 U15863 ( .A1(n12663), .A2(n12662), .ZN(n12670) );
  INV_X1 U15864 ( .A(n12670), .ZN(n12664) );
  XNOR2_X1 U15865 ( .A(n12671), .B(n12664), .ZN(n12665) );
  NAND2_X1 U15866 ( .A1(n12666), .A2(n12665), .ZN(n12667) );
  NAND2_X1 U15867 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  OR2_X1 U15868 ( .A1(n12669), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16035) );
  NAND2_X1 U15869 ( .A1(n12669), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16034) );
  NAND2_X1 U15870 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NOR2_X1 U15871 ( .A1(n13541), .A2(n12672), .ZN(n12673) );
  NAND2_X1 U15872 ( .A1(n13836), .A2(n13835), .ZN(n12674) );
  INV_X1 U15873 ( .A(n13836), .ZN(n12675) );
  NAND2_X1 U15874 ( .A1(n12675), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12676) );
  INV_X2 U15875 ( .A(n16008), .ZN(n16009) );
  INV_X1 U15876 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12679) );
  AOI21_X1 U15877 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16009), .ZN(n16018) );
  NAND2_X1 U15878 ( .A1(n14647), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16005) );
  OAI21_X1 U15879 ( .B1(n16009), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16005), .ZN(n14745) );
  NOR3_X1 U15880 ( .A1(n16018), .A2(n14743), .A3(n14745), .ZN(n16004) );
  OR2_X1 U15881 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12680) );
  NAND2_X1 U15882 ( .A1(n16004), .A2(n12680), .ZN(n14835) );
  NAND2_X1 U15883 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12681) );
  NAND2_X1 U15884 ( .A1(n16005), .A2(n12681), .ZN(n14832) );
  AND2_X1 U15885 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14836) );
  NOR2_X1 U15886 ( .A1(n14832), .A2(n14836), .ZN(n14731) );
  NAND2_X1 U15887 ( .A1(n14835), .A2(n14731), .ZN(n12683) );
  NOR2_X1 U15888 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15994) );
  XNOR2_X1 U15889 ( .A(n16009), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14838) );
  NOR2_X1 U15890 ( .A1(n15994), .A2(n14838), .ZN(n12682) );
  NAND2_X1 U15891 ( .A1(n12683), .A2(n12682), .ZN(n14730) );
  INV_X1 U15892 ( .A(n14730), .ZN(n12684) );
  NAND2_X1 U15893 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16016) );
  INV_X1 U15894 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15895 ( .A1(n12685), .A2(n12742), .ZN(n12686) );
  NAND2_X1 U15896 ( .A1(n16009), .A2(n12686), .ZN(n16017) );
  XNOR2_X1 U15897 ( .A(n16009), .B(n14825), .ZN(n14719) );
  NAND3_X1 U15898 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14623) );
  NAND2_X1 U15899 ( .A1(n12688), .A2(n10154), .ZN(n14655) );
  NAND3_X1 U15900 ( .A1(n14673), .A2(n14794), .A3(n16049), .ZN(n14624) );
  AND2_X1 U15901 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14769) );
  NOR2_X1 U15902 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14768) );
  NAND2_X1 U15903 ( .A1(n12695), .A2(n11634), .ZN(n12704) );
  AND2_X1 U15904 ( .A1(n14846), .A2(n12696), .ZN(n12697) );
  NOR2_X1 U15905 ( .A1(n12698), .A2(n12697), .ZN(n12713) );
  AND2_X1 U15906 ( .A1(n12704), .A2(n11627), .ZN(n12699) );
  NAND2_X1 U15907 ( .A1(n11637), .A2(n12699), .ZN(n12732) );
  NAND2_X1 U15908 ( .A1(n12713), .A2(n12732), .ZN(n12700) );
  NAND2_X1 U15909 ( .A1(n12700), .A2(n12313), .ZN(n13323) );
  NAND2_X1 U15910 ( .A1(n11616), .A2(n20879), .ZN(n12702) );
  NAND3_X1 U15911 ( .A1(n12702), .A2(n12701), .A3(n11618), .ZN(n12703) );
  OAI211_X1 U15912 ( .C1(n12704), .C2(n15882), .A(n13323), .B(n12703), .ZN(
        n12706) );
  NAND2_X1 U15913 ( .A1(n12706), .A2(n12705), .ZN(n12711) );
  NAND2_X1 U15914 ( .A1(n13327), .A2(n12707), .ZN(n12708) );
  NAND3_X1 U15915 ( .A1(n12708), .A2(n11627), .A3(n11647), .ZN(n12709) );
  NAND3_X1 U15916 ( .A1(n12709), .A2(n13224), .A3(n11625), .ZN(n12710) );
  INV_X1 U15917 ( .A(n12712), .ZN(n12730) );
  INV_X1 U15918 ( .A(n13386), .ZN(n12714) );
  NOR2_X1 U15919 ( .A1(n15862), .A2(n12714), .ZN(n14308) );
  NAND2_X1 U15920 ( .A1(n11650), .A2(n11609), .ZN(n12715) );
  NAND3_X1 U15921 ( .A1(n11645), .A2(n14308), .A3(n12715), .ZN(n12716) );
  AOI22_X1 U15922 ( .A1(n12717), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n12341), .ZN(n12722) );
  OR2_X1 U15923 ( .A1(n12718), .A2(n12690), .ZN(n12720) );
  NAND2_X1 U15924 ( .A1(n12341), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15925 ( .A1(n12720), .A2(n12719), .ZN(n12865) );
  INV_X1 U15926 ( .A(n14504), .ZN(n12725) );
  OR2_X1 U15927 ( .A1(n12259), .A2(n11616), .ZN(n15876) );
  OAI21_X1 U15928 ( .B1(n12723), .B2(n11609), .A(n15876), .ZN(n12724) );
  INV_X1 U15929 ( .A(n13778), .ZN(n12726) );
  NAND2_X1 U15930 ( .A1(n12743), .A2(n13403), .ZN(n14810) );
  OAI21_X1 U15931 ( .B1(n12575), .B2(n12727), .A(n11616), .ZN(n12734) );
  OAI211_X1 U15932 ( .C1(n12730), .C2(n13778), .A(n12728), .B(n12729), .ZN(
        n12731) );
  INV_X1 U15933 ( .A(n12731), .ZN(n12733) );
  AND3_X1 U15934 ( .A1(n12734), .A2(n12733), .A3(n12732), .ZN(n12735) );
  OAI21_X1 U15935 ( .B1(n12736), .B2(n13777), .A(n12735), .ZN(n13314) );
  OAI21_X1 U15936 ( .B1(n12737), .B2(n11627), .A(n12738), .ZN(n12739) );
  OR2_X1 U15937 ( .A1(n13314), .A2(n12739), .ZN(n12740) );
  NAND2_X1 U15938 ( .A1(n12743), .A2(n12740), .ZN(n20161) );
  INV_X1 U15939 ( .A(n14306), .ZN(n12741) );
  INV_X1 U15940 ( .A(n20162), .ZN(n13349) );
  NOR2_X1 U15941 ( .A1(n15889), .A2(n14804), .ZN(n14803) );
  INV_X1 U15942 ( .A(n20157), .ZN(n12749) );
  NAND2_X1 U15943 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U15944 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14824) );
  NOR3_X1 U15945 ( .A1(n14825), .A2(n14821), .A3(n14824), .ZN(n14800) );
  INV_X1 U15946 ( .A(n14800), .ZN(n12747) );
  NOR2_X1 U15947 ( .A1(n13835), .A2(n16168), .ZN(n16143) );
  NAND4_X1 U15948 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16143), .ZN(n16119) );
  NOR2_X1 U15949 ( .A1(n12742), .A2(n16119), .ZN(n16127) );
  NAND2_X1 U15950 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16127), .ZN(
        n14822) );
  NAND2_X1 U15951 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13623) );
  INV_X1 U15952 ( .A(n13623), .ZN(n12745) );
  NAND3_X1 U15953 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n12745), .ZN(n13622) );
  NOR2_X1 U15954 ( .A1(n16179), .A2(n13622), .ZN(n16139) );
  INV_X1 U15955 ( .A(n16139), .ZN(n16118) );
  NOR2_X1 U15956 ( .A1(n14822), .A2(n16118), .ZN(n12759) );
  INV_X1 U15957 ( .A(n12759), .ZN(n12757) );
  NOR2_X1 U15958 ( .A1(n12747), .A2(n12757), .ZN(n16080) );
  NOR2_X1 U15959 ( .A1(n20161), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12744) );
  NOR2_X1 U15960 ( .A1(n12743), .A2(n20149), .ZN(n20171) );
  INV_X1 U15961 ( .A(n13352), .ZN(n13621) );
  AOI21_X1 U15962 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13468) );
  INV_X1 U15963 ( .A(n13468), .ZN(n13466) );
  NAND2_X1 U15964 ( .A1(n12745), .A2(n13466), .ZN(n16175) );
  NOR2_X1 U15965 ( .A1(n16179), .A2(n16175), .ZN(n13626) );
  INV_X1 U15966 ( .A(n14822), .ZN(n12746) );
  NAND2_X1 U15967 ( .A1(n13626), .A2(n12746), .ZN(n12758) );
  OAI21_X1 U15968 ( .B1(n12747), .B2(n12758), .A(n13349), .ZN(n12748) );
  OAI211_X1 U15969 ( .C1(n16140), .C2(n16080), .A(n13621), .B(n12748), .ZN(
        n16073) );
  OAI22_X1 U15970 ( .A1(n12754), .A2(n16073), .B1(n20157), .B2(n13352), .ZN(
        n15888) );
  OAI21_X1 U15971 ( .B1(n14803), .B2(n12749), .A(n15888), .ZN(n16065) );
  AOI21_X1 U15972 ( .B1(n13349), .B2(n14673), .A(n16065), .ZN(n14787) );
  AOI22_X1 U15973 ( .A1(n14794), .A2(n20157), .B1(n16117), .B2(n14673), .ZN(
        n12750) );
  NAND2_X1 U15974 ( .A1(n14787), .A2(n12750), .ZN(n16057) );
  NOR2_X1 U15975 ( .A1(n16049), .A2(n12408), .ZN(n16048) );
  INV_X1 U15976 ( .A(n16048), .ZN(n12761) );
  AND2_X1 U15977 ( .A1(n20157), .A2(n12761), .ZN(n12751) );
  NOR2_X1 U15978 ( .A1(n16057), .A2(n12751), .ZN(n14778) );
  INV_X1 U15979 ( .A(n14769), .ZN(n14759) );
  NAND2_X1 U15980 ( .A1(n20157), .A2(n14759), .ZN(n12752) );
  NAND2_X1 U15981 ( .A1(n14778), .A2(n12752), .ZN(n14765) );
  AOI211_X1 U15982 ( .C1(n12843), .C2(n20157), .A(n12690), .B(n14765), .ZN(
        n14752) );
  OAI21_X1 U15983 ( .B1(n16057), .B2(n20157), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U15984 ( .A1(n20149), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n12889) );
  OAI21_X1 U15985 ( .B1(n14752), .B2(n12753), .A(n12889), .ZN(n12763) );
  INV_X1 U15986 ( .A(n12754), .ZN(n12760) );
  INV_X1 U15987 ( .A(n14810), .ZN(n20172) );
  INV_X1 U15988 ( .A(n20161), .ZN(n12755) );
  NAND2_X1 U15989 ( .A1(n12755), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12756) );
  OAI22_X1 U15990 ( .A1(n20162), .A2(n12758), .B1(n12757), .B2(n12756), .ZN(
        n14799) );
  AOI21_X1 U15991 ( .B1(n20172), .B2(n12759), .A(n14799), .ZN(n16115) );
  INV_X1 U15992 ( .A(n16115), .ZN(n16100) );
  NAND4_X1 U15993 ( .A1(n12760), .A2(n16100), .A3(n14800), .A4(n14803), .ZN(
        n16072) );
  NOR2_X1 U15994 ( .A1(n14673), .A2(n16072), .ZN(n14795) );
  NAND2_X1 U15995 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14795), .ZN(
        n16064) );
  NOR2_X1 U15996 ( .A1(n16064), .A2(n12761), .ZN(n14784) );
  NAND3_X1 U15997 ( .A1(n14784), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14769), .ZN(n14753) );
  NOR3_X1 U15998 ( .A1(n14753), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12690), .ZN(n12762) );
  INV_X1 U15999 ( .A(n12768), .ZN(n12765) );
  NAND2_X1 U16000 ( .A1(n15137), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15138) );
  OAI21_X1 U16001 ( .B1(n12769), .B2(n12768), .A(n12767), .ZN(n12770) );
  NAND2_X1 U16002 ( .A1(n15138), .A2(n12770), .ZN(n12773) );
  XNOR2_X1 U16003 ( .A(n12771), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12772) );
  XNOR2_X1 U16004 ( .A(n12773), .B(n12772), .ZN(n12802) );
  OR2_X2 U16005 ( .A1(n12775), .A2(n12774), .ZN(n15276) );
  AOI21_X2 U16006 ( .B1(n12776), .B2(n15276), .A(n15123), .ZN(n12808) );
  NOR2_X1 U16007 ( .A1(n15031), .A2(n12777), .ZN(n12778) );
  NOR2_X1 U16008 ( .A1(n15328), .A2(n15340), .ZN(n15323) );
  AND2_X1 U16009 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15323), .ZN(
        n12779) );
  AND2_X1 U16010 ( .A1(n12780), .A2(n12779), .ZN(n15287) );
  NAND2_X1 U16011 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12791) );
  INV_X1 U16012 ( .A(n12791), .ZN(n12781) );
  NAND2_X1 U16013 ( .A1(n15287), .A2(n12781), .ZN(n12782) );
  NAND2_X1 U16014 ( .A1(n12782), .A2(n15424), .ZN(n15280) );
  INV_X1 U16015 ( .A(n15280), .ZN(n12788) );
  NOR2_X1 U16016 ( .A1(n12785), .A2(n12784), .ZN(n12786) );
  OR2_X2 U16017 ( .A1(n12783), .A2(n12786), .ZN(n16231) );
  NAND2_X1 U16018 ( .A1(n19286), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12803) );
  OAI21_X1 U16019 ( .B1(n16231), .B2(n19305), .A(n12803), .ZN(n12787) );
  AOI21_X1 U16020 ( .B1(n12788), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12787), .ZN(n12798) );
  INV_X1 U16021 ( .A(n15323), .ZN(n12789) );
  NAND3_X1 U16022 ( .A1(n15364), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15349), .ZN(n15335) );
  NOR2_X1 U16023 ( .A1(n12789), .A2(n15335), .ZN(n15313) );
  NOR2_X1 U16024 ( .A1(n12791), .A2(n12790), .ZN(n12792) );
  NAND2_X1 U16025 ( .A1(n15313), .A2(n12792), .ZN(n15277) );
  INV_X1 U16026 ( .A(n12793), .ZN(n12795) );
  NAND2_X1 U16027 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  OR2_X1 U16028 ( .A1(n15277), .A2(n12796), .ZN(n12797) );
  OAI211_X1 U16029 ( .C1(n16222), .C2(n16400), .A(n12798), .B(n12797), .ZN(
        n12799) );
  AOI21_X1 U16030 ( .B1(n12808), .B2(n16388), .A(n12799), .ZN(n12800) );
  NAND2_X1 U16031 ( .A1(n12801), .A2(n12800), .ZN(P2_U3018) );
  INV_X1 U16032 ( .A(n16228), .ZN(n12805) );
  OAI21_X1 U16033 ( .B1(n16365), .B2(n10219), .A(n12803), .ZN(n12804) );
  AOI21_X1 U16034 ( .B1(n16355), .B2(n12805), .A(n12804), .ZN(n12806) );
  OAI21_X1 U16035 ( .B1(n16231), .B2(n15258), .A(n12806), .ZN(n12807) );
  AOI21_X1 U16036 ( .B1(n12808), .B2(n10925), .A(n12807), .ZN(n12809) );
  NAND2_X1 U16037 ( .A1(n12810), .A2(n12809), .ZN(P2_U2986) );
  AND3_X1 U16038 ( .A1(n16196), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n12811) );
  NAND2_X1 U16039 ( .A1(n12812), .A2(n20178), .ZN(n12825) );
  XNOR2_X1 U16040 ( .A(n16009), .B(n12843), .ZN(n12813) );
  OR2_X1 U16041 ( .A1(n12815), .A2(n20858), .ZN(n20873) );
  NAND2_X1 U16042 ( .A1(n20873), .A2(n16196), .ZN(n12816) );
  NAND2_X1 U16043 ( .A1(n16196), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U16044 ( .A1(n12818), .A2(n12817), .ZN(n20151) );
  OAI22_X1 U16045 ( .A1(n16047), .A2(n12819), .B1(n20140), .B2(n21187), .ZN(
        n12820) );
  AOI21_X1 U16046 ( .B1(n16043), .B2(n12821), .A(n12820), .ZN(n12822) );
  NAND2_X1 U16047 ( .A1(n12825), .A2(n12824), .ZN(P1_U2970) );
  NAND2_X1 U16048 ( .A1(n12826), .A2(n16391), .ZN(n12836) );
  AOI222_X1 U16049 ( .A1(n11327), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12478), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11291), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12828) );
  NOR4_X1 U16050 ( .A1(n15277), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12851), .A4(n15262), .ZN(n12829) );
  AOI21_X1 U16051 ( .B1(n19302), .B2(n15262), .A(n12851), .ZN(n12831) );
  NAND2_X1 U16052 ( .A1(n15280), .A2(n12831), .ZN(n12854) );
  NAND3_X1 U16053 ( .A1(n12854), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15424), .ZN(n12832) );
  OAI211_X1 U16054 ( .C1(n16204), .C2(n16400), .A(n12833), .B(n12832), .ZN(
        n12834) );
  INV_X1 U16055 ( .A(n12834), .ZN(n12835) );
  OAI211_X1 U16056 ( .C1(n12837), .C2(n19311), .A(n12836), .B(n12835), .ZN(
        P2_U3015) );
  INV_X1 U16057 ( .A(n12839), .ZN(n12840) );
  NAND2_X1 U16058 ( .A1(n12256), .A2(n12840), .ZN(n12842) );
  NAND2_X1 U16059 ( .A1(n12842), .A2(n12841), .ZN(n14048) );
  INV_X1 U16060 ( .A(n14048), .ZN(n12862) );
  INV_X2 U16061 ( .A(n20142), .ZN(n20178) );
  NAND2_X1 U16062 ( .A1(n12862), .A2(n20178), .ZN(n12850) );
  NAND2_X1 U16063 ( .A1(n12844), .A2(n12843), .ZN(n12846) );
  NOR2_X1 U16064 ( .A1(n20141), .A2(n12866), .ZN(n12848) );
  NAND2_X1 U16065 ( .A1(n20149), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14751) );
  OAI21_X1 U16066 ( .B1(n16047), .B2(n12867), .A(n14751), .ZN(n12847) );
  OAI21_X1 U16067 ( .B1(n15277), .B2(n15262), .A(n12851), .ZN(n12855) );
  OAI21_X1 U16068 ( .B1(n14292), .B2(n19305), .A(n12852), .ZN(n12853) );
  AOI21_X1 U16069 ( .B1(n12855), .B2(n12854), .A(n12853), .ZN(n12856) );
  OAI21_X1 U16070 ( .B1(n14289), .B2(n16400), .A(n12856), .ZN(n12857) );
  NAND2_X1 U16071 ( .A1(n12862), .A2(n20047), .ZN(n12878) );
  OAI22_X1 U16072 ( .A1(n12867), .A2(n20057), .B1(n20059), .B2(n12866), .ZN(
        n12874) );
  INV_X1 U16073 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n12872) );
  NOR2_X1 U16074 ( .A1(n21187), .A2(n12868), .ZN(n12879) );
  INV_X1 U16075 ( .A(n12879), .ZN(n12871) );
  NAND2_X1 U16076 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n12870) );
  OAI21_X1 U16077 ( .B1(n12870), .B2(n12869), .A(n20029), .ZN(n12881) );
  AOI21_X1 U16078 ( .B1(n12872), .B2(n12871), .A(n12881), .ZN(n12873) );
  AOI211_X1 U16079 ( .C1(n20043), .C2(P1_EBX_REG_30__SCAN_IN), .A(n12874), .B(
        n12873), .ZN(n12875) );
  OAI21_X1 U16080 ( .B1(n14750), .B2(n15963), .A(n12875), .ZN(n12876) );
  INV_X1 U16081 ( .A(n12876), .ZN(n12877) );
  NAND2_X1 U16082 ( .A1(n12878), .A2(n12877), .ZN(P1_U2810) );
  NAND2_X1 U16083 ( .A1(n12888), .A2(n20047), .ZN(n12887) );
  INV_X1 U16084 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U16085 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n12879), .ZN(n12880) );
  OAI22_X1 U16086 ( .A1(n20057), .A2(n12890), .B1(P1_REIP_REG_31__SCAN_IN), 
        .B2(n12880), .ZN(n12883) );
  INV_X1 U16087 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21184) );
  NOR2_X1 U16088 ( .A1(n12881), .A2(n21184), .ZN(n12882) );
  AOI211_X1 U16089 ( .C1(P1_EBX_REG_31__SCAN_IN), .C2(n20043), .A(n12883), .B(
        n12882), .ZN(n12884) );
  NAND2_X1 U16090 ( .A1(n12887), .A2(n12886), .ZN(P1_U2809) );
  NAND2_X1 U16091 ( .A1(n12888), .A2(n20178), .ZN(n12895) );
  OAI21_X1 U16092 ( .B1(n16047), .B2(n12890), .A(n12889), .ZN(n12891) );
  AOI21_X1 U16093 ( .B1(n16043), .B2(n12892), .A(n12891), .ZN(n12894) );
  NOR2_X1 U16094 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12897) );
  NOR4_X1 U16095 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12896) );
  NAND4_X1 U16096 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12897), .A4(n12896), .ZN(n12909) );
  INV_X1 U16097 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21056) );
  NOR3_X1 U16098 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21056), .ZN(n12899) );
  NOR4_X1 U16099 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12898)
         );
  NAND4_X1 U16100 ( .A1(n20177), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12899), .A4(
        n12898), .ZN(U214) );
  NOR4_X1 U16101 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12903) );
  NOR4_X1 U16102 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12902) );
  NOR4_X1 U16103 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12901) );
  NOR4_X1 U16104 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12900) );
  NAND4_X1 U16105 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        n12908) );
  NOR4_X1 U16106 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12906) );
  NOR4_X1 U16107 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12905) );
  NOR4_X1 U16108 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12904) );
  NAND4_X1 U16109 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n19895), .ZN(
        n12907) );
  NOR2_X1 U16110 ( .A1(n13930), .A2(n12909), .ZN(n16547) );
  NAND2_X1 U16111 ( .A1(n16547), .A2(U214), .ZN(U212) );
  INV_X1 U16112 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16688) );
  NOR2_X1 U16113 ( .A1(n17954), .A2(n17956), .ZN(n17939) );
  NAND2_X1 U16114 ( .A1(n17939), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16678) );
  INV_X1 U16115 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17897) );
  NOR2_X1 U16116 ( .A1(n17912), .A2(n17897), .ZN(n17895) );
  INV_X1 U16117 ( .A(n17895), .ZN(n16924) );
  NAND2_X1 U16118 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17864) );
  NOR2_X1 U16119 ( .A1(n17848), .A2(n16885), .ZN(n16863) );
  INV_X1 U16120 ( .A(n16863), .ZN(n17834) );
  NAND3_X1 U16121 ( .A1(n17751), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17737) );
  NAND2_X1 U16122 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17671) );
  NAND2_X1 U16123 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17635) );
  NAND2_X1 U16124 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16510), .ZN(
        n16483) );
  NAND2_X1 U16125 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16507), .ZN(
        n12910) );
  XOR2_X2 U16126 ( .A(n16688), .B(n12910), .Z(n17001) );
  NAND2_X1 U16127 ( .A1(n17001), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13028) );
  INV_X1 U16128 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18877) );
  NOR2_X2 U16129 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18975), .ZN(n18745) );
  NAND2_X1 U16130 ( .A1(n18745), .A2(n18985), .ZN(n18870) );
  NAND2_X1 U16131 ( .A1(n18985), .A2(n18975), .ZN(n18979) );
  NAND2_X2 U16132 ( .A1(n18877), .A2(n19037), .ZN(n18216) );
  NOR3_X1 U16133 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18882) );
  NOR2_X1 U16134 ( .A1(n18330), .A2(n18878), .ZN(n13027) );
  INV_X2 U16135 ( .A(n17304), .ZN(n15676) );
  AOI22_X1 U16136 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12914) );
  OAI21_X1 U16137 ( .B1(n17283), .B2(n18354), .A(n12914), .ZN(n12929) );
  NOR2_X2 U16138 ( .A1(n18828), .A2(n12921), .ZN(n12915) );
  AOI22_X1 U16139 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12927) );
  INV_X1 U16140 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18608) );
  OR2_X2 U16141 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12918), .ZN(
        n17186) );
  AOI22_X1 U16142 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12919) );
  OAI21_X1 U16143 ( .B1(n9844), .B2(n18608), .A(n12919), .ZN(n12925) );
  AOI22_X1 U16144 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U16145 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12922) );
  OAI211_X1 U16146 ( .C1(n15691), .C2(n15602), .A(n12923), .B(n12922), .ZN(
        n12924) );
  AOI211_X1 U16147 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n12925), .B(n12924), .ZN(n12926) );
  OAI211_X1 U16148 ( .C1(n10447), .C2(n17185), .A(n12927), .B(n12926), .ZN(
        n12928) );
  AOI211_X4 U16149 ( .C1(n15676), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n12929), .B(n12928), .ZN(n19025) );
  INV_X1 U16150 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18392) );
  AOI22_X1 U16151 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16152 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12930) );
  OAI211_X1 U16153 ( .C1(n17306), .C2(n18392), .A(n12931), .B(n12930), .ZN(
        n12937) );
  AOI22_X1 U16154 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15714), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16155 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16156 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12933) );
  NAND2_X1 U16157 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12932) );
  NAND4_X1 U16158 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n12936) );
  AOI22_X1 U16159 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12940) );
  OAI21_X1 U16160 ( .B1(n9846), .B2(n17051), .A(n12940), .ZN(n12949) );
  AOI22_X1 U16161 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12947) );
  INV_X1 U16162 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U16163 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12941) );
  OAI21_X1 U16164 ( .B1(n15691), .B2(n17215), .A(n12941), .ZN(n12945) );
  INV_X1 U16165 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17057) );
  BUF_X2 U16166 ( .A(n15715), .Z(n17325) );
  AOI22_X1 U16167 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16168 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15714), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12942) );
  OAI211_X1 U16169 ( .C1(n17161), .C2(n17057), .A(n12943), .B(n12942), .ZN(
        n12944) );
  AOI211_X1 U16170 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n12945), .B(n12944), .ZN(n12946) );
  OAI211_X1 U16171 ( .C1(n17186), .C2(n18507), .A(n12947), .B(n12946), .ZN(
        n12948) );
  INV_X1 U16172 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18696) );
  INV_X2 U16173 ( .A(n9846), .ZN(n15654) );
  AOI22_X1 U16174 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12959) );
  INV_X1 U16175 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U16176 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16177 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12950) );
  OAI211_X1 U16178 ( .C1(n15691), .C2(n17156), .A(n12951), .B(n12950), .ZN(
        n12957) );
  AOI22_X1 U16179 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16180 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U16181 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U16182 ( .A1(n15686), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12952) );
  NAND4_X1 U16183 ( .A1(n12955), .A2(n12954), .A3(n12953), .A4(n12952), .ZN(
        n12956) );
  AOI211_X1 U16184 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n12957), .B(n12956), .ZN(n12958) );
  AOI22_X1 U16185 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12969) );
  INV_X1 U16186 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15633) );
  AOI22_X1 U16187 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16188 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12960) );
  OAI211_X1 U16189 ( .C1(n15691), .C2(n15633), .A(n12961), .B(n12960), .ZN(
        n12967) );
  AOI22_X1 U16190 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16191 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16192 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12963) );
  NAND2_X1 U16193 ( .A1(n15686), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12962) );
  NAND4_X1 U16194 ( .A1(n12965), .A2(n12964), .A3(n12963), .A4(n12962), .ZN(
        n12966) );
  INV_X1 U16195 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U16196 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12970) );
  OAI21_X1 U16197 ( .B1(n17304), .B2(n17259), .A(n12970), .ZN(n12980) );
  INV_X1 U16198 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U16199 ( .A1(n15607), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12977) );
  INV_X1 U16200 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17140) );
  OAI22_X1 U16201 ( .A1(n17161), .A2(n17140), .B1(n17283), .B2(n18368), .ZN(
        n12975) );
  AOI22_X1 U16202 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16203 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16204 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12971) );
  NAND3_X1 U16205 ( .A1(n12973), .A2(n12972), .A3(n12971), .ZN(n12974) );
  AOI211_X1 U16206 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n12975), .B(n12974), .ZN(n12976) );
  OAI211_X1 U16207 ( .C1(n17158), .C2(n12978), .A(n12977), .B(n12976), .ZN(
        n12979) );
  AOI22_X1 U16208 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12981) );
  OAI21_X1 U16209 ( .B1(n15688), .B2(n17235), .A(n12981), .ZN(n12988) );
  AOI22_X1 U16210 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12987) );
  INV_X1 U16211 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17111) );
  OAI22_X1 U16212 ( .A1(n17161), .A2(n17111), .B1(n17304), .B2(n17121), .ZN(
        n12986) );
  AOI22_X1 U16213 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16214 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U16215 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12982) );
  NAND3_X1 U16216 ( .A1(n12984), .A2(n12983), .A3(n12982), .ZN(n12985) );
  NAND2_X1 U16217 ( .A1(n18365), .A2(n9849), .ZN(n18819) );
  AOI22_X1 U16218 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12998) );
  INV_X1 U16219 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U16220 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16221 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12989) );
  OAI211_X1 U16222 ( .C1(n17161), .C2(n15566), .A(n12990), .B(n12989), .ZN(
        n12996) );
  AOI22_X1 U16223 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16224 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16225 ( .A1(n15607), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U16226 ( .A1(n15686), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12991) );
  NAND4_X1 U16227 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n12995) );
  NOR2_X1 U16228 ( .A1(n18355), .A2(n13000), .ZN(n14012) );
  INV_X1 U16229 ( .A(n18867), .ZN(n17561) );
  INV_X1 U16230 ( .A(n9849), .ZN(n18376) );
  NAND2_X1 U16231 ( .A1(n13012), .A2(n18355), .ZN(n14017) );
  NAND2_X1 U16232 ( .A1(n18867), .A2(n18350), .ZN(n13014) );
  NAND2_X1 U16233 ( .A1(n13000), .A2(n18821), .ZN(n15550) );
  INV_X1 U16234 ( .A(n18355), .ZN(n15773) );
  NAND2_X1 U16235 ( .A1(n18371), .A2(n15773), .ZN(n15772) );
  NAND2_X1 U16236 ( .A1(n9849), .A2(n18371), .ZN(n15919) );
  INV_X1 U16237 ( .A(n15919), .ZN(n18842) );
  NOR2_X1 U16238 ( .A1(n17371), .A2(n18842), .ZN(n15918) );
  NOR3_X1 U16239 ( .A1(n18350), .A2(n15915), .A3(n15918), .ZN(n14015) );
  AOI21_X1 U16240 ( .B1(n15772), .B2(n13010), .A(n14015), .ZN(n13002) );
  INV_X1 U16241 ( .A(n13002), .ZN(n13011) );
  NAND2_X1 U16242 ( .A1(n18384), .A2(n15778), .ZN(n13006) );
  NOR2_X1 U16243 ( .A1(n13003), .A2(n18360), .ZN(n13005) );
  NOR2_X1 U16244 ( .A1(n15919), .A2(n18365), .ZN(n13004) );
  AOI211_X1 U16245 ( .C1(n18365), .C2(n13006), .A(n13005), .B(n13004), .ZN(
        n13009) );
  NAND2_X1 U16246 ( .A1(n18350), .A2(n15915), .ZN(n14011) );
  INV_X1 U16247 ( .A(n14011), .ZN(n13007) );
  OAI21_X1 U16248 ( .B1(n13007), .B2(n18355), .A(n15778), .ZN(n13008) );
  OAI211_X1 U16249 ( .C1(n13010), .C2(n18345), .A(n13009), .B(n13008), .ZN(
        n14014) );
  NAND2_X1 U16250 ( .A1(n13012), .A2(n15765), .ZN(n15768) );
  INV_X1 U16251 ( .A(n14010), .ZN(n18834) );
  INV_X1 U16252 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18869) );
  OAI22_X1 U16253 ( .A1(n18999), .A2(n18847), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14020) );
  AND2_X1 U16254 ( .A1(n14020), .A2(n14018), .ZN(n13015) );
  AOI22_X1 U16255 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18852), .B2(n18992), .ZN(
        n13020) );
  OAI22_X1 U16256 ( .A1(n18856), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n13017), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13022) );
  NOR2_X1 U16257 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18856), .ZN(
        n13018) );
  NAND2_X1 U16258 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13017), .ZN(
        n13023) );
  AOI22_X1 U16259 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13022), .B1(
        n13018), .B2(n13023), .ZN(n14019) );
  NAND2_X1 U16260 ( .A1(n13021), .A2(n13020), .ZN(n13019) );
  OAI211_X1 U16261 ( .C1(n13021), .C2(n13020), .A(n14019), .B(n13019), .ZN(
        n14021) );
  XNOR2_X1 U16262 ( .A(n14018), .B(n14020), .ZN(n13026) );
  INV_X1 U16263 ( .A(n13022), .ZN(n13025) );
  NAND2_X1 U16264 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13023), .ZN(
        n13024) );
  AOI221_X1 U16265 ( .B1(n13028), .B2(n17003), .C1(n17019), .C2(n17003), .A(
        n17987), .ZN(n13036) );
  NAND2_X1 U16266 ( .A1(n18878), .A2(n13028), .ZN(n16960) );
  INV_X1 U16267 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19008) );
  OAI22_X1 U16268 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16960), .B1(
        n19008), .B2(n17017), .ZN(n13035) );
  INV_X1 U16269 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18897) );
  NAND2_X1 U16270 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18897), .ZN(n19033) );
  NOR2_X1 U16271 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18885) );
  NAND2_X1 U16272 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19026) );
  INV_X1 U16273 ( .A(n19026), .ZN(n18884) );
  AOI211_X1 U16274 ( .C1(n19025), .C2(n19023), .A(n18884), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18866) );
  INV_X1 U16275 ( .A(n13030), .ZN(n19038) );
  AOI211_X4 U16276 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18350), .A(n18866), .B(
        n19038), .ZN(n17014) );
  INV_X1 U16277 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17361) );
  NAND2_X1 U16278 ( .A1(n18828), .A2(n13029), .ZN(n18993) );
  NOR2_X1 U16279 ( .A1(n18345), .A2(n19036), .ZN(n17013) );
  INV_X1 U16280 ( .A(n17013), .ZN(n17042) );
  OAI22_X1 U16281 ( .A1(n17037), .A2(n17361), .B1(n18993), .B2(n17042), .ZN(
        n13034) );
  INV_X1 U16282 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19024) );
  NAND2_X1 U16283 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18350), .ZN(n13031) );
  AOI211_X4 U16284 ( .C1(n19026), .C2(n19024), .A(n19038), .B(n13031), .ZN(
        n17007) );
  INV_X1 U16285 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17367) );
  NAND2_X1 U16286 ( .A1(n17367), .A2(n17361), .ZN(n17025) );
  NOR2_X1 U16287 ( .A1(n17367), .A2(n17361), .ZN(n17357) );
  INV_X1 U16288 ( .A(n17357), .ZN(n13032) );
  NAND2_X1 U16289 ( .A1(n17025), .A2(n13032), .ZN(n17362) );
  OAI22_X1 U16290 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17026), .B1(n17036), 
        .B2(n17362), .ZN(n13033) );
  INV_X1 U16291 ( .A(n13145), .ZN(n13037) );
  AND2_X1 U16292 ( .A1(n13038), .A2(n13037), .ZN(n19213) );
  INV_X1 U16293 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13041) );
  NOR2_X1 U16294 ( .A1(n19756), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19042) );
  INV_X1 U16295 ( .A(n19042), .ZN(n13039) );
  OAI211_X1 U16296 ( .C1(n19213), .C2(n13041), .A(n13040), .B(n13039), .ZN(
        P2_U2814) );
  NOR2_X1 U16297 ( .A1(n14043), .A2(n19872), .ZN(n13083) );
  INV_X1 U16298 ( .A(n13083), .ZN(n13043) );
  INV_X1 U16299 ( .A(n13042), .ZN(n13081) );
  NOR2_X1 U16300 ( .A1(n16430), .A2(n13044), .ZN(n16439) );
  NOR2_X1 U16301 ( .A1(n16439), .A2(n13144), .ZN(n20003) );
  OAI21_X1 U16302 ( .B1(n13089), .B2(n20003), .A(n13045), .ZN(P2_U2819) );
  INV_X1 U16303 ( .A(n13148), .ZN(n13141) );
  AOI22_X1 U16304 ( .A1(n13118), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n13141), .ZN(n13048) );
  AOI22_X1 U16305 ( .A1(n19315), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19313), .ZN(n19322) );
  INV_X1 U16306 ( .A(n19322), .ZN(n13047) );
  NAND2_X1 U16307 ( .A1(n13077), .A2(n13047), .ZN(n13125) );
  NAND2_X1 U16308 ( .A1(n13048), .A2(n13125), .ZN(P2_U2952) );
  AOI22_X1 U16309 ( .A1(n13118), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13141), .ZN(n13050) );
  AOI22_X1 U16310 ( .A1(n19315), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13930), .ZN(n15017) );
  INV_X1 U16311 ( .A(n15017), .ZN(n13049) );
  NAND2_X1 U16312 ( .A1(n13077), .A2(n13049), .ZN(n13066) );
  NAND2_X1 U16313 ( .A1(n13050), .A2(n13066), .ZN(P2_U2980) );
  AOI22_X1 U16314 ( .A1(n13118), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16315 ( .A1(n19315), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13930), .ZN(n19354) );
  INV_X1 U16316 ( .A(n19354), .ZN(n13051) );
  NAND2_X1 U16317 ( .A1(n13077), .A2(n13051), .ZN(n13129) );
  NAND2_X1 U16318 ( .A1(n13052), .A2(n13129), .ZN(P2_U2974) );
  AOI22_X1 U16319 ( .A1(n13118), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16320 ( .A1(n19315), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13930), .ZN(n19340) );
  INV_X1 U16321 ( .A(n19340), .ZN(n13053) );
  NAND2_X1 U16322 ( .A1(n13077), .A2(n13053), .ZN(n13121) );
  NAND2_X1 U16323 ( .A1(n13054), .A2(n13121), .ZN(P2_U2971) );
  AOI22_X1 U16324 ( .A1(n13118), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16325 ( .A1(n19315), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19313), .ZN(n13477) );
  INV_X1 U16326 ( .A(n13477), .ZN(n15037) );
  NAND2_X1 U16327 ( .A1(n13077), .A2(n15037), .ZN(n13068) );
  NAND2_X1 U16328 ( .A1(n13055), .A2(n13068), .ZN(P2_U2977) );
  AOI22_X1 U16329 ( .A1(n13118), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16330 ( .A1(n19315), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13930), .ZN(n19333) );
  INV_X1 U16331 ( .A(n19333), .ZN(n19244) );
  NAND2_X1 U16332 ( .A1(n13077), .A2(n19244), .ZN(n13119) );
  NAND2_X1 U16333 ( .A1(n13056), .A2(n13119), .ZN(P2_U2969) );
  AOI22_X1 U16334 ( .A1(n13118), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16335 ( .A1(n19315), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13930), .ZN(n19336) );
  INV_X1 U16336 ( .A(n19336), .ZN(n13506) );
  NAND2_X1 U16337 ( .A1(n13077), .A2(n13506), .ZN(n13131) );
  NAND2_X1 U16338 ( .A1(n13057), .A2(n13131), .ZN(P2_U2970) );
  AOI22_X1 U16339 ( .A1(n13118), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16340 ( .A1(n19315), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13930), .ZN(n19346) );
  INV_X1 U16341 ( .A(n19346), .ZN(n13058) );
  NAND2_X1 U16342 ( .A1(n13077), .A2(n13058), .ZN(n13123) );
  NAND2_X1 U16343 ( .A1(n13059), .A2(n13123), .ZN(P2_U2973) );
  AOI22_X1 U16344 ( .A1(n13118), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16345 ( .A1(n19315), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19313), .ZN(n13540) );
  INV_X1 U16346 ( .A(n13540), .ZN(n15028) );
  NAND2_X1 U16347 ( .A1(n13077), .A2(n15028), .ZN(n13140) );
  NAND2_X1 U16348 ( .A1(n13060), .A2(n13140), .ZN(P2_U2978) );
  AOI22_X1 U16349 ( .A1(n13118), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16350 ( .A1(n19315), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19313), .ZN(n19329) );
  INV_X1 U16351 ( .A(n19329), .ZN(n13061) );
  NAND2_X1 U16352 ( .A1(n13077), .A2(n13061), .ZN(n13133) );
  NAND2_X1 U16353 ( .A1(n13062), .A2(n13133), .ZN(P2_U2968) );
  AOI22_X1 U16354 ( .A1(n13118), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16355 ( .A1(n19315), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13930), .ZN(n19343) );
  INV_X1 U16356 ( .A(n19343), .ZN(n19232) );
  NAND2_X1 U16357 ( .A1(n13077), .A2(n19232), .ZN(n13127) );
  NAND2_X1 U16358 ( .A1(n13063), .A2(n13127), .ZN(P2_U2972) );
  AOI22_X1 U16359 ( .A1(n13118), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16360 ( .A1(n19315), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19313), .ZN(n13445) );
  INV_X1 U16361 ( .A(n13445), .ZN(n15046) );
  NAND2_X1 U16362 ( .A1(n13077), .A2(n15046), .ZN(n13136) );
  NAND2_X1 U16363 ( .A1(n13064), .A2(n13136), .ZN(P2_U2976) );
  INV_X1 U16364 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U16365 ( .A1(n13118), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13065) );
  OAI211_X1 U16366 ( .C1(n13148), .C2(n13255), .A(n13066), .B(n13065), .ZN(
        P2_U2965) );
  INV_X1 U16367 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13252) );
  NAND2_X1 U16368 ( .A1(n13118), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13067) );
  OAI211_X1 U16369 ( .C1(n13148), .C2(n13252), .A(n13068), .B(n13067), .ZN(
        P2_U2962) );
  INV_X1 U16370 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19258) );
  INV_X1 U16371 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16576) );
  OR2_X1 U16372 ( .A1(n19313), .A2(n16576), .ZN(n13070) );
  NAND2_X1 U16373 ( .A1(n19313), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U16374 ( .A1(n13070), .A2(n13069), .ZN(n19224) );
  NAND2_X1 U16375 ( .A1(n13077), .A2(n19224), .ZN(n13074) );
  NAND2_X1 U16376 ( .A1(n13118), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13071) );
  OAI211_X1 U16377 ( .C1(n19258), .C2(n13148), .A(n13074), .B(n13071), .ZN(
        P2_U2979) );
  INV_X1 U16378 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19266) );
  INV_X1 U16379 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16584) );
  INV_X1 U16380 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17490) );
  AOI22_X1 U16381 ( .A1(n19315), .A2(n16584), .B1(n17490), .B2(n19313), .ZN(
        n19228) );
  NAND2_X1 U16382 ( .A1(n13077), .A2(n19228), .ZN(n13080) );
  NAND2_X1 U16383 ( .A1(n13118), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13072) );
  OAI211_X1 U16384 ( .C1(n19266), .C2(n13148), .A(n13080), .B(n13072), .ZN(
        P2_U2975) );
  INV_X1 U16385 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13158) );
  NAND2_X1 U16386 ( .A1(n13118), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13073) );
  OAI211_X1 U16387 ( .C1(n13158), .C2(n13148), .A(n13074), .B(n13073), .ZN(
        P2_U2964) );
  INV_X1 U16388 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19254) );
  INV_X1 U16389 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16572) );
  OR2_X1 U16390 ( .A1(n19313), .A2(n16572), .ZN(n13076) );
  NAND2_X1 U16391 ( .A1(n19313), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U16392 ( .A1(n13076), .A2(n13075), .ZN(n19221) );
  NAND2_X1 U16393 ( .A1(n13077), .A2(n19221), .ZN(n13138) );
  NAND2_X1 U16394 ( .A1(n13118), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13078) );
  OAI211_X1 U16395 ( .C1(n19254), .C2(n13148), .A(n13138), .B(n13078), .ZN(
        P2_U2981) );
  INV_X1 U16396 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U16397 ( .A1(n13118), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13079) );
  OAI211_X1 U16398 ( .C1(n13250), .C2(n13148), .A(n13080), .B(n13079), .ZN(
        P2_U2960) );
  NOR2_X1 U16399 ( .A1(n13145), .A2(n13081), .ZN(n13082) );
  NAND2_X1 U16400 ( .A1(n13147), .A2(n13082), .ZN(n13088) );
  NOR2_X1 U16401 ( .A1(n16430), .A2(n13084), .ZN(n13085) );
  AOI21_X1 U16402 ( .B1(n16432), .B2(n16433), .A(n13085), .ZN(n13180) );
  INV_X1 U16403 ( .A(n16432), .ZN(n16434) );
  INV_X1 U16404 ( .A(n13086), .ZN(n16431) );
  NAND2_X1 U16405 ( .A1(n16434), .A2(n16431), .ZN(n13169) );
  AND4_X1 U16406 ( .A1(n13088), .A2(n13180), .A3(n13087), .A4(n13169), .ZN(
        n16427) );
  OR2_X1 U16407 ( .A1(n16427), .A2(n13144), .ZN(n13092) );
  NOR2_X1 U16408 ( .A1(n19798), .A2(n15506), .ZN(n19991) );
  NAND2_X1 U16409 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19991), .ZN(n16469) );
  NOR2_X1 U16410 ( .A1(n13089), .A2(n16469), .ZN(n13090) );
  AOI21_X1 U16411 ( .B1(n19863), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13090), 
        .ZN(n13091) );
  AND2_X1 U16412 ( .A1(n13092), .A2(n13091), .ZN(n15546) );
  INV_X1 U16413 ( .A(n15546), .ZN(n13100) );
  INV_X1 U16414 ( .A(n13093), .ZN(n13094) );
  NOR2_X1 U16415 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  NAND2_X1 U16416 ( .A1(n13097), .A2(n13096), .ZN(n16440) );
  OR3_X1 U16417 ( .A1(n15546), .A2(n16440), .A3(n19958), .ZN(n13098) );
  OAI21_X1 U16418 ( .B1(n13100), .B2(n13099), .A(n13098), .ZN(P2_U3595) );
  OAI21_X1 U16419 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19204), .A(
        n13113), .ZN(n16404) );
  INV_X1 U16420 ( .A(n16404), .ZN(n13104) );
  NOR2_X1 U16421 ( .A1(n19170), .A2(n19060), .ZN(n16406) );
  OAI21_X1 U16422 ( .B1(n13102), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13101), .ZN(n16402) );
  NOR2_X1 U16423 ( .A1(n16358), .A2(n16402), .ZN(n13103) );
  AOI211_X1 U16424 ( .C1(n19291), .C2(n13104), .A(n16406), .B(n13103), .ZN(
        n13107) );
  OAI21_X1 U16425 ( .B1(n19287), .B2(n13105), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13106) );
  OAI211_X1 U16426 ( .C1(n15258), .C2(n19208), .A(n13107), .B(n13106), .ZN(
        P2_U3014) );
  INV_X1 U16427 ( .A(n13108), .ZN(n13109) );
  INV_X1 U16428 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21205) );
  NAND2_X1 U16429 ( .A1(n20858), .A2(n16195), .ZN(n13738) );
  OAI211_X1 U16430 ( .C1(n13109), .C2(n21205), .A(n13543), .B(n13738), .ZN(
        P1_U2801) );
  OAI21_X1 U16431 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13111), .A(
        n13110), .ZN(n19312) );
  NAND2_X1 U16432 ( .A1(n19286), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19309) );
  OAI21_X1 U16433 ( .B1(n16358), .B2(n19312), .A(n19309), .ZN(n13116) );
  OAI21_X1 U16434 ( .B1(n13113), .B2(n19182), .A(n13112), .ZN(n13114) );
  XOR2_X1 U16435 ( .A(n13114), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n19299) );
  OAI22_X1 U16436 ( .A1(n19299), .A2(n16356), .B1(n19180), .B2(n16365), .ZN(
        n13115) );
  AOI211_X1 U16437 ( .C1(n16355), .C2(n19180), .A(n13116), .B(n13115), .ZN(
        n13117) );
  OAI21_X1 U16438 ( .B1(n19304), .B2(n15258), .A(n13117), .ZN(P2_U3013) );
  AOI22_X1 U16439 ( .A1(n13118), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13141), .ZN(n13120) );
  NAND2_X1 U16440 ( .A1(n13120), .A2(n13119), .ZN(P2_U2954) );
  AOI22_X1 U16441 ( .A1(n13118), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13141), .ZN(n13122) );
  NAND2_X1 U16442 ( .A1(n13122), .A2(n13121), .ZN(P2_U2956) );
  AOI22_X1 U16443 ( .A1(n13118), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13141), .ZN(n13124) );
  NAND2_X1 U16444 ( .A1(n13124), .A2(n13123), .ZN(P2_U2958) );
  AOI22_X1 U16445 ( .A1(n13118), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U16446 ( .A1(n13126), .A2(n13125), .ZN(P2_U2967) );
  AOI22_X1 U16447 ( .A1(n13118), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U16448 ( .A1(n13128), .A2(n13127), .ZN(P2_U2957) );
  AOI22_X1 U16449 ( .A1(n13118), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16450 ( .A1(n13130), .A2(n13129), .ZN(P2_U2959) );
  AOI22_X1 U16451 ( .A1(n13118), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13132) );
  NAND2_X1 U16452 ( .A1(n13132), .A2(n13131), .ZN(P2_U2955) );
  AOI22_X1 U16453 ( .A1(n13118), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13134) );
  NAND2_X1 U16454 ( .A1(n13134), .A2(n13133), .ZN(P2_U2953) );
  INV_X1 U16455 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13156) );
  NAND2_X1 U16456 ( .A1(n13118), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13135) );
  OAI211_X1 U16457 ( .C1(n13148), .C2(n13156), .A(n13136), .B(n13135), .ZN(
        P2_U2961) );
  INV_X1 U16458 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U16459 ( .A1(n13118), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13137) );
  OAI211_X1 U16460 ( .C1(n13152), .C2(n13148), .A(n13138), .B(n13137), .ZN(
        P2_U2966) );
  INV_X1 U16461 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13154) );
  NAND2_X1 U16462 ( .A1(n13118), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13139) );
  OAI211_X1 U16463 ( .C1(n13148), .C2(n13154), .A(n13140), .B(n13139), .ZN(
        P2_U2963) );
  AOI22_X1 U16464 ( .A1(n19315), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19313), .ZN(n13833) );
  AOI22_X1 U16465 ( .A1(n13118), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n13141), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n13142) );
  OAI21_X1 U16466 ( .B1(n13833), .B2(n13143), .A(n13142), .ZN(P2_U2982) );
  NOR2_X1 U16467 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  NAND2_X1 U16468 ( .A1(n13147), .A2(n13146), .ZN(n13149) );
  NAND2_X1 U16469 ( .A1(n19250), .A2(n13150), .ZN(n13254) );
  NAND2_X1 U16470 ( .A1(n19863), .A2(n19991), .ZN(n14861) );
  INV_X2 U16471 ( .A(n14861), .ZN(n19282) );
  NOR2_X4 U16472 ( .A1(n19250), .A2(n19282), .ZN(n19267) );
  AOI22_X1 U16473 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19267), .B1(n19282), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13151) );
  OAI21_X1 U16474 ( .B1(n13152), .B2(n13254), .A(n13151), .ZN(P2_U2921) );
  AOI22_X1 U16475 ( .A1(n19282), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13153) );
  OAI21_X1 U16476 ( .B1(n13154), .B2(n13254), .A(n13153), .ZN(P2_U2924) );
  AOI22_X1 U16477 ( .A1(n19282), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13155) );
  OAI21_X1 U16478 ( .B1(n13156), .B2(n13254), .A(n13155), .ZN(P2_U2926) );
  AOI22_X1 U16479 ( .A1(n19282), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13157) );
  OAI21_X1 U16480 ( .B1(n13158), .B2(n13254), .A(n13157), .ZN(P2_U2923) );
  INV_X1 U16481 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U16482 ( .A1(n19282), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13159) );
  OAI21_X1 U16483 ( .B1(n15055), .B2(n13254), .A(n13159), .ZN(P2_U2928) );
  NAND2_X1 U16484 ( .A1(n13291), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13160) );
  NOR2_X1 U16485 ( .A1(n19756), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13161) );
  AOI21_X1 U16486 ( .B1(n13287), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13161), .ZN(n13162) );
  AOI21_X4 U16487 ( .B1(n13164), .B2(n13284), .A(n13163), .ZN(n15501) );
  NAND2_X1 U16488 ( .A1(n14957), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13166) );
  NAND4_X1 U16489 ( .A1(n13165), .A2(n13166), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19809), .ZN(n13167) );
  INV_X1 U16490 ( .A(n13168), .ZN(n15519) );
  NAND2_X1 U16491 ( .A1(n13169), .A2(n15519), .ZN(n13170) );
  NAND2_X1 U16492 ( .A1(n13170), .A2(n19866), .ZN(n13301) );
  MUX2_X1 U16493 ( .A(n19208), .B(n19201), .S(n15010), .Z(n13171) );
  OAI21_X1 U16494 ( .B1(n19988), .B2(n15012), .A(n13171), .ZN(P2_U2887) );
  NOR2_X1 U16495 ( .A1(n14313), .A2(n13172), .ZN(n13175) );
  INV_X1 U16496 ( .A(n13738), .ZN(n13173) );
  OAI21_X1 U16497 ( .B1(n13173), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20875), 
        .ZN(n13174) );
  OAI21_X1 U16498 ( .B1(n20875), .B2(n13175), .A(n13174), .ZN(P1_U3487) );
  INV_X1 U16499 ( .A(n13176), .ZN(n13178) );
  NAND2_X1 U16500 ( .A1(n13178), .A2(n13177), .ZN(n13179) );
  NAND2_X1 U16501 ( .A1(n13180), .A2(n13179), .ZN(n13181) );
  AND2_X1 U16502 ( .A1(n13182), .A2(n13925), .ZN(n13183) );
  NOR2_X1 U16503 ( .A1(n13186), .A2(n13185), .ZN(n13187) );
  NOR2_X1 U16504 ( .A1(n13188), .A2(n13187), .ZN(n19198) );
  NOR3_X1 U16505 ( .A1(n19988), .A2(n15120), .A3(n19198), .ZN(n13189) );
  AOI21_X1 U16506 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19231), .A(n13189), .ZN(
        n13192) );
  NAND2_X1 U16507 ( .A1(n19249), .A2(n19352), .ZN(n15023) );
  OAI21_X1 U16508 ( .B1(n15120), .B2(n19316), .A(n15023), .ZN(n13190) );
  NAND2_X1 U16509 ( .A1(n13190), .A2(n19198), .ZN(n13191) );
  OAI211_X1 U16510 ( .C1(n19322), .C2(n13834), .A(n13192), .B(n13191), .ZN(
        P2_U2919) );
  NAND2_X1 U16511 ( .A1(n13194), .A2(n13193), .ZN(n13196) );
  AND2_X1 U16512 ( .A1(n13196), .A2(n10260), .ZN(n14911) );
  INV_X1 U16513 ( .A(n14911), .ZN(n19971) );
  OAI21_X1 U16514 ( .B1(n13199), .B2(n13198), .A(n13197), .ZN(n14298) );
  NAND2_X1 U16515 ( .A1(n13201), .A2(n13200), .ZN(n14301) );
  NAND3_X1 U16516 ( .A1(n16391), .A2(n14302), .A3(n14301), .ZN(n13202) );
  OAI21_X1 U16517 ( .B1(n14298), .B2(n19311), .A(n13202), .ZN(n13203) );
  AOI21_X1 U16518 ( .B1(n19971), .B2(n19308), .A(n13203), .ZN(n13212) );
  INV_X1 U16519 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19892) );
  NOR2_X1 U16520 ( .A1(n19170), .A2(n19892), .ZN(n14296) );
  AOI21_X1 U16521 ( .B1(n16390), .B2(n15526), .A(n14296), .ZN(n13208) );
  NAND2_X1 U16522 ( .A1(n13205), .A2(n13204), .ZN(n13206) );
  NAND2_X1 U16523 ( .A1(n15381), .A2(n13206), .ZN(n13207) );
  OAI211_X1 U16524 ( .C1(n13209), .C2(n19301), .A(n13208), .B(n13207), .ZN(
        n13210) );
  INV_X1 U16525 ( .A(n13210), .ZN(n13211) );
  OAI211_X1 U16526 ( .C1(n13214), .C2(n13213), .A(n13212), .B(n13211), .ZN(
        P2_U3044) );
  NAND2_X1 U16527 ( .A1(n14174), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13216) );
  NAND2_X1 U16528 ( .A1(n15501), .A2(n13216), .ZN(n13269) );
  INV_X1 U16529 ( .A(n15501), .ZN(n13218) );
  INV_X1 U16530 ( .A(n13216), .ZN(n13217) );
  NAND2_X1 U16531 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  NAND2_X1 U16532 ( .A1(n13287), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13220) );
  XNOR2_X1 U16533 ( .A(n19984), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19451) );
  NAND2_X1 U16534 ( .A1(n19451), .A2(n19961), .ZN(n19632) );
  NAND2_X1 U16535 ( .A1(n13220), .A2(n19632), .ZN(n13221) );
  MUX2_X1 U16536 ( .A(n19304), .B(n10929), .S(n15010), .Z(n13223) );
  OAI21_X1 U16537 ( .B1(n19447), .B2(n15012), .A(n13223), .ZN(P2_U2886) );
  INV_X1 U16538 ( .A(n13403), .ZN(n14845) );
  NAND2_X1 U16539 ( .A1(n15876), .A2(n14845), .ZN(n13226) );
  INV_X1 U16540 ( .A(n20879), .ZN(n13225) );
  NAND2_X1 U16541 ( .A1(n16196), .A2(n15874), .ZN(n20877) );
  INV_X2 U16542 ( .A(n20877), .ZN(n20120) );
  NOR2_X4 U16543 ( .A1(n20095), .A2(n20120), .ZN(n15907) );
  AOI22_X1 U16544 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U16545 ( .B1(n12248), .B2(n13375), .A(n13227), .ZN(P1_U2907) );
  INV_X1 U16546 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21201) );
  AOI22_X1 U16547 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13228) );
  OAI21_X1 U16548 ( .B1(n21201), .B2(n13375), .A(n13228), .ZN(P1_U2908) );
  AOI22_X1 U16549 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13229) );
  OAI21_X1 U16550 ( .B1(n12211), .B2(n13375), .A(n13229), .ZN(P1_U2909) );
  AOI22_X1 U16551 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13230) );
  OAI21_X1 U16552 ( .B1(n12074), .B2(n13375), .A(n13230), .ZN(P1_U2916) );
  AOI22_X1 U16553 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16554 ( .B1(n21019), .B2(n13375), .A(n13231), .ZN(P1_U2912) );
  INV_X1 U16555 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21178) );
  AOI22_X1 U16556 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13232) );
  OAI21_X1 U16557 ( .B1(n21178), .B2(n13375), .A(n13232), .ZN(P1_U2914) );
  INV_X1 U16558 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21157) );
  AOI22_X1 U16559 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16560 ( .B1(n21157), .B2(n13375), .A(n13233), .ZN(P1_U2915) );
  AOI22_X1 U16561 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13234) );
  OAI21_X1 U16562 ( .B1(n12176), .B2(n13375), .A(n13234), .ZN(P1_U2911) );
  AOI22_X1 U16563 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16564 ( .B1(n12010), .B2(n13375), .A(n13235), .ZN(P1_U2920) );
  AOI22_X1 U16565 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13236) );
  OAI21_X1 U16566 ( .B1(n12136), .B2(n13375), .A(n13236), .ZN(P1_U2913) );
  OR3_X1 U16567 ( .A1(n13239), .A2(n13238), .A3(n13237), .ZN(n13240) );
  NAND2_X1 U16568 ( .A1(n13241), .A2(n13240), .ZN(n13965) );
  INV_X1 U16569 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19271) );
  OAI222_X1 U16570 ( .A1(n13834), .A2(n19346), .B1(n13965), .B2(n19239), .C1(
        n19271), .C2(n19249), .ZN(P2_U2913) );
  INV_X1 U16571 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U16572 ( .A1(n19282), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13242) );
  OAI21_X1 U16573 ( .B1(n15066), .B2(n13254), .A(n13242), .ZN(P2_U2929) );
  INV_X1 U16574 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15073) );
  AOI22_X1 U16575 ( .A1(n19282), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13243) );
  OAI21_X1 U16576 ( .B1(n15073), .B2(n13254), .A(n13243), .ZN(P2_U2930) );
  INV_X1 U16577 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15085) );
  AOI22_X1 U16578 ( .A1(n19282), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13244) );
  OAI21_X1 U16579 ( .B1(n15085), .B2(n13254), .A(n13244), .ZN(P2_U2931) );
  INV_X1 U16580 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U16581 ( .A1(n19282), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13245) );
  OAI21_X1 U16582 ( .B1(n15092), .B2(n13254), .A(n13245), .ZN(P2_U2932) );
  INV_X1 U16583 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U16584 ( .A1(n19282), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13246) );
  OAI21_X1 U16585 ( .B1(n15103), .B2(n13254), .A(n13246), .ZN(P2_U2933) );
  INV_X1 U16586 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U16587 ( .A1(n19282), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13247) );
  OAI21_X1 U16588 ( .B1(n15109), .B2(n13254), .A(n13247), .ZN(P2_U2934) );
  INV_X1 U16589 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U16590 ( .A1(n19282), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13248) );
  OAI21_X1 U16591 ( .B1(n13928), .B2(n13254), .A(n13248), .ZN(P2_U2935) );
  AOI22_X1 U16592 ( .A1(n19282), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U16593 ( .B1(n13250), .B2(n13254), .A(n13249), .ZN(P2_U2927) );
  AOI22_X1 U16594 ( .A1(n19282), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13251) );
  OAI21_X1 U16595 ( .B1(n13252), .B2(n13254), .A(n13251), .ZN(P2_U2925) );
  AOI22_X1 U16596 ( .A1(n19282), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U16597 ( .B1(n13255), .B2(n13254), .A(n13253), .ZN(P2_U2922) );
  OAI21_X1 U16598 ( .B1(n13258), .B2(n13257), .A(n13256), .ZN(n20148) );
  NAND2_X1 U16599 ( .A1(n11608), .A2(n11554), .ZN(n13259) );
  NAND2_X1 U16600 ( .A1(n20179), .A2(DATAI_0_), .ZN(n13261) );
  NAND2_X1 U16601 ( .A1(n20177), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13260) );
  AND2_X1 U16602 ( .A1(n13261), .A2(n13260), .ZN(n20187) );
  INV_X1 U16603 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20123) );
  OAI222_X1 U16604 ( .A1(n20148), .A2(n14622), .B1(n14604), .B2(n20187), .C1(
        n14602), .C2(n20123), .ZN(P1_U2904) );
  OAI21_X1 U16605 ( .B1(n13264), .B2(n13263), .A(n13262), .ZN(n20143) );
  NAND2_X1 U16606 ( .A1(n20179), .A2(DATAI_1_), .ZN(n13266) );
  NAND2_X1 U16607 ( .A1(n20177), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13265) );
  AND2_X1 U16608 ( .A1(n13266), .A2(n13265), .ZN(n20196) );
  INV_X1 U16609 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20119) );
  OAI222_X1 U16610 ( .A1(n20143), .A2(n14622), .B1(n14604), .B2(n20196), .C1(
        n14602), .C2(n20119), .ZN(P1_U2903) );
  OAI21_X1 U16611 ( .B1(n13268), .B2(n13267), .A(n16384), .ZN(n19159) );
  OAI222_X1 U16612 ( .A1(n13834), .A2(n19354), .B1(n19159), .B2(n19239), .C1(
        n19269), .C2(n19249), .ZN(P2_U2912) );
  INV_X1 U16613 ( .A(n13269), .ZN(n13270) );
  AOI21_X2 U16614 ( .B1(n13272), .B2(n13271), .A(n13270), .ZN(n13497) );
  NAND2_X1 U16615 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19662) );
  NAND2_X1 U16616 ( .A1(n19662), .A2(n19973), .ZN(n13274) );
  NOR2_X1 U16617 ( .A1(n19973), .A2(n19984), .ZN(n19797) );
  INV_X1 U16618 ( .A(n13285), .ZN(n13273) );
  NAND2_X1 U16619 ( .A1(n13274), .A2(n13273), .ZN(n19450) );
  NOR2_X1 U16620 ( .A1(n19450), .A2(n19756), .ZN(n13275) );
  AOI21_X1 U16621 ( .B1(n13287), .B2(n15529), .A(n13275), .ZN(n13276) );
  OAI21_X2 U16622 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n13281) );
  NAND2_X1 U16623 ( .A1(n14174), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13279) );
  XNOR2_X1 U16624 ( .A(n13281), .B(n13279), .ZN(n13496) );
  NAND2_X1 U16625 ( .A1(n13497), .A2(n13496), .ZN(n13283) );
  INV_X1 U16626 ( .A(n13279), .ZN(n13280) );
  NAND2_X1 U16627 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  OAI21_X1 U16628 ( .B1(n13285), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19961), .ZN(n13286) );
  NOR2_X1 U16629 ( .A1(n13286), .A2(n19851), .ZN(n19691) );
  AOI21_X1 U16630 ( .B1(n13287), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19691), .ZN(n13288) );
  NAND2_X1 U16631 ( .A1(n14174), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13290) );
  NAND2_X1 U16632 ( .A1(n13337), .A2(n13338), .ZN(n13295) );
  INV_X1 U16633 ( .A(n13290), .ZN(n13292) );
  AOI22_X1 U16634 ( .A1(n13293), .A2(n13292), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13291), .ZN(n13294) );
  INV_X1 U16635 ( .A(n14174), .ZN(n14222) );
  INV_X1 U16636 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13296) );
  XOR2_X1 U16637 ( .A(n13358), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13305)
         );
  NAND2_X1 U16638 ( .A1(n13298), .A2(n13297), .ZN(n13300) );
  AND2_X1 U16639 ( .A1(n13300), .A2(n10344), .ZN(n16361) );
  NOR2_X1 U16640 ( .A1(n15000), .A2(n13302), .ZN(n13303) );
  AOI21_X1 U16641 ( .B1(n16361), .B2(n15000), .A(n13303), .ZN(n13304) );
  OAI21_X1 U16642 ( .B1(n13305), .B2(n15012), .A(n13304), .ZN(P2_U2882) );
  XNOR2_X1 U16643 ( .A(n13307), .B(n13306), .ZN(n19977) );
  XNOR2_X1 U16644 ( .A(n19447), .B(n19977), .ZN(n13309) );
  NAND2_X1 U16645 ( .A1(n19316), .A2(n19198), .ZN(n13308) );
  NAND2_X1 U16646 ( .A1(n13309), .A2(n13308), .ZN(n13500) );
  OAI21_X1 U16647 ( .B1(n13309), .B2(n13308), .A(n13500), .ZN(n13310) );
  NAND2_X1 U16648 ( .A1(n13310), .A2(n19246), .ZN(n13312) );
  AOI22_X1 U16649 ( .A1(n19245), .A2(n19977), .B1(n19231), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13311) );
  OAI211_X1 U16650 ( .C1(n19329), .C2(n13834), .A(n13312), .B(n13311), .ZN(
        P2_U2918) );
  XNOR2_X1 U16651 ( .A(n13780), .B(n12718), .ZN(n20160) );
  INV_X1 U16652 ( .A(n20092), .ZN(n14537) );
  AOI22_X1 U16653 ( .A1(n20088), .A2(n20160), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14537), .ZN(n13313) );
  OAI21_X1 U16654 ( .B1(n20143), .B2(n14539), .A(n13313), .ZN(P1_U2871) );
  INV_X1 U16655 ( .A(n20861), .ZN(n13320) );
  INV_X1 U16656 ( .A(n13314), .ZN(n13319) );
  NAND2_X1 U16657 ( .A1(n13316), .A2(n12737), .ZN(n13317) );
  NOR2_X1 U16658 ( .A1(n13315), .A2(n13317), .ZN(n13318) );
  NAND3_X1 U16659 ( .A1(n13319), .A2(n13318), .A3(n12572), .ZN(n14849) );
  INV_X1 U16660 ( .A(n14849), .ZN(n13399) );
  OAI22_X1 U16661 ( .A1(n13320), .A2(n13399), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14846), .ZN(n15849) );
  OAI22_X1 U16662 ( .A1(n16195), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20841), .ZN(n13321) );
  AOI21_X1 U16663 ( .B1(n15849), .B2(n16188), .A(n13321), .ZN(n13336) );
  OAI211_X1 U16664 ( .C1(n13778), .C2(n11618), .A(n13323), .B(n13322), .ZN(
        n13324) );
  INV_X1 U16665 ( .A(n13324), .ZN(n13326) );
  AND2_X1 U16666 ( .A1(n13326), .A2(n13325), .ZN(n13333) );
  NAND2_X1 U16667 ( .A1(n13403), .A2(n20880), .ZN(n13329) );
  INV_X1 U16668 ( .A(n13327), .ZN(n13328) );
  AOI21_X1 U16669 ( .B1(n13329), .B2(n13328), .A(n20879), .ZN(n13331) );
  OAI21_X1 U16670 ( .B1(n13331), .B2(n13330), .A(n15882), .ZN(n13332) );
  NAND2_X1 U16671 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15874), .ZN(n16198) );
  INV_X1 U16672 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20014) );
  OAI22_X1 U16673 ( .A1(n15852), .A2(n20008), .B1(n16198), .B2(n20014), .ZN(
        n16186) );
  AOI21_X1 U16674 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n16196), .A(n16186), 
        .ZN(n20842) );
  NOR2_X1 U16675 ( .A1(n14845), .A2(n13334), .ZN(n15850) );
  AOI22_X1 U16676 ( .A1(n15850), .A2(n16188), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20842), .ZN(n13335) );
  OAI21_X1 U16677 ( .B1(n13336), .B2(n20842), .A(n13335), .ZN(P1_U3474) );
  INV_X1 U16678 ( .A(n19963), .ZN(n19360) );
  NOR2_X1 U16679 ( .A1(n13340), .A2(n13301), .ZN(n13341) );
  AOI21_X1 U16680 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n13301), .A(n13341), .ZN(
        n13342) );
  OAI21_X1 U16681 ( .B1(n19360), .B2(n15012), .A(n13342), .ZN(P2_U2884) );
  OAI21_X1 U16682 ( .B1(n12341), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13343), .ZN(n20166) );
  OAI222_X1 U16683 ( .A1(n20166), .A2(n14546), .B1(n20995), .B2(n20092), .C1(
        n20148), .C2(n14539), .ZN(P1_U2872) );
  XNOR2_X1 U16684 ( .A(n13345), .B(n13344), .ZN(n13442) );
  INV_X1 U16685 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14850) );
  NAND2_X1 U16686 ( .A1(n14850), .A2(n14810), .ZN(n20156) );
  NAND2_X1 U16687 ( .A1(n20156), .A2(n16117), .ZN(n14788) );
  NOR2_X1 U16688 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  OR2_X1 U16689 ( .A1(n13471), .A2(n13348), .ZN(n13818) );
  NAND2_X1 U16690 ( .A1(n20149), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13438) );
  NOR2_X1 U16691 ( .A1(n14850), .A2(n12328), .ZN(n13350) );
  OAI221_X1 U16692 ( .B1(n13468), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n13468), .C2(n13350), .A(n13349), .ZN(n13351) );
  OAI211_X1 U16693 ( .C1(n16151), .C2(n13818), .A(n13438), .B(n13351), .ZN(
        n13355) );
  NAND2_X1 U16694 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13353) );
  AOI21_X1 U16695 ( .B1(n16117), .B2(n13353), .A(n13352), .ZN(n13465) );
  NOR2_X1 U16696 ( .A1(n13465), .A2(n13356), .ZN(n13354) );
  AOI211_X1 U16697 ( .C1(n13467), .C2(n13356), .A(n13355), .B(n13354), .ZN(
        n13357) );
  OAI21_X1 U16698 ( .B1(n20176), .B2(n13442), .A(n13357), .ZN(P1_U3029) );
  INV_X1 U16699 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13360) );
  NOR2_X1 U16700 ( .A1(n13358), .A2(n13360), .ZN(n13362) );
  INV_X1 U16701 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13359) );
  OAI211_X1 U16702 ( .C1(n13362), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14961), .B(n13479), .ZN(n13367) );
  NOR2_X1 U16703 ( .A1(n13364), .A2(n13299), .ZN(n13365) );
  OR2_X1 U16704 ( .A1(n13363), .A2(n13365), .ZN(n13969) );
  INV_X1 U16705 ( .A(n13969), .ZN(n16348) );
  NAND2_X1 U16706 ( .A1(n15000), .A2(n16348), .ZN(n13366) );
  OAI211_X1 U16707 ( .C1(n15000), .C2(n13368), .A(n13367), .B(n13366), .ZN(
        P2_U2881) );
  INV_X1 U16708 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21250) );
  AOI22_X1 U16709 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20120), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15907), .ZN(n13369) );
  OAI21_X1 U16710 ( .B1(n21250), .B2(n13375), .A(n13369), .ZN(P1_U2906) );
  INV_X1 U16711 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U16712 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U16713 ( .B1(n13371), .B2(n13375), .A(n13370), .ZN(P1_U2918) );
  AOI22_X1 U16714 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13372) );
  OAI21_X1 U16715 ( .B1(n12026), .B2(n13375), .A(n13372), .ZN(P1_U2919) );
  AOI22_X1 U16716 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13373) );
  OAI21_X1 U16717 ( .B1(n12054), .B2(n13375), .A(n13373), .ZN(P1_U2917) );
  INV_X1 U16718 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U16719 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13374) );
  OAI21_X1 U16720 ( .B1(n20990), .B2(n13375), .A(n13374), .ZN(P1_U2910) );
  NAND2_X1 U16721 ( .A1(n20850), .A2(n14849), .ZN(n13392) );
  OR2_X1 U16722 ( .A1(n14849), .A2(n13376), .ZN(n13405) );
  AOI21_X1 U16723 ( .B1(n13377), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11795), .ZN(n13378) );
  NOR2_X1 U16724 ( .A1(n13379), .A2(n13378), .ZN(n20831) );
  INV_X1 U16725 ( .A(n13380), .ZN(n13381) );
  MUX2_X1 U16726 ( .A(n13381), .B(n11795), .S(n13400), .Z(n13383) );
  INV_X1 U16727 ( .A(n13382), .ZN(n13385) );
  NAND2_X1 U16728 ( .A1(n13383), .A2(n13385), .ZN(n13388) );
  OAI21_X1 U16729 ( .B1(n13377), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11795), .ZN(n13384) );
  AOI22_X1 U16730 ( .A1(n13385), .A2(n13384), .B1(n13377), .B2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U16731 ( .A1(n14306), .A2(n13386), .ZN(n13401) );
  AOI22_X1 U16732 ( .A1(n13403), .A2(n13388), .B1(n13387), .B2(n13401), .ZN(
        n13389) );
  OAI21_X1 U16733 ( .B1(n13405), .B2(n20831), .A(n13389), .ZN(n13390) );
  INV_X1 U16734 ( .A(n13390), .ZN(n13391) );
  NAND2_X1 U16735 ( .A1(n13392), .A2(n13391), .ZN(n20830) );
  INV_X1 U16736 ( .A(n15852), .ZN(n13409) );
  NAND2_X1 U16737 ( .A1(n20830), .A2(n13409), .ZN(n13394) );
  NAND2_X1 U16738 ( .A1(n15852), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13393) );
  NAND2_X1 U16739 ( .A1(n13394), .A2(n13393), .ZN(n15861) );
  NAND2_X1 U16740 ( .A1(n15861), .A2(n16195), .ZN(n13396) );
  AND2_X1 U16741 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20014), .ZN(n13412) );
  NAND2_X1 U16742 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13412), .ZN(
        n13395) );
  NAND2_X1 U16743 ( .A1(n13396), .A2(n13395), .ZN(n15873) );
  INV_X1 U16744 ( .A(n13397), .ZN(n13415) );
  OR2_X1 U16745 ( .A1(n13398), .A2(n13399), .ZN(n13408) );
  XNOR2_X1 U16746 ( .A(n13377), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n20840) );
  XNOR2_X1 U16747 ( .A(n13400), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13402) );
  AOI22_X1 U16748 ( .A1(n13403), .A2(n13402), .B1(n13401), .B2(n20840), .ZN(
        n13404) );
  OAI21_X1 U16749 ( .B1(n13405), .B2(n20840), .A(n13404), .ZN(n13406) );
  INV_X1 U16750 ( .A(n13406), .ZN(n13407) );
  NAND2_X1 U16751 ( .A1(n13408), .A2(n13407), .ZN(n20835) );
  NAND2_X1 U16752 ( .A1(n20835), .A2(n13409), .ZN(n13411) );
  NAND2_X1 U16753 ( .A1(n15852), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13410) );
  NAND2_X1 U16754 ( .A1(n13411), .A2(n13410), .ZN(n15857) );
  NAND2_X1 U16755 ( .A1(n15857), .A2(n16195), .ZN(n13414) );
  NAND2_X1 U16756 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13412), .ZN(
        n13413) );
  NAND2_X1 U16757 ( .A1(n13414), .A2(n13413), .ZN(n15872) );
  NAND3_X1 U16758 ( .A1(n15873), .A2(n13415), .A3(n15872), .ZN(n13423) );
  OR2_X1 U16759 ( .A1(n13416), .A2(n10037), .ZN(n13417) );
  XNOR2_X1 U16760 ( .A(n13417), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16189) );
  NAND2_X1 U16761 ( .A1(n16189), .A2(n16187), .ZN(n13419) );
  OR2_X1 U16762 ( .A1(n15852), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13420) );
  INV_X1 U16763 ( .A(n13420), .ZN(n13418) );
  NAND2_X1 U16764 ( .A1(n13419), .A2(n13418), .ZN(n13422) );
  OAI21_X1 U16765 ( .B1(n11821), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13420), .ZN(
        n13421) );
  NAND2_X1 U16766 ( .A1(n13422), .A2(n13421), .ZN(n15870) );
  NAND2_X1 U16767 ( .A1(n13423), .A2(n15870), .ZN(n15875) );
  INV_X1 U16768 ( .A(n16198), .ZN(n13424) );
  OAI21_X1 U16769 ( .B1(n15875), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13424), .ZN(
        n13425) );
  OAI21_X1 U16770 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n16196), .ZN(n20884) );
  NAND2_X1 U16771 ( .A1(n13425), .A2(n20236), .ZN(n20857) );
  NAND2_X1 U16772 ( .A1(n20466), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20860) );
  INV_X1 U16773 ( .A(n20860), .ZN(n13431) );
  NAND2_X1 U16774 ( .A1(n13427), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20708) );
  OAI211_X1 U16775 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n13427), .A(n20708), 
        .B(n20858), .ZN(n13428) );
  OAI21_X1 U16776 ( .B1(n20586), .B2(n13431), .A(n13428), .ZN(n13429) );
  NAND2_X1 U16777 ( .A1(n20857), .A2(n13429), .ZN(n13430) );
  OAI21_X1 U16778 ( .B1(n20857), .B2(n20514), .A(n13430), .ZN(P1_U3477) );
  XNOR2_X1 U16779 ( .A(n20456), .B(n20708), .ZN(n13432) );
  OAI22_X1 U16780 ( .A1(n13432), .A2(n20852), .B1(n13398), .B2(n13431), .ZN(
        n13433) );
  NAND2_X1 U16781 ( .A1(n20857), .A2(n13433), .ZN(n13434) );
  OAI21_X1 U16782 ( .B1(n20857), .B2(n15856), .A(n13434), .ZN(P1_U3476) );
  INV_X1 U16783 ( .A(n13436), .ZN(n13437) );
  AOI21_X1 U16784 ( .B1(n13435), .B2(n13262), .A(n13437), .ZN(n13452) );
  NOR2_X1 U16785 ( .A1(n20141), .A2(n13816), .ZN(n13440) );
  INV_X1 U16786 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13815) );
  OAI21_X1 U16787 ( .B1(n16047), .B2(n13815), .A(n13438), .ZN(n13439) );
  AOI211_X1 U16788 ( .C1(n13452), .C2(n20178), .A(n13440), .B(n13439), .ZN(
        n13441) );
  OAI21_X1 U16789 ( .B1(n20155), .B2(n13442), .A(n13441), .ZN(P1_U2997) );
  OR2_X1 U16790 ( .A1(n13443), .A2(n16383), .ZN(n13444) );
  NAND2_X1 U16791 ( .A1(n13444), .A2(n13475), .ZN(n15491) );
  INV_X1 U16792 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19264) );
  OAI222_X1 U16793 ( .A1(n13834), .A2(n13445), .B1(n15491), .B2(n19239), .C1(
        n19264), .C2(n19249), .ZN(P2_U2910) );
  XOR2_X1 U16794 ( .A(n13479), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13451)
         );
  NOR2_X1 U16795 ( .A1(n13363), .A2(n13447), .ZN(n13448) );
  OR2_X1 U16796 ( .A1(n13446), .A2(n13448), .ZN(n19157) );
  MUX2_X1 U16797 ( .A(n19157), .B(n13449), .S(n15010), .Z(n13450) );
  OAI21_X1 U16798 ( .B1(n13451), .B2(n15012), .A(n13450), .ZN(P2_U2880) );
  INV_X1 U16799 ( .A(n13452), .ZN(n13826) );
  NAND2_X1 U16800 ( .A1(n20179), .A2(DATAI_2_), .ZN(n13454) );
  NAND2_X1 U16801 ( .A1(n20177), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13453) );
  AND2_X1 U16802 ( .A1(n13454), .A2(n13453), .ZN(n20201) );
  INV_X1 U16803 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20117) );
  OAI222_X1 U16804 ( .A1(n13826), .A2(n14622), .B1(n14604), .B2(n20201), .C1(
        n14602), .C2(n20117), .ZN(P1_U2902) );
  OAI222_X1 U16805 ( .A1(n13826), .A2(n14539), .B1(n20092), .B2(n10158), .C1(
        n13818), .C2(n14546), .ZN(P1_U2870) );
  OAI21_X1 U16806 ( .B1(n13456), .B2(n13457), .A(n13459), .ZN(n13487) );
  NAND2_X1 U16807 ( .A1(n20179), .A2(DATAI_3_), .ZN(n13461) );
  NAND2_X1 U16808 ( .A1(n20177), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13460) );
  AND2_X1 U16809 ( .A1(n13461), .A2(n13460), .ZN(n20206) );
  INV_X1 U16810 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13462) );
  OAI222_X1 U16811 ( .A1(n13487), .A2(n14622), .B1(n14604), .B2(n20206), .C1(
        n13462), .C2(n14602), .ZN(P1_U2901) );
  XNOR2_X1 U16812 ( .A(n13464), .B(n13463), .ZN(n13492) );
  OAI21_X1 U16813 ( .B1(n20162), .B2(n13466), .A(n13465), .ZN(n13515) );
  NAND2_X1 U16814 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13467), .ZN(
        n16116) );
  AOI22_X1 U16815 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13515), .B1(
        n13625), .B2(n13469), .ZN(n13474) );
  OAI21_X1 U16816 ( .B1(n13471), .B2(n13470), .A(n13512), .ZN(n13472) );
  INV_X1 U16817 ( .A(n13472), .ZN(n20087) );
  AND2_X1 U16818 ( .A1(n20149), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13488) );
  AOI21_X1 U16819 ( .B1(n20087), .B2(n20169), .A(n13488), .ZN(n13473) );
  OAI211_X1 U16820 ( .C1(n20176), .C2(n13492), .A(n13474), .B(n13473), .ZN(
        P1_U3028) );
  XNOR2_X1 U16821 ( .A(n13476), .B(n13475), .ZN(n15476) );
  INV_X1 U16822 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19262) );
  OAI222_X1 U16823 ( .A1(n13834), .A2(n13477), .B1(n15476), .B2(n19239), .C1(
        n19262), .C2(n19249), .ZN(P2_U2909) );
  INV_X1 U16824 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U16825 ( .A1(n13480), .A2(n13482), .ZN(n13529) );
  OAI211_X1 U16826 ( .C1(n13480), .C2(n13482), .A(n13481), .B(n14961), .ZN(
        n13486) );
  OAI21_X1 U16827 ( .B1(n13446), .B2(n13484), .A(n13483), .ZN(n19150) );
  INV_X1 U16828 ( .A(n19150), .ZN(n16389) );
  NAND2_X1 U16829 ( .A1(n15000), .A2(n16389), .ZN(n13485) );
  OAI211_X1 U16830 ( .C1(n15000), .C2(n11111), .A(n13486), .B(n13485), .ZN(
        P2_U2879) );
  INV_X1 U16831 ( .A(n13487), .ZN(n20090) );
  AOI21_X1 U16832 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13488), .ZN(n13489) );
  OAI21_X1 U16833 ( .B1(n20072), .B2(n20141), .A(n13489), .ZN(n13490) );
  AOI21_X1 U16834 ( .B1(n20090), .B2(n20178), .A(n13490), .ZN(n13491) );
  OAI21_X1 U16835 ( .B1(n20155), .B2(n13492), .A(n13491), .ZN(P1_U2996) );
  OR2_X1 U16836 ( .A1(n13494), .A2(n13493), .ZN(n13495) );
  NAND2_X1 U16837 ( .A1(n13495), .A2(n13590), .ZN(n13719) );
  XNOR2_X1 U16838 ( .A(n19963), .B(n13719), .ZN(n13504) );
  INV_X1 U16839 ( .A(n13497), .ZN(n13498) );
  INV_X1 U16840 ( .A(n19448), .ZN(n19969) );
  NAND2_X1 U16841 ( .A1(n19969), .A2(n14911), .ZN(n13502) );
  XNOR2_X1 U16842 ( .A(n19448), .B(n14911), .ZN(n19242) );
  INV_X1 U16843 ( .A(n19977), .ZN(n13499) );
  NAND2_X1 U16844 ( .A1(n19447), .A2(n13499), .ZN(n13501) );
  NAND2_X1 U16845 ( .A1(n13501), .A2(n13500), .ZN(n19241) );
  NAND2_X1 U16846 ( .A1(n19242), .A2(n19241), .ZN(n19240) );
  NAND2_X1 U16847 ( .A1(n13502), .A2(n19240), .ZN(n13503) );
  NAND2_X1 U16848 ( .A1(n13504), .A2(n13503), .ZN(n13589) );
  OAI21_X1 U16849 ( .B1(n13504), .B2(n13503), .A(n13589), .ZN(n13505) );
  NAND2_X1 U16850 ( .A1(n13505), .A2(n19246), .ZN(n13508) );
  AOI22_X1 U16851 ( .A1(n19243), .A2(n13506), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19231), .ZN(n13507) );
  OAI211_X1 U16852 ( .C1(n13719), .C2(n15023), .A(n13508), .B(n13507), .ZN(
        P2_U2916) );
  XNOR2_X1 U16853 ( .A(n13510), .B(n13509), .ZN(n13525) );
  OAI211_X1 U16854 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13623), .B(n13625), .ZN(n13517) );
  INV_X1 U16855 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21170) );
  NOR2_X1 U16856 ( .A1(n20140), .A2(n21170), .ZN(n13521) );
  NAND2_X1 U16857 ( .A1(n13512), .A2(n13511), .ZN(n13513) );
  NAND2_X1 U16858 ( .A1(n16171), .A2(n13513), .ZN(n14494) );
  NOR2_X1 U16859 ( .A1(n14494), .A2(n16151), .ZN(n13514) );
  AOI211_X1 U16860 ( .C1(n13515), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13521), .B(n13514), .ZN(n13516) );
  OAI211_X1 U16861 ( .C1(n13525), .C2(n20176), .A(n13517), .B(n13516), .ZN(
        P1_U3027) );
  AOI21_X1 U16862 ( .B1(n13520), .B2(n13459), .A(n11853), .ZN(n13526) );
  AOI21_X1 U16863 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13521), .ZN(n13522) );
  OAI21_X1 U16864 ( .B1(n14493), .B2(n20141), .A(n13522), .ZN(n13523) );
  AOI21_X1 U16865 ( .B1(n13526), .B2(n20178), .A(n13523), .ZN(n13524) );
  OAI21_X1 U16866 ( .B1(n20155), .B2(n13525), .A(n13524), .ZN(P1_U2995) );
  INV_X1 U16867 ( .A(n13526), .ZN(n14502) );
  NAND2_X1 U16868 ( .A1(n20179), .A2(DATAI_4_), .ZN(n13528) );
  NAND2_X1 U16869 ( .A1(n20177), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13527) );
  AND2_X1 U16870 ( .A1(n13528), .A2(n13527), .ZN(n20210) );
  INV_X1 U16871 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20114) );
  OAI222_X1 U16872 ( .A1(n14502), .A2(n14622), .B1(n14604), .B2(n20210), .C1(
        n14602), .C2(n20114), .ZN(P1_U2900) );
  INV_X1 U16873 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20982) );
  OAI222_X1 U16874 ( .A1(n14502), .A2(n14539), .B1(n20092), .B2(n20982), .C1(
        n14494), .C2(n14546), .ZN(P1_U2868) );
  INV_X2 U16875 ( .A(n13529), .ZN(n13532) );
  OAI211_X1 U16876 ( .C1(n13532), .C2(n13531), .A(n14961), .B(n13634), .ZN(
        n13537) );
  NAND2_X1 U16877 ( .A1(n13533), .A2(n13483), .ZN(n13535) );
  INV_X1 U16878 ( .A(n13600), .ZN(n13534) );
  AND2_X1 U16879 ( .A1(n13535), .A2(n13534), .ZN(n16332) );
  NAND2_X1 U16880 ( .A1(n15000), .A2(n16332), .ZN(n13536) );
  OAI211_X1 U16881 ( .C1(n15000), .C2(n11114), .A(n13537), .B(n13536), .ZN(
        P2_U2878) );
  INV_X1 U16882 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19260) );
  OAI21_X1 U16883 ( .B1(n13539), .B2(n13538), .A(n15441), .ZN(n19130) );
  OAI222_X1 U16884 ( .A1(n13834), .A2(n13540), .B1(n19249), .B2(n19260), .C1(
        n19239), .C2(n19130), .ZN(P2_U2908) );
  NAND2_X1 U16885 ( .A1(n13587), .A2(n11616), .ZN(n13588) );
  INV_X1 U16886 ( .A(DATAI_14_), .ZN(n21245) );
  NAND2_X1 U16887 ( .A1(n20177), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13544) );
  OAI21_X1 U16888 ( .B1(n20177), .B2(n21245), .A(n13544), .ZN(n14606) );
  NAND2_X1 U16889 ( .A1(n13766), .A2(n14606), .ZN(n20136) );
  NAND2_X1 U16890 ( .A1(n20134), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13545) );
  OAI211_X1 U16891 ( .C1(n21250), .C2(n13748), .A(n20136), .B(n13545), .ZN(
        P1_U2951) );
  INV_X1 U16892 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20108) );
  INV_X1 U16893 ( .A(DATAI_8_), .ZN(n21188) );
  NAND2_X1 U16894 ( .A1(n20177), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13546) );
  OAI21_X1 U16895 ( .B1(n20177), .B2(n21188), .A(n13546), .ZN(n14567) );
  NAND2_X1 U16896 ( .A1(n13766), .A2(n14567), .ZN(n13751) );
  NAND2_X1 U16897 ( .A1(n20134), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13547) );
  OAI211_X1 U16898 ( .C1(n20108), .C2(n13748), .A(n13751), .B(n13547), .ZN(
        P1_U2960) );
  INV_X1 U16899 ( .A(DATAI_12_), .ZN(n13549) );
  NAND2_X1 U16900 ( .A1(n20177), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13548) );
  OAI21_X1 U16901 ( .B1(n20177), .B2(n13549), .A(n13548), .ZN(n14611) );
  NAND2_X1 U16902 ( .A1(n13766), .A2(n14611), .ZN(n20130) );
  NAND2_X1 U16903 ( .A1(n20134), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13550) );
  OAI211_X1 U16904 ( .C1(n21201), .C2(n13748), .A(n20130), .B(n13550), .ZN(
        P1_U2949) );
  INV_X1 U16905 ( .A(DATAI_11_), .ZN(n21182) );
  NAND2_X1 U16906 ( .A1(n20177), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13551) );
  OAI21_X1 U16907 ( .B1(n20177), .B2(n21182), .A(n13551), .ZN(n14619) );
  NAND2_X1 U16908 ( .A1(n13766), .A2(n14619), .ZN(n20128) );
  NAND2_X1 U16909 ( .A1(n20134), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13552) );
  OAI211_X1 U16910 ( .C1(n12211), .C2(n13748), .A(n20128), .B(n13552), .ZN(
        P1_U2948) );
  INV_X1 U16911 ( .A(DATAI_10_), .ZN(n21234) );
  INV_X1 U16912 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16580) );
  MUX2_X1 U16913 ( .A(n21234), .B(n16580), .S(n20177), .Z(n14555) );
  INV_X1 U16914 ( .A(n14555), .ZN(n13553) );
  NAND2_X1 U16915 ( .A1(n13766), .A2(n13553), .ZN(n20126) );
  NAND2_X1 U16916 ( .A1(n20134), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13554) );
  OAI211_X1 U16917 ( .C1(n20990), .C2(n13748), .A(n20126), .B(n13554), .ZN(
        P1_U2947) );
  INV_X1 U16918 ( .A(DATAI_13_), .ZN(n21047) );
  NAND2_X1 U16919 ( .A1(n20177), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16920 ( .B1(n20177), .B2(n21047), .A(n13555), .ZN(n14609) );
  NAND2_X1 U16921 ( .A1(n13766), .A2(n14609), .ZN(n20132) );
  NAND2_X1 U16922 ( .A1(n20134), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13556) );
  OAI211_X1 U16923 ( .C1(n12248), .C2(n13748), .A(n20132), .B(n13556), .ZN(
        P1_U2950) );
  INV_X1 U16924 ( .A(DATAI_9_), .ZN(n21022) );
  NAND2_X1 U16925 ( .A1(n20177), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13557) );
  OAI21_X1 U16926 ( .B1(n20177), .B2(n21022), .A(n13557), .ZN(n14560) );
  NAND2_X1 U16927 ( .A1(n13766), .A2(n14560), .ZN(n20124) );
  NAND2_X1 U16928 ( .A1(n20134), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13558) );
  OAI211_X1 U16929 ( .C1(n12176), .C2(n13748), .A(n20124), .B(n13558), .ZN(
        P1_U2946) );
  INV_X1 U16930 ( .A(n13561), .ZN(n13562) );
  NAND2_X1 U16931 ( .A1(n13562), .A2(n13519), .ZN(n13563) );
  AND2_X1 U16932 ( .A1(n13560), .A2(n13563), .ZN(n20085) );
  INV_X1 U16933 ( .A(n20085), .ZN(n13567) );
  NAND2_X1 U16934 ( .A1(n20179), .A2(DATAI_5_), .ZN(n13565) );
  NAND2_X1 U16935 ( .A1(n20177), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13564) );
  AND2_X1 U16936 ( .A1(n13565), .A2(n13564), .ZN(n20215) );
  OAI222_X1 U16937 ( .A1(n13567), .A2(n14622), .B1(n14604), .B2(n20215), .C1(
        n13566), .C2(n14602), .ZN(P1_U2899) );
  NAND2_X1 U16938 ( .A1(n13569), .A2(n13568), .ZN(n13571) );
  XNOR2_X1 U16939 ( .A(n13571), .B(n13570), .ZN(n14031) );
  INV_X1 U16940 ( .A(n13572), .ZN(n13573) );
  XNOR2_X1 U16941 ( .A(n13574), .B(n13573), .ZN(n14032) );
  AOI21_X1 U16942 ( .B1(n15381), .B2(n13576), .A(n13575), .ZN(n13989) );
  INV_X1 U16943 ( .A(n13662), .ZN(n13578) );
  MUX2_X1 U16944 ( .A(n13989), .B(n13578), .S(n13577), .Z(n13582) );
  INV_X1 U16945 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19894) );
  NOR2_X1 U16946 ( .A1(n19894), .A2(n19170), .ZN(n13580) );
  AOI21_X1 U16947 ( .B1(n16390), .B2(n15545), .A(n13580), .ZN(n13581) );
  OAI211_X1 U16948 ( .C1(n16400), .C2(n13719), .A(n13582), .B(n13581), .ZN(
        n13583) );
  AOI21_X1 U16949 ( .B1(n16388), .B2(n14032), .A(n13583), .ZN(n13584) );
  OAI21_X1 U16950 ( .B1(n14031), .B2(n19300), .A(n13584), .ZN(P2_U3043) );
  INV_X1 U16951 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14601) );
  INV_X1 U16952 ( .A(DATAI_15_), .ZN(n13586) );
  INV_X1 U16953 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13585) );
  MUX2_X1 U16954 ( .A(n13586), .B(n13585), .S(n20177), .Z(n14603) );
  INV_X1 U16955 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20094) );
  OAI222_X1 U16956 ( .A1(n13748), .A2(n14601), .B1(n13588), .B2(n14603), .C1(
        n13587), .C2(n20094), .ZN(P1_U2967) );
  INV_X1 U16957 ( .A(n13719), .ZN(n19962) );
  OAI21_X1 U16958 ( .B1(n19963), .B2(n19962), .A(n13589), .ZN(n13592) );
  XNOR2_X1 U16959 ( .A(n13591), .B(n13590), .ZN(n13665) );
  NAND2_X1 U16960 ( .A1(n13592), .A2(n13665), .ZN(n19235) );
  OAI21_X1 U16961 ( .B1(n13594), .B2(n13593), .A(n13358), .ZN(n19233) );
  XNOR2_X1 U16962 ( .A(n19235), .B(n19233), .ZN(n13595) );
  NAND2_X1 U16963 ( .A1(n13595), .A2(n19246), .ZN(n13597) );
  INV_X1 U16964 ( .A(n13665), .ZN(n19168) );
  AOI22_X1 U16965 ( .A1(n19245), .A2(n19168), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19231), .ZN(n13596) );
  OAI211_X1 U16966 ( .C1(n19340), .C2(n13834), .A(n13597), .B(n13596), .ZN(
        P2_U2915) );
  INV_X1 U16967 ( .A(n13634), .ZN(n13599) );
  OR2_X1 U16968 ( .A1(n13634), .A2(n13631), .ZN(n13637) );
  OAI211_X1 U16969 ( .C1(n13599), .C2(n13598), .A(n14961), .B(n13637), .ZN(
        n13604) );
  OR2_X1 U16970 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  NAND2_X1 U16971 ( .A1(n13602), .A2(n13605), .ZN(n15471) );
  INV_X1 U16972 ( .A(n15471), .ZN(n16323) );
  NAND2_X1 U16973 ( .A1(n15000), .A2(n16323), .ZN(n13603) );
  OAI211_X1 U16974 ( .C1(n14983), .C2(n11118), .A(n13604), .B(n13603), .ZN(
        P2_U2877) );
  INV_X1 U16975 ( .A(n13630), .ZN(n13636) );
  XNOR2_X1 U16976 ( .A(n13637), .B(n13636), .ZN(n13610) );
  NAND2_X1 U16977 ( .A1(n13606), .A2(n13605), .ZN(n13607) );
  INV_X1 U16978 ( .A(n16319), .ZN(n19139) );
  MUX2_X1 U16979 ( .A(n19139), .B(n13608), .S(n15010), .Z(n13609) );
  OAI21_X1 U16980 ( .B1(n13610), .B2(n15012), .A(n13609), .ZN(P2_U2876) );
  OAI21_X1 U16981 ( .B1(n13612), .B2(n13615), .A(n13614), .ZN(n16038) );
  INV_X1 U16982 ( .A(DATAI_7_), .ZN(n13617) );
  NAND2_X1 U16983 ( .A1(n20177), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13616) );
  OAI21_X1 U16984 ( .B1(n20177), .B2(n13617), .A(n13616), .ZN(n20229) );
  AOI22_X1 U16985 ( .A1(n14620), .A2(n20229), .B1(P1_EAX_REG_7__SCAN_IN), .B2(
        n14618), .ZN(n13618) );
  OAI21_X1 U16986 ( .B1(n16038), .B2(n14622), .A(n13618), .ZN(P1_U2897) );
  XNOR2_X1 U16987 ( .A(n13620), .B(n13619), .ZN(n13653) );
  OR2_X1 U16988 ( .A1(n13626), .A2(n20162), .ZN(n16176) );
  NAND2_X1 U16989 ( .A1(n16176), .A2(n13621), .ZN(n16141) );
  AOI21_X1 U16990 ( .B1(n13622), .B2(n16117), .A(n16141), .ZN(n16180) );
  NOR2_X1 U16991 ( .A1(n16116), .A2(n13623), .ZN(n13624) );
  NAND2_X1 U16992 ( .A1(n13624), .A2(n16179), .ZN(n16184) );
  NAND2_X1 U16993 ( .A1(n16180), .A2(n16184), .ZN(n13840) );
  INV_X1 U16994 ( .A(n16138), .ZN(n16128) );
  AOI22_X1 U16995 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13840), .B1(
        n16128), .B2(n13841), .ZN(n13628) );
  XNOR2_X1 U16996 ( .A(n16173), .B(n16160), .ZN(n20040) );
  AND2_X1 U16997 ( .A1(n20149), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n13649) );
  AOI21_X1 U16998 ( .B1(n20040), .B2(n20169), .A(n13649), .ZN(n13627) );
  OAI211_X1 U16999 ( .C1(n13653), .C2(n20176), .A(n13628), .B(n13627), .ZN(
        P1_U3025) );
  NAND2_X1 U17000 ( .A1(n13630), .A2(n13629), .ZN(n13632) );
  INV_X1 U17001 ( .A(n13677), .ZN(n13639) );
  OAI21_X1 U17002 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13638) );
  NAND3_X1 U17003 ( .A1(n13639), .A2(n14961), .A3(n13638), .ZN(n13644) );
  OR2_X1 U17004 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  AND2_X1 U17005 ( .A1(n13642), .A2(n13673), .ZN(n19117) );
  NAND2_X1 U17006 ( .A1(n15000), .A2(n19117), .ZN(n13643) );
  OAI211_X1 U17007 ( .C1(n15000), .C2(n11124), .A(n13644), .B(n13643), .ZN(
        P2_U2875) );
  AOI21_X1 U17008 ( .B1(n13645), .B2(n13560), .A(n13612), .ZN(n20048) );
  INV_X1 U17009 ( .A(n20048), .ZN(n13656) );
  AOI22_X1 U17010 ( .A1(n20040), .A2(n20088), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14537), .ZN(n13646) );
  OAI21_X1 U17011 ( .B1(n13656), .B2(n14539), .A(n13646), .ZN(P1_U2866) );
  OAI21_X1 U17012 ( .B1(n13648), .B2(n13647), .A(n16367), .ZN(n15428) );
  INV_X1 U17013 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19256) );
  OAI222_X1 U17014 ( .A1(n13834), .A2(n15017), .B1(n15428), .B2(n19239), .C1(
        n19256), .C2(n19249), .ZN(P2_U2906) );
  AOI21_X1 U17015 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13649), .ZN(n13650) );
  OAI21_X1 U17016 ( .B1(n20041), .B2(n20141), .A(n13650), .ZN(n13651) );
  AOI21_X1 U17017 ( .B1(n20048), .B2(n20178), .A(n13651), .ZN(n13652) );
  OAI21_X1 U17018 ( .B1(n20155), .B2(n13653), .A(n13652), .ZN(P1_U2993) );
  INV_X1 U17019 ( .A(DATAI_6_), .ZN(n13655) );
  NAND2_X1 U17020 ( .A1(n20177), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13654) );
  OAI21_X1 U17021 ( .B1(n20177), .B2(n13655), .A(n13654), .ZN(n14572) );
  INV_X1 U17022 ( .A(n14572), .ZN(n20221) );
  OAI222_X1 U17023 ( .A1(n13656), .A2(n14622), .B1(n14604), .B2(n20221), .C1(
        n14602), .C2(n11870), .ZN(P1_U2898) );
  XOR2_X1 U17024 ( .A(n13658), .B(n13657), .Z(n19292) );
  INV_X1 U17025 ( .A(n19292), .ZN(n13672) );
  NAND2_X1 U17026 ( .A1(n13660), .A2(n13659), .ZN(n13661) );
  XNOR2_X1 U17027 ( .A(n13661), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19288) );
  NAND2_X1 U17028 ( .A1(n13662), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13967) );
  OAI21_X1 U17029 ( .B1(n13664), .B2(n13663), .A(n13297), .ZN(n19173) );
  INV_X1 U17030 ( .A(n19173), .ZN(n19289) );
  NAND2_X1 U17031 ( .A1(n19289), .A2(n16390), .ZN(n13669) );
  OAI21_X1 U17032 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16410), .A(
        n13989), .ZN(n13966) );
  INV_X1 U17033 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19896) );
  NOR2_X1 U17034 ( .A1(n19896), .A2(n19170), .ZN(n13667) );
  NOR2_X1 U17035 ( .A1(n16400), .A2(n13665), .ZN(n13666) );
  AOI211_X1 U17036 ( .C1(n13966), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13667), .B(n13666), .ZN(n13668) );
  OAI211_X1 U17037 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13967), .A(
        n13669), .B(n13668), .ZN(n13670) );
  AOI21_X1 U17038 ( .B1(n19288), .B2(n16388), .A(n13670), .ZN(n13671) );
  OAI21_X1 U17039 ( .B1(n13672), .B2(n19300), .A(n13671), .ZN(P2_U3042) );
  AOI21_X1 U17040 ( .B1(n13674), .B2(n13673), .A(n10347), .ZN(n16308) );
  INV_X1 U17041 ( .A(n16308), .ZN(n13680) );
  INV_X1 U17042 ( .A(n13723), .ZN(n13675) );
  OAI211_X1 U17043 ( .C1(n13677), .C2(n13676), .A(n13675), .B(n14961), .ZN(
        n13679) );
  NAND2_X1 U17044 ( .A1(n15010), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13678) );
  OAI211_X1 U17045 ( .C1(n13680), .C2(n15010), .A(n13679), .B(n13678), .ZN(
        P2_U2874) );
  NOR2_X1 U17046 ( .A1(n19165), .A2(n13681), .ZN(n13682) );
  XNOR2_X1 U17047 ( .A(n13682), .B(n16353), .ZN(n13689) );
  INV_X1 U17048 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19900) );
  OAI21_X1 U17049 ( .B1(n19900), .B2(n19179), .A(n19170), .ZN(n13685) );
  OAI22_X1 U17050 ( .A1(n19202), .A2(n13368), .B1(n13683), .B2(n19141), .ZN(
        n13684) );
  AOI211_X1 U17051 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19167), .A(
        n13685), .B(n13684), .ZN(n13687) );
  NAND2_X1 U17052 ( .A1(n19185), .A2(n16348), .ZN(n13686) );
  OAI211_X1 U17053 ( .C1(n13965), .C2(n19158), .A(n13687), .B(n13686), .ZN(
        n13688) );
  AOI21_X1 U17054 ( .B1(n13689), .B2(n19108), .A(n13688), .ZN(n13690) );
  INV_X1 U17055 ( .A(n13690), .ZN(P2_U2849) );
  NOR2_X1 U17056 ( .A1(n19165), .A2(n13691), .ZN(n13692) );
  XNOR2_X1 U17057 ( .A(n13692), .B(n16327), .ZN(n13699) );
  INV_X1 U17058 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19908) );
  OAI21_X1 U17059 ( .B1(n19908), .B2(n19179), .A(n19170), .ZN(n13695) );
  OAI22_X1 U17060 ( .A1(n19202), .A2(n11118), .B1(n13693), .B2(n19141), .ZN(
        n13694) );
  AOI211_X1 U17061 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19167), .A(
        n13695), .B(n13694), .ZN(n13697) );
  NAND2_X1 U17062 ( .A1(n19185), .A2(n16323), .ZN(n13696) );
  OAI211_X1 U17063 ( .C1(n15476), .C2(n19158), .A(n13697), .B(n13696), .ZN(
        n13698) );
  AOI21_X1 U17064 ( .B1(n13699), .B2(n19108), .A(n13698), .ZN(n13700) );
  INV_X1 U17065 ( .A(n13700), .ZN(P2_U2845) );
  NAND2_X1 U17066 ( .A1(n19152), .A2(n13701), .ZN(n13702) );
  XNOR2_X1 U17067 ( .A(n16328), .B(n13702), .ZN(n13709) );
  INV_X1 U17068 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U17069 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n19183), .B1(n19205), .B2(
        n13703), .ZN(n13704) );
  OAI211_X1 U17070 ( .C1(n19906), .C2(n19179), .A(n13704), .B(n19170), .ZN(
        n13705) );
  AOI21_X1 U17071 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19167), .A(
        n13705), .ZN(n13707) );
  NAND2_X1 U17072 ( .A1(n19185), .A2(n16332), .ZN(n13706) );
  OAI211_X1 U17073 ( .C1(n15491), .C2(n19158), .A(n13707), .B(n13706), .ZN(
        n13708) );
  AOI21_X1 U17074 ( .B1(n13709), .B2(n19108), .A(n13708), .ZN(n13710) );
  INV_X1 U17075 ( .A(n13710), .ZN(P2_U2846) );
  NAND2_X1 U17076 ( .A1(n19152), .A2(n13711), .ZN(n13712) );
  XNOR2_X1 U17077 ( .A(n14035), .B(n13712), .ZN(n13721) );
  NAND2_X1 U17078 ( .A1(n19963), .A2(n19213), .ZN(n13718) );
  OAI22_X1 U17079 ( .A1(n19202), .A2(n13714), .B1(n13713), .B2(n19141), .ZN(
        n13716) );
  OAI22_X1 U17080 ( .A1(n14033), .A2(n19210), .B1(n19894), .B2(n19179), .ZN(
        n13715) );
  AOI211_X1 U17081 ( .C1(n19185), .C2(n15545), .A(n13716), .B(n13715), .ZN(
        n13717) );
  OAI211_X1 U17082 ( .C1(n13719), .C2(n19158), .A(n13718), .B(n13717), .ZN(
        n13720) );
  AOI21_X1 U17083 ( .B1(n13721), .B2(n19108), .A(n13720), .ZN(n13722) );
  INV_X1 U17084 ( .A(n13722), .ZN(P2_U2852) );
  OAI211_X1 U17085 ( .C1(n13723), .C2(n13724), .A(n13806), .B(n14961), .ZN(
        n13729) );
  AND2_X1 U17086 ( .A1(n13726), .A2(n13725), .ZN(n13727) );
  OR2_X1 U17087 ( .A1(n13727), .A2(n13804), .ZN(n19112) );
  NAND2_X1 U17088 ( .A1(n15000), .A2(n16371), .ZN(n13728) );
  OAI211_X1 U17089 ( .C1(n14983), .C2(n11136), .A(n13729), .B(n13728), .ZN(
        P2_U2873) );
  NAND2_X1 U17090 ( .A1(n13614), .A2(n13731), .ZN(n13732) );
  NAND2_X1 U17091 ( .A1(n13730), .A2(n13732), .ZN(n13863) );
  AOI22_X1 U17092 ( .A1(n14620), .A2(n14567), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14618), .ZN(n13733) );
  OAI21_X1 U17093 ( .B1(n13863), .B2(n14622), .A(n13733), .ZN(P1_U2896) );
  AOI21_X1 U17094 ( .B1(n13734), .B2(n20077), .A(n20030), .ZN(n14488) );
  INV_X1 U17095 ( .A(n14488), .ZN(n13746) );
  NAND2_X1 U17096 ( .A1(n20077), .A2(n13735), .ZN(n13939) );
  NAND2_X1 U17097 ( .A1(n13839), .A2(n13939), .ZN(n13745) );
  OR2_X1 U17098 ( .A1(n16162), .A2(n13736), .ZN(n13737) );
  AND2_X1 U17099 ( .A1(n13883), .A2(n13737), .ZN(n13844) );
  NAND2_X1 U17100 ( .A1(n13844), .A2(n20070), .ZN(n13743) );
  OAI21_X1 U17101 ( .B1(n20057), .B2(n13739), .A(n20055), .ZN(n13741) );
  NOR2_X1 U17102 ( .A1(n20059), .A2(n13858), .ZN(n13740) );
  NOR2_X1 U17103 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  OAI211_X1 U17104 ( .C1(n14471), .C2(n10164), .A(n13743), .B(n13742), .ZN(
        n13744) );
  AOI21_X1 U17105 ( .B1(n13746), .B2(n13745), .A(n13744), .ZN(n13747) );
  OAI21_X1 U17106 ( .B1(n13863), .B2(n15978), .A(n13747), .ZN(P1_U2832) );
  AOI22_X1 U17107 ( .A1(n20135), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20134), .ZN(n13749) );
  INV_X1 U17108 ( .A(n20215), .ZN(n14575) );
  NAND2_X1 U17109 ( .A1(n13766), .A2(n14575), .ZN(n13758) );
  NAND2_X1 U17110 ( .A1(n13749), .A2(n13758), .ZN(P1_U2942) );
  AOI22_X1 U17111 ( .A1(n20135), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20134), .ZN(n13750) );
  INV_X1 U17112 ( .A(n20206), .ZN(n14582) );
  NAND2_X1 U17113 ( .A1(n13766), .A2(n14582), .ZN(n13764) );
  NAND2_X1 U17114 ( .A1(n13750), .A2(n13764), .ZN(P1_U2940) );
  AOI22_X1 U17115 ( .A1(n20135), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20134), .ZN(n13752) );
  NAND2_X1 U17116 ( .A1(n13752), .A2(n13751), .ZN(P1_U2945) );
  AOI22_X1 U17117 ( .A1(n20135), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20134), .ZN(n13753) );
  INV_X1 U17118 ( .A(n20210), .ZN(n14578) );
  NAND2_X1 U17119 ( .A1(n13766), .A2(n14578), .ZN(n13760) );
  NAND2_X1 U17120 ( .A1(n13753), .A2(n13760), .ZN(P1_U2941) );
  AOI22_X1 U17121 ( .A1(n20135), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20134), .ZN(n13754) );
  NAND2_X1 U17122 ( .A1(n13766), .A2(n14572), .ZN(n13768) );
  NAND2_X1 U17123 ( .A1(n13754), .A2(n13768), .ZN(P1_U2943) );
  AOI22_X1 U17124 ( .A1(n20135), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20134), .ZN(n13755) );
  INV_X1 U17125 ( .A(n20201), .ZN(n14586) );
  NAND2_X1 U17126 ( .A1(n13766), .A2(n14586), .ZN(n13762) );
  NAND2_X1 U17127 ( .A1(n13755), .A2(n13762), .ZN(P1_U2954) );
  AOI22_X1 U17128 ( .A1(n20135), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20134), .ZN(n13756) );
  NAND2_X1 U17129 ( .A1(n13766), .A2(n20229), .ZN(n13770) );
  NAND2_X1 U17130 ( .A1(n13756), .A2(n13770), .ZN(P1_U2944) );
  AOI22_X1 U17131 ( .A1(n20135), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20134), .ZN(n13757) );
  INV_X1 U17132 ( .A(n20187), .ZN(n14594) );
  NAND2_X1 U17133 ( .A1(n13766), .A2(n14594), .ZN(n13774) );
  NAND2_X1 U17134 ( .A1(n13757), .A2(n13774), .ZN(P1_U2952) );
  AOI22_X1 U17135 ( .A1(n20135), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20134), .ZN(n13759) );
  NAND2_X1 U17136 ( .A1(n13759), .A2(n13758), .ZN(P1_U2957) );
  AOI22_X1 U17137 ( .A1(n20135), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20134), .ZN(n13761) );
  NAND2_X1 U17138 ( .A1(n13761), .A2(n13760), .ZN(P1_U2956) );
  AOI22_X1 U17139 ( .A1(n20135), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20134), .ZN(n13763) );
  NAND2_X1 U17140 ( .A1(n13763), .A2(n13762), .ZN(P1_U2939) );
  AOI22_X1 U17141 ( .A1(n20135), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20134), .ZN(n13765) );
  NAND2_X1 U17142 ( .A1(n13765), .A2(n13764), .ZN(P1_U2955) );
  AOI22_X1 U17143 ( .A1(n20135), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20134), .ZN(n13767) );
  INV_X1 U17144 ( .A(n20196), .ZN(n14589) );
  NAND2_X1 U17145 ( .A1(n13766), .A2(n14589), .ZN(n13772) );
  NAND2_X1 U17146 ( .A1(n13767), .A2(n13772), .ZN(P1_U2938) );
  AOI22_X1 U17147 ( .A1(n20135), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20134), .ZN(n13769) );
  NAND2_X1 U17148 ( .A1(n13769), .A2(n13768), .ZN(P1_U2958) );
  AOI22_X1 U17149 ( .A1(n20135), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20134), .ZN(n13771) );
  NAND2_X1 U17150 ( .A1(n13771), .A2(n13770), .ZN(P1_U2959) );
  AOI22_X1 U17151 ( .A1(n20135), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20134), .ZN(n13773) );
  NAND2_X1 U17152 ( .A1(n13773), .A2(n13772), .ZN(P1_U2953) );
  AOI22_X1 U17153 ( .A1(n20135), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20134), .ZN(n13775) );
  NAND2_X1 U17154 ( .A1(n13775), .A2(n13774), .ZN(P1_U2937) );
  INV_X1 U17155 ( .A(n13844), .ZN(n13776) );
  OAI222_X1 U17156 ( .A1(n13863), .A2(n14539), .B1(n20092), .B2(n10164), .C1(
        n13776), .C2(n14546), .ZN(P1_U2864) );
  OAI21_X1 U17157 ( .B1(n13779), .B2(n13777), .A(n15978), .ZN(n20076) );
  INV_X1 U17158 ( .A(n20076), .ZN(n14503) );
  NOR2_X1 U17159 ( .A1(n13779), .A2(n13778), .ZN(n20071) );
  INV_X1 U17160 ( .A(n20071), .ZN(n13788) );
  AOI22_X1 U17161 ( .A1(n20070), .A2(n13780), .B1(n20043), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13787) );
  NAND2_X1 U17162 ( .A1(n20030), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13781) );
  OAI21_X1 U17163 ( .B1(n20059), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13781), .ZN(n13782) );
  INV_X1 U17164 ( .A(n13782), .ZN(n13784) );
  NAND2_X1 U17165 ( .A1(n20069), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13783) );
  OAI211_X1 U17166 ( .C1(n20032), .C2(P1_REIP_REG_1__SCAN_IN), .A(n13784), .B(
        n13783), .ZN(n13785) );
  INV_X1 U17167 ( .A(n13785), .ZN(n13786) );
  OAI211_X1 U17168 ( .C1(n20586), .C2(n13788), .A(n13787), .B(n13786), .ZN(
        n13789) );
  INV_X1 U17169 ( .A(n13789), .ZN(n13790) );
  OAI21_X1 U17170 ( .B1(n20143), .B2(n14503), .A(n13790), .ZN(P1_U2839) );
  NAND2_X1 U17171 ( .A1(n19152), .A2(n13791), .ZN(n13792) );
  XNOR2_X1 U17172 ( .A(n16354), .B(n13792), .ZN(n13801) );
  OAI21_X1 U17173 ( .B1(n9916), .B2(n13794), .A(n13793), .ZN(n19238) );
  INV_X1 U17174 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19898) );
  OAI21_X1 U17175 ( .B1(n19898), .B2(n19179), .A(n19170), .ZN(n13797) );
  OAI22_X1 U17176 ( .A1(n13795), .A2(n19141), .B1(n16364), .B2(n19210), .ZN(
        n13796) );
  AOI211_X1 U17177 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19183), .A(n13797), .B(
        n13796), .ZN(n13799) );
  NAND2_X1 U17178 ( .A1(n19185), .A2(n16361), .ZN(n13798) );
  OAI211_X1 U17179 ( .C1(n19238), .C2(n19158), .A(n13799), .B(n13798), .ZN(
        n13800) );
  AOI21_X1 U17180 ( .B1(n13801), .B2(n19108), .A(n13800), .ZN(n13802) );
  INV_X1 U17181 ( .A(n13802), .ZN(P2_U2850) );
  OR2_X1 U17182 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  NAND2_X1 U17183 ( .A1(n13910), .A2(n13805), .ZN(n15410) );
  INV_X1 U17184 ( .A(n13806), .ZN(n13810) );
  INV_X1 U17185 ( .A(n13907), .ZN(n13904) );
  OAI211_X1 U17186 ( .C1(n13810), .C2(n13809), .A(n14961), .B(n13904), .ZN(
        n13812) );
  NAND2_X1 U17187 ( .A1(n13301), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13811) );
  OAI211_X1 U17188 ( .C1(n15410), .C2(n15010), .A(n13812), .B(n13811), .ZN(
        P2_U2872) );
  NAND2_X1 U17189 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13813) );
  NAND2_X1 U17190 ( .A1(n20077), .A2(n13813), .ZN(n13822) );
  NAND2_X1 U17191 ( .A1(n13822), .A2(n13814), .ZN(n20075) );
  INV_X1 U17192 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20867) );
  OAI22_X1 U17193 ( .A1(n13816), .A2(n20059), .B1(n20057), .B2(n13815), .ZN(
        n13817) );
  AOI21_X1 U17194 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(n20043), .A(n13817), .ZN(
        n13821) );
  INV_X1 U17195 ( .A(n13818), .ZN(n13819) );
  NAND2_X1 U17196 ( .A1(n20070), .A2(n13819), .ZN(n13820) );
  OAI211_X1 U17197 ( .C1(n13822), .C2(n20867), .A(n13821), .B(n13820), .ZN(
        n13823) );
  AOI21_X1 U17198 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n20075), .A(n13823), .ZN(
        n13825) );
  INV_X1 U17199 ( .A(n13398), .ZN(n20459) );
  NAND2_X1 U17200 ( .A1(n20459), .A2(n20071), .ZN(n13824) );
  OAI211_X1 U17201 ( .C1(n13826), .C2(n14503), .A(n13825), .B(n13824), .ZN(
        P1_U2838) );
  NAND2_X1 U17202 ( .A1(n20057), .A2(n20059), .ZN(n13827) );
  AOI22_X1 U17203 ( .A1(n20043), .A2(P1_EBX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13827), .ZN(n13829) );
  NAND2_X1 U17204 ( .A1(n20029), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13828) );
  OAI211_X1 U17205 ( .C1(n20166), .C2(n15963), .A(n13829), .B(n13828), .ZN(
        n13830) );
  AOI21_X1 U17206 ( .B1(n20861), .B2(n20071), .A(n13830), .ZN(n13831) );
  OAI21_X1 U17207 ( .B1(n20148), .B2(n14503), .A(n13831), .ZN(P1_U2840) );
  OAI21_X1 U17208 ( .B1(n16366), .B2(n13832), .A(n13923), .ZN(n15408) );
  INV_X1 U17209 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19252) );
  OAI222_X1 U17210 ( .A1(n13834), .A2(n13833), .B1(n15408), .B2(n19239), .C1(
        n19252), .C2(n19249), .ZN(P2_U2904) );
  XNOR2_X1 U17211 ( .A(n13836), .B(n13835), .ZN(n13837) );
  XNOR2_X1 U17212 ( .A(n13838), .B(n13837), .ZN(n13857) );
  INV_X1 U17213 ( .A(n13857), .ZN(n13846) );
  INV_X1 U17214 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13839) );
  NOR2_X1 U17215 ( .A1(n20140), .A2(n13839), .ZN(n13860) );
  NOR2_X1 U17216 ( .A1(n13841), .A2(n16138), .ZN(n16164) );
  OAI21_X1 U17217 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16164), .ZN(n13842) );
  AOI21_X1 U17218 ( .B1(n13841), .B2(n20157), .A(n13840), .ZN(n16169) );
  OAI22_X1 U17219 ( .A1(n16143), .A2(n13842), .B1(n16169), .B2(n13835), .ZN(
        n13843) );
  AOI211_X1 U17220 ( .C1(n20169), .C2(n13844), .A(n13860), .B(n13843), .ZN(
        n13845) );
  OAI21_X1 U17221 ( .B1(n13846), .B2(n20176), .A(n13845), .ZN(P1_U3023) );
  NAND2_X1 U17222 ( .A1(n19152), .A2(n13847), .ZN(n13848) );
  XNOR2_X1 U17223 ( .A(n16304), .B(n13848), .ZN(n13849) );
  NAND2_X1 U17224 ( .A1(n13849), .A2(n19108), .ZN(n13856) );
  NAND2_X1 U17225 ( .A1(n19197), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13850) );
  OAI211_X1 U17226 ( .C1(n19158), .C2(n15428), .A(n13850), .B(n19170), .ZN(
        n13854) );
  AOI22_X1 U17227 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19183), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19167), .ZN(n13851) );
  OAI21_X1 U17228 ( .B1(n13852), .B2(n19141), .A(n13851), .ZN(n13853) );
  AOI211_X1 U17229 ( .C1(n16308), .C2(n19185), .A(n13854), .B(n13853), .ZN(
        n13855) );
  NAND2_X1 U17230 ( .A1(n13856), .A2(n13855), .ZN(P2_U2842) );
  INV_X1 U17231 ( .A(n20155), .ZN(n16045) );
  NAND2_X1 U17232 ( .A1(n13857), .A2(n16045), .ZN(n13862) );
  NOR2_X1 U17233 ( .A1(n20141), .A2(n13858), .ZN(n13859) );
  AOI211_X1 U17234 ( .C1(n20152), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13860), .B(n13859), .ZN(n13861) );
  OAI211_X1 U17235 ( .C1(n20142), .C2(n13863), .A(n13862), .B(n13861), .ZN(
        P1_U2991) );
  AOI21_X1 U17236 ( .B1(n13864), .B2(n13730), .A(n13916), .ZN(n14490) );
  INV_X1 U17237 ( .A(n14490), .ZN(n13885) );
  AOI22_X1 U17238 ( .A1(n14620), .A2(n14560), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14618), .ZN(n13865) );
  OAI21_X1 U17239 ( .B1(n13885), .B2(n14622), .A(n13865), .ZN(P1_U2895) );
  XNOR2_X1 U17240 ( .A(n13867), .B(n13866), .ZN(n16357) );
  AND2_X1 U17241 ( .A1(n13868), .A2(n10860), .ZN(n13869) );
  INV_X1 U17242 ( .A(n16359), .ZN(n13880) );
  NOR2_X1 U17243 ( .A1(n19898), .A2(n19170), .ZN(n13876) );
  AOI211_X1 U17244 ( .C1(n13874), .C2(n13873), .A(n13872), .B(n13967), .ZN(
        n13875) );
  AOI211_X1 U17245 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13966), .A(
        n13876), .B(n13875), .ZN(n13878) );
  NAND2_X1 U17246 ( .A1(n16390), .A2(n16361), .ZN(n13877) );
  OAI211_X1 U17247 ( .C1(n19238), .C2(n16400), .A(n13878), .B(n13877), .ZN(
        n13879) );
  AOI21_X1 U17248 ( .B1(n13880), .B2(n16388), .A(n13879), .ZN(n13881) );
  OAI21_X1 U17249 ( .B1(n19300), .B2(n16357), .A(n13881), .ZN(P2_U3041) );
  NAND2_X1 U17250 ( .A1(n13883), .A2(n13882), .ZN(n13884) );
  NAND2_X1 U17251 ( .A1(n13918), .A2(n13884), .ZN(n16152) );
  OAI222_X1 U17252 ( .A1(n13885), .A2(n14539), .B1(n21227), .B2(n20092), .C1(
        n16152), .C2(n14546), .ZN(P1_U2863) );
  NOR2_X1 U17253 ( .A1(n10155), .A2(n13887), .ZN(n13888) );
  XNOR2_X1 U17254 ( .A(n13889), .B(n13888), .ZN(n16149) );
  AOI22_X1 U17255 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13890) );
  OAI21_X1 U17256 ( .B1(n20141), .B2(n13891), .A(n13890), .ZN(n13892) );
  AOI21_X1 U17257 ( .B1(n14490), .B2(n20178), .A(n13892), .ZN(n13893) );
  OAI21_X1 U17258 ( .B1(n16149), .B2(n20155), .A(n13893), .ZN(P1_U2990) );
  AOI22_X1 U17259 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17260 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17261 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17262 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13894) );
  NAND4_X1 U17263 ( .A1(n13897), .A2(n13896), .A3(n13895), .A4(n13894), .ZN(
        n13903) );
  AOI22_X1 U17264 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17265 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17266 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U17267 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13898) );
  NAND4_X1 U17268 ( .A1(n13901), .A2(n13900), .A3(n13899), .A4(n13898), .ZN(
        n13902) );
  NOR2_X1 U17269 ( .A1(n13903), .A2(n13902), .ZN(n13905) );
  AND2_X1 U17270 ( .A1(n13904), .A2(n13905), .ZN(n13908) );
  INV_X1 U17271 ( .A(n13905), .ZN(n13906) );
  OR2_X1 U17272 ( .A1(n13908), .A2(n13955), .ZN(n13937) );
  NAND2_X1 U17273 ( .A1(n13910), .A2(n13909), .ZN(n13911) );
  AND2_X1 U17274 ( .A1(n13958), .A2(n13911), .ZN(n19097) );
  NOR2_X1 U17275 ( .A1(n15000), .A2(n13912), .ZN(n13913) );
  AOI21_X1 U17276 ( .B1(n19097), .B2(n15000), .A(n13913), .ZN(n13914) );
  OAI21_X1 U17277 ( .B1(n13937), .B2(n15012), .A(n13914), .ZN(P2_U2871) );
  XOR2_X1 U17278 ( .A(n13916), .B(n13915), .Z(n14006) );
  NAND2_X1 U17279 ( .A1(n13918), .A2(n13917), .ZN(n13919) );
  NAND2_X1 U17280 ( .A1(n15972), .A2(n13919), .ZN(n16144) );
  OAI22_X1 U17281 ( .A1(n16144), .A2(n14546), .B1(n20979), .B2(n20092), .ZN(
        n13920) );
  AOI21_X1 U17282 ( .B1(n14006), .B2(n20089), .A(n13920), .ZN(n13921) );
  INV_X1 U17283 ( .A(n13921), .ZN(P1_U2862) );
  AND2_X1 U17284 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  OR2_X1 U17285 ( .A1(n13924), .A2(n14885), .ZN(n15403) );
  INV_X1 U17286 ( .A(n15403), .ZN(n19098) );
  AND2_X1 U17287 ( .A1(n13926), .A2(n13925), .ZN(n13927) );
  INV_X1 U17288 ( .A(n16286), .ZN(n15110) );
  OAI22_X1 U17289 ( .A1(n15110), .A2(n19322), .B1(n19249), .B2(n13928), .ZN(
        n13935) );
  INV_X1 U17290 ( .A(n19215), .ZN(n15114) );
  INV_X1 U17291 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n13933) );
  INV_X1 U17292 ( .A(n19217), .ZN(n15112) );
  INV_X1 U17293 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n13932) );
  OAI22_X1 U17294 ( .A1(n15114), .A2(n13933), .B1(n15112), .B2(n13932), .ZN(
        n13934) );
  AOI211_X1 U17295 ( .C1(n19098), .C2(n19245), .A(n13935), .B(n13934), .ZN(
        n13936) );
  OAI21_X1 U17296 ( .B1(n15120), .B2(n13937), .A(n13936), .ZN(P2_U2903) );
  INV_X1 U17297 ( .A(n14006), .ZN(n14000) );
  INV_X1 U17298 ( .A(n14004), .ZN(n13938) );
  AOI22_X1 U17299 ( .A1(n13938), .A2(n20073), .B1(n20069), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13941) );
  INV_X1 U17300 ( .A(n20029), .ZN(n15930) );
  OAI21_X1 U17301 ( .B1(n14421), .B2(n15930), .A(n14488), .ZN(n15950) );
  OAI221_X1 U17302 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n14479), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(P1_REIP_REG_9__SCAN_IN), .A(n15950), 
        .ZN(n13940) );
  NAND3_X1 U17303 ( .A1(n13941), .A2(n13940), .A3(n20055), .ZN(n13943) );
  NOR2_X1 U17304 ( .A1(n16144), .A2(n15963), .ZN(n13942) );
  AOI211_X1 U17305 ( .C1(n20043), .C2(P1_EBX_REG_10__SCAN_IN), .A(n13943), .B(
        n13942), .ZN(n13944) );
  OAI21_X1 U17306 ( .B1(n14000), .B2(n15978), .A(n13944), .ZN(P1_U2830) );
  AOI22_X1 U17307 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U17308 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U17309 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13946) );
  AOI22_X1 U17310 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10762), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13945) );
  NAND4_X1 U17311 ( .A1(n13948), .A2(n13947), .A3(n13946), .A4(n13945), .ZN(
        n13954) );
  AOI22_X1 U17312 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17313 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17314 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13950) );
  AOI22_X1 U17315 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n14108), .ZN(n13949) );
  NAND4_X1 U17316 ( .A1(n13952), .A2(n13951), .A3(n13950), .A4(n13949), .ZN(
        n13953) );
  OAI21_X1 U17317 ( .B1(n13955), .B2(n13956), .A(n14049), .ZN(n15119) );
  AND2_X1 U17318 ( .A1(n13958), .A2(n13957), .ZN(n13959) );
  OR2_X1 U17319 ( .A1(n13959), .A2(n15006), .ZN(n15391) );
  MUX2_X1 U17320 ( .A(n15391), .B(n11146), .S(n15010), .Z(n13960) );
  OAI21_X1 U17321 ( .B1(n15119), .B2(n15012), .A(n13960), .ZN(P2_U2870) );
  OAI21_X1 U17322 ( .B1(n13961), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13962), .ZN(n16347) );
  XOR2_X1 U17323 ( .A(n13964), .B(n13963), .Z(n16349) );
  NOR2_X1 U17324 ( .A1(n13965), .A2(n16400), .ZN(n13976) );
  AOI21_X1 U17325 ( .B1(n19302), .B2(n13968), .A(n13966), .ZN(n13974) );
  NOR3_X1 U17326 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13968), .A3(
        n13967), .ZN(n13971) );
  NOR2_X1 U17327 ( .A1(n19305), .A2(n13969), .ZN(n13970) );
  AOI211_X1 U17328 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19286), .A(n13971), .B(
        n13970), .ZN(n13972) );
  OAI21_X1 U17329 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13975) );
  AOI211_X1 U17330 ( .C1(n16349), .C2(n16391), .A(n13976), .B(n13975), .ZN(
        n13977) );
  OAI21_X1 U17331 ( .B1(n19311), .B2(n16347), .A(n13977), .ZN(P2_U3040) );
  NOR2_X1 U17332 ( .A1(n10371), .A2(n13980), .ZN(n13981) );
  XNOR2_X1 U17333 ( .A(n13978), .B(n13981), .ZN(n13999) );
  NAND2_X1 U17334 ( .A1(n16340), .A2(n16338), .ZN(n13983) );
  XNOR2_X1 U17335 ( .A(n13982), .B(n13983), .ZN(n13996) );
  OAI22_X1 U17336 ( .A1(n16365), .A2(n13984), .B1(n19902), .B2(n19170), .ZN(
        n13985) );
  AOI21_X1 U17337 ( .B1(n16355), .B2(n19153), .A(n13985), .ZN(n13986) );
  OAI21_X1 U17338 ( .B1(n15258), .B2(n19157), .A(n13986), .ZN(n13987) );
  AOI21_X1 U17339 ( .B1(n13996), .B2(n19291), .A(n13987), .ZN(n13988) );
  OAI21_X1 U17340 ( .B1(n13999), .B2(n16358), .A(n13988), .ZN(P2_U3007) );
  OAI21_X1 U17341 ( .B1(n16410), .B2(n13990), .A(n13989), .ZN(n16386) );
  INV_X1 U17342 ( .A(n13991), .ZN(n16394) );
  AOI22_X1 U17343 ( .A1(n19286), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n13992), 
        .B2(n16394), .ZN(n13993) );
  OAI21_X1 U17344 ( .B1(n19305), .B2(n19157), .A(n13993), .ZN(n13995) );
  NOR2_X1 U17345 ( .A1(n19159), .A2(n16400), .ZN(n13994) );
  AOI211_X1 U17346 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16386), .A(
        n13995), .B(n13994), .ZN(n13998) );
  NAND2_X1 U17347 ( .A1(n13996), .A2(n16391), .ZN(n13997) );
  OAI211_X1 U17348 ( .C1(n13999), .C2(n19311), .A(n13998), .B(n13997), .ZN(
        P2_U3039) );
  INV_X1 U17349 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14001) );
  OAI222_X1 U17350 ( .A1(n14602), .A2(n14001), .B1(n14604), .B2(n14555), .C1(
        n14622), .C2(n14000), .ZN(P1_U2894) );
  MUX2_X1 U17351 ( .A(n16025), .B(n16026), .S(n10154), .Z(n14002) );
  XOR2_X1 U17352 ( .A(n12685), .B(n14002), .Z(n16147) );
  INV_X1 U17353 ( .A(n16147), .ZN(n14008) );
  AOI22_X1 U17354 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14003) );
  OAI21_X1 U17355 ( .B1(n14004), .B2(n20141), .A(n14003), .ZN(n14005) );
  AOI21_X1 U17356 ( .B1(n14006), .B2(n20178), .A(n14005), .ZN(n14007) );
  OAI21_X1 U17357 ( .B1(n14008), .B2(n20155), .A(n14007), .ZN(P1_U2989) );
  INV_X1 U17358 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18863) );
  OAI21_X1 U17359 ( .B1(n15645), .B2(n18999), .A(n18863), .ZN(n14009) );
  NAND2_X1 U17360 ( .A1(n14010), .A2(n14009), .ZN(n18814) );
  NOR2_X1 U17361 ( .A1(n18979), .A2(n18814), .ZN(n14028) );
  NAND2_X1 U17362 ( .A1(n18877), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18344) );
  NAND2_X1 U17363 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  INV_X1 U17364 ( .A(n15784), .ZN(n14016) );
  AOI211_X1 U17365 ( .C1(n14017), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        n15783) );
  AOI21_X1 U17366 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19006), .A(
        n14018), .ZN(n15770) );
  AND2_X1 U17367 ( .A1(n14020), .A2(n14019), .ZN(n14023) );
  NAND2_X1 U17368 ( .A1(n14022), .A2(n14021), .ZN(n15769) );
  NAND2_X1 U17369 ( .A1(n15767), .A2(n18812), .ZN(n15548) );
  NAND4_X1 U17370 ( .A1(n18806), .A2(n14025), .A3(n15775), .A4(n19026), .ZN(
        n14026) );
  NAND4_X1 U17371 ( .A1(n15783), .A2(n15548), .A3(n15917), .A4(n14026), .ZN(
        n18840) );
  NOR3_X1 U17372 ( .A1(n18877), .A2(n18869), .A3(n18985), .ZN(n18972) );
  AOI22_X1 U17373 ( .A1(n18840), .A2(n19020), .B1(P3_FLUSH_REG_SCAN_IN), .B2(
        n18972), .ZN(n14027) );
  NAND2_X1 U17374 ( .A1(n18344), .A2(n14027), .ZN(n19004) );
  MUX2_X1 U17375 ( .A(n14028), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19007), .Z(P3_U3284) );
  INV_X1 U17376 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14029) );
  OAI222_X1 U17377 ( .A1(n14539), .A2(n14048), .B1(n14029), .B2(n20092), .C1(
        n14750), .C2(n14546), .ZN(P1_U2842) );
  MUX2_X1 U17378 ( .A(n14305), .B(n14907), .S(n15010), .Z(n14030) );
  OAI21_X1 U17379 ( .B1(n19969), .B2(n15012), .A(n14030), .ZN(P2_U2885) );
  NOR2_X1 U17380 ( .A1(n14031), .A2(n16356), .ZN(n14039) );
  NAND2_X1 U17381 ( .A1(n14032), .A2(n10925), .ZN(n14037) );
  OAI22_X1 U17382 ( .A1(n16365), .A2(n14033), .B1(n19894), .B2(n19170), .ZN(
        n14034) );
  AOI21_X1 U17383 ( .B1(n16355), .B2(n14035), .A(n14034), .ZN(n14036) );
  OAI211_X1 U17384 ( .C1(n13340), .C2(n15258), .A(n14037), .B(n14036), .ZN(
        n14038) );
  OR2_X1 U17385 ( .A1(n14039), .A2(n14038), .ZN(P2_U3011) );
  MUX2_X1 U17386 ( .A(n14040), .B(n19173), .S(n15000), .Z(n14041) );
  OAI21_X1 U17387 ( .B1(n19233), .B2(n15012), .A(n14041), .ZN(P2_U2883) );
  OAI21_X1 U17388 ( .B1(n19042), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19043), 
        .ZN(n14042) );
  OAI21_X1 U17389 ( .B1(n14043), .B2(n19043), .A(n14042), .ZN(P2_U3612) );
  AOI22_X1 U17390 ( .A1(n14592), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14618), .ZN(n14047) );
  NOR3_X1 U17391 ( .A1(n14618), .A2(n14044), .A3(n20213), .ZN(n14045) );
  AOI22_X1 U17392 ( .A1(n14595), .A2(n14606), .B1(n14593), .B2(DATAI_30_), 
        .ZN(n14046) );
  OAI211_X1 U17393 ( .C1(n14048), .C2(n14622), .A(n14047), .B(n14046), .ZN(
        P1_U2874) );
  AOI22_X1 U17394 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14053) );
  AOI22_X1 U17395 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U17396 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17397 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10762), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14050) );
  NAND4_X1 U17398 ( .A1(n14053), .A2(n14052), .A3(n14051), .A4(n14050), .ZN(
        n14059) );
  AOI22_X1 U17399 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17400 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14056) );
  AOI22_X1 U17401 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17402 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n14108), .ZN(n14054) );
  NAND4_X1 U17403 ( .A1(n14057), .A2(n14056), .A3(n14055), .A4(n14054), .ZN(
        n14058) );
  NOR2_X1 U17404 ( .A1(n14059), .A2(n14058), .ZN(n15003) );
  INV_X1 U17405 ( .A(n15003), .ZN(n14060) );
  AOI22_X1 U17406 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U17407 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U17408 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U17409 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10762), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14061) );
  NAND4_X1 U17410 ( .A1(n14064), .A2(n14063), .A3(n14062), .A4(n14061), .ZN(
        n14070) );
  AOI22_X1 U17411 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17412 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14067) );
  AOI22_X1 U17413 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U17414 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14065) );
  NAND4_X1 U17415 ( .A1(n14068), .A2(n14067), .A3(n14066), .A4(n14065), .ZN(
        n14069) );
  NOR2_X1 U17416 ( .A1(n14070), .A2(n14069), .ZN(n14998) );
  AOI22_X1 U17417 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U17418 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U17419 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10742), .B1(
        n15540), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U17420 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10762), .B1(
        n10761), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14071) );
  NAND4_X1 U17421 ( .A1(n14074), .A2(n14073), .A3(n14072), .A4(n14071), .ZN(
        n14080) );
  AOI22_X1 U17422 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17423 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17424 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U17425 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n14108), .ZN(n14075) );
  NAND4_X1 U17426 ( .A1(n14078), .A2(n14077), .A3(n14076), .A4(n14075), .ZN(
        n14079) );
  NOR2_X1 U17427 ( .A1(n14080), .A2(n14079), .ZN(n14991) );
  AOI22_X1 U17428 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U17429 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U17430 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17431 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14082) );
  NAND4_X1 U17432 ( .A1(n14085), .A2(n14084), .A3(n14083), .A4(n14082), .ZN(
        n14091) );
  AOI22_X1 U17433 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U17434 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14088) );
  AOI22_X1 U17435 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U17436 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14086) );
  NAND4_X1 U17437 ( .A1(n14089), .A2(n14088), .A3(n14087), .A4(n14086), .ZN(
        n14090) );
  OR2_X1 U17438 ( .A1(n14091), .A2(n14090), .ZN(n14987) );
  NAND2_X1 U17439 ( .A1(n14986), .A2(n14987), .ZN(n14974) );
  AOI22_X1 U17440 ( .A1(n10760), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17441 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17442 ( .A1(n15540), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U17443 ( .A1(n10761), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14092) );
  NAND4_X1 U17444 ( .A1(n14095), .A2(n14094), .A3(n14093), .A4(n14092), .ZN(
        n14102) );
  AOI22_X1 U17445 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14100) );
  AOI22_X1 U17446 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U17447 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17448 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14108), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14097) );
  NAND4_X1 U17449 ( .A1(n14100), .A2(n14099), .A3(n14098), .A4(n14097), .ZN(
        n14101) );
  NOR2_X1 U17450 ( .A1(n14102), .A2(n14101), .ZN(n14975) );
  AOI22_X1 U17451 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10760), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U17452 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U17453 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n15540), .B1(
        n10742), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17454 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10761), .B1(
        n10762), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14103) );
  NAND4_X1 U17455 ( .A1(n14106), .A2(n14105), .A3(n14104), .A4(n14103), .ZN(
        n14115) );
  AOI22_X1 U17456 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17457 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10748), .B1(
        n10734), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17458 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14096), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U17459 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14108), .ZN(n14110) );
  NAND4_X1 U17460 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        n14114) );
  NAND2_X1 U17461 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14119) );
  NAND2_X1 U17462 ( .A1(n14270), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14118) );
  NAND2_X1 U17463 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14117) );
  NAND2_X1 U17464 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14116) );
  AND4_X1 U17465 ( .A1(n14119), .A2(n14118), .A3(n14117), .A4(n14116), .ZN(
        n14122) );
  AOI22_X1 U17466 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17467 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14120) );
  XNOR2_X1 U17468 ( .A(n15529), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14277) );
  NAND4_X1 U17469 ( .A1(n14122), .A2(n14121), .A3(n14120), .A4(n14277), .ZN(
        n14131) );
  NAND2_X1 U17470 ( .A1(n9806), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14126) );
  NAND2_X1 U17471 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14125) );
  NAND2_X1 U17472 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14124) );
  NAND2_X1 U17473 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14123) );
  AND4_X1 U17474 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        n14129) );
  AOI22_X1 U17475 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14128) );
  AOI22_X1 U17476 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14127) );
  NAND4_X1 U17477 ( .A1(n14129), .A2(n14268), .A3(n14128), .A4(n14127), .ZN(
        n14130) );
  AND2_X1 U17478 ( .A1(n14131), .A2(n14130), .ZN(n14132) );
  AND2_X1 U17479 ( .A1(n14133), .A2(n14132), .ZN(n14155) );
  NAND2_X1 U17480 ( .A1(n14155), .A2(n14957), .ZN(n14136) );
  INV_X1 U17481 ( .A(n14132), .ZN(n14137) );
  INV_X1 U17482 ( .A(n14133), .ZN(n14134) );
  OAI21_X1 U17483 ( .B1(n9992), .B2(n14137), .A(n14134), .ZN(n14135) );
  NOR2_X1 U17484 ( .A1(n14957), .A2(n14137), .ZN(n14970) );
  NAND2_X1 U17485 ( .A1(n9804), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14142) );
  NAND2_X1 U17486 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14141) );
  NAND2_X1 U17487 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14140) );
  NAND2_X1 U17488 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14139) );
  AND4_X1 U17489 ( .A1(n14142), .A2(n14141), .A3(n14140), .A4(n14139), .ZN(
        n14145) );
  AOI22_X1 U17490 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U17491 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14143) );
  NAND4_X1 U17492 ( .A1(n14145), .A2(n14144), .A3(n14143), .A4(n14277), .ZN(
        n14154) );
  NAND2_X1 U17493 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n14149) );
  NAND2_X1 U17494 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14148) );
  NAND2_X1 U17495 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14147) );
  NAND2_X1 U17496 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14146) );
  AND4_X1 U17497 ( .A1(n14149), .A2(n14148), .A3(n14147), .A4(n14146), .ZN(
        n14152) );
  AOI22_X1 U17498 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17499 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14150) );
  NAND4_X1 U17500 ( .A1(n14152), .A2(n14268), .A3(n14151), .A4(n14150), .ZN(
        n14153) );
  NAND2_X1 U17501 ( .A1(n14154), .A2(n14153), .ZN(n14956) );
  INV_X1 U17502 ( .A(n14155), .ZN(n14156) );
  NOR2_X1 U17503 ( .A1(n14156), .A2(n14956), .ZN(n14175) );
  AOI211_X1 U17504 ( .C1(n14956), .C2(n14156), .A(n14222), .B(n14175), .ZN(
        n14959) );
  INV_X1 U17505 ( .A(n14970), .ZN(n14157) );
  NAND2_X1 U17506 ( .A1(n9806), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14161) );
  NAND2_X1 U17507 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14160) );
  NAND2_X1 U17508 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14159) );
  NAND2_X1 U17509 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14158) );
  AND4_X1 U17510 ( .A1(n14161), .A2(n14160), .A3(n14159), .A4(n14158), .ZN(
        n14164) );
  AOI22_X1 U17511 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14163) );
  AOI22_X1 U17512 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14162) );
  NAND4_X1 U17513 ( .A1(n14164), .A2(n14163), .A3(n14162), .A4(n14277), .ZN(
        n14173) );
  NAND2_X1 U17514 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14168) );
  NAND2_X1 U17515 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14167) );
  NAND2_X1 U17516 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14166) );
  NAND2_X1 U17517 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14165) );
  AND4_X1 U17518 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n14171) );
  AOI22_X1 U17519 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17520 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14169) );
  NAND4_X1 U17521 ( .A1(n14171), .A2(n14268), .A3(n14170), .A4(n14169), .ZN(
        n14172) );
  AND2_X1 U17522 ( .A1(n14173), .A2(n14172), .ZN(n14176) );
  NAND2_X1 U17523 ( .A1(n14175), .A2(n14176), .ZN(n14199) );
  OAI211_X1 U17524 ( .C1(n14175), .C2(n14176), .A(n14199), .B(n14174), .ZN(
        n14179) );
  XNOR2_X2 U17525 ( .A(n14178), .B(n14180), .ZN(n14948) );
  INV_X1 U17526 ( .A(n14176), .ZN(n14177) );
  NOR2_X1 U17527 ( .A1(n14957), .A2(n14177), .ZN(n14947) );
  NAND2_X2 U17528 ( .A1(n14948), .A2(n14947), .ZN(n14946) );
  NAND2_X1 U17529 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14186) );
  NAND2_X1 U17530 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14185) );
  NAND2_X1 U17531 ( .A1(n14254), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14184) );
  NAND2_X1 U17532 ( .A1(n14276), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14183) );
  AND4_X1 U17533 ( .A1(n14186), .A2(n14185), .A3(n14184), .A4(n14183), .ZN(
        n14189) );
  AOI22_X1 U17534 ( .A1(n9809), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14273), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14188) );
  AOI22_X1 U17535 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14187) );
  NAND4_X1 U17536 ( .A1(n14189), .A2(n14188), .A3(n14187), .A4(n14277), .ZN(
        n14198) );
  NAND2_X1 U17537 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n14193) );
  NAND2_X1 U17538 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14192) );
  NAND2_X1 U17539 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14191) );
  NAND2_X1 U17540 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14190) );
  AND4_X1 U17541 ( .A1(n14193), .A2(n14192), .A3(n14191), .A4(n14190), .ZN(
        n14196) );
  AOI22_X1 U17542 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14195) );
  AOI22_X1 U17543 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14194) );
  NAND4_X1 U17544 ( .A1(n14196), .A2(n14268), .A3(n14195), .A4(n14194), .ZN(
        n14197) );
  NAND2_X1 U17545 ( .A1(n14198), .A2(n14197), .ZN(n14201) );
  AOI21_X1 U17546 ( .B1(n14199), .B2(n14201), .A(n14222), .ZN(n14200) );
  NAND2_X1 U17547 ( .A1(n14200), .A2(n14223), .ZN(n14202) );
  NOR2_X1 U17548 ( .A1(n14957), .A2(n14201), .ZN(n14940) );
  INV_X1 U17549 ( .A(n14202), .ZN(n14203) );
  AOI21_X2 U17550 ( .B1(n14939), .B2(n14940), .A(n14205), .ZN(n14228) );
  NAND2_X1 U17551 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14209) );
  NAND2_X1 U17552 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14208) );
  NAND2_X1 U17553 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14207) );
  NAND2_X1 U17554 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14206) );
  AND4_X1 U17555 ( .A1(n14209), .A2(n14208), .A3(n14207), .A4(n14206), .ZN(
        n14212) );
  AOI22_X1 U17556 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14211) );
  AOI22_X1 U17557 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14210) );
  NAND4_X1 U17558 ( .A1(n14212), .A2(n14211), .A3(n14210), .A4(n14277), .ZN(
        n14221) );
  NAND2_X1 U17559 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14216) );
  NAND2_X1 U17560 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14215) );
  NAND2_X1 U17561 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14214) );
  NAND2_X1 U17562 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14213) );
  AND4_X1 U17563 ( .A1(n14216), .A2(n14215), .A3(n14214), .A4(n14213), .ZN(
        n14219) );
  AOI22_X1 U17564 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14218) );
  AOI22_X1 U17565 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14217) );
  NAND4_X1 U17566 ( .A1(n14219), .A2(n14268), .A3(n14218), .A4(n14217), .ZN(
        n14220) );
  NAND2_X1 U17567 ( .A1(n14221), .A2(n14220), .ZN(n14225) );
  AOI21_X1 U17568 ( .B1(n14223), .B2(n14225), .A(n14222), .ZN(n14224) );
  OR2_X1 U17569 ( .A1(n14223), .A2(n14225), .ZN(n14246) );
  NAND2_X1 U17570 ( .A1(n14224), .A2(n14246), .ZN(n14229) );
  INV_X1 U17571 ( .A(n14225), .ZN(n14226) );
  NAND2_X1 U17572 ( .A1(n14227), .A2(n14226), .ZN(n14934) );
  NAND2_X1 U17573 ( .A1(n9804), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14233) );
  NAND2_X1 U17574 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14232) );
  NAND2_X1 U17575 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14231) );
  NAND2_X1 U17576 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14230) );
  AND4_X1 U17577 ( .A1(n14233), .A2(n14232), .A3(n14231), .A4(n14230), .ZN(
        n14236) );
  AOI22_X1 U17578 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14235) );
  AOI22_X1 U17579 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14234) );
  NAND4_X1 U17580 ( .A1(n14236), .A2(n14235), .A3(n14234), .A4(n14277), .ZN(
        n14245) );
  NAND2_X1 U17581 ( .A1(n9804), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n14240) );
  NAND2_X1 U17582 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14239) );
  NAND2_X1 U17583 ( .A1(n15518), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14238) );
  NAND2_X1 U17584 ( .A1(n14272), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14237) );
  AND4_X1 U17585 ( .A1(n14240), .A2(n14239), .A3(n14238), .A4(n14237), .ZN(
        n14243) );
  AOI22_X1 U17586 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U17587 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14241) );
  NAND4_X1 U17588 ( .A1(n14243), .A2(n14268), .A3(n14242), .A4(n14241), .ZN(
        n14244) );
  AND2_X1 U17589 ( .A1(n14245), .A2(n14244), .ZN(n14929) );
  INV_X1 U17590 ( .A(n14246), .ZN(n14927) );
  NAND3_X1 U17591 ( .A1(n14927), .A2(n14929), .A3(n14957), .ZN(n14263) );
  AOI22_X1 U17592 ( .A1(n9806), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U17593 ( .A1(n14247), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U17594 ( .A1(n14249), .A2(n14248), .ZN(n14261) );
  AOI22_X1 U17595 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14251) );
  AOI22_X1 U17596 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14250) );
  NAND3_X1 U17597 ( .A1(n14251), .A2(n14250), .A3(n14277), .ZN(n14260) );
  AOI22_X1 U17598 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14253) );
  AOI22_X1 U17599 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14252) );
  NAND2_X1 U17600 ( .A1(n14253), .A2(n14252), .ZN(n14259) );
  AOI22_X1 U17601 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14257) );
  AOI22_X1 U17602 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14256) );
  NAND3_X1 U17603 ( .A1(n14257), .A2(n14256), .A3(n14268), .ZN(n14258) );
  OAI22_X1 U17604 ( .A1(n14261), .A2(n14260), .B1(n14259), .B2(n14258), .ZN(
        n14262) );
  XNOR2_X1 U17605 ( .A(n14263), .B(n14262), .ZN(n14922) );
  AOI22_X1 U17606 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17607 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14265) );
  NAND2_X1 U17608 ( .A1(n14266), .A2(n14265), .ZN(n14283) );
  AOI22_X1 U17609 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14269) );
  AOI22_X1 U17610 ( .A1(n14276), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14267) );
  NAND3_X1 U17611 ( .A1(n14269), .A2(n14268), .A3(n14267), .ZN(n14282) );
  AOI22_X1 U17612 ( .A1(n14271), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14270), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U17613 ( .A1(n14273), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14274) );
  NAND2_X1 U17614 ( .A1(n14275), .A2(n14274), .ZN(n14281) );
  AOI22_X1 U17615 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14276), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14279) );
  AOI22_X1 U17616 ( .A1(n9822), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14254), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14278) );
  NAND3_X1 U17617 ( .A1(n14279), .A2(n14278), .A3(n14277), .ZN(n14280) );
  OAI22_X1 U17618 ( .A1(n14283), .A2(n14282), .B1(n14281), .B2(n14280), .ZN(
        n14284) );
  INV_X1 U17619 ( .A(n14284), .ZN(n14285) );
  XNOR2_X1 U17620 ( .A(n14286), .B(n14285), .ZN(n14295) );
  AOI22_X1 U17621 ( .A1(n16286), .A2(n19221), .B1(n19231), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U17622 ( .A1(n19215), .A2(BUF2_REG_30__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14287) );
  OAI211_X1 U17623 ( .C1(n14289), .C2(n15023), .A(n14288), .B(n14287), .ZN(
        n14290) );
  INV_X1 U17624 ( .A(n14290), .ZN(n14291) );
  OAI21_X1 U17625 ( .B1(n14295), .B2(n15120), .A(n14291), .ZN(P2_U2889) );
  NOR2_X1 U17626 ( .A1(n14292), .A2(n13301), .ZN(n14293) );
  AOI21_X1 U17627 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15010), .A(n14293), .ZN(
        n14294) );
  OAI21_X1 U17628 ( .B1(n14295), .B2(n15012), .A(n14294), .ZN(P2_U2857) );
  INV_X1 U17629 ( .A(n14296), .ZN(n14297) );
  OAI21_X1 U17630 ( .B1(n14298), .B2(n16358), .A(n14297), .ZN(n14300) );
  NOR2_X1 U17631 ( .A1(n19296), .A2(n14914), .ZN(n14299) );
  AOI211_X1 U17632 ( .C1(n19287), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14300), .B(n14299), .ZN(n14304) );
  NAND3_X1 U17633 ( .A1(n14302), .A2(n19291), .A3(n14301), .ZN(n14303) );
  OAI211_X1 U17634 ( .C1(n15258), .C2(n14305), .A(n14304), .B(n14303), .ZN(
        P2_U3012) );
  NOR2_X1 U17635 ( .A1(n14307), .A2(n14306), .ZN(n14310) );
  AOI21_X1 U17636 ( .B1(n14308), .B2(n12259), .A(n15882), .ZN(n14309) );
  AOI211_X1 U17637 ( .C1(n11607), .C2(n14311), .A(n14310), .B(n14309), .ZN(
        n15864) );
  INV_X1 U17638 ( .A(n15864), .ZN(n14315) );
  OAI21_X1 U17639 ( .B1(n12313), .B2(n14311), .A(n12259), .ZN(n14312) );
  OAI21_X1 U17640 ( .B1(n14313), .B2(n15882), .A(n14312), .ZN(n20009) );
  NOR2_X1 U17641 ( .A1(n12718), .A2(n14313), .ZN(n20878) );
  AOI21_X1 U17642 ( .B1(n20878), .B2(n20879), .A(n20876), .ZN(n14314) );
  NOR2_X1 U17643 ( .A1(n20009), .A2(n14314), .ZN(n15868) );
  NOR2_X1 U17644 ( .A1(n15868), .A2(n20008), .ZN(n20015) );
  MUX2_X1 U17645 ( .A(P1_MORE_REG_SCAN_IN), .B(n14315), .S(n20015), .Z(
        P1_U3484) );
  OAI21_X1 U17646 ( .B1(n14319), .B2(n14318), .A(n14317), .ZN(n14773) );
  INV_X1 U17647 ( .A(n14773), .ZN(n14327) );
  INV_X1 U17648 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21153) );
  OAI22_X1 U17649 ( .A1(n14320), .A2(n20057), .B1(n20059), .B2(n14631), .ZN(
        n14323) );
  INV_X1 U17650 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21220) );
  NOR4_X1 U17651 ( .A1(n14369), .A2(n14321), .A3(P1_REIP_REG_28__SCAN_IN), 
        .A4(n21220), .ZN(n14322) );
  AOI211_X1 U17652 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n20043), .A(n14323), .B(
        n14322), .ZN(n14324) );
  OAI21_X1 U17653 ( .B1(n21153), .B2(n14325), .A(n14324), .ZN(n14326) );
  AOI21_X1 U17654 ( .B1(n14327), .B2(n20070), .A(n14326), .ZN(n14328) );
  OAI21_X1 U17655 ( .B1(n14629), .B2(n15978), .A(n14328), .ZN(P1_U2812) );
  NAND2_X1 U17656 ( .A1(n14643), .A2(n20047), .ZN(n14336) );
  NOR2_X1 U17657 ( .A1(n15930), .A2(n14329), .ZN(n14348) );
  AOI22_X1 U17658 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20069), .B1(
        n20073), .B2(n14639), .ZN(n14330) );
  OAI21_X1 U17659 ( .B1(n14471), .B2(n14331), .A(n14330), .ZN(n14334) );
  NOR2_X1 U17660 ( .A1(n14332), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14333) );
  AOI211_X1 U17661 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14348), .A(n14334), 
        .B(n14333), .ZN(n14335) );
  OAI211_X1 U17662 ( .C1(n14780), .C2(n15963), .A(n14336), .B(n14335), .ZN(
        P1_U2813) );
  BUF_X1 U17663 ( .A(n14337), .Z(n14338) );
  OAI21_X1 U17664 ( .B1(n14338), .B2(n14339), .A(n12440), .ZN(n14649) );
  INV_X1 U17665 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21212) );
  INV_X1 U17666 ( .A(n14369), .ZN(n14340) );
  INV_X1 U17667 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21199) );
  NAND4_X1 U17668 ( .A1(n14340), .A2(P1_REIP_REG_24__SCAN_IN), .A3(
        P1_REIP_REG_25__SCAN_IN), .A4(n21199), .ZN(n14343) );
  INV_X1 U17669 ( .A(n14651), .ZN(n14341) );
  AOI22_X1 U17670 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20069), .B1(
        n20073), .B2(n14341), .ZN(n14342) );
  OAI211_X1 U17671 ( .C1(n21212), .C2(n14471), .A(n14343), .B(n14342), .ZN(
        n14347) );
  XNOR2_X1 U17672 ( .A(n14345), .B(n14344), .ZN(n16052) );
  NOR2_X1 U17673 ( .A1(n16052), .A2(n15963), .ZN(n14346) );
  AOI211_X1 U17674 ( .C1(n14348), .C2(P1_REIP_REG_26__SCAN_IN), .A(n14347), 
        .B(n14346), .ZN(n14349) );
  OAI21_X1 U17675 ( .B1(n14649), .B2(n15978), .A(n14349), .ZN(P1_U2814) );
  AOI21_X1 U17676 ( .B1(n14352), .B2(n14351), .A(n14338), .ZN(n14662) );
  INV_X1 U17677 ( .A(n14662), .ZN(n14563) );
  AND2_X1 U17678 ( .A1(n20029), .A2(n14353), .ZN(n14391) );
  XNOR2_X1 U17679 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14357) );
  OAI22_X1 U17680 ( .A1(n14354), .A2(n20057), .B1(n20059), .B2(n14660), .ZN(
        n14355) );
  AOI21_X1 U17681 ( .B1(n20043), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14355), .ZN(
        n14356) );
  OAI21_X1 U17682 ( .B1(n14369), .B2(n14357), .A(n14356), .ZN(n14362) );
  NAND2_X1 U17683 ( .A1(n14371), .A2(n14358), .ZN(n14359) );
  NAND2_X1 U17684 ( .A1(n14360), .A2(n14359), .ZN(n16059) );
  NOR2_X1 U17685 ( .A1(n16059), .A2(n15963), .ZN(n14361) );
  AOI211_X1 U17686 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14391), .A(n14362), 
        .B(n14361), .ZN(n14363) );
  OAI21_X1 U17687 ( .B1(n14563), .B2(n15978), .A(n14363), .ZN(P1_U2815) );
  OAI21_X1 U17689 ( .B1(n14378), .B2(n14365), .A(n14351), .ZN(n14668) );
  INV_X1 U17690 ( .A(n14671), .ZN(n14366) );
  OAI22_X1 U17691 ( .A1(n14667), .A2(n20057), .B1(n20059), .B2(n14366), .ZN(
        n14367) );
  AOI21_X1 U17692 ( .B1(n20043), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14367), .ZN(
        n14368) );
  OAI21_X1 U17693 ( .B1(n14369), .B2(P1_REIP_REG_24__SCAN_IN), .A(n14368), 
        .ZN(n14375) );
  INV_X1 U17694 ( .A(n14387), .ZN(n14373) );
  INV_X1 U17695 ( .A(n14370), .ZN(n14372) );
  OAI21_X1 U17696 ( .B1(n14373), .B2(n14372), .A(n14371), .ZN(n14792) );
  NOR2_X1 U17697 ( .A1(n14792), .A2(n15963), .ZN(n14374) );
  AOI211_X1 U17698 ( .C1(n14391), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14375), 
        .B(n14374), .ZN(n14376) );
  OAI21_X1 U17699 ( .B1(n14668), .B2(n15978), .A(n14376), .ZN(P1_U2816) );
  AOI21_X1 U17700 ( .B1(n14379), .B2(n14377), .A(n14378), .ZN(n14380) );
  INV_X1 U17701 ( .A(n14380), .ZN(n14678) );
  INV_X1 U17702 ( .A(n14381), .ZN(n14383) );
  OAI21_X1 U17703 ( .B1(n14383), .B2(n14382), .A(n14676), .ZN(n14390) );
  AOI22_X1 U17704 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20069), .B1(
        n20073), .B2(n14681), .ZN(n14384) );
  OAI21_X1 U17705 ( .B1(n14471), .B2(n21214), .A(n14384), .ZN(n14389) );
  OR2_X1 U17706 ( .A1(n14396), .A2(n14385), .ZN(n14386) );
  NAND2_X1 U17707 ( .A1(n14387), .A2(n14386), .ZN(n16067) );
  NOR2_X1 U17708 ( .A1(n16067), .A2(n15963), .ZN(n14388) );
  AOI211_X1 U17709 ( .C1(n14391), .C2(n14390), .A(n14389), .B(n14388), .ZN(
        n14392) );
  OAI21_X1 U17710 ( .B1(n14678), .B2(n15978), .A(n14392), .ZN(P1_U2817) );
  OAI21_X1 U17711 ( .B1(n14393), .B2(n14394), .A(n14377), .ZN(n14686) );
  INV_X1 U17712 ( .A(n14395), .ZN(n14398) );
  INV_X1 U17713 ( .A(n14416), .ZN(n14397) );
  AOI21_X1 U17714 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14807) );
  INV_X1 U17715 ( .A(n14399), .ZN(n14400) );
  NAND2_X1 U17716 ( .A1(n20029), .A2(n14400), .ZN(n14434) );
  INV_X1 U17717 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14798) );
  OAI22_X1 U17718 ( .A1(n14401), .A2(n20057), .B1(n20059), .B2(n14688), .ZN(
        n14402) );
  AOI21_X1 U17719 ( .B1(n20043), .B2(P1_EBX_REG_22__SCAN_IN), .A(n14402), .ZN(
        n14406) );
  OAI21_X1 U17720 ( .B1(n14403), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14404) );
  OAI211_X1 U17721 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(P1_REIP_REG_22__SCAN_IN), .A(n20077), .B(n14404), .ZN(n14405) );
  OAI211_X1 U17722 ( .C1(n14434), .C2(n14798), .A(n14406), .B(n14405), .ZN(
        n14407) );
  AOI21_X1 U17723 ( .B1(n14807), .B2(n20070), .A(n14407), .ZN(n14408) );
  OAI21_X1 U17724 ( .B1(n14686), .B2(n15978), .A(n14408), .ZN(P1_U2818) );
  INV_X1 U17725 ( .A(n14393), .ZN(n14410) );
  OAI21_X1 U17726 ( .B1(n14411), .B2(n14409), .A(n14410), .ZN(n14696) );
  NOR2_X1 U17727 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20032), .ZN(n14412) );
  AOI22_X1 U17728 ( .A1(n14699), .A2(n20073), .B1(n14413), .B2(n14412), .ZN(
        n14420) );
  AND2_X1 U17729 ( .A1(n14427), .A2(n14414), .ZN(n14415) );
  NOR2_X1 U17730 ( .A1(n14416), .A2(n14415), .ZN(n15892) );
  INV_X1 U17731 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15887) );
  AOI22_X1 U17732 ( .A1(n20043), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20069), .ZN(n14417) );
  OAI21_X1 U17733 ( .B1(n14434), .B2(n15887), .A(n14417), .ZN(n14418) );
  AOI21_X1 U17734 ( .B1(n15892), .B2(n20070), .A(n14418), .ZN(n14419) );
  OAI211_X1 U17735 ( .C1(n14696), .C2(n15978), .A(n14420), .B(n14419), .ZN(
        P1_U2819) );
  INV_X1 U17736 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20966) );
  INV_X1 U17737 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21229) );
  NOR2_X1 U17738 ( .A1(n20966), .A2(n21229), .ZN(n14422) );
  NAND2_X1 U17739 ( .A1(n14421), .A2(n14479), .ZN(n15985) );
  NOR2_X1 U17740 ( .A1(n14444), .A2(n15985), .ZN(n14443) );
  AOI21_X1 U17741 ( .B1(n14422), .B2(n14443), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14435) );
  AOI21_X1 U17742 ( .B1(n14424), .B2(n14423), .A(n14409), .ZN(n14709) );
  NAND2_X1 U17743 ( .A1(n14709), .A2(n20047), .ZN(n14433) );
  OAI22_X1 U17744 ( .A1(n14425), .A2(n20057), .B1(n20059), .B2(n14707), .ZN(
        n14431) );
  INV_X1 U17745 ( .A(n14442), .ZN(n14429) );
  INV_X1 U17746 ( .A(n14426), .ZN(n14428) );
  OAI21_X1 U17747 ( .B1(n14429), .B2(n14428), .A(n14427), .ZN(n14813) );
  NOR2_X1 U17748 ( .A1(n14813), .A2(n15963), .ZN(n14430) );
  AOI211_X1 U17749 ( .C1(n20043), .C2(P1_EBX_REG_20__SCAN_IN), .A(n14431), .B(
        n14430), .ZN(n14432) );
  OAI211_X1 U17750 ( .C1(n14435), .C2(n14434), .A(n14433), .B(n14432), .ZN(
        P1_U2820) );
  INV_X1 U17751 ( .A(n14423), .ZN(n14438) );
  AOI21_X1 U17752 ( .B1(n14439), .B2(n14437), .A(n14438), .ZN(n14713) );
  INV_X1 U17753 ( .A(n14713), .ZN(n14585) );
  OR2_X1 U17754 ( .A1(n14457), .A2(n14440), .ZN(n14441) );
  AND2_X1 U17755 ( .A1(n14442), .A2(n14441), .ZN(n16075) );
  AOI22_X1 U17756 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20069), .B1(
        n20073), .B2(n14716), .ZN(n14448) );
  INV_X1 U17757 ( .A(n14443), .ZN(n14449) );
  NOR2_X1 U17758 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14449), .ZN(n14461) );
  INV_X1 U17759 ( .A(n14444), .ZN(n14445) );
  INV_X1 U17760 ( .A(n15950), .ZN(n15983) );
  OAI21_X1 U17761 ( .B1(n15930), .B2(n14445), .A(n15983), .ZN(n14477) );
  OAI21_X1 U17762 ( .B1(n14461), .B2(n14477), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14447) );
  NAND2_X1 U17763 ( .A1(n20043), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14446) );
  NAND4_X1 U17764 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n20055), .ZN(
        n14451) );
  NOR3_X1 U17765 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n21229), .A3(n14449), 
        .ZN(n14450) );
  AOI211_X1 U17766 ( .C1(n16075), .C2(n20070), .A(n14451), .B(n14450), .ZN(
        n14452) );
  OAI21_X1 U17767 ( .B1(n14585), .B2(n15978), .A(n14452), .ZN(P1_U2821) );
  OAI21_X1 U17768 ( .B1(n9858), .B2(n14453), .A(n14437), .ZN(n14721) );
  NAND2_X1 U17769 ( .A1(n20069), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14454) );
  OAI211_X1 U17770 ( .C1(n20059), .C2(n14722), .A(n14454), .B(n20055), .ZN(
        n14459) );
  NOR2_X1 U17771 ( .A1(n14469), .A2(n14455), .ZN(n14456) );
  OR2_X1 U17772 ( .A1(n14457), .A2(n14456), .ZN(n14819) );
  NOR2_X1 U17773 ( .A1(n14819), .A2(n15963), .ZN(n14458) );
  AOI211_X1 U17774 ( .C1(n20043), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14459), .B(
        n14458), .ZN(n14460) );
  INV_X1 U17775 ( .A(n14460), .ZN(n14462) );
  AOI211_X1 U17776 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14477), .A(n14462), 
        .B(n14461), .ZN(n14463) );
  OAI21_X1 U17777 ( .B1(n14721), .B2(n15978), .A(n14463), .ZN(P1_U2822) );
  AND2_X1 U17778 ( .A1(n14464), .A2(n14465), .ZN(n14466) );
  OR2_X1 U17779 ( .A1(n14466), .A2(n9858), .ZN(n14740) );
  NAND2_X1 U17780 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15922) );
  INV_X1 U17781 ( .A(n15985), .ZN(n15961) );
  NAND2_X1 U17782 ( .A1(n15929), .A2(n15961), .ZN(n15944) );
  INV_X1 U17783 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21244) );
  OAI21_X1 U17784 ( .B1(n15922), .B2(n15944), .A(n21244), .ZN(n14476) );
  AND2_X1 U17785 ( .A1(n14515), .A2(n14467), .ZN(n14468) );
  NOR2_X1 U17786 ( .A1(n14469), .A2(n14468), .ZN(n16085) );
  INV_X1 U17787 ( .A(n16085), .ZN(n14513) );
  INV_X1 U17788 ( .A(n14470), .ZN(n14738) );
  OAI21_X1 U17789 ( .B1(n20057), .B2(n14736), .A(n20055), .ZN(n14473) );
  NOR2_X1 U17790 ( .A1(n14471), .A2(n12380), .ZN(n14472) );
  AOI211_X1 U17791 ( .C1(n20073), .C2(n14738), .A(n14473), .B(n14472), .ZN(
        n14474) );
  OAI21_X1 U17792 ( .B1(n14513), .B2(n15963), .A(n14474), .ZN(n14475) );
  AOI21_X1 U17793 ( .B1(n14477), .B2(n14476), .A(n14475), .ZN(n14478) );
  OAI21_X1 U17794 ( .B1(n14740), .B2(n15978), .A(n14478), .ZN(P1_U2823) );
  NAND2_X1 U17795 ( .A1(n14479), .A2(n21251), .ZN(n14487) );
  INV_X1 U17796 ( .A(n16152), .ZN(n14485) );
  NAND2_X1 U17797 ( .A1(n20043), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U17798 ( .A1(n20069), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14482) );
  NAND2_X1 U17799 ( .A1(n20073), .A2(n14480), .ZN(n14481) );
  NAND4_X1 U17800 ( .A1(n14483), .A2(n20055), .A3(n14482), .A4(n14481), .ZN(
        n14484) );
  AOI21_X1 U17801 ( .B1(n14485), .B2(n20070), .A(n14484), .ZN(n14486) );
  OAI211_X1 U17802 ( .C1(n14488), .C2(n21251), .A(n14487), .B(n14486), .ZN(
        n14489) );
  AOI21_X1 U17803 ( .B1(n14490), .B2(n20047), .A(n14489), .ZN(n14491) );
  INV_X1 U17804 ( .A(n14491), .ZN(P1_U2831) );
  OAI21_X1 U17805 ( .B1(n20032), .B2(n20053), .A(n20029), .ZN(n20068) );
  NAND2_X1 U17806 ( .A1(n20069), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14492) );
  OAI211_X1 U17807 ( .C1(n20059), .C2(n14493), .A(n14492), .B(n20055), .ZN(
        n14496) );
  NOR2_X1 U17808 ( .A1(n15963), .A2(n14494), .ZN(n14495) );
  AOI211_X1 U17809 ( .C1(n20043), .C2(P1_EBX_REG_4__SCAN_IN), .A(n14496), .B(
        n14495), .ZN(n14497) );
  OAI21_X1 U17810 ( .B1(n21170), .B2(n20068), .A(n14497), .ZN(n14500) );
  NAND3_X1 U17811 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14498) );
  NOR3_X1 U17812 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20032), .A3(n14498), .ZN(
        n14499) );
  AOI211_X1 U17813 ( .C1(n20071), .C2(n16189), .A(n14500), .B(n14499), .ZN(
        n14501) );
  OAI21_X1 U17814 ( .B1(n14503), .B2(n14502), .A(n14501), .ZN(P1_U2836) );
  OAI22_X1 U17815 ( .A1(n14504), .A2(n14546), .B1(n20092), .B2(n21167), .ZN(
        P1_U2841) );
  OAI222_X1 U17816 ( .A1(n14539), .A2(n14505), .B1(n21165), .B2(n20092), .C1(
        n14762), .C2(n14546), .ZN(P1_U2843) );
  OAI222_X1 U17817 ( .A1(n14629), .A2(n14539), .B1(n14506), .B2(n20092), .C1(
        n14773), .C2(n14546), .ZN(P1_U2844) );
  OAI222_X1 U17818 ( .A1(n14539), .A2(n14649), .B1(n21212), .B2(n20092), .C1(
        n14546), .C2(n16052), .ZN(P1_U2846) );
  OAI222_X1 U17819 ( .A1(n14539), .A2(n14563), .B1(n21211), .B2(n20092), .C1(
        n16059), .C2(n14546), .ZN(P1_U2847) );
  INV_X1 U17820 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n20955) );
  OAI222_X1 U17821 ( .A1(n14539), .A2(n14668), .B1(n20955), .B2(n20092), .C1(
        n14792), .C2(n14546), .ZN(P1_U2848) );
  OAI222_X1 U17822 ( .A1(n14678), .A2(n14539), .B1(n21214), .B2(n20092), .C1(
        n16067), .C2(n14546), .ZN(P1_U2849) );
  INV_X1 U17823 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21168) );
  INV_X1 U17824 ( .A(n14807), .ZN(n14507) );
  OAI222_X1 U17825 ( .A1(n14686), .A2(n14539), .B1(n21168), .B2(n20092), .C1(
        n14507), .C2(n14546), .ZN(P1_U2850) );
  AOI22_X1 U17826 ( .A1(n15892), .A2(n20088), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14537), .ZN(n14508) );
  OAI21_X1 U17827 ( .B1(n14696), .B2(n14539), .A(n14508), .ZN(P1_U2851) );
  INV_X1 U17828 ( .A(n14709), .ZN(n14581) );
  INV_X1 U17829 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14509) );
  OAI222_X1 U17830 ( .A1(n14581), .A2(n14539), .B1(n20092), .B2(n14509), .C1(
        n14813), .C2(n14546), .ZN(P1_U2852) );
  AOI22_X1 U17831 ( .A1(n16075), .A2(n20088), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14537), .ZN(n14510) );
  OAI21_X1 U17832 ( .B1(n14585), .B2(n14539), .A(n14510), .ZN(P1_U2853) );
  OAI22_X1 U17833 ( .A1(n14819), .A2(n14546), .B1(n21043), .B2(n20092), .ZN(
        n14511) );
  INV_X1 U17834 ( .A(n14511), .ZN(n14512) );
  OAI21_X1 U17835 ( .B1(n14721), .B2(n14539), .A(n14512), .ZN(P1_U2854) );
  OAI222_X1 U17836 ( .A1(n14740), .A2(n14539), .B1(n20092), .B2(n12380), .C1(
        n14513), .C2(n14546), .ZN(P1_U2855) );
  INV_X1 U17837 ( .A(n15937), .ZN(n14517) );
  INV_X1 U17838 ( .A(n14514), .ZN(n14516) );
  OAI21_X1 U17839 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n15926) );
  INV_X1 U17840 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21248) );
  INV_X1 U17841 ( .A(n14464), .ZN(n14519) );
  AOI21_X1 U17842 ( .B1(n14520), .B2(n14518), .A(n14519), .ZN(n15990) );
  INV_X1 U17843 ( .A(n15990), .ZN(n14598) );
  OAI222_X1 U17844 ( .A1(n15926), .A2(n14546), .B1(n20092), .B2(n21248), .C1(
        n14598), .C2(n14539), .ZN(P1_U2856) );
  OAI21_X1 U17845 ( .B1(n14522), .B2(n14525), .A(n14524), .ZN(n14608) );
  INV_X1 U17846 ( .A(n14608), .ZN(n16013) );
  NAND2_X1 U17847 ( .A1(n16013), .A2(n20089), .ZN(n14529) );
  AND2_X1 U17848 ( .A1(n14535), .A2(n14526), .ZN(n14527) );
  NOR2_X1 U17849 ( .A1(n15935), .A2(n14527), .ZN(n16101) );
  NAND2_X1 U17850 ( .A1(n16101), .A2(n20088), .ZN(n14528) );
  OAI211_X1 U17851 ( .C1(n14530), .C2(n20092), .A(n14529), .B(n14528), .ZN(
        P1_U2858) );
  AND2_X1 U17852 ( .A1(n14532), .A2(n14533), .ZN(n14534) );
  OR2_X1 U17853 ( .A1(n14534), .A2(n14522), .ZN(n15955) );
  AOI21_X1 U17854 ( .B1(n14536), .B2(n14542), .A(n12370), .ZN(n16110) );
  AOI22_X1 U17855 ( .A1(n16110), .A2(n20088), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14537), .ZN(n14538) );
  OAI21_X1 U17856 ( .B1(n15955), .B2(n14539), .A(n14538), .ZN(P1_U2859) );
  OR2_X1 U17857 ( .A1(n15974), .A2(n14540), .ZN(n14541) );
  NAND2_X1 U17858 ( .A1(n14542), .A2(n14541), .ZN(n16123) );
  OAI21_X1 U17859 ( .B1(n14544), .B2(n14545), .A(n14532), .ZN(n15962) );
  OAI222_X1 U17860 ( .A1(n16123), .A2(n14546), .B1(n20092), .B2(n10167), .C1(
        n15962), .C2(n14539), .ZN(P1_U2860) );
  AOI22_X1 U17861 ( .A1(n14592), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14618), .ZN(n14548) );
  AOI22_X1 U17862 ( .A1(n14595), .A2(n14609), .B1(n14593), .B2(DATAI_29_), 
        .ZN(n14547) );
  OAI211_X1 U17863 ( .C1(n14505), .C2(n14622), .A(n14548), .B(n14547), .ZN(
        P1_U2875) );
  AOI22_X1 U17864 ( .A1(n14592), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14618), .ZN(n14550) );
  AOI22_X1 U17865 ( .A1(n14595), .A2(n14611), .B1(n14593), .B2(DATAI_28_), 
        .ZN(n14549) );
  OAI211_X1 U17866 ( .C1(n14629), .C2(n14622), .A(n14550), .B(n14549), .ZN(
        P1_U2876) );
  AOI22_X1 U17867 ( .A1(n14592), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14618), .ZN(n14552) );
  AOI22_X1 U17868 ( .A1(n14595), .A2(n14619), .B1(n14593), .B2(DATAI_27_), 
        .ZN(n14551) );
  OAI211_X1 U17869 ( .C1(n14553), .C2(n14622), .A(n14552), .B(n14551), .ZN(
        P1_U2877) );
  INV_X1 U17870 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16558) );
  NOR2_X1 U17871 ( .A1(n14565), .A2(n16558), .ZN(n14558) );
  INV_X1 U17872 ( .A(n14595), .ZN(n14556) );
  INV_X1 U17873 ( .A(n14593), .ZN(n14554) );
  OAI22_X1 U17874 ( .A1(n14556), .A2(n14555), .B1(n14554), .B2(n20984), .ZN(
        n14557) );
  AOI211_X1 U17875 ( .C1(n14618), .C2(P1_EAX_REG_26__SCAN_IN), .A(n14558), .B(
        n14557), .ZN(n14559) );
  OAI21_X1 U17876 ( .B1(n14649), .B2(n14622), .A(n14559), .ZN(P1_U2878) );
  AOI22_X1 U17877 ( .A1(n14592), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14618), .ZN(n14562) );
  AOI22_X1 U17878 ( .A1(n14595), .A2(n14560), .B1(n14593), .B2(DATAI_25_), 
        .ZN(n14561) );
  OAI211_X1 U17879 ( .C1(n14563), .C2(n14622), .A(n14562), .B(n14561), .ZN(
        P1_U2879) );
  INV_X1 U17880 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14564) );
  OAI22_X1 U17881 ( .A1(n14565), .A2(n14564), .B1(n21019), .B2(n14602), .ZN(
        n14566) );
  INV_X1 U17882 ( .A(n14566), .ZN(n14569) );
  AOI22_X1 U17883 ( .A1(n14595), .A2(n14567), .B1(n14593), .B2(DATAI_24_), 
        .ZN(n14568) );
  OAI211_X1 U17884 ( .C1(n14668), .C2(n14622), .A(n14569), .B(n14568), .ZN(
        P1_U2880) );
  AOI22_X1 U17885 ( .A1(n14592), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14618), .ZN(n14571) );
  AOI22_X1 U17886 ( .A1(n14595), .A2(n20229), .B1(n14593), .B2(DATAI_23_), 
        .ZN(n14570) );
  OAI211_X1 U17887 ( .C1(n14678), .C2(n14622), .A(n14571), .B(n14570), .ZN(
        P1_U2881) );
  AOI22_X1 U17888 ( .A1(n14592), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14618), .ZN(n14574) );
  AOI22_X1 U17889 ( .A1(n14595), .A2(n14572), .B1(n14593), .B2(DATAI_22_), 
        .ZN(n14573) );
  OAI211_X1 U17890 ( .C1(n14686), .C2(n14622), .A(n14574), .B(n14573), .ZN(
        P1_U2882) );
  AOI22_X1 U17891 ( .A1(n14592), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14618), .ZN(n14577) );
  AOI22_X1 U17892 ( .A1(n14595), .A2(n14575), .B1(n14593), .B2(DATAI_21_), 
        .ZN(n14576) );
  OAI211_X1 U17893 ( .C1(n14696), .C2(n14622), .A(n14577), .B(n14576), .ZN(
        P1_U2883) );
  AOI22_X1 U17894 ( .A1(n14592), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14618), .ZN(n14580) );
  AOI22_X1 U17895 ( .A1(n14595), .A2(n14578), .B1(n14593), .B2(DATAI_20_), 
        .ZN(n14579) );
  OAI211_X1 U17896 ( .C1(n14581), .C2(n14622), .A(n14580), .B(n14579), .ZN(
        P1_U2884) );
  AOI22_X1 U17897 ( .A1(n14592), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14618), .ZN(n14584) );
  AOI22_X1 U17898 ( .A1(n14595), .A2(n14582), .B1(n14593), .B2(DATAI_19_), 
        .ZN(n14583) );
  OAI211_X1 U17899 ( .C1(n14585), .C2(n14622), .A(n14584), .B(n14583), .ZN(
        P1_U2885) );
  AOI22_X1 U17900 ( .A1(n14592), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14618), .ZN(n14588) );
  AOI22_X1 U17901 ( .A1(n14595), .A2(n14586), .B1(n14593), .B2(DATAI_18_), 
        .ZN(n14587) );
  OAI211_X1 U17902 ( .C1(n14721), .C2(n14622), .A(n14588), .B(n14587), .ZN(
        P1_U2886) );
  AOI22_X1 U17903 ( .A1(n14592), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14618), .ZN(n14591) );
  AOI22_X1 U17904 ( .A1(n14595), .A2(n14589), .B1(n14593), .B2(DATAI_17_), 
        .ZN(n14590) );
  OAI211_X1 U17905 ( .C1(n14740), .C2(n14622), .A(n14591), .B(n14590), .ZN(
        P1_U2887) );
  AOI22_X1 U17906 ( .A1(n14592), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14618), .ZN(n14597) );
  AOI22_X1 U17907 ( .A1(n14595), .A2(n14594), .B1(n14593), .B2(DATAI_16_), 
        .ZN(n14596) );
  OAI211_X1 U17908 ( .C1(n14598), .C2(n14622), .A(n14597), .B(n14596), .ZN(
        P1_U2888) );
  INV_X1 U17909 ( .A(n14518), .ZN(n14599) );
  AOI21_X1 U17910 ( .B1(n14600), .B2(n14524), .A(n14599), .ZN(n16001) );
  INV_X1 U17911 ( .A(n16001), .ZN(n14605) );
  OAI222_X1 U17912 ( .A1(n14605), .A2(n14622), .B1(n14604), .B2(n14603), .C1(
        n14602), .C2(n14601), .ZN(P1_U2889) );
  AOI22_X1 U17913 ( .A1(n14620), .A2(n14606), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14618), .ZN(n14607) );
  OAI21_X1 U17914 ( .B1(n14608), .B2(n14622), .A(n14607), .ZN(P1_U2890) );
  AOI22_X1 U17915 ( .A1(n14620), .A2(n14609), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14618), .ZN(n14610) );
  OAI21_X1 U17916 ( .B1(n15955), .B2(n14622), .A(n14610), .ZN(P1_U2891) );
  AOI22_X1 U17917 ( .A1(n14620), .A2(n14611), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14618), .ZN(n14612) );
  OAI21_X1 U17918 ( .B1(n15962), .B2(n14622), .A(n14612), .ZN(P1_U2892) );
  INV_X1 U17919 ( .A(n14614), .ZN(n14615) );
  AOI21_X1 U17920 ( .B1(n14617), .B2(n14616), .A(n14615), .ZN(n16030) );
  INV_X1 U17921 ( .A(n16030), .ZN(n15979) );
  AOI22_X1 U17922 ( .A1(n14620), .A2(n14619), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14618), .ZN(n14621) );
  OAI21_X1 U17923 ( .B1(n15979), .B2(n14622), .A(n14621), .ZN(P1_U2893) );
  NAND2_X1 U17924 ( .A1(n10154), .A2(n14623), .ZN(n14645) );
  NAND2_X1 U17925 ( .A1(n14675), .A2(n14645), .ZN(n14627) );
  OAI21_X1 U17926 ( .B1(n14624), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14627), .ZN(n14626) );
  MUX2_X1 U17927 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14783), .S(
        n16009), .Z(n14625) );
  OAI211_X1 U17928 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14627), .A(
        n14626), .B(n14625), .ZN(n14628) );
  XOR2_X1 U17929 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14628), .Z(
        n14777) );
  INV_X1 U17930 ( .A(n14629), .ZN(n14633) );
  NAND2_X1 U17931 ( .A1(n20149), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14772) );
  NAND2_X1 U17932 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14630) );
  OAI211_X1 U17933 ( .C1(n20141), .C2(n14631), .A(n14772), .B(n14630), .ZN(
        n14632) );
  AOI21_X1 U17934 ( .B1(n14633), .B2(n20178), .A(n14632), .ZN(n14634) );
  OAI21_X1 U17935 ( .B1(n20155), .B2(n14777), .A(n14634), .ZN(P1_U2971) );
  INV_X1 U17936 ( .A(n14635), .ZN(n14637) );
  MUX2_X1 U17937 ( .A(n14637), .B(n14636), .S(n14647), .Z(n14638) );
  XNOR2_X1 U17938 ( .A(n14638), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14786) );
  NAND2_X1 U17939 ( .A1(n16043), .A2(n14639), .ZN(n14640) );
  NAND2_X1 U17940 ( .A1(n20149), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14779) );
  OAI211_X1 U17941 ( .C1(n16047), .C2(n14641), .A(n14640), .B(n14779), .ZN(
        n14642) );
  AOI21_X1 U17942 ( .B1(n14643), .B2(n20178), .A(n14642), .ZN(n14644) );
  OAI21_X1 U17943 ( .B1(n20155), .B2(n14786), .A(n14644), .ZN(P1_U2972) );
  OAI211_X1 U17944 ( .C1(n14647), .C2(n14675), .A(n14646), .B(n14645), .ZN(
        n14648) );
  XOR2_X1 U17945 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14648), .Z(
        n16056) );
  INV_X1 U17946 ( .A(n14649), .ZN(n14653) );
  NOR2_X1 U17947 ( .A1(n20140), .A2(n21199), .ZN(n16050) );
  AOI21_X1 U17948 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16050), .ZN(n14650) );
  OAI21_X1 U17949 ( .B1(n14651), .B2(n20141), .A(n14650), .ZN(n14652) );
  AOI21_X1 U17950 ( .B1(n14653), .B2(n20178), .A(n14652), .ZN(n14654) );
  OAI21_X1 U17951 ( .B1(n20155), .B2(n16056), .A(n14654), .ZN(P1_U2973) );
  NOR3_X1 U17952 ( .A1(n14675), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14657) );
  NAND2_X1 U17953 ( .A1(n14655), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14664) );
  NOR2_X1 U17954 ( .A1(n14664), .A2(n14794), .ZN(n14656) );
  MUX2_X1 U17955 ( .A(n14657), .B(n14656), .S(n10154), .Z(n14658) );
  XNOR2_X1 U17956 ( .A(n14658), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16058) );
  AOI22_X1 U17957 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14659) );
  OAI21_X1 U17958 ( .B1(n14660), .B2(n20141), .A(n14659), .ZN(n14661) );
  AOI21_X1 U17959 ( .B1(n14662), .B2(n20178), .A(n14661), .ZN(n14663) );
  OAI21_X1 U17960 ( .B1(n20155), .B2(n16058), .A(n14663), .ZN(P1_U2974) );
  NOR2_X1 U17961 ( .A1(n14675), .A2(n10154), .ZN(n14665) );
  MUX2_X1 U17962 ( .A(n16008), .B(n14665), .S(n14664), .Z(n14666) );
  XNOR2_X1 U17963 ( .A(n14666), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14797) );
  NAND2_X1 U17964 ( .A1(n20149), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14791) );
  OAI21_X1 U17965 ( .B1(n16047), .B2(n14667), .A(n14791), .ZN(n14670) );
  NOR2_X1 U17966 ( .A1(n14668), .A2(n20142), .ZN(n14669) );
  OAI21_X1 U17967 ( .B1(n14797), .B2(n20155), .A(n14672), .ZN(P1_U2975) );
  XNOR2_X1 U17968 ( .A(n14647), .B(n14673), .ZN(n14674) );
  XNOR2_X1 U17969 ( .A(n14675), .B(n14674), .ZN(n16066) );
  OAI22_X1 U17970 ( .A1(n16047), .A2(n14677), .B1(n20140), .B2(n14676), .ZN(
        n14680) );
  NOR2_X1 U17971 ( .A1(n14678), .A2(n20142), .ZN(n14679) );
  AOI211_X1 U17972 ( .C1(n16043), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        n14682) );
  OAI21_X1 U17973 ( .B1(n16066), .B2(n20155), .A(n14682), .ZN(P1_U2976) );
  NAND2_X1 U17974 ( .A1(n14684), .A2(n14683), .ZN(n14685) );
  XOR2_X1 U17975 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14685), .Z(
        n14809) );
  INV_X1 U17976 ( .A(n14686), .ZN(n14690) );
  AOI22_X1 U17977 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14687) );
  OAI21_X1 U17978 ( .B1(n14688), .B2(n20141), .A(n14687), .ZN(n14689) );
  AOI21_X1 U17979 ( .B1(n14690), .B2(n20178), .A(n14689), .ZN(n14691) );
  OAI21_X1 U17980 ( .B1(n20155), .B2(n14809), .A(n14691), .ZN(P1_U2977) );
  MUX2_X1 U17981 ( .A(n14693), .B(n14692), .S(n10154), .Z(n14694) );
  XNOR2_X1 U17982 ( .A(n14694), .B(n15889), .ZN(n15891) );
  OAI22_X1 U17983 ( .A1(n16047), .A2(n14695), .B1(n20140), .B2(n15887), .ZN(
        n14698) );
  NOR2_X1 U17984 ( .A1(n14696), .A2(n20142), .ZN(n14697) );
  AOI211_X1 U17985 ( .C1(n16043), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14700) );
  OAI21_X1 U17986 ( .B1(n20155), .B2(n15891), .A(n14700), .ZN(P1_U2978) );
  INV_X1 U17987 ( .A(n14701), .ZN(n14702) );
  NAND2_X1 U17988 ( .A1(n14702), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14703) );
  MUX2_X1 U17989 ( .A(n14704), .B(n14703), .S(n10154), .Z(n14705) );
  XOR2_X1 U17990 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n14705), .Z(
        n14818) );
  AOI22_X1 U17991 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n14706) );
  OAI21_X1 U17992 ( .B1(n14707), .B2(n20141), .A(n14706), .ZN(n14708) );
  AOI21_X1 U17993 ( .B1(n14709), .B2(n20178), .A(n14708), .ZN(n14710) );
  OAI21_X1 U17994 ( .B1(n20155), .B2(n14818), .A(n14710), .ZN(P1_U2979) );
  NOR2_X1 U17995 ( .A1(n10154), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14711) );
  MUX2_X1 U17996 ( .A(n16008), .B(n14711), .S(n14701), .Z(n14712) );
  XNOR2_X1 U17997 ( .A(n14712), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16074) );
  NAND2_X1 U17998 ( .A1(n14713), .A2(n20178), .ZN(n14718) );
  OAI22_X1 U17999 ( .A1(n16047), .A2(n14714), .B1(n20140), .B2(n20966), .ZN(
        n14715) );
  AOI21_X1 U18000 ( .B1(n16043), .B2(n14716), .A(n14715), .ZN(n14717) );
  OAI211_X1 U18001 ( .C1(n16074), .C2(n20155), .A(n14718), .B(n14717), .ZN(
        P1_U2980) );
  OAI21_X1 U18002 ( .B1(n14720), .B2(n14719), .A(n14701), .ZN(n14831) );
  INV_X1 U18003 ( .A(n14721), .ZN(n14726) );
  NOR2_X1 U18004 ( .A1(n20141), .A2(n14722), .ZN(n14725) );
  INV_X1 U18005 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U18006 ( .A1(n20149), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14820) );
  OAI21_X1 U18007 ( .B1(n16047), .B2(n14723), .A(n14820), .ZN(n14724) );
  AOI211_X1 U18008 ( .C1(n14726), .C2(n20178), .A(n14725), .B(n14724), .ZN(
        n14727) );
  OAI21_X1 U18009 ( .B1(n20155), .B2(n14831), .A(n14727), .ZN(P1_U2981) );
  INV_X1 U18010 ( .A(n16026), .ZN(n14729) );
  INV_X1 U18011 ( .A(n14833), .ZN(n14728) );
  NOR2_X1 U18012 ( .A1(n14729), .A2(n14728), .ZN(n16006) );
  AOI21_X1 U18013 ( .B1(n14731), .B2(n16006), .A(n14730), .ZN(n14734) );
  NOR2_X1 U18014 ( .A1(n10154), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14733) );
  NAND2_X1 U18015 ( .A1(n14734), .A2(n16009), .ZN(n14732) );
  OAI21_X1 U18016 ( .B1(n14734), .B2(n14733), .A(n14732), .ZN(n14735) );
  XOR2_X1 U18017 ( .A(n12679), .B(n14735), .Z(n16086) );
  OAI22_X1 U18018 ( .A1(n16047), .A2(n14736), .B1(n20140), .B2(n21244), .ZN(
        n14737) );
  AOI21_X1 U18019 ( .B1(n16043), .B2(n14738), .A(n14737), .ZN(n14739) );
  OAI21_X1 U18020 ( .B1(n14740), .B2(n20142), .A(n14739), .ZN(n14741) );
  AOI21_X1 U18021 ( .B1(n16086), .B2(n16045), .A(n14741), .ZN(n14742) );
  INV_X1 U18022 ( .A(n14742), .ZN(P1_U2982) );
  OR3_X1 U18023 ( .A1(n16006), .A2(n16018), .A3(n14743), .ZN(n14744) );
  XOR2_X1 U18024 ( .A(n14745), .B(n14744), .Z(n16111) );
  NAND2_X1 U18025 ( .A1(n20149), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16108) );
  OAI21_X1 U18026 ( .B1(n16047), .B2(n15953), .A(n16108), .ZN(n14746) );
  AOI21_X1 U18027 ( .B1(n16043), .B2(n15958), .A(n14746), .ZN(n14747) );
  OAI21_X1 U18028 ( .B1(n15955), .B2(n20142), .A(n14747), .ZN(n14748) );
  AOI21_X1 U18029 ( .B1(n16111), .B2(n16045), .A(n14748), .ZN(n14749) );
  INV_X1 U18030 ( .A(n14749), .ZN(P1_U2986) );
  INV_X1 U18031 ( .A(n14751), .ZN(n14755) );
  AOI21_X1 U18032 ( .B1(n12690), .B2(n14753), .A(n14752), .ZN(n14754) );
  AOI211_X1 U18033 ( .C1(n20169), .C2(n14756), .A(n14755), .B(n14754), .ZN(
        n14757) );
  OAI21_X1 U18034 ( .B1(n14758), .B2(n20176), .A(n14757), .ZN(P1_U3001) );
  INV_X1 U18035 ( .A(n14784), .ZN(n14760) );
  NOR3_X1 U18036 ( .A1(n14760), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14759), .ZN(n14764) );
  NAND2_X1 U18037 ( .A1(n20149), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14761) );
  OAI21_X1 U18038 ( .B1(n14762), .B2(n16151), .A(n14761), .ZN(n14763) );
  AOI211_X1 U18039 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14765), .A(
        n14764), .B(n14763), .ZN(n14766) );
  OAI21_X1 U18040 ( .B1(n14767), .B2(n20176), .A(n14766), .ZN(P1_U3002) );
  NOR2_X1 U18041 ( .A1(n14769), .A2(n14768), .ZN(n14775) );
  INV_X1 U18042 ( .A(n14778), .ZN(n14770) );
  NAND2_X1 U18043 ( .A1(n14770), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14771) );
  OAI211_X1 U18044 ( .C1(n14773), .C2(n16151), .A(n14772), .B(n14771), .ZN(
        n14774) );
  AOI21_X1 U18045 ( .B1(n14784), .B2(n14775), .A(n14774), .ZN(n14776) );
  OAI21_X1 U18046 ( .B1(n14777), .B2(n20176), .A(n14776), .ZN(P1_U3003) );
  NOR2_X1 U18047 ( .A1(n14778), .A2(n14783), .ZN(n14782) );
  OAI21_X1 U18048 ( .B1(n14780), .B2(n16151), .A(n14779), .ZN(n14781) );
  AOI211_X1 U18049 ( .C1(n14784), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14785) );
  OAI21_X1 U18050 ( .B1(n14786), .B2(n20176), .A(n14785), .ZN(P1_U3004) );
  OAI21_X1 U18051 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14788), .A(
        n14787), .ZN(n14789) );
  NAND2_X1 U18052 ( .A1(n14789), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14790) );
  OAI211_X1 U18053 ( .C1(n14792), .C2(n16151), .A(n14791), .B(n14790), .ZN(
        n14793) );
  AOI21_X1 U18054 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14796) );
  OAI21_X1 U18055 ( .B1(n14797), .B2(n20176), .A(n14796), .ZN(P1_U3007) );
  OAI22_X1 U18056 ( .A1(n14804), .A2(n15888), .B1(n20140), .B2(n14798), .ZN(
        n14806) );
  INV_X1 U18057 ( .A(n16080), .ZN(n14802) );
  NAND2_X1 U18058 ( .A1(n14800), .A2(n14799), .ZN(n16077) );
  AOI221_X1 U18059 ( .B1(n14802), .B2(n16077), .C1(n14810), .C2(n16077), .A(
        n14801), .ZN(n14816) );
  NAND2_X1 U18060 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14816), .ZN(
        n15896) );
  AOI211_X1 U18061 ( .C1(n15889), .C2(n14804), .A(n14803), .B(n15896), .ZN(
        n14805) );
  AOI211_X1 U18062 ( .C1(n20169), .C2(n14807), .A(n14806), .B(n14805), .ZN(
        n14808) );
  OAI21_X1 U18063 ( .B1(n14809), .B2(n20176), .A(n14808), .ZN(P1_U3009) );
  AOI21_X1 U18064 ( .B1(n14810), .B2(n16077), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16078) );
  INV_X1 U18065 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21172) );
  NOR2_X1 U18066 ( .A1(n20140), .A2(n21172), .ZN(n14811) );
  AOI221_X1 U18067 ( .B1(n16078), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), 
        .C1(n16073), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n14811), .ZN(
        n14812) );
  OAI21_X1 U18068 ( .B1(n16151), .B2(n14813), .A(n14812), .ZN(n14814) );
  AOI21_X1 U18069 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14817) );
  OAI21_X1 U18070 ( .B1(n14818), .B2(n20176), .A(n14817), .ZN(P1_U3011) );
  NAND2_X1 U18071 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14840) );
  NAND3_X1 U18072 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n16100), .ZN(n16091) );
  NOR2_X1 U18073 ( .A1(n14840), .A2(n16091), .ZN(n16084) );
  NAND3_X1 U18074 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16084), .A3(
        n14825), .ZN(n14830) );
  INV_X1 U18075 ( .A(n14819), .ZN(n14828) );
  INV_X1 U18076 ( .A(n14820), .ZN(n14827) );
  INV_X1 U18077 ( .A(n16141), .ZN(n16121) );
  OAI21_X1 U18078 ( .B1(n14822), .B2(n14821), .A(n20157), .ZN(n14823) );
  OAI211_X1 U18079 ( .C1(n16140), .C2(n16139), .A(n16121), .B(n14823), .ZN(
        n16112) );
  AOI21_X1 U18080 ( .B1(n14824), .B2(n20157), .A(n16112), .ZN(n16090) );
  NOR2_X1 U18081 ( .A1(n16090), .A2(n14825), .ZN(n14826) );
  AOI211_X1 U18082 ( .C1(n20169), .C2(n14828), .A(n14827), .B(n14826), .ZN(
        n14829) );
  OAI211_X1 U18083 ( .C1(n14831), .C2(n20176), .A(n14830), .B(n14829), .ZN(
        P1_U3013) );
  INV_X1 U18084 ( .A(n14832), .ZN(n14834) );
  OAI211_X1 U18085 ( .C1(n14835), .C2(n16026), .A(n14834), .B(n14833), .ZN(
        n15998) );
  NOR3_X1 U18086 ( .A1(n15998), .A2(n14836), .A3(n15994), .ZN(n15996) );
  NOR2_X1 U18087 ( .A1(n15994), .A2(n15996), .ZN(n14837) );
  XNOR2_X1 U18088 ( .A(n14838), .B(n14837), .ZN(n15989) );
  INV_X1 U18089 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14839) );
  OAI22_X1 U18090 ( .A1(n15926), .A2(n16151), .B1(n20140), .B2(n14839), .ZN(
        n14843) );
  INV_X1 U18091 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16104) );
  AOI21_X1 U18092 ( .B1(n16104), .B2(n20157), .A(n16112), .ZN(n16099) );
  OAI21_X1 U18093 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n14840), .ZN(n14841) );
  OAI22_X1 U18094 ( .A1(n16099), .A2(n12377), .B1(n16091), .B2(n14841), .ZN(
        n14842) );
  AOI211_X1 U18095 ( .C1(n15989), .C2(n16182), .A(n14843), .B(n14842), .ZN(
        n14844) );
  INV_X1 U18096 ( .A(n14844), .ZN(P1_U3015) );
  NOR2_X1 U18097 ( .A1(n14845), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14848) );
  NOR3_X1 U18098 ( .A1(n14846), .A2(n13377), .A3(n13397), .ZN(n14847) );
  AOI211_X1 U18099 ( .C1(n20660), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n15851) );
  INV_X1 U18100 ( .A(n16188), .ZN(n20837) );
  NOR2_X1 U18101 ( .A1(n16195), .A2(n14850), .ZN(n20834) );
  OAI22_X1 U18102 ( .A1(n12328), .A2(n12694), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20838) );
  NOR3_X1 U18103 ( .A1(n13397), .A2(n13377), .A3(n20841), .ZN(n14851) );
  AOI21_X1 U18104 ( .B1(n20834), .B2(n20838), .A(n14851), .ZN(n14852) );
  OAI21_X1 U18105 ( .B1(n15851), .B2(n20837), .A(n14852), .ZN(n14853) );
  MUX2_X1 U18106 ( .A(n14853), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20842), .Z(P1_U3473) );
  NOR2_X1 U18107 ( .A1(n9992), .A2(n16437), .ZN(n14857) );
  INV_X1 U18108 ( .A(n19877), .ZN(n14855) );
  AOI21_X1 U18109 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n14855), .A(n14854), 
        .ZN(n14856) );
  AOI21_X1 U18110 ( .B1(n14857), .B2(n19877), .A(n14856), .ZN(n14859) );
  OAI22_X1 U18111 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15910), .B1(n19872), 
        .B2(n19798), .ZN(n14858) );
  OAI21_X1 U18112 ( .B1(n14859), .B2(n19863), .A(n14858), .ZN(n14863) );
  OAI21_X1 U18113 ( .B1(n16452), .B2(n19798), .A(n19809), .ZN(n14860) );
  OAI211_X1 U18114 ( .C1(n19872), .C2(n14861), .A(n19043), .B(n14860), .ZN(
        n14862) );
  MUX2_X1 U18115 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n14863), .S(n14862), 
        .Z(P2_U3610) );
  OAI22_X1 U18116 ( .A1(n11084), .A2(n19210), .B1(n19929), .B2(n19179), .ZN(
        n14866) );
  OAI22_X1 U18117 ( .A1(n19202), .A2(n11160), .B1(n14864), .B2(n19141), .ZN(
        n14865) );
  AOI211_X1 U18118 ( .C1(n15199), .C2(n19185), .A(n14866), .B(n14865), .ZN(
        n14870) );
  OAI211_X1 U18119 ( .C1(n14868), .C2(n15195), .A(n19108), .B(n14867), .ZN(
        n14869) );
  OAI211_X1 U18120 ( .C1(n14871), .C2(n19158), .A(n14870), .B(n14869), .ZN(
        P2_U2834) );
  AND2_X1 U18121 ( .A1(n15100), .A2(n14872), .ZN(n14873) );
  OR2_X1 U18122 ( .A1(n14873), .A2(n15082), .ZN(n15366) );
  INV_X1 U18123 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19925) );
  AOI22_X1 U18124 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19183), .B1(n14874), 
        .B2(n19205), .ZN(n14875) );
  OAI211_X1 U18125 ( .C1(n19925), .C2(n19179), .A(n14875), .B(n19170), .ZN(
        n14876) );
  AOI21_X1 U18126 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19167), .A(
        n14876), .ZN(n14883) );
  NAND2_X1 U18127 ( .A1(n19152), .A2(n14877), .ZN(n14878) );
  XNOR2_X1 U18128 ( .A(n15221), .B(n14878), .ZN(n14881) );
  OAI21_X1 U18129 ( .B1(n15008), .B2(n14879), .A(n14993), .ZN(n15361) );
  INV_X1 U18130 ( .A(n15361), .ZN(n14880) );
  AOI22_X1 U18131 ( .A1(n14881), .A2(n19108), .B1(n14880), .B2(n19185), .ZN(
        n14882) );
  OAI211_X1 U18132 ( .C1(n15366), .C2(n19158), .A(n14883), .B(n14882), .ZN(
        P2_U2836) );
  OAI21_X1 U18133 ( .B1(n14885), .B2(n14884), .A(n15101), .ZN(n15389) );
  INV_X1 U18134 ( .A(n15389), .ZN(n15117) );
  NOR2_X1 U18135 ( .A1(n19152), .A2(n19869), .ZN(n19135) );
  INV_X1 U18136 ( .A(n19135), .ZN(n19195) );
  AOI22_X1 U18137 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19197), .ZN(n14886) );
  OAI211_X1 U18138 ( .C1(n15238), .C2(n19195), .A(n14886), .B(n19170), .ZN(
        n14894) );
  NOR2_X1 U18139 ( .A1(n19165), .A2(n14887), .ZN(n19080) );
  OAI211_X1 U18140 ( .C1(n14888), .C2(n15238), .A(n19108), .B(n19080), .ZN(
        n14892) );
  OAI22_X1 U18141 ( .A1(n19202), .A2(n11146), .B1(n14889), .B2(n19141), .ZN(
        n14890) );
  INV_X1 U18142 ( .A(n14890), .ZN(n14891) );
  OAI211_X1 U18143 ( .C1(n19207), .C2(n15391), .A(n14892), .B(n14891), .ZN(
        n14893) );
  AOI211_X1 U18144 ( .C1(n15117), .C2(n19199), .A(n14894), .B(n14893), .ZN(
        n14895) );
  INV_X1 U18145 ( .A(n14895), .ZN(P2_U2838) );
  INV_X1 U18146 ( .A(n14896), .ZN(n15256) );
  NAND2_X1 U18147 ( .A1(n19152), .A2(n14897), .ZN(n14898) );
  XOR2_X1 U18148 ( .A(n15256), .B(n14898), .Z(n14904) );
  INV_X1 U18149 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19917) );
  OAI21_X1 U18150 ( .B1(n19917), .B2(n19179), .A(n19170), .ZN(n14901) );
  OAI22_X1 U18151 ( .A1(n14899), .A2(n19141), .B1(n15257), .B2(n19210), .ZN(
        n14900) );
  AOI211_X1 U18152 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19183), .A(n14901), .B(
        n14900), .ZN(n14902) );
  OAI21_X1 U18153 ( .B1(n15410), .B2(n19207), .A(n14902), .ZN(n14903) );
  AOI21_X1 U18154 ( .B1(n14904), .B2(n19108), .A(n14903), .ZN(n14905) );
  OAI21_X1 U18155 ( .B1(n15408), .B2(n19158), .A(n14905), .ZN(P2_U2840) );
  AOI22_X1 U18156 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19197), .ZN(n14910) );
  OAI22_X1 U18157 ( .A1(n19202), .A2(n14907), .B1(n14906), .B2(n19141), .ZN(
        n14908) );
  AOI21_X1 U18158 ( .B1(n15526), .B2(n19185), .A(n14908), .ZN(n14909) );
  OAI211_X1 U18159 ( .C1(n14911), .C2(n19158), .A(n14910), .B(n14909), .ZN(
        n14917) );
  INV_X1 U18160 ( .A(n14914), .ZN(n14915) );
  NOR2_X1 U18161 ( .A1(n19165), .A2(n14912), .ZN(n15508) );
  INV_X1 U18162 ( .A(n15508), .ZN(n14913) );
  AOI221_X1 U18163 ( .B1(n14915), .B2(n15508), .C1(n14914), .C2(n14913), .A(
        n19869), .ZN(n14916) );
  AOI211_X1 U18164 ( .C1(n19213), .C2(n19448), .A(n14917), .B(n14916), .ZN(
        n14918) );
  INV_X1 U18165 ( .A(n14918), .ZN(P2_U2853) );
  NAND2_X1 U18166 ( .A1(n16205), .A2(n14983), .ZN(n14919) );
  OAI21_X1 U18167 ( .B1(n14983), .B2(n14920), .A(n14919), .ZN(P2_U2856) );
  XNOR2_X1 U18168 ( .A(n14921), .B(n14922), .ZN(n15020) );
  OAI21_X1 U18169 ( .B1(n12783), .B2(n14924), .A(n14923), .ZN(n15265) );
  NOR2_X1 U18170 ( .A1(n15265), .A2(n13301), .ZN(n14925) );
  AOI21_X1 U18171 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n13301), .A(n14925), .ZN(
        n14926) );
  OAI21_X1 U18172 ( .B1(n15020), .B2(n15012), .A(n14926), .ZN(P2_U2858) );
  NOR2_X1 U18173 ( .A1(n10306), .A2(n14927), .ZN(n14928) );
  XOR2_X1 U18174 ( .A(n14929), .B(n14928), .Z(n15026) );
  NOR2_X1 U18175 ( .A1(n16231), .A2(n13301), .ZN(n14930) );
  AOI21_X1 U18176 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15010), .A(n14930), .ZN(
        n14931) );
  OAI21_X1 U18177 ( .B1(n15026), .B2(n15012), .A(n14931), .ZN(P2_U2859) );
  XOR2_X1 U18178 ( .A(n14932), .B(n14943), .Z(n16233) );
  INV_X1 U18179 ( .A(n16233), .ZN(n14938) );
  NAND2_X1 U18180 ( .A1(n15027), .A2(n14961), .ZN(n14937) );
  NAND2_X1 U18181 ( .A1(n15010), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14936) );
  OAI211_X1 U18182 ( .C1(n14938), .C2(n15010), .A(n14937), .B(n14936), .ZN(
        P2_U2860) );
  XNOR2_X1 U18183 ( .A(n14939), .B(n14940), .ZN(n15036) );
  NAND2_X1 U18184 ( .A1(n14952), .A2(n14941), .ZN(n14942) );
  NAND2_X1 U18185 ( .A1(n14943), .A2(n14942), .ZN(n16243) );
  NOR2_X1 U18186 ( .A1(n16243), .A2(n13301), .ZN(n14944) );
  AOI21_X1 U18187 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15010), .A(n14944), .ZN(
        n14945) );
  OAI21_X1 U18188 ( .B1(n15036), .B2(n15012), .A(n14945), .ZN(P2_U2861) );
  OAI21_X1 U18189 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n15045) );
  OR2_X1 U18190 ( .A1(n14949), .A2(n14950), .ZN(n14951) );
  NAND2_X1 U18191 ( .A1(n14952), .A2(n14951), .ZN(n16255) );
  NOR2_X1 U18192 ( .A1(n16255), .A2(n13301), .ZN(n14953) );
  AOI21_X1 U18193 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15010), .A(n14953), .ZN(
        n14954) );
  OAI21_X1 U18194 ( .B1(n15045), .B2(n15012), .A(n14954), .ZN(P2_U2862) );
  INV_X1 U18195 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16267) );
  NOR2_X1 U18196 ( .A1(n14957), .A2(n14956), .ZN(n14958) );
  XNOR2_X1 U18197 ( .A(n14959), .B(n14958), .ZN(n14960) );
  XNOR2_X1 U18198 ( .A(n14955), .B(n14960), .ZN(n16287) );
  NAND2_X1 U18199 ( .A1(n16287), .A2(n14961), .ZN(n14967) );
  NOR2_X1 U18200 ( .A1(n14963), .A2(n14962), .ZN(n14964) );
  OR2_X1 U18201 ( .A1(n14949), .A2(n14964), .ZN(n16275) );
  INV_X1 U18202 ( .A(n16275), .ZN(n14965) );
  NAND2_X1 U18203 ( .A1(n14965), .A2(n15000), .ZN(n14966) );
  OAI211_X1 U18204 ( .C1(n14983), .C2(n16267), .A(n14967), .B(n14966), .ZN(
        P2_U2863) );
  OAI21_X1 U18205 ( .B1(n14968), .B2(n14970), .A(n14969), .ZN(n15061) );
  NAND2_X1 U18206 ( .A1(n13301), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14973) );
  XOR2_X1 U18207 ( .A(n14971), .B(n14982), .Z(n16277) );
  NAND2_X1 U18208 ( .A1(n16277), .A2(n15000), .ZN(n14972) );
  OAI211_X1 U18209 ( .C1(n15061), .C2(n15012), .A(n14973), .B(n14972), .ZN(
        P2_U2864) );
  INV_X1 U18210 ( .A(n14974), .ZN(n14978) );
  INV_X1 U18211 ( .A(n14975), .ZN(n14977) );
  OAI21_X1 U18212 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n15072) );
  NAND2_X1 U18213 ( .A1(n15010), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14985) );
  AND2_X1 U18214 ( .A1(n14980), .A2(n14979), .ZN(n14981) );
  NOR2_X1 U18215 ( .A1(n14982), .A2(n14981), .ZN(n15841) );
  NAND2_X1 U18216 ( .A1(n15841), .A2(n14983), .ZN(n14984) );
  OAI211_X1 U18217 ( .C1(n15072), .C2(n15012), .A(n14985), .B(n14984), .ZN(
        P2_U2865) );
  OR2_X1 U18218 ( .A1(n14986), .A2(n14987), .ZN(n14988) );
  NAND2_X1 U18219 ( .A1(n14974), .A2(n14988), .ZN(n15080) );
  NOR2_X1 U18220 ( .A1(n15000), .A2(n11160), .ZN(n14989) );
  AOI21_X1 U18221 ( .B1(n15199), .B2(n15000), .A(n14989), .ZN(n14990) );
  OAI21_X1 U18222 ( .B1(n15080), .B2(n15012), .A(n14990), .ZN(P2_U2866) );
  AOI21_X1 U18223 ( .B1(n14991), .B2(n9836), .A(n14986), .ZN(n14992) );
  INV_X1 U18224 ( .A(n14992), .ZN(n15091) );
  OAI21_X1 U18225 ( .B1(n9810), .B2(n10335), .A(n14995), .ZN(n19078) );
  MUX2_X1 U18226 ( .A(n11156), .B(n19078), .S(n15000), .Z(n14996) );
  OAI21_X1 U18227 ( .B1(n15091), .B2(n15012), .A(n14996), .ZN(P2_U2867) );
  NAND2_X1 U18228 ( .A1(n14997), .A2(n14998), .ZN(n14999) );
  NAND2_X1 U18229 ( .A1(n9836), .A2(n14999), .ZN(n15099) );
  INV_X1 U18230 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n15001) );
  MUX2_X1 U18231 ( .A(n15001), .B(n15361), .S(n15000), .Z(n15002) );
  OAI21_X1 U18232 ( .B1(n15099), .B2(n15012), .A(n15002), .ZN(P2_U2868) );
  NAND2_X1 U18233 ( .A1(n14049), .A2(n15003), .ZN(n15004) );
  NAND2_X1 U18234 ( .A1(n14997), .A2(n15004), .ZN(n15108) );
  NOR2_X1 U18235 ( .A1(n15006), .A2(n15005), .ZN(n15007) );
  OR2_X1 U18236 ( .A1(n15008), .A2(n15007), .ZN(n19084) );
  NOR2_X1 U18237 ( .A1(n19084), .A2(n13301), .ZN(n15009) );
  AOI21_X1 U18238 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n15010), .A(n15009), .ZN(
        n15011) );
  OAI21_X1 U18239 ( .B1(n15108), .B2(n15012), .A(n15011), .ZN(P2_U2869) );
  XOR2_X1 U18240 ( .A(n15014), .B(n15013), .Z(n16212) );
  AOI22_X1 U18241 ( .A1(n19215), .A2(BUF2_REG_29__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U18242 ( .A1(n19231), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n15015) );
  OAI211_X1 U18243 ( .C1(n15017), .C2(n15110), .A(n15016), .B(n15015), .ZN(
        n15018) );
  AOI21_X1 U18244 ( .B1(n16212), .B2(n19245), .A(n15018), .ZN(n15019) );
  OAI21_X1 U18245 ( .B1(n15020), .B2(n15120), .A(n15019), .ZN(P2_U2890) );
  AOI22_X1 U18246 ( .A1(n16286), .A2(n19224), .B1(n19231), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U18247 ( .A1(n19215), .A2(BUF2_REG_28__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15021) );
  OAI211_X1 U18248 ( .C1(n16222), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15024) );
  INV_X1 U18249 ( .A(n15024), .ZN(n15025) );
  OAI21_X1 U18250 ( .B1(n15026), .B2(n15120), .A(n15025), .ZN(P2_U2891) );
  NAND2_X1 U18251 ( .A1(n15027), .A2(n19246), .ZN(n15035) );
  AOI22_X1 U18252 ( .A1(n16286), .A2(n15028), .B1(n19231), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15034) );
  AOI22_X1 U18253 ( .A1(n19215), .A2(BUF2_REG_27__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15033) );
  AND2_X1 U18254 ( .A1(n9845), .A2(n15029), .ZN(n15030) );
  NOR2_X1 U18255 ( .A1(n15031), .A2(n15030), .ZN(n16234) );
  NAND2_X1 U18256 ( .A1(n16234), .A2(n19245), .ZN(n15032) );
  NAND4_X1 U18257 ( .A1(n15035), .A2(n15034), .A3(n15033), .A4(n15032), .ZN(
        P2_U2892) );
  OR2_X1 U18258 ( .A1(n15036), .A2(n15120), .ZN(n15044) );
  AOI22_X1 U18259 ( .A1(n16286), .A2(n15037), .B1(n19231), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U18260 ( .A1(n19215), .A2(BUF2_REG_26__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15042) );
  NAND2_X1 U18261 ( .A1(n15039), .A2(n15038), .ZN(n15040) );
  AND2_X1 U18262 ( .A1(n9845), .A2(n15040), .ZN(n16245) );
  NAND2_X1 U18263 ( .A1(n16245), .A2(n19245), .ZN(n15041) );
  NAND4_X1 U18264 ( .A1(n15044), .A2(n15043), .A3(n15042), .A4(n15041), .ZN(
        P2_U2893) );
  OR2_X1 U18265 ( .A1(n15045), .A2(n15120), .ZN(n15052) );
  AOI22_X1 U18266 ( .A1(n16286), .A2(n15046), .B1(n19231), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15051) );
  AOI22_X1 U18267 ( .A1(n19215), .A2(BUF2_REG_25__SCAN_IN), .B1(n19217), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15050) );
  INV_X1 U18268 ( .A(n15047), .ZN(n15048) );
  XNOR2_X1 U18269 ( .A(n15309), .B(n15048), .ZN(n16257) );
  NAND2_X1 U18270 ( .A1(n16257), .A2(n19245), .ZN(n15049) );
  NAND4_X1 U18271 ( .A1(n15052), .A2(n15051), .A3(n15050), .A4(n15049), .ZN(
        P2_U2894) );
  INV_X1 U18272 ( .A(n15310), .ZN(n15053) );
  AOI21_X1 U18273 ( .B1(n15054), .B2(n15062), .A(n15053), .ZN(n16278) );
  OAI22_X1 U18274 ( .A1(n15110), .A2(n19354), .B1(n19249), .B2(n15055), .ZN(
        n15059) );
  INV_X1 U18275 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15057) );
  INV_X1 U18276 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n15056) );
  OAI22_X1 U18277 ( .A1(n15114), .A2(n15057), .B1(n15112), .B2(n15056), .ZN(
        n15058) );
  AOI211_X1 U18278 ( .C1(n16278), .C2(n19245), .A(n15059), .B(n15058), .ZN(
        n15060) );
  OAI21_X1 U18279 ( .B1(n15120), .B2(n15061), .A(n15060), .ZN(P2_U2896) );
  INV_X1 U18280 ( .A(n15062), .ZN(n15063) );
  AOI21_X1 U18281 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15842) );
  OAI22_X1 U18282 ( .A1(n15110), .A2(n19346), .B1(n19249), .B2(n15066), .ZN(
        n15070) );
  INV_X1 U18283 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15068) );
  INV_X1 U18284 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n15067) );
  OAI22_X1 U18285 ( .A1(n15114), .A2(n15068), .B1(n15112), .B2(n15067), .ZN(
        n15069) );
  AOI211_X1 U18286 ( .C1(n15842), .C2(n19245), .A(n15070), .B(n15069), .ZN(
        n15071) );
  OAI21_X1 U18287 ( .B1(n15120), .B2(n15072), .A(n15071), .ZN(P2_U2897) );
  OAI22_X1 U18288 ( .A1(n15110), .A2(n19343), .B1(n19249), .B2(n15073), .ZN(
        n15077) );
  INV_X1 U18289 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15075) );
  INV_X1 U18290 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15074) );
  OAI22_X1 U18291 ( .A1(n15114), .A2(n15075), .B1(n15112), .B2(n15074), .ZN(
        n15076) );
  AOI211_X1 U18292 ( .C1(n15078), .C2(n19245), .A(n15077), .B(n15076), .ZN(
        n15079) );
  OAI21_X1 U18293 ( .B1(n15120), .B2(n15080), .A(n15079), .ZN(P2_U2898) );
  NOR2_X1 U18294 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  OR2_X1 U18295 ( .A1(n15084), .A2(n15083), .ZN(n15353) );
  INV_X1 U18296 ( .A(n15353), .ZN(n19072) );
  OAI22_X1 U18297 ( .A1(n15110), .A2(n19340), .B1(n19249), .B2(n15085), .ZN(
        n15089) );
  INV_X1 U18298 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15087) );
  INV_X1 U18299 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n15086) );
  OAI22_X1 U18300 ( .A1(n15114), .A2(n15087), .B1(n15112), .B2(n15086), .ZN(
        n15088) );
  AOI211_X1 U18301 ( .C1(n19072), .C2(n19245), .A(n15089), .B(n15088), .ZN(
        n15090) );
  OAI21_X1 U18302 ( .B1(n15120), .B2(n15091), .A(n15090), .ZN(P2_U2899) );
  INV_X1 U18303 ( .A(n15366), .ZN(n15097) );
  OAI22_X1 U18304 ( .A1(n15110), .A2(n19336), .B1(n19249), .B2(n15092), .ZN(
        n15096) );
  INV_X1 U18305 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15094) );
  INV_X1 U18306 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15093) );
  OAI22_X1 U18307 ( .A1(n15114), .A2(n15094), .B1(n15112), .B2(n15093), .ZN(
        n15095) );
  AOI211_X1 U18308 ( .C1(n15097), .C2(n19245), .A(n15096), .B(n15095), .ZN(
        n15098) );
  OAI21_X1 U18309 ( .B1(n15120), .B2(n15099), .A(n15098), .ZN(P2_U2900) );
  AOI21_X1 U18310 ( .B1(n15102), .B2(n15101), .A(n11425), .ZN(n19086) );
  OAI22_X1 U18311 ( .A1(n15110), .A2(n19333), .B1(n19249), .B2(n15103), .ZN(
        n15106) );
  INV_X1 U18312 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15104) );
  OAI22_X1 U18313 ( .A1(n15114), .A2(n15104), .B1(n15112), .B2(n20199), .ZN(
        n15105) );
  AOI211_X1 U18314 ( .C1(n19086), .C2(n19245), .A(n15106), .B(n15105), .ZN(
        n15107) );
  OAI21_X1 U18315 ( .B1(n15120), .B2(n15108), .A(n15107), .ZN(P2_U2901) );
  OAI22_X1 U18316 ( .A1(n15110), .A2(n19329), .B1(n19249), .B2(n15109), .ZN(
        n15116) );
  INV_X1 U18317 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15113) );
  INV_X1 U18318 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n15111) );
  OAI22_X1 U18319 ( .A1(n15114), .A2(n15113), .B1(n15112), .B2(n15111), .ZN(
        n15115) );
  AOI211_X1 U18320 ( .C1(n15117), .C2(n19245), .A(n15116), .B(n15115), .ZN(
        n15118) );
  OAI21_X1 U18321 ( .B1(n15120), .B2(n15119), .A(n15118), .ZN(P2_U2902) );
  INV_X1 U18322 ( .A(n15121), .ZN(n15122) );
  OAI21_X1 U18323 ( .B1(n15123), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15122), .ZN(n15274) );
  NAND2_X1 U18324 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  XNOR2_X1 U18325 ( .A(n15127), .B(n15126), .ZN(n15271) );
  NOR2_X1 U18326 ( .A1(n19170), .A2(n19944), .ZN(n15266) );
  AOI21_X1 U18327 ( .B1(n19287), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15266), .ZN(n15130) );
  NAND2_X1 U18328 ( .A1(n16355), .A2(n15128), .ZN(n15129) );
  OAI211_X1 U18329 ( .C1(n15265), .C2(n15258), .A(n15130), .B(n15129), .ZN(
        n15131) );
  AOI21_X1 U18330 ( .B1(n15271), .B2(n19291), .A(n15131), .ZN(n15132) );
  OAI21_X1 U18331 ( .B1(n15274), .B2(n16358), .A(n15132), .ZN(P2_U2985) );
  NAND2_X1 U18332 ( .A1(n12775), .A2(n12774), .ZN(n15275) );
  NAND3_X1 U18333 ( .A1(n15276), .A2(n10925), .A3(n15275), .ZN(n15141) );
  NAND2_X1 U18334 ( .A1(n16355), .A2(n15133), .ZN(n15134) );
  NAND2_X1 U18335 ( .A1(n19286), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15279) );
  OAI211_X1 U18336 ( .C1(n16365), .C2(n15135), .A(n15134), .B(n15279), .ZN(
        n15136) );
  AOI21_X1 U18337 ( .B1(n16233), .B2(n19290), .A(n15136), .ZN(n15140) );
  OR2_X1 U18338 ( .A1(n15137), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15283) );
  NAND3_X1 U18339 ( .A1(n15283), .A2(n15138), .A3(n19291), .ZN(n15139) );
  NAND3_X1 U18340 ( .A1(n15141), .A2(n15140), .A3(n15139), .ZN(P2_U2987) );
  OAI21_X1 U18341 ( .B1(n15142), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12775), .ZN(n15297) );
  NAND2_X1 U18342 ( .A1(n15153), .A2(n15150), .ZN(n15143) );
  NAND2_X1 U18343 ( .A1(n15143), .A2(n15151), .ZN(n15145) );
  XNOR2_X1 U18344 ( .A(n15145), .B(n15144), .ZN(n15294) );
  INV_X1 U18345 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19938) );
  NOR2_X1 U18346 ( .A1(n19170), .A2(n19938), .ZN(n15290) );
  NOR2_X1 U18347 ( .A1(n19296), .A2(n16248), .ZN(n15146) );
  AOI211_X1 U18348 ( .C1(n19287), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15290), .B(n15146), .ZN(n15147) );
  OAI21_X1 U18349 ( .B1(n16243), .B2(n15258), .A(n15147), .ZN(n15148) );
  AOI21_X1 U18350 ( .B1(n15294), .B2(n19291), .A(n15148), .ZN(n15149) );
  OAI21_X1 U18351 ( .B1(n15297), .B2(n16358), .A(n15149), .ZN(P2_U2988) );
  NAND2_X1 U18352 ( .A1(n15151), .A2(n15150), .ZN(n15152) );
  XNOR2_X1 U18353 ( .A(n15153), .B(n15152), .ZN(n15308) );
  INV_X1 U18354 ( .A(n15154), .ZN(n15163) );
  AOI21_X1 U18355 ( .B1(n15155), .B2(n15163), .A(n15142), .ZN(n15298) );
  NAND2_X1 U18356 ( .A1(n15298), .A2(n10925), .ZN(n15161) );
  NAND2_X1 U18357 ( .A1(n19286), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15299) );
  OAI21_X1 U18358 ( .B1(n16365), .B2(n15156), .A(n15299), .ZN(n15158) );
  NOR2_X1 U18359 ( .A1(n16255), .A2(n15258), .ZN(n15157) );
  AOI211_X1 U18360 ( .C1(n16355), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15160) );
  OAI211_X1 U18361 ( .C1(n16356), .C2(n15308), .A(n15161), .B(n15160), .ZN(
        P2_U2989) );
  INV_X1 U18362 ( .A(n15162), .ZN(n15164) );
  OAI21_X1 U18363 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15164), .A(
        n15163), .ZN(n15321) );
  NAND2_X1 U18364 ( .A1(n9890), .A2(n15165), .ZN(n15166) );
  XNOR2_X1 U18365 ( .A(n15167), .B(n15166), .ZN(n15318) );
  INV_X1 U18366 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19934) );
  NOR2_X1 U18367 ( .A1(n19170), .A2(n19934), .ZN(n15314) );
  NOR2_X1 U18368 ( .A1(n19296), .A2(n16272), .ZN(n15168) );
  AOI211_X1 U18369 ( .C1(n19287), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15314), .B(n15168), .ZN(n15169) );
  OAI21_X1 U18370 ( .B1(n16275), .B2(n15258), .A(n15169), .ZN(n15170) );
  AOI21_X1 U18371 ( .B1(n15318), .B2(n19291), .A(n15170), .ZN(n15171) );
  OAI21_X1 U18372 ( .B1(n15321), .B2(n16358), .A(n15171), .ZN(P2_U2990) );
  OAI21_X1 U18373 ( .B1(n15172), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15162), .ZN(n15334) );
  NAND2_X1 U18374 ( .A1(n16355), .A2(n15173), .ZN(n15174) );
  NAND2_X1 U18375 ( .A1(n19286), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15322) );
  OAI211_X1 U18376 ( .C1(n16365), .C2(n15175), .A(n15174), .B(n15322), .ZN(
        n15183) );
  NAND2_X1 U18377 ( .A1(n15176), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15177) );
  XNOR2_X1 U18378 ( .A(n15178), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15180) );
  NOR2_X1 U18379 ( .A1(n15179), .A2(n15180), .ZN(n15330) );
  INV_X1 U18380 ( .A(n15180), .ZN(n15181) );
  NOR3_X1 U18381 ( .A1(n15330), .A2(n15329), .A3(n16356), .ZN(n15182) );
  AOI211_X1 U18382 ( .C1(n19290), .C2(n16277), .A(n15183), .B(n15182), .ZN(
        n15184) );
  OAI21_X1 U18383 ( .B1(n15334), .B2(n16358), .A(n15184), .ZN(P2_U2991) );
  INV_X1 U18384 ( .A(n15172), .ZN(n15185) );
  OAI21_X1 U18385 ( .B1(n11473), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15185), .ZN(n15345) );
  XNOR2_X1 U18386 ( .A(n15186), .B(n15340), .ZN(n15187) );
  XNOR2_X1 U18387 ( .A(n15176), .B(n15187), .ZN(n15343) );
  NAND2_X1 U18388 ( .A1(n15841), .A2(n19290), .ZN(n15190) );
  INV_X1 U18389 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15188) );
  NOR2_X1 U18390 ( .A1(n19170), .A2(n15188), .ZN(n15337) );
  AOI21_X1 U18391 ( .B1(n19287), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15337), .ZN(n15189) );
  OAI211_X1 U18392 ( .C1(n19296), .C2(n15844), .A(n15190), .B(n15189), .ZN(
        n15191) );
  AOI21_X1 U18393 ( .B1(n15343), .B2(n19291), .A(n15191), .ZN(n15192) );
  OAI21_X1 U18394 ( .B1(n15345), .B2(n16358), .A(n15192), .ZN(P2_U2992) );
  NAND2_X1 U18395 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15193) );
  OAI211_X1 U18396 ( .C1(n19296), .C2(n15195), .A(n15194), .B(n15193), .ZN(
        n15198) );
  NOR3_X1 U18397 ( .A1(n15196), .A2(n11473), .A3(n16358), .ZN(n15197) );
  AOI211_X1 U18398 ( .C1(n19290), .C2(n15199), .A(n15198), .B(n15197), .ZN(
        n15200) );
  OAI21_X1 U18399 ( .B1(n15201), .B2(n16356), .A(n15200), .ZN(P2_U2993) );
  NAND2_X1 U18400 ( .A1(n15203), .A2(n15202), .ZN(n15207) );
  NAND2_X1 U18401 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  XNOR2_X1 U18402 ( .A(n15207), .B(n15206), .ZN(n15357) );
  AOI21_X1 U18403 ( .B1(n15208), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15209) );
  NOR2_X1 U18404 ( .A1(n15209), .A2(n9854), .ZN(n15355) );
  NOR2_X1 U18405 ( .A1(n19170), .A2(n19927), .ZN(n15347) );
  NOR2_X1 U18406 ( .A1(n19296), .A2(n19075), .ZN(n15210) );
  AOI211_X1 U18407 ( .C1(n19287), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15347), .B(n15210), .ZN(n15211) );
  OAI21_X1 U18408 ( .B1(n19078), .B2(n15258), .A(n15211), .ZN(n15212) );
  AOI21_X1 U18409 ( .B1(n15355), .B2(n10925), .A(n15212), .ZN(n15213) );
  OAI21_X1 U18410 ( .B1(n15357), .B2(n16356), .A(n15213), .ZN(P2_U2994) );
  NAND2_X1 U18411 ( .A1(n15215), .A2(n15214), .ZN(n15218) );
  INV_X1 U18412 ( .A(n15226), .ZN(n15216) );
  AOI21_X1 U18413 ( .B1(n15228), .B2(n15225), .A(n15216), .ZN(n15217) );
  XOR2_X1 U18414 ( .A(n15218), .B(n15217), .Z(n15370) );
  XNOR2_X1 U18415 ( .A(n15208), .B(n15363), .ZN(n15368) );
  NAND2_X1 U18416 ( .A1(n19286), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15359) );
  OAI21_X1 U18417 ( .B1(n16365), .B2(n15219), .A(n15359), .ZN(n15220) );
  AOI21_X1 U18418 ( .B1(n15221), .B2(n16355), .A(n15220), .ZN(n15222) );
  OAI21_X1 U18419 ( .B1(n15361), .B2(n15258), .A(n15222), .ZN(n15223) );
  AOI21_X1 U18420 ( .B1(n15368), .B2(n10925), .A(n15223), .ZN(n15224) );
  OAI21_X1 U18421 ( .B1(n15370), .B2(n16356), .A(n15224), .ZN(P2_U2995) );
  NAND2_X1 U18422 ( .A1(n15226), .A2(n15225), .ZN(n15227) );
  XNOR2_X1 U18423 ( .A(n15228), .B(n15227), .ZN(n15379) );
  AOI21_X1 U18424 ( .B1(n15382), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15230) );
  NOR2_X1 U18425 ( .A1(n15230), .A2(n15208), .ZN(n15376) );
  NOR2_X1 U18426 ( .A1(n19084), .A2(n15258), .ZN(n15233) );
  NAND2_X1 U18427 ( .A1(n19286), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15372) );
  NAND2_X1 U18428 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15231) );
  OAI211_X1 U18429 ( .C1(n19296), .C2(n19079), .A(n15372), .B(n15231), .ZN(
        n15232) );
  AOI211_X1 U18430 ( .C1(n15376), .C2(n10925), .A(n15233), .B(n15232), .ZN(
        n15234) );
  OAI21_X1 U18431 ( .B1(n15379), .B2(n16356), .A(n15234), .ZN(P2_U2996) );
  XOR2_X1 U18432 ( .A(n15236), .B(n15235), .Z(n15398) );
  NOR2_X1 U18433 ( .A1(n15391), .A2(n15258), .ZN(n15240) );
  NAND2_X1 U18434 ( .A1(n19286), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15390) );
  NAND2_X1 U18435 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15237) );
  OAI211_X1 U18436 ( .C1(n19296), .C2(n15238), .A(n15390), .B(n15237), .ZN(
        n15239) );
  AOI211_X1 U18437 ( .C1(n15241), .C2(n10925), .A(n15240), .B(n15239), .ZN(
        n15242) );
  OAI21_X1 U18438 ( .B1(n15398), .B2(n16356), .A(n15242), .ZN(P2_U2997) );
  XNOR2_X1 U18439 ( .A(n15244), .B(n15243), .ZN(n15407) );
  INV_X1 U18440 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19919) );
  NOR2_X1 U18441 ( .A1(n19919), .A2(n19170), .ZN(n15246) );
  INV_X1 U18442 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19093) );
  OAI22_X1 U18443 ( .A1(n16365), .A2(n19093), .B1(n19296), .B2(n19091), .ZN(
        n15245) );
  AOI211_X1 U18444 ( .C1(n19290), .C2(n19097), .A(n15246), .B(n15245), .ZN(
        n15249) );
  INV_X1 U18445 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15399) );
  OAI21_X1 U18446 ( .B1(n9852), .B2(n15385), .A(n15399), .ZN(n15247) );
  OAI211_X1 U18447 ( .C1(n15407), .C2(n16356), .A(n15249), .B(n15248), .ZN(
        P2_U2998) );
  XNOR2_X1 U18448 ( .A(n9852), .B(n15385), .ZN(n15420) );
  NAND2_X1 U18449 ( .A1(n15251), .A2(n15250), .ZN(n15255) );
  INV_X1 U18450 ( .A(n16295), .ZN(n15252) );
  NOR2_X1 U18451 ( .A1(n15253), .A2(n15252), .ZN(n15254) );
  XOR2_X1 U18452 ( .A(n15255), .B(n15254), .Z(n15418) );
  OAI22_X1 U18453 ( .A1(n16365), .A2(n15257), .B1(n19296), .B2(n15256), .ZN(
        n15260) );
  OAI22_X1 U18454 ( .A1(n15258), .A2(n15410), .B1(n19917), .B2(n19170), .ZN(
        n15259) );
  AOI211_X1 U18455 ( .C1(n15418), .C2(n19291), .A(n15260), .B(n15259), .ZN(
        n15261) );
  OAI21_X1 U18456 ( .B1(n16358), .B2(n15420), .A(n15261), .ZN(P2_U2999) );
  INV_X1 U18457 ( .A(n15277), .ZN(n15263) );
  OAI211_X1 U18458 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15264), .A(
        n15263), .B(n15262), .ZN(n15268) );
  INV_X1 U18459 ( .A(n15265), .ZN(n16211) );
  AOI21_X1 U18460 ( .B1(n16211), .B2(n16390), .A(n15266), .ZN(n15267) );
  OAI211_X1 U18461 ( .C1(n15280), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        n15270) );
  AOI21_X1 U18462 ( .B1(n16212), .B2(n19308), .A(n15270), .ZN(n15273) );
  NAND2_X1 U18463 ( .A1(n15271), .A2(n16391), .ZN(n15272) );
  OAI211_X1 U18464 ( .C1(n15274), .C2(n19311), .A(n15273), .B(n15272), .ZN(
        P2_U3017) );
  NAND3_X1 U18465 ( .A1(n15276), .A2(n16388), .A3(n15275), .ZN(n15286) );
  NOR2_X1 U18466 ( .A1(n15277), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15282) );
  NAND2_X1 U18467 ( .A1(n16233), .A2(n16390), .ZN(n15278) );
  OAI211_X1 U18468 ( .C1(n15280), .C2(n12774), .A(n15279), .B(n15278), .ZN(
        n15281) );
  AOI211_X1 U18469 ( .C1(n16234), .C2(n19308), .A(n15282), .B(n15281), .ZN(
        n15285) );
  NAND3_X1 U18470 ( .A1(n15283), .A2(n15138), .A3(n16391), .ZN(n15284) );
  NAND3_X1 U18471 ( .A1(n15286), .A2(n15285), .A3(n15284), .ZN(P2_U3019) );
  NOR2_X1 U18472 ( .A1(n15287), .A2(n15452), .ZN(n15312) );
  NAND2_X1 U18473 ( .A1(n15312), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15292) );
  XNOR2_X1 U18474 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15288) );
  NAND2_X1 U18475 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15313), .ZN(
        n15300) );
  NOR2_X1 U18476 ( .A1(n15288), .A2(n15300), .ZN(n15289) );
  NOR2_X1 U18477 ( .A1(n15290), .A2(n15289), .ZN(n15291) );
  OAI211_X1 U18478 ( .C1(n16243), .C2(n19305), .A(n15292), .B(n15291), .ZN(
        n15293) );
  AOI21_X1 U18479 ( .B1(n16245), .B2(n19308), .A(n15293), .ZN(n15296) );
  NAND2_X1 U18480 ( .A1(n15294), .A2(n16391), .ZN(n15295) );
  OAI211_X1 U18481 ( .C1(n15297), .C2(n19311), .A(n15296), .B(n15295), .ZN(
        P2_U3020) );
  NAND2_X1 U18482 ( .A1(n15298), .A2(n16388), .ZN(n15307) );
  NAND2_X1 U18483 ( .A1(n15312), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15304) );
  INV_X1 U18484 ( .A(n16255), .ZN(n15302) );
  OAI21_X1 U18485 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15300), .A(
        n15299), .ZN(n15301) );
  AOI21_X1 U18486 ( .B1(n15302), .B2(n16390), .A(n15301), .ZN(n15303) );
  NAND2_X1 U18487 ( .A1(n15304), .A2(n15303), .ZN(n15305) );
  AOI21_X1 U18488 ( .B1(n16257), .B2(n19308), .A(n15305), .ZN(n15306) );
  OAI211_X1 U18489 ( .C1(n15308), .C2(n19300), .A(n15307), .B(n15306), .ZN(
        P2_U3021) );
  AOI21_X1 U18490 ( .B1(n15311), .B2(n15310), .A(n15309), .ZN(n16288) );
  OAI21_X1 U18491 ( .B1(n15313), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15312), .ZN(n15316) );
  INV_X1 U18492 ( .A(n15314), .ZN(n15315) );
  OAI211_X1 U18493 ( .C1(n16275), .C2(n19305), .A(n15316), .B(n15315), .ZN(
        n15317) );
  AOI21_X1 U18494 ( .B1(n16288), .B2(n19308), .A(n15317), .ZN(n15320) );
  NAND2_X1 U18495 ( .A1(n15318), .A2(n16391), .ZN(n15319) );
  OAI211_X1 U18496 ( .C1(n15321), .C2(n19311), .A(n15320), .B(n15319), .ZN(
        P2_U3022) );
  INV_X1 U18497 ( .A(n15322), .ZN(n15326) );
  NOR3_X1 U18498 ( .A1(n15335), .A2(n15324), .A3(n15323), .ZN(n15325) );
  AOI211_X1 U18499 ( .C1(n16390), .C2(n16277), .A(n15326), .B(n15325), .ZN(
        n15327) );
  OAI21_X1 U18500 ( .B1(n15328), .B2(n15341), .A(n15327), .ZN(n15332) );
  NOR3_X1 U18501 ( .A1(n15330), .A2(n15329), .A3(n19300), .ZN(n15331) );
  AOI211_X1 U18502 ( .C1(n19308), .C2(n16278), .A(n15332), .B(n15331), .ZN(
        n15333) );
  OAI21_X1 U18503 ( .B1(n15334), .B2(n19311), .A(n15333), .ZN(P2_U3023) );
  NAND2_X1 U18504 ( .A1(n15842), .A2(n19308), .ZN(n15339) );
  NOR2_X1 U18505 ( .A1(n15335), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15336) );
  AOI211_X1 U18506 ( .C1(n15841), .C2(n16390), .A(n15337), .B(n15336), .ZN(
        n15338) );
  OAI211_X1 U18507 ( .C1(n15341), .C2(n15340), .A(n15339), .B(n15338), .ZN(
        n15342) );
  AOI21_X1 U18508 ( .B1(n16391), .B2(n15343), .A(n15342), .ZN(n15344) );
  OAI21_X1 U18509 ( .B1(n15345), .B2(n19311), .A(n15344), .ZN(P2_U3024) );
  INV_X1 U18510 ( .A(n19078), .ZN(n15348) );
  AND3_X1 U18511 ( .A1(n15358), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15424), .ZN(n15346) );
  AOI211_X1 U18512 ( .C1(n15348), .C2(n16390), .A(n15347), .B(n15346), .ZN(
        n15352) );
  INV_X1 U18513 ( .A(n15349), .ZN(n15350) );
  OAI211_X1 U18514 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15364), .B(n15350), .ZN(
        n15351) );
  OAI211_X1 U18515 ( .C1(n15353), .C2(n16400), .A(n15352), .B(n15351), .ZN(
        n15354) );
  AOI21_X1 U18516 ( .B1(n15355), .B2(n16388), .A(n15354), .ZN(n15356) );
  OAI21_X1 U18517 ( .B1(n15357), .B2(n19300), .A(n15356), .ZN(P2_U3026) );
  NAND3_X1 U18518 ( .A1(n15358), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15424), .ZN(n15360) );
  OAI211_X1 U18519 ( .C1(n15361), .C2(n19305), .A(n15360), .B(n15359), .ZN(
        n15362) );
  AOI21_X1 U18520 ( .B1(n15364), .B2(n15363), .A(n15362), .ZN(n15365) );
  OAI21_X1 U18521 ( .B1(n15366), .B2(n16400), .A(n15365), .ZN(n15367) );
  AOI21_X1 U18522 ( .B1(n15368), .B2(n16388), .A(n15367), .ZN(n15369) );
  OAI21_X1 U18523 ( .B1(n15370), .B2(n19300), .A(n15369), .ZN(P2_U3027) );
  NOR4_X1 U18524 ( .A1(n15415), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15394), .A4(n15388), .ZN(n15375) );
  NAND3_X1 U18525 ( .A1(n15380), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n10890), .ZN(n15371) );
  NAND3_X1 U18526 ( .A1(n15371), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15424), .ZN(n15373) );
  OAI211_X1 U18527 ( .C1(n19084), .C2(n19305), .A(n15373), .B(n15372), .ZN(
        n15374) );
  AOI211_X1 U18528 ( .C1(n19086), .C2(n19308), .A(n15375), .B(n15374), .ZN(
        n15378) );
  NAND2_X1 U18529 ( .A1(n15376), .A2(n16388), .ZN(n15377) );
  OAI211_X1 U18530 ( .C1(n15379), .C2(n19300), .A(n15378), .B(n15377), .ZN(
        P2_U3028) );
  NOR2_X1 U18531 ( .A1(n15380), .A2(n15452), .ZN(n15409) );
  INV_X1 U18532 ( .A(n15381), .ZN(n15383) );
  AOI21_X1 U18533 ( .B1(n19311), .B2(n15383), .A(n15382), .ZN(n15384) );
  NAND2_X1 U18534 ( .A1(n15387), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15397) );
  NOR2_X1 U18535 ( .A1(n15389), .A2(n16400), .ZN(n15393) );
  OAI21_X1 U18536 ( .B1(n19305), .B2(n15391), .A(n15390), .ZN(n15392) );
  AOI211_X1 U18537 ( .C1(n15395), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15396) );
  OAI211_X1 U18538 ( .C1(n15398), .C2(n19300), .A(n15397), .B(n15396), .ZN(
        P2_U3029) );
  OAI21_X1 U18539 ( .B1(n9852), .B2(n19311), .A(n15415), .ZN(n15400) );
  NAND3_X1 U18540 ( .A1(n15400), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15399), .ZN(n15402) );
  AOI22_X1 U18541 ( .A1(n16390), .A2(n19097), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19286), .ZN(n15401) );
  OAI211_X1 U18542 ( .C1(n16400), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        n15404) );
  AOI21_X1 U18543 ( .B1(n15405), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15404), .ZN(n15406) );
  OAI21_X1 U18544 ( .B1(n19300), .B2(n15407), .A(n15406), .ZN(P2_U3030) );
  NOR2_X1 U18545 ( .A1(n15408), .A2(n16400), .ZN(n15417) );
  NAND2_X1 U18546 ( .A1(n15409), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15414) );
  INV_X1 U18547 ( .A(n15410), .ZN(n15412) );
  NOR2_X1 U18548 ( .A1(n19917), .A2(n19170), .ZN(n15411) );
  AOI21_X1 U18549 ( .B1(n16390), .B2(n15412), .A(n15411), .ZN(n15413) );
  OAI211_X1 U18550 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15415), .A(
        n15414), .B(n15413), .ZN(n15416) );
  AOI211_X1 U18551 ( .C1(n15418), .C2(n16391), .A(n15417), .B(n15416), .ZN(
        n15419) );
  OAI21_X1 U18552 ( .B1(n19311), .B2(n15420), .A(n15419), .ZN(P2_U3031) );
  OAI21_X1 U18553 ( .B1(n15421), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16293), .ZN(n16306) );
  XNOR2_X1 U18554 ( .A(n15423), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15433) );
  AND2_X1 U18555 ( .A1(n15425), .A2(n15424), .ZN(n16369) );
  NAND2_X1 U18556 ( .A1(n16369), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15427) );
  AOI22_X1 U18557 ( .A1(n16390), .A2(n16308), .B1(P2_REIP_REG_13__SCAN_IN), 
        .B2(n19286), .ZN(n15426) );
  OAI211_X1 U18558 ( .C1(n16400), .C2(n15428), .A(n15427), .B(n15426), .ZN(
        n15432) );
  OAI22_X1 U18559 ( .A1(n15430), .A2(n16298), .B1(n9871), .B2(n15429), .ZN(
        n16305) );
  NOR2_X1 U18560 ( .A1(n16305), .A2(n19300), .ZN(n15431) );
  AOI211_X1 U18561 ( .C1(n16377), .C2(n15433), .A(n15432), .B(n15431), .ZN(
        n15434) );
  OAI21_X1 U18562 ( .B1(n19311), .B2(n16306), .A(n15434), .ZN(P2_U3033) );
  AOI21_X1 U18563 ( .B1(n15443), .B2(n9855), .A(n15421), .ZN(n16313) );
  INV_X1 U18564 ( .A(n16313), .ZN(n15448) );
  INV_X1 U18565 ( .A(n15435), .ZN(n15436) );
  NOR2_X1 U18566 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  XNOR2_X1 U18567 ( .A(n15439), .B(n15438), .ZN(n16312) );
  XNOR2_X1 U18568 ( .A(n15441), .B(n15440), .ZN(n19226) );
  INV_X1 U18569 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19912) );
  NOR2_X1 U18570 ( .A1(n19912), .A2(n19170), .ZN(n15442) );
  AOI221_X1 U18571 ( .B1(n16369), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C1(n16377), .C2(n15443), .A(n15442), .ZN(n15445) );
  NAND2_X1 U18572 ( .A1(n16390), .A2(n19117), .ZN(n15444) );
  OAI211_X1 U18573 ( .C1(n19226), .C2(n16400), .A(n15445), .B(n15444), .ZN(
        n15446) );
  AOI21_X1 U18574 ( .B1(n16312), .B2(n16391), .A(n15446), .ZN(n15447) );
  OAI21_X1 U18575 ( .B1(n15448), .B2(n19311), .A(n15447), .ZN(P2_U3034) );
  OAI21_X1 U18576 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n9829), .A(
        n9855), .ZN(n16317) );
  XNOR2_X1 U18577 ( .A(n15449), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15450) );
  XNOR2_X1 U18578 ( .A(n15451), .B(n15450), .ZN(n16316) );
  NOR2_X1 U18579 ( .A1(n15452), .A2(n15487), .ZN(n15474) );
  AOI211_X1 U18580 ( .C1(n15454), .C2(n15462), .A(n15453), .B(n15470), .ZN(
        n15456) );
  INV_X1 U18581 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19910) );
  NOR2_X1 U18582 ( .A1(n19910), .A2(n19170), .ZN(n15455) );
  AOI211_X1 U18583 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15474), .A(
        n15456), .B(n15455), .ZN(n15459) );
  INV_X1 U18584 ( .A(n19130), .ZN(n15457) );
  AOI22_X1 U18585 ( .A1(n15457), .A2(n19308), .B1(n16390), .B2(n16319), .ZN(
        n15458) );
  OAI211_X1 U18586 ( .C1(n16316), .C2(n19300), .A(n15459), .B(n15458), .ZN(
        n15460) );
  INV_X1 U18587 ( .A(n15460), .ZN(n15461) );
  OAI21_X1 U18588 ( .B1(n16317), .B2(n19311), .A(n15461), .ZN(P2_U3035) );
  AOI21_X1 U18589 ( .B1(n15462), .B2(n10381), .A(n9829), .ZN(n16322) );
  INV_X1 U18590 ( .A(n16322), .ZN(n15480) );
  AOI21_X1 U18591 ( .B1(n15486), .B2(n15483), .A(n15482), .ZN(n15469) );
  INV_X1 U18592 ( .A(n15465), .ZN(n15467) );
  NOR2_X1 U18593 ( .A1(n15467), .A2(n15466), .ZN(n15468) );
  XNOR2_X1 U18594 ( .A(n15469), .B(n15468), .ZN(n16324) );
  NOR2_X1 U18595 ( .A1(n15470), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15478) );
  NOR2_X1 U18596 ( .A1(n19908), .A2(n19170), .ZN(n15473) );
  NOR2_X1 U18597 ( .A1(n19305), .A2(n15471), .ZN(n15472) );
  AOI211_X1 U18598 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n15474), .A(
        n15473), .B(n15472), .ZN(n15475) );
  OAI21_X1 U18599 ( .B1(n16400), .B2(n15476), .A(n15475), .ZN(n15477) );
  AOI211_X1 U18600 ( .C1(n16324), .C2(n16391), .A(n15478), .B(n15477), .ZN(
        n15479) );
  OAI21_X1 U18601 ( .B1(n15480), .B2(n19311), .A(n15479), .ZN(P2_U3036) );
  OAI21_X1 U18602 ( .B1(n15481), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10381), .ZN(n16330) );
  INV_X1 U18603 ( .A(n15482), .ZN(n15484) );
  AND2_X1 U18604 ( .A1(n15484), .A2(n15483), .ZN(n15485) );
  XNOR2_X1 U18605 ( .A(n15486), .B(n15485), .ZN(n16329) );
  INV_X1 U18606 ( .A(n15487), .ZN(n15490) );
  NOR2_X1 U18607 ( .A1(n19906), .A2(n19170), .ZN(n15488) );
  AOI221_X1 U18608 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15490), .C1(
        n15489), .C2(n15490), .A(n15488), .ZN(n15494) );
  INV_X1 U18609 ( .A(n15491), .ZN(n15492) );
  AOI22_X1 U18610 ( .A1(n19308), .A2(n15492), .B1(n16390), .B2(n16332), .ZN(
        n15493) );
  OAI211_X1 U18611 ( .C1(n16329), .C2(n19300), .A(n15494), .B(n15493), .ZN(
        n15495) );
  INV_X1 U18612 ( .A(n15495), .ZN(n15496) );
  OAI21_X1 U18613 ( .B1(n16330), .B2(n19311), .A(n15496), .ZN(P2_U3037) );
  INV_X1 U18614 ( .A(n15544), .ZN(n15499) );
  INV_X1 U18615 ( .A(n15497), .ZN(n15498) );
  NOR2_X1 U18616 ( .A1(n15498), .A2(n11260), .ZN(n15512) );
  OAI22_X1 U18617 ( .A1(n19208), .A2(n15499), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15512), .ZN(n16415) );
  INV_X1 U18618 ( .A(n19958), .ZN(n15502) );
  INV_X1 U18619 ( .A(n16457), .ZN(n15500) );
  AOI22_X1 U18620 ( .A1(n19165), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19196), .B2(n19152), .ZN(n15507) );
  AOI222_X1 U18621 ( .A1(n16415), .A2(n15502), .B1(n15501), .B2(n15500), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15507), .ZN(n15505) );
  AOI21_X1 U18622 ( .B1(n15502), .B2(n16416), .A(n15546), .ZN(n15504) );
  OAI22_X1 U18623 ( .A1(n15505), .A2(n15546), .B1(n15504), .B2(n15503), .ZN(
        P2_U3601) );
  OR2_X1 U18624 ( .A1(n15507), .A2(n15506), .ZN(n15527) );
  OAI21_X1 U18625 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(n19192) );
  OAI21_X1 U18626 ( .B1(n19152), .B2(n19298), .A(n19192), .ZN(n15516) );
  INV_X1 U18627 ( .A(n16416), .ZN(n15536) );
  NOR2_X1 U18628 ( .A1(n15536), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15514) );
  NOR3_X1 U18629 ( .A1(n15512), .A2(n15521), .A3(n15511), .ZN(n15513) );
  AOI211_X1 U18630 ( .C1(n13222), .C2(n15544), .A(n15514), .B(n15513), .ZN(
        n16421) );
  OAI222_X1 U18631 ( .A1(n16457), .A2(n19447), .B1(n15527), .B2(n15516), .C1(
        n19958), .C2(n16421), .ZN(n15515) );
  MUX2_X1 U18632 ( .A(n15515), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15546), .Z(P2_U3600) );
  INV_X1 U18633 ( .A(n15516), .ZN(n15528) );
  OR2_X1 U18634 ( .A1(n16431), .A2(n16433), .ZN(n15532) );
  AOI22_X1 U18635 ( .A1(n15532), .A2(n15518), .B1(n15517), .B2(n16416), .ZN(
        n15524) );
  AOI21_X1 U18636 ( .B1(n15520), .B2(n15519), .A(n15518), .ZN(n15533) );
  NOR2_X1 U18637 ( .A1(n15521), .A2(n15529), .ZN(n15522) );
  INV_X1 U18638 ( .A(n15522), .ZN(n15531) );
  NAND2_X1 U18639 ( .A1(n15533), .A2(n15531), .ZN(n15523) );
  NAND2_X1 U18640 ( .A1(n15532), .A2(n15522), .ZN(n15535) );
  NAND3_X1 U18641 ( .A1(n15524), .A2(n15523), .A3(n15535), .ZN(n15525) );
  AOI21_X1 U18642 ( .B1(n15526), .B2(n15544), .A(n15525), .ZN(n16413) );
  OAI222_X1 U18643 ( .A1(n15528), .A2(n15527), .B1(n19958), .B2(n16413), .C1(
        n16457), .C2(n19969), .ZN(n15530) );
  MUX2_X1 U18644 ( .A(n15530), .B(n15529), .S(n15546), .Z(P2_U3599) );
  AOI22_X1 U18645 ( .A1(n15532), .A2(n15531), .B1(n10721), .B2(n16416), .ZN(
        n15539) );
  INV_X1 U18646 ( .A(n15533), .ZN(n15534) );
  OAI211_X1 U18647 ( .C1(n10721), .C2(n15536), .A(n15535), .B(n15534), .ZN(
        n15537) );
  INV_X1 U18648 ( .A(n15537), .ZN(n15538) );
  MUX2_X1 U18649 ( .A(n15539), .B(n15538), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15542) );
  INV_X1 U18650 ( .A(n15540), .ZN(n15541) );
  NAND2_X1 U18651 ( .A1(n15542), .A2(n15541), .ZN(n15543) );
  AOI21_X1 U18652 ( .B1(n15545), .B2(n15544), .A(n15543), .ZN(n16414) );
  OAI22_X1 U18653 ( .A1(n19360), .A2(n16457), .B1(n16414), .B2(n19958), .ZN(
        n15547) );
  MUX2_X1 U18654 ( .A(n15547), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15546), .Z(P2_U3596) );
  INV_X1 U18655 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16729) );
  INV_X1 U18656 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16750) );
  INV_X1 U18657 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16791) );
  INV_X1 U18658 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17170) );
  INV_X1 U18659 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17211) );
  INV_X1 U18660 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17248) );
  NAND2_X1 U18661 ( .A1(n17371), .A2(n15779), .ZN(n15549) );
  INV_X1 U18662 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17008) );
  NAND3_X1 U18663 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17354) );
  NOR2_X1 U18664 ( .A1(n17008), .A2(n17354), .ZN(n17353) );
  INV_X1 U18665 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17344) );
  INV_X1 U18666 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16972) );
  INV_X1 U18667 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16985) );
  NOR3_X1 U18668 ( .A1(n17344), .A2(n16972), .A3(n16985), .ZN(n17323) );
  INV_X1 U18669 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17299) );
  INV_X1 U18670 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16940) );
  NOR4_X1 U18671 ( .A1(n17277), .A2(n17299), .A3(n16933), .A4(n16940), .ZN(
        n15551) );
  NAND4_X1 U18672 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17323), .A4(n15551), .ZN(n17243) );
  NAND2_X1 U18673 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17183), .ZN(n17168) );
  NAND2_X1 U18674 ( .A1(n17371), .A2(n17125), .ZN(n17139) );
  NAND4_X1 U18675 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(n17105), .ZN(n17092) );
  NAND2_X1 U18676 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17097), .ZN(n17082) );
  NAND2_X1 U18677 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17087), .ZN(n17081) );
  INV_X1 U18678 ( .A(n17081), .ZN(n15630) );
  AOI21_X1 U18679 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17360), .A(n17087), .ZN(
        n15629) );
  AOI22_X1 U18680 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15553) );
  OAI21_X1 U18681 ( .B1(n17317), .B2(n18368), .A(n15553), .ZN(n15563) );
  AOI22_X1 U18682 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15561) );
  INV_X1 U18683 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18404) );
  INV_X1 U18684 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18701) );
  OAI22_X1 U18685 ( .A1(n17287), .A2(n18404), .B1(n17161), .B2(n18701), .ZN(
        n15559) );
  AOI22_X1 U18686 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U18687 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15556) );
  AOI22_X1 U18688 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15555) );
  NAND3_X1 U18689 ( .A1(n15557), .A2(n15556), .A3(n15555), .ZN(n15558) );
  AOI211_X1 U18690 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15559), .B(n15558), .ZN(n15560) );
  OAI211_X1 U18691 ( .C1(n17186), .C2(n17140), .A(n15561), .B(n15560), .ZN(
        n15562) );
  AOI211_X1 U18692 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n15563), .B(n15562), .ZN(n17084) );
  AOI22_X1 U18693 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15564) );
  OAI21_X1 U18694 ( .B1(n9848), .B2(n17282), .A(n15564), .ZN(n15575) );
  INV_X1 U18695 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U18696 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15607), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18697 ( .A1(n15686), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15565) );
  OAI21_X1 U18698 ( .B1(n17186), .B2(n15566), .A(n15565), .ZN(n15570) );
  AOI22_X1 U18699 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18700 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15567) );
  OAI211_X1 U18701 ( .C1(n15691), .C2(n17285), .A(n15568), .B(n15567), .ZN(
        n15569) );
  AOI211_X1 U18702 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n15570), .B(n15569), .ZN(n15571) );
  OAI211_X1 U18703 ( .C1(n15688), .C2(n15573), .A(n15572), .B(n15571), .ZN(
        n15574) );
  AOI211_X1 U18704 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n15575), .B(n15574), .ZN(n17094) );
  INV_X1 U18705 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U18706 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15576) );
  OAI21_X1 U18707 ( .B1(n17283), .B2(n17200), .A(n15576), .ZN(n15585) );
  AOI22_X1 U18708 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15583) );
  INV_X1 U18709 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U18710 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15577) );
  OAI21_X1 U18711 ( .B1(n17306), .B2(n18487), .A(n15577), .ZN(n15581) );
  AOI22_X1 U18712 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15579) );
  AOI22_X1 U18713 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15578) );
  OAI211_X1 U18714 ( .C1(n17161), .C2(n18685), .A(n15579), .B(n15578), .ZN(
        n15580) );
  AOI211_X1 U18715 ( .C1(n15554), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n15581), .B(n15580), .ZN(n15582) );
  OAI211_X1 U18716 ( .C1(n17287), .C2(n18392), .A(n15583), .B(n15582), .ZN(
        n15584) );
  AOI211_X1 U18717 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n15585), .B(n15584), .ZN(n17107) );
  AOI22_X1 U18718 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15586) );
  OAI21_X1 U18719 ( .B1(n9827), .B2(n18507), .A(n15586), .ZN(n15595) );
  INV_X1 U18720 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18716) );
  AOI22_X1 U18721 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15593) );
  INV_X1 U18722 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18388) );
  OAI22_X1 U18723 ( .A1(n17287), .A2(n18388), .B1(n17306), .B2(n17051), .ZN(
        n15591) );
  AOI22_X1 U18724 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15735), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U18725 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U18726 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15587) );
  NAND3_X1 U18727 ( .A1(n15589), .A2(n15588), .A3(n15587), .ZN(n15590) );
  AOI211_X1 U18728 ( .C1(n15676), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n15591), .B(n15590), .ZN(n15592) );
  OAI211_X1 U18729 ( .C1(n9844), .C2(n18716), .A(n15593), .B(n15592), .ZN(
        n15594) );
  AOI211_X1 U18730 ( .C1(n15714), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n15595), .B(n15594), .ZN(n17106) );
  NOR2_X1 U18731 ( .A1(n17107), .A2(n17106), .ZN(n17102) );
  AOI22_X1 U18732 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15606) );
  INV_X1 U18733 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U18734 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15596) );
  OAI21_X1 U18735 ( .B1(n9844), .B2(n17316), .A(n15596), .ZN(n15604) );
  AOI22_X1 U18736 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15601) );
  INV_X1 U18737 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U18738 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U18739 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15597) );
  OAI211_X1 U18740 ( .C1(n15691), .C2(n17305), .A(n15598), .B(n15597), .ZN(
        n15599) );
  AOI21_X1 U18741 ( .B1(n15694), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n15599), .ZN(n15600) );
  OAI211_X1 U18742 ( .C1(n10447), .C2(n15602), .A(n15601), .B(n15600), .ZN(
        n15603) );
  AOI211_X1 U18743 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n15604), .B(n15603), .ZN(n15605) );
  OAI211_X1 U18744 ( .C1(n17317), .C2(n18354), .A(n15606), .B(n15605), .ZN(
        n17101) );
  NAND2_X1 U18745 ( .A1(n17102), .A2(n17101), .ZN(n17100) );
  NOR2_X1 U18746 ( .A1(n17094), .A2(n17100), .ZN(n17093) );
  INV_X1 U18747 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U18748 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18749 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15735), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15608) );
  OAI21_X1 U18750 ( .B1(n17304), .B2(n17273), .A(n15608), .ZN(n15615) );
  INV_X1 U18751 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U18752 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15613) );
  AOI22_X1 U18753 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15610) );
  AOI22_X1 U18754 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15609) );
  OAI211_X1 U18755 ( .C1(n17161), .C2(n18696), .A(n15610), .B(n15609), .ZN(
        n15611) );
  AOI21_X1 U18756 ( .B1(n15686), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15611), .ZN(n15612) );
  OAI211_X1 U18757 ( .C1(n15691), .C2(n17268), .A(n15613), .B(n15612), .ZN(
        n15614) );
  AOI211_X1 U18758 ( .C1(n15714), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15615), .B(n15614), .ZN(n15616) );
  OAI211_X1 U18759 ( .C1(n17317), .C2(n18363), .A(n15617), .B(n15616), .ZN(
        n17089) );
  NAND2_X1 U18760 ( .A1(n17093), .A2(n17089), .ZN(n17088) );
  NOR2_X1 U18761 ( .A1(n17084), .A2(n17088), .ZN(n17083) );
  INV_X1 U18762 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18407) );
  AOI22_X1 U18763 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15627) );
  INV_X1 U18764 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U18765 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15619) );
  AOI22_X1 U18766 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17280), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15618) );
  OAI211_X1 U18767 ( .C1(n15691), .C2(n15631), .A(n15619), .B(n15618), .ZN(
        n15625) );
  AOI22_X1 U18768 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15623) );
  AOI22_X1 U18769 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U18770 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15621) );
  NAND2_X1 U18771 ( .A1(n15686), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n15620) );
  NAND4_X1 U18772 ( .A1(n15623), .A2(n15622), .A3(n15621), .A4(n15620), .ZN(
        n15624) );
  AOI211_X1 U18773 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15625), .B(n15624), .ZN(n15626) );
  OAI211_X1 U18774 ( .C1(n17287), .C2(n18407), .A(n15627), .B(n15626), .ZN(
        n15628) );
  NAND2_X1 U18775 ( .A1(n17083), .A2(n15628), .ZN(n17077) );
  OAI21_X1 U18776 ( .B1(n17083), .B2(n15628), .A(n17077), .ZN(n17388) );
  OAI22_X1 U18777 ( .A1(n15630), .A2(n15629), .B1(n17388), .B2(n17360), .ZN(
        P3_U2675) );
  INV_X1 U18778 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17137) );
  OAI22_X1 U18779 ( .A1(n17306), .A2(n15631), .B1(n17317), .B2(n17137), .ZN(
        n15642) );
  AOI22_X1 U18780 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15640) );
  AOI22_X1 U18781 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15735), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15639) );
  AOI22_X1 U18782 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15632) );
  OAI21_X1 U18783 ( .B1(n17287), .B2(n15633), .A(n15632), .ZN(n15637) );
  AOI22_X1 U18784 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U18785 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15634) );
  OAI211_X1 U18786 ( .C1(n15691), .C2(n18407), .A(n15635), .B(n15634), .ZN(
        n15636) );
  AOI211_X1 U18787 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15637), .B(n15636), .ZN(n15638) );
  NAND3_X1 U18788 ( .A1(n15640), .A2(n15639), .A3(n15638), .ZN(n15641) );
  AOI211_X1 U18789 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15642), .B(n15641), .ZN(n17462) );
  INV_X1 U18790 ( .A(n15643), .ZN(n17349) );
  NAND2_X1 U18791 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17321), .ZN(n17320) );
  NOR3_X1 U18792 ( .A1(n17277), .A2(n17299), .A3(n17320), .ZN(n17276) );
  AND2_X1 U18793 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17276), .ZN(n17263) );
  NOR2_X1 U18794 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17263), .ZN(n15644) );
  NOR2_X1 U18795 ( .A1(n18384), .A2(n15643), .ZN(n17352) );
  INV_X1 U18796 ( .A(n17352), .ZN(n17242) );
  OAI21_X1 U18797 ( .B1(n17243), .B2(n17242), .A(n17360), .ZN(n17247) );
  OAI22_X1 U18798 ( .A1(n17462), .A2(n17360), .B1(n15644), .B2(n17247), .ZN(
        P3_U2690) );
  NOR2_X1 U18799 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18975), .ZN(
        n18389) );
  OAI211_X1 U18800 ( .C1(n18999), .C2(n15645), .A(n17287), .B(n18863), .ZN(
        n18336) );
  AOI221_X1 U18801 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18972), .C1(n18336), .C2(
        n18972), .A(n18511), .ZN(n15646) );
  NOR2_X1 U18802 ( .A1(n18389), .A2(n15646), .ZN(n15648) );
  NAND3_X1 U18803 ( .A1(n18869), .A2(n18975), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18720) );
  INV_X1 U18804 ( .A(n15646), .ZN(n18342) );
  NAND2_X1 U18805 ( .A1(n18869), .A2(n18975), .ZN(n16647) );
  NOR2_X1 U18806 ( .A1(n18985), .A2(n19024), .ZN(n17955) );
  INV_X1 U18807 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18845) );
  OAI22_X1 U18808 ( .A1(n19019), .A2(n17955), .B1(n18975), .B2(n18845), .ZN(
        n15651) );
  NAND3_X1 U18809 ( .A1(n18847), .A2(n18342), .A3(n15651), .ZN(n15647) );
  OAI221_X1 U18810 ( .B1(n18847), .B2(n15648), .C1(n18847), .C2(n18720), .A(
        n15647), .ZN(P3_U2864) );
  NOR2_X1 U18811 ( .A1(n18847), .A2(n18852), .ZN(n18532) );
  OR2_X1 U18812 ( .A1(n19019), .A2(n17955), .ZN(n15649) );
  OAI221_X1 U18813 ( .B1(n18975), .B2(n18532), .C1(n15649), .C2(n18532), .A(
        n15648), .ZN(n15650) );
  INV_X1 U18814 ( .A(n15650), .ZN(n18341) );
  INV_X1 U18815 ( .A(n18720), .ZN(n15652) );
  OAI221_X1 U18816 ( .B1(n15652), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n15652), .C2(n15651), .A(n18342), .ZN(n18339) );
  AOI22_X1 U18817 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18341), .B1(
        n18339), .B2(n18852), .ZN(P3_U2865) );
  NAND2_X1 U18818 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15836) );
  NAND2_X1 U18819 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18006) );
  NAND2_X1 U18820 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18204) );
  NOR2_X1 U18821 ( .A1(n18204), .A2(n17857), .ZN(n18178) );
  NAND2_X1 U18822 ( .A1(n18178), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17839) );
  INV_X1 U18823 ( .A(n17839), .ZN(n18162) );
  NAND2_X1 U18824 ( .A1(n18162), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17820) );
  NOR2_X1 U18825 ( .A1(n18170), .A2(n17820), .ZN(n18151) );
  NAND2_X1 U18826 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18151), .ZN(
        n17791) );
  AOI22_X1 U18827 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15653) );
  OAI21_X1 U18828 ( .B1(n17283), .B2(n18415), .A(n15653), .ZN(n15663) );
  AOI22_X1 U18829 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18830 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15655) );
  OAI21_X1 U18831 ( .B1(n15691), .B2(n18388), .A(n15655), .ZN(n15659) );
  INV_X1 U18832 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18627) );
  AOI22_X1 U18833 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18834 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15656) );
  OAI211_X1 U18835 ( .C1(n17161), .C2(n18627), .A(n15657), .B(n15656), .ZN(
        n15658) );
  AOI211_X1 U18836 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15659), .B(n15658), .ZN(n15660) );
  OAI211_X1 U18837 ( .C1(n17317), .C2(n18716), .A(n15661), .B(n15660), .ZN(
        n15662) );
  AOI211_X4 U18838 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15663), .B(n15662), .ZN(n17494) );
  INV_X1 U18839 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U18840 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15664) );
  OAI21_X1 U18841 ( .B1(n9850), .B2(n15665), .A(n15664), .ZN(n15674) );
  INV_X1 U18842 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U18843 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15672) );
  OAI22_X1 U18844 ( .A1(n17287), .A2(n17137), .B1(n15691), .B2(n18374), .ZN(
        n15670) );
  AOI22_X1 U18845 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15668) );
  AOI22_X1 U18846 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U18847 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15666) );
  NAND3_X1 U18848 ( .A1(n15668), .A2(n15667), .A3(n15666), .ZN(n15669) );
  AOI211_X1 U18849 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15670), .B(n15669), .ZN(n15671) );
  OAI211_X1 U18850 ( .C1(n15688), .C2(n17128), .A(n15672), .B(n15671), .ZN(
        n15673) );
  AOI22_X1 U18851 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15675) );
  OAI21_X1 U18852 ( .B1(n9827), .B2(n17268), .A(n15675), .ZN(n15685) );
  AOI22_X1 U18853 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15683) );
  INV_X1 U18854 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18613) );
  AOI22_X1 U18855 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15676), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15677) );
  OAI21_X1 U18856 ( .B1(n17161), .B2(n18613), .A(n15677), .ZN(n15681) );
  AOI22_X1 U18857 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U18858 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15735), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15678) );
  OAI211_X1 U18859 ( .C1(n15691), .C2(n18363), .A(n15679), .B(n15678), .ZN(
        n15680) );
  OAI211_X1 U18860 ( .C1(n10447), .C2(n17273), .A(n15683), .B(n15682), .ZN(
        n15684) );
  AOI22_X1 U18861 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15687) );
  OAI21_X1 U18862 ( .B1(n9844), .B2(n17185), .A(n15687), .ZN(n15693) );
  AOI22_X1 U18863 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U18864 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15689) );
  OAI211_X1 U18865 ( .C1(n15691), .C2(n18354), .A(n15690), .B(n15689), .ZN(
        n15692) );
  AOI211_X1 U18866 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n15693), .B(n15692), .ZN(n15701) );
  INV_X1 U18867 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U18868 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15695) );
  OAI21_X1 U18869 ( .B1(n17158), .B2(n17307), .A(n15695), .ZN(n15699) );
  AOI22_X1 U18870 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15697) );
  NAND3_X1 U18871 ( .A1(n15697), .A2(n10456), .A3(n15696), .ZN(n15698) );
  AOI22_X1 U18872 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15702) );
  OAI21_X1 U18873 ( .B1(n9846), .B2(n18487), .A(n15702), .ZN(n15711) );
  AOI22_X1 U18874 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15709) );
  INV_X1 U18875 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18605) );
  AOI22_X1 U18876 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15703) );
  OAI21_X1 U18877 ( .B1(n17161), .B2(n18605), .A(n15703), .ZN(n15707) );
  INV_X1 U18878 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18349) );
  AOI22_X1 U18879 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15705) );
  AOI22_X1 U18880 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15704) );
  OAI211_X1 U18881 ( .C1(n15691), .C2(n18349), .A(n15705), .B(n15704), .ZN(
        n15706) );
  AOI211_X1 U18882 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n15707), .B(n15706), .ZN(n15708) );
  OAI211_X1 U18883 ( .C1(n15688), .C2(n17200), .A(n15709), .B(n15708), .ZN(
        n15710) );
  INV_X1 U18884 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18358) );
  AOI22_X1 U18885 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15722) );
  AOI22_X1 U18886 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U18887 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17308), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15712) );
  OAI211_X1 U18888 ( .C1(n17306), .C2(n17282), .A(n15713), .B(n15712), .ZN(
        n15720) );
  AOI22_X1 U18889 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18890 ( .A1(n15716), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15715), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U18891 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n15717) );
  OAI211_X1 U18892 ( .C1(n15691), .C2(n18358), .A(n15722), .B(n15721), .ZN(
        n17514) );
  NOR2_X1 U18893 ( .A1(n15789), .A2(n9859), .ZN(n15746) );
  INV_X1 U18894 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U18895 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U18896 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U18897 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15723) );
  OAI211_X1 U18898 ( .C1(n15691), .C2(n18368), .A(n15724), .B(n15723), .ZN(
        n15730) );
  AOI22_X1 U18899 ( .A1(n17280), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U18900 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15727) );
  AOI22_X1 U18901 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15726) );
  NAND2_X1 U18902 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n15725) );
  NAND4_X1 U18903 ( .A1(n15728), .A2(n15727), .A3(n15726), .A4(n15725), .ZN(
        n15729) );
  AOI211_X1 U18904 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15730), .B(n15729), .ZN(n15731) );
  OAI211_X1 U18905 ( .C1(n10447), .C2(n17250), .A(n15732), .B(n15731), .ZN(
        n15787) );
  NAND2_X1 U18906 ( .A1(n15746), .A2(n15787), .ZN(n15745) );
  AOI22_X1 U18907 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n9811), .ZN(n15743) );
  INV_X1 U18908 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U18909 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n17330), .B1(
        n17280), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U18910 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15714), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15733) );
  OAI211_X1 U18911 ( .C1(n17306), .C2(n17230), .A(n15734), .B(n15733), .ZN(
        n15741) );
  AOI22_X1 U18912 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n15676), .ZN(n15739) );
  AOI22_X1 U18913 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n17308), .B1(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n17326), .ZN(n15738) );
  AOI22_X1 U18914 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n15735), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n17325), .ZN(n15737) );
  NAND2_X1 U18915 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n17231), .ZN(
        n15736) );
  NAND4_X1 U18916 ( .A1(n15739), .A2(n15738), .A3(n15737), .A4(n15736), .ZN(
        n15740) );
  AOI211_X1 U18917 ( .C1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .C2(n15694), .A(
        n15741), .B(n15740), .ZN(n15742) );
  OAI211_X1 U18918 ( .C1(n15691), .C2(n18379), .A(n15743), .B(n15742), .ZN(
        n15808) );
  NAND2_X1 U18919 ( .A1(n17925), .A2(n15808), .ZN(n15744) );
  NOR2_X1 U18920 ( .A1(n17494), .A2(n15744), .ZN(n15762) );
  XOR2_X1 U18921 ( .A(n17494), .B(n15744), .Z(n15758) );
  XOR2_X1 U18922 ( .A(n17501), .B(n15745), .Z(n15754) );
  AND2_X1 U18923 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15754), .ZN(
        n15755) );
  INV_X1 U18924 ( .A(n15787), .ZN(n17505) );
  XNOR2_X1 U18925 ( .A(n17505), .B(n15746), .ZN(n15752) );
  AND2_X1 U18926 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15752), .ZN(
        n15753) );
  XOR2_X1 U18927 ( .A(n9859), .B(n15789), .Z(n15750) );
  AND2_X1 U18928 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15750), .ZN(
        n15751) );
  AOI21_X1 U18929 ( .B1(n15790), .B2(n15920), .A(n9859), .ZN(n15748) );
  INV_X1 U18930 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18304) );
  NOR2_X1 U18931 ( .A1(n15748), .A2(n18304), .ZN(n15749) );
  NOR2_X1 U18932 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15920), .ZN(
        n17992) );
  INV_X1 U18933 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18987) );
  XNOR2_X1 U18934 ( .A(n18987), .B(n15793), .ZN(n17983) );
  INV_X1 U18935 ( .A(n17983), .ZN(n17985) );
  NAND2_X1 U18936 ( .A1(n17992), .A2(n17985), .ZN(n17984) );
  OAI211_X1 U18937 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n10112), .A(
        n15747), .B(n17984), .ZN(n17975) );
  INV_X1 U18938 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18291) );
  XOR2_X1 U18939 ( .A(n18291), .B(n15750), .Z(n17962) );
  NOR2_X1 U18940 ( .A1(n15751), .A2(n17961), .ZN(n17947) );
  INV_X1 U18941 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18274) );
  XOR2_X1 U18942 ( .A(n18274), .B(n15752), .Z(n17946) );
  INV_X1 U18943 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18270) );
  XOR2_X1 U18944 ( .A(n18270), .B(n15754), .Z(n17937) );
  INV_X1 U18945 ( .A(n15808), .ZN(n17498) );
  INV_X1 U18946 ( .A(n17925), .ZN(n17923) );
  XNOR2_X1 U18947 ( .A(n17498), .B(n17923), .ZN(n15756) );
  AOI222_X1 U18948 ( .A1(n17924), .A2(n15813), .B1(n17924), .B2(n15756), .C1(
        n15813), .C2(n15756), .ZN(n15759) );
  INV_X1 U18949 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18250) );
  NAND2_X1 U18950 ( .A1(n15762), .A2(n15757), .ZN(n15763) );
  AND2_X1 U18951 ( .A1(n15759), .A2(n15758), .ZN(n17915) );
  AOI21_X1 U18952 ( .B1(n15762), .B2(n15761), .A(n17915), .ZN(n15760) );
  NAND2_X1 U18953 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17900), .ZN(
        n17899) );
  NOR2_X1 U18954 ( .A1(n18142), .A2(n18129), .ZN(n18120) );
  NAND2_X1 U18955 ( .A1(n18120), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18083) );
  NAND2_X1 U18956 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18087) );
  NOR2_X1 U18957 ( .A1(n18088), .A2(n18087), .ZN(n15831) );
  INV_X1 U18958 ( .A(n15831), .ZN(n18072) );
  NOR2_X1 U18959 ( .A1(n18083), .A2(n18072), .ZN(n18071) );
  NAND2_X1 U18960 ( .A1(n18071), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18073) );
  INV_X1 U18961 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18002) );
  NOR2_X1 U18962 ( .A1(n18073), .A2(n18002), .ZN(n17686) );
  NAND2_X1 U18963 ( .A1(n17686), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18029) );
  INV_X1 U18964 ( .A(n17641), .ZN(n18011) );
  NOR2_X1 U18965 ( .A1(n15836), .A2(n18011), .ZN(n16535) );
  NAND3_X1 U18966 ( .A1(n15764), .A2(n17524), .A3(n18350), .ZN(n15766) );
  NAND2_X1 U18967 ( .A1(n15766), .A2(n15765), .ZN(n18820) );
  AOI21_X1 U18968 ( .B1(n15770), .B2(n15769), .A(n15776), .ZN(n16471) );
  NAND2_X1 U18969 ( .A1(n15773), .A2(n18350), .ZN(n15771) );
  NOR2_X1 U18970 ( .A1(n9849), .A2(n15771), .ZN(n15785) );
  INV_X1 U18971 ( .A(n15772), .ZN(n15777) );
  XNOR2_X1 U18972 ( .A(n15773), .B(n18350), .ZN(n15774) );
  OAI21_X1 U18973 ( .B1(n15775), .B2(n15774), .A(n19026), .ZN(n16649) );
  NOR3_X1 U18974 ( .A1(n15777), .A2(n15776), .A3(n16649), .ZN(n15781) );
  INV_X1 U18975 ( .A(n18812), .ZN(n16472) );
  AOI211_X1 U18976 ( .C1(n15779), .C2(n15778), .A(n18355), .B(n16472), .ZN(
        n15780) );
  AOI211_X1 U18977 ( .C1(n16471), .C2(n15785), .A(n15781), .B(n15780), .ZN(
        n15782) );
  NAND2_X1 U18978 ( .A1(n18197), .A2(n18315), .ZN(n18334) );
  INV_X1 U18979 ( .A(n17494), .ZN(n15786) );
  NAND2_X1 U18980 ( .A1(n15785), .A2(n15784), .ZN(n16473) );
  INV_X1 U18981 ( .A(n16473), .ZN(n18809) );
  NOR2_X1 U18982 ( .A1(n15786), .A2(n18332), .ZN(n18242) );
  INV_X1 U18983 ( .A(n18242), .ZN(n18042) );
  XOR2_X1 U18984 ( .A(n15805), .B(n17501), .Z(n15801) );
  XNOR2_X1 U18985 ( .A(n15788), .B(n17505), .ZN(n15799) );
  XOR2_X1 U18986 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15799), .Z(
        n17952) );
  XNOR2_X1 U18987 ( .A(n15790), .B(n15789), .ZN(n15797) );
  NAND2_X1 U18988 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15797), .ZN(
        n15798) );
  OR2_X1 U18989 ( .A1(n18304), .A2(n15792), .ZN(n15796) );
  NAND2_X1 U18990 ( .A1(n15793), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15795) );
  INV_X1 U18991 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19003) );
  NOR2_X1 U18992 ( .A1(n15794), .A2(n19003), .ZN(n17993) );
  NAND2_X1 U18993 ( .A1(n15795), .A2(n17982), .ZN(n18293) );
  NAND2_X1 U18994 ( .A1(n15796), .A2(n18292), .ZN(n17965) );
  NAND2_X1 U18995 ( .A1(n15798), .A2(n17964), .ZN(n17951) );
  NAND2_X1 U18996 ( .A1(n17952), .A2(n17951), .ZN(n17950) );
  NAND2_X1 U18997 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15799), .ZN(
        n15800) );
  NAND2_X1 U18998 ( .A1(n17950), .A2(n15800), .ZN(n15803) );
  NAND2_X1 U18999 ( .A1(n15801), .A2(n15803), .ZN(n15804) );
  INV_X1 U19000 ( .A(n15801), .ZN(n15802) );
  XNOR2_X1 U19001 ( .A(n15803), .B(n15802), .ZN(n17935) );
  NAND2_X1 U19002 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17935), .ZN(
        n17934) );
  NAND2_X1 U19003 ( .A1(n15804), .A2(n17934), .ZN(n17921) );
  XNOR2_X1 U19004 ( .A(n15813), .B(n15808), .ZN(n17926) );
  XOR2_X1 U19005 ( .A(n15809), .B(n17926), .Z(n17922) );
  AOI21_X1 U19006 ( .B1(n17494), .B2(n16533), .A(n17793), .ZN(n15811) );
  NAND2_X1 U19007 ( .A1(n15811), .A2(n17790), .ZN(n15812) );
  NAND2_X1 U19008 ( .A1(n17862), .A2(n18115), .ZN(n18067) );
  INV_X1 U19009 ( .A(n17686), .ZN(n17685) );
  NAND2_X1 U19010 ( .A1(n18044), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17674) );
  NAND3_X1 U19011 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18009), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16528) );
  INV_X1 U19012 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18016) );
  NOR2_X1 U19013 ( .A1(n18006), .A2(n18029), .ZN(n15834) );
  INV_X1 U19014 ( .A(n15834), .ZN(n18001) );
  NOR2_X1 U19015 ( .A1(n18016), .A2(n18001), .ZN(n16539) );
  NAND3_X1 U19016 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18259) );
  NOR2_X1 U19017 ( .A1(n15813), .A2(n18259), .ZN(n18254) );
  NAND3_X1 U19018 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18254), .ZN(n15830) );
  INV_X1 U19019 ( .A(n15830), .ZN(n18112) );
  AOI21_X1 U19020 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18111) );
  INV_X1 U19021 ( .A(n18111), .ZN(n18300) );
  NAND2_X1 U19022 ( .A1(n18112), .A2(n18300), .ZN(n18138) );
  NOR2_X1 U19023 ( .A1(n17791), .A2(n18138), .ZN(n18116) );
  INV_X1 U19024 ( .A(n18116), .ZN(n18028) );
  NAND2_X1 U19025 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18232) );
  NAND2_X1 U19026 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18254), .ZN(
        n18234) );
  OR3_X1 U19027 ( .A1(n18237), .A2(n18232), .A3(n18234), .ZN(n18139) );
  NOR2_X1 U19028 ( .A1(n17791), .A2(n18139), .ZN(n18066) );
  INV_X1 U19029 ( .A(n18066), .ZN(n18117) );
  NAND2_X1 U19030 ( .A1(n10247), .A2(n19003), .ZN(n18314) );
  NAND2_X1 U19031 ( .A1(n18314), .A2(n18231), .ZN(n18298) );
  OAI22_X1 U19032 ( .A1(n18835), .A2(n18028), .B1(n18117), .B2(n18298), .ZN(
        n18025) );
  NAND4_X1 U19033 ( .A1(n18315), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16539), .A4(n18025), .ZN(n16516) );
  OAI21_X1 U19034 ( .B1(n18042), .B2(n16528), .A(n16516), .ZN(n15814) );
  AOI21_X1 U19035 ( .B1(n16535), .B2(n18322), .A(n15814), .ZN(n15901) );
  NOR2_X1 U19036 ( .A1(n17494), .A2(n16473), .ZN(n16531) );
  INV_X1 U19037 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16518) );
  NOR2_X1 U19038 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17793), .ZN(
        n16529) );
  INV_X1 U19039 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18034) );
  NOR2_X1 U19040 ( .A1(n17793), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17768) );
  INV_X1 U19041 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18109) );
  NAND2_X1 U19042 ( .A1(n17768), .A2(n18109), .ZN(n15815) );
  NOR2_X1 U19043 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15815), .ZN(
        n17730) );
  NAND2_X1 U19044 ( .A1(n17730), .A2(n18088), .ZN(n17717) );
  NAND2_X1 U19045 ( .A1(n15816), .A2(n18237), .ZN(n17883) );
  INV_X1 U19046 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18195) );
  NAND2_X1 U19047 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15818), .ZN(
        n15819) );
  NAND2_X1 U19048 ( .A1(n18243), .A2(n17902), .ZN(n17901) );
  NAND2_X1 U19049 ( .A1(n15819), .A2(n17901), .ZN(n17874) );
  NAND2_X1 U19050 ( .A1(n18115), .A2(n17874), .ZN(n15820) );
  NAND2_X1 U19051 ( .A1(n10446), .A2(n18129), .ZN(n17779) );
  OR2_X1 U19052 ( .A1(n17793), .A2(n17688), .ZN(n17675) );
  OAI221_X1 U19053 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17902), 
        .C1(n18034), .C2(n17676), .A(n17675), .ZN(n17657) );
  NOR2_X1 U19054 ( .A1(n17676), .A2(n17902), .ZN(n15825) );
  NOR2_X1 U19055 ( .A1(n17902), .A2(n15823), .ZN(n15824) );
  NOR2_X1 U19056 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15827), .ZN(
        n16530) );
  NAND2_X1 U19057 ( .A1(n16529), .A2(n16530), .ZN(n15900) );
  INV_X1 U19058 ( .A(n15900), .ZN(n15828) );
  INV_X1 U19059 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16538) );
  NOR2_X1 U19060 ( .A1(n15828), .A2(n15899), .ZN(n15829) );
  XOR2_X1 U19061 ( .A(n16518), .B(n15829), .Z(n16506) );
  NOR2_X1 U19062 ( .A1(n10244), .A2(n18826), .ZN(n18214) );
  OR2_X1 U19063 ( .A1(n19003), .A2(n18232), .ZN(n18299) );
  NOR2_X1 U19064 ( .A1(n15830), .A2(n18299), .ZN(n18222) );
  NAND2_X1 U19065 ( .A1(n18115), .A2(n18222), .ZN(n18137) );
  INV_X1 U19066 ( .A(n16539), .ZN(n17633) );
  NAND2_X1 U19067 ( .A1(n15831), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15832) );
  INV_X1 U19068 ( .A(n18083), .ZN(n18065) );
  NAND2_X1 U19069 ( .A1(n18065), .A2(n18116), .ZN(n18070) );
  NOR2_X1 U19070 ( .A1(n15832), .A2(n18070), .ZN(n18047) );
  NAND3_X1 U19071 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n18047), .ZN(n15833) );
  OAI21_X1 U19072 ( .B1(n18006), .B2(n15833), .A(n10244), .ZN(n18008) );
  OAI221_X1 U19073 ( .B1(n10247), .B2(n15834), .C1(n10247), .C2(n18066), .A(
        n18008), .ZN(n15835) );
  AOI221_X1 U19074 ( .B1(n18137), .B2(n18841), .C1(n17633), .C2(n18841), .A(
        n15835), .ZN(n15897) );
  OAI21_X1 U19075 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18214), .A(
        n15897), .ZN(n16527) );
  AOI21_X1 U19076 ( .B1(n16538), .B2(n18249), .A(n16527), .ZN(n15837) );
  NOR2_X1 U19077 ( .A1(n15836), .A2(n16518), .ZN(n16493) );
  NAND2_X1 U19078 ( .A1(n17641), .A2(n16493), .ZN(n16492) );
  NAND2_X1 U19079 ( .A1(n18009), .A2(n16493), .ZN(n16491) );
  AOI22_X1 U19080 ( .A1(n18322), .A2(n16492), .B1(n18242), .B2(n16491), .ZN(
        n15904) );
  OAI211_X1 U19081 ( .C1(n15837), .C2(n18305), .A(n15904), .B(n18317), .ZN(
        n15838) );
  AOI22_X1 U19082 ( .A1(n18241), .A2(n16506), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15838), .ZN(n15839) );
  NAND2_X1 U19083 ( .A1(n18330), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16513) );
  OAI211_X1 U19084 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15901), .A(
        n15839), .B(n16513), .ZN(P3_U2833) );
  AOI22_X1 U19085 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19197), .ZN(n15848) );
  AOI22_X1 U19086 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19183), .B1(n15840), 
        .B2(n19205), .ZN(n15847) );
  AOI22_X1 U19087 ( .A1(n15842), .A2(n19199), .B1(n15841), .B2(n19185), .ZN(
        n15846) );
  NAND4_X1 U19088 ( .A1(n15848), .A2(n15847), .A3(n15846), .A4(n15845), .ZN(
        P2_U2833) );
  INV_X1 U19089 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21041) );
  NAND2_X1 U19090 ( .A1(n21041), .A2(n20014), .ZN(n15867) );
  INV_X1 U19091 ( .A(n15857), .ZN(n15859) );
  NOR3_X1 U19092 ( .A1(n15850), .A2(n15849), .A3(n20866), .ZN(n15853) );
  NAND2_X1 U19093 ( .A1(n15853), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15855) );
  OAI22_X1 U19094 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15853), .B1(
        n15852), .B2(n15851), .ZN(n15854) );
  OAI211_X1 U19095 ( .C1(n15857), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        n15858) );
  OAI21_X1 U19096 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15859), .A(
        n15858), .ZN(n15860) );
  AOI222_X1 U19097 ( .A1(n20856), .A2(n15861), .B1(n20856), .B2(n15860), .C1(
        n15861), .C2(n15860), .ZN(n15865) );
  INV_X1 U19098 ( .A(n15862), .ZN(n15863) );
  OAI211_X1 U19099 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15865), .A(
        n15864), .B(n15863), .ZN(n15866) );
  AOI21_X1 U19100 ( .B1(n15868), .B2(n15867), .A(n15866), .ZN(n15869) );
  NAND2_X1 U19101 ( .A1(n15870), .A2(n15869), .ZN(n15871) );
  AOI21_X1 U19102 ( .B1(n15873), .B2(n15872), .A(n15871), .ZN(n15886) );
  INV_X1 U19103 ( .A(n15874), .ZN(n16192) );
  NOR2_X1 U19104 ( .A1(n15875), .A2(n16192), .ZN(n20862) );
  NOR2_X1 U19105 ( .A1(n15883), .A2(n16196), .ZN(n15880) );
  NOR2_X1 U19106 ( .A1(n15876), .A2(n20879), .ZN(n15879) );
  NAND3_X1 U19107 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20876), .A3(n16196), 
        .ZN(n15877) );
  AOI22_X1 U19108 ( .A1(n15879), .A2(n15878), .B1(n20766), .B2(n15877), .ZN(
        n16191) );
  OAI221_X1 U19109 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15886), 
        .A(n16191), .ZN(n15881) );
  OAI211_X1 U19110 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20880), .A(n15880), 
        .B(n15881), .ZN(n16194) );
  INV_X1 U19111 ( .A(n15881), .ZN(n16197) );
  AOI21_X1 U19112 ( .B1(n15883), .B2(n15882), .A(n16197), .ZN(n15884) );
  OAI22_X1 U19113 ( .A1(n20862), .A2(n16194), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15884), .ZN(n15885) );
  OAI21_X1 U19114 ( .B1(n15886), .B2(n20008), .A(n15885), .ZN(P1_U3161) );
  OAI22_X1 U19115 ( .A1(n15889), .A2(n15888), .B1(n20140), .B2(n15887), .ZN(
        n15890) );
  INV_X1 U19116 ( .A(n15890), .ZN(n15895) );
  INV_X1 U19117 ( .A(n15891), .ZN(n15893) );
  AOI22_X1 U19118 ( .A1(n15893), .A2(n16182), .B1(n20169), .B2(n15892), .ZN(
        n15894) );
  OAI211_X1 U19119 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15896), .A(
        n15895), .B(n15894), .ZN(P1_U3010) );
  INV_X1 U19120 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16517) );
  INV_X1 U19121 ( .A(n18317), .ZN(n18056) );
  OAI21_X1 U19122 ( .B1(n18826), .B2(n18316), .A(n18315), .ZN(n18312) );
  OAI22_X1 U19123 ( .A1(n15897), .A2(n18305), .B1(n16493), .B2(n18312), .ZN(
        n15898) );
  NOR2_X1 U19124 ( .A1(n18056), .A2(n15898), .ZN(n16515) );
  INV_X1 U19125 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18959) );
  NOR2_X1 U19126 ( .A1(n18216), .A2(n18959), .ZN(n16494) );
  NOR3_X1 U19127 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15901), .A3(
        n16518), .ZN(n15902) );
  OAI221_X1 U19128 ( .B1(n16517), .B2(n16515), .C1(n16517), .C2(n15904), .A(
        n15903), .ZN(P3_U2832) );
  INV_X1 U19129 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20773) );
  INV_X1 U19130 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20971) );
  NOR2_X1 U19131 ( .A1(n20776), .A2(n20971), .ZN(n15905) );
  INV_X1 U19132 ( .A(HOLD), .ZN(n21001) );
  INV_X1 U19133 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U19134 ( .A1(n15905), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n15905), 
        .B2(HOLD), .C1(n21001), .C2(n20782), .ZN(n15906) );
  OAI211_X1 U19135 ( .C1(n20880), .C2(n20773), .A(n15906), .B(n20879), .ZN(
        P1_U3195) );
  AND2_X1 U19136 ( .A1(n15907), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U19137 ( .A1(n19872), .A2(n19862), .ZN(n16464) );
  NAND2_X1 U19138 ( .A1(n16469), .A2(n16464), .ZN(n15908) );
  AOI211_X1 U19139 ( .C1(n15909), .C2(n19633), .A(n15910), .B(n15908), .ZN(
        P2_U3178) );
  INV_X1 U19140 ( .A(n16469), .ZN(n16449) );
  INV_X1 U19141 ( .A(n15910), .ZN(n16456) );
  INV_X1 U19142 ( .A(n19991), .ZN(n15911) );
  NAND2_X1 U19143 ( .A1(n16456), .A2(n15911), .ZN(n15912) );
  AOI221_X1 U19144 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16449), .C1(n19998), .C2(
        n16449), .A(n19807), .ZN(n19995) );
  INV_X1 U19145 ( .A(n19995), .ZN(n19992) );
  NOR2_X1 U19146 ( .A1(n16426), .A2(n19992), .ZN(P2_U3047) );
  NAND3_X1 U19147 ( .A1(n15915), .A2(n19025), .A3(n15914), .ZN(n15916) );
  INV_X1 U19148 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17592) );
  NOR2_X1 U19149 ( .A1(n17372), .A2(n17592), .ZN(n17521) );
  NAND2_X1 U19150 ( .A1(n17371), .A2(n17513), .ZN(n17491) );
  NAND2_X1 U19151 ( .A1(n15918), .A2(n17513), .ZN(n17509) );
  AOI22_X1 U19152 ( .A1(n17518), .A2(BUF2_REG_0__SCAN_IN), .B1(n17517), .B2(
        n15920), .ZN(n15921) );
  OAI221_X1 U19153 ( .B1(n17521), .B2(n17592), .C1(n17521), .C2(n17491), .A(
        n15921), .ZN(P3_U2735) );
  OAI21_X1 U19154 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15922), .ZN(n15933) );
  INV_X1 U19155 ( .A(n20055), .ZN(n15975) );
  AOI21_X1 U19156 ( .B1(n20073), .B2(n15923), .A(n15975), .ZN(n15924) );
  OAI21_X1 U19157 ( .B1(n15925), .B2(n20057), .A(n15924), .ZN(n15928) );
  NOR2_X1 U19158 ( .A1(n15926), .A2(n15963), .ZN(n15927) );
  AOI211_X1 U19159 ( .C1(n20043), .C2(P1_EBX_REG_16__SCAN_IN), .A(n15928), .B(
        n15927), .ZN(n15932) );
  OAI21_X1 U19160 ( .B1(n15930), .B2(n15929), .A(n15983), .ZN(n15945) );
  AOI22_X1 U19161 ( .A1(n15990), .A2(n20047), .B1(P1_REIP_REG_16__SCAN_IN), 
        .B2(n15945), .ZN(n15931) );
  OAI211_X1 U19162 ( .C1(n15944), .C2(n15933), .A(n15932), .B(n15931), .ZN(
        P1_U2824) );
  OR2_X1 U19163 ( .A1(n15935), .A2(n15934), .ZN(n15936) );
  NAND2_X1 U19164 ( .A1(n15937), .A2(n15936), .ZN(n16092) );
  INV_X1 U19165 ( .A(n16092), .ZN(n15986) );
  OAI21_X1 U19166 ( .B1(n20057), .B2(n15938), .A(n20055), .ZN(n15939) );
  AOI21_X1 U19167 ( .B1(n20043), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15939), .ZN(
        n15940) );
  OAI21_X1 U19168 ( .B1(n15999), .B2(n20059), .A(n15940), .ZN(n15941) );
  AOI21_X1 U19169 ( .B1(n15986), .B2(n20070), .A(n15941), .ZN(n15943) );
  AOI22_X1 U19170 ( .A1(n16001), .A2(n20047), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15945), .ZN(n15942) );
  OAI211_X1 U19171 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15944), .A(n15943), 
        .B(n15942), .ZN(P1_U2825) );
  AOI22_X1 U19172 ( .A1(n16101), .A2(n20070), .B1(n20073), .B2(n16012), .ZN(
        n15949) );
  AOI22_X1 U19173 ( .A1(n20043), .A2(P1_EBX_REG_14__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20069), .ZN(n15948) );
  NAND3_X1 U19174 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15961), .ZN(n15954) );
  OAI21_X1 U19175 ( .B1(n15960), .B2(n15954), .A(n21232), .ZN(n15946) );
  AOI22_X1 U19176 ( .A1(n16013), .A2(n20047), .B1(n15946), .B2(n15945), .ZN(
        n15947) );
  NAND4_X1 U19177 ( .A1(n15949), .A2(n15948), .A3(n15947), .A4(n20055), .ZN(
        P1_U2826) );
  NAND2_X1 U19178 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15951) );
  AOI21_X1 U19179 ( .B1(n15951), .B2(n20029), .A(n15950), .ZN(n15970) );
  AOI22_X1 U19180 ( .A1(n16110), .A2(n20070), .B1(n20043), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15952) );
  OAI211_X1 U19181 ( .C1(n20057), .C2(n15953), .A(n15952), .B(n20055), .ZN(
        n15957) );
  OAI22_X1 U19182 ( .A1(n15955), .A2(n15978), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15954), .ZN(n15956) );
  AOI211_X1 U19183 ( .C1(n15958), .C2(n20073), .A(n15957), .B(n15956), .ZN(
        n15959) );
  OAI21_X1 U19184 ( .B1(n15970), .B2(n15960), .A(n15959), .ZN(P1_U2827) );
  AOI21_X1 U19185 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15961), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19186 ( .A1(n20043), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n20073), 
        .B2(n16021), .ZN(n15968) );
  INV_X1 U19187 ( .A(n15962), .ZN(n16022) );
  NOR2_X1 U19188 ( .A1(n16123), .A2(n15963), .ZN(n15966) );
  OAI21_X1 U19189 ( .B1(n20057), .B2(n15964), .A(n20055), .ZN(n15965) );
  AOI211_X1 U19190 ( .C1(n16022), .C2(n20047), .A(n15966), .B(n15965), .ZN(
        n15967) );
  OAI211_X1 U19191 ( .C1(n15970), .C2(n15969), .A(n15968), .B(n15967), .ZN(
        P1_U2828) );
  AND2_X1 U19192 ( .A1(n15972), .A2(n15971), .ZN(n15973) );
  NOR2_X1 U19193 ( .A1(n15974), .A2(n15973), .ZN(n16132) );
  NAND2_X1 U19194 ( .A1(n20043), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n15977) );
  AOI21_X1 U19195 ( .B1(n20069), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15975), .ZN(n15976) );
  OAI211_X1 U19196 ( .C1(n20059), .C2(n16033), .A(n15977), .B(n15976), .ZN(
        n15981) );
  NOR2_X1 U19197 ( .A1(n15979), .A2(n15978), .ZN(n15980) );
  AOI211_X1 U19198 ( .C1(n16132), .C2(n20070), .A(n15981), .B(n15980), .ZN(
        n15982) );
  OAI221_X1 U19199 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15985), .C1(n15984), 
        .C2(n15983), .A(n15982), .ZN(P1_U2829) );
  AOI22_X1 U19200 ( .A1(n16001), .A2(n20089), .B1(n20088), .B2(n15986), .ZN(
        n15987) );
  OAI21_X1 U19201 ( .B1(n20092), .B2(n12374), .A(n15987), .ZN(P1_U2857) );
  AOI22_X1 U19202 ( .A1(n16030), .A2(n20089), .B1(n20088), .B2(n16132), .ZN(
        n15988) );
  OAI21_X1 U19203 ( .B1(n20092), .B2(n21230), .A(n15988), .ZN(P1_U2861) );
  AOI22_X1 U19204 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15992) );
  AOI22_X1 U19205 ( .A1(n15990), .A2(n20178), .B1(n16045), .B2(n15989), .ZN(
        n15991) );
  OAI211_X1 U19206 ( .C1(n20141), .C2(n15993), .A(n15992), .B(n15991), .ZN(
        P1_U2983) );
  INV_X1 U19207 ( .A(n15994), .ZN(n15995) );
  OAI21_X1 U19208 ( .B1(n16098), .B2(n10154), .A(n15995), .ZN(n15997) );
  AOI21_X1 U19209 ( .B1(n15998), .B2(n15997), .A(n15996), .ZN(n16093) );
  AOI22_X1 U19210 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16003) );
  INV_X1 U19211 ( .A(n15999), .ZN(n16000) );
  AOI22_X1 U19212 ( .A1(n16001), .A2(n20178), .B1(n16043), .B2(n16000), .ZN(
        n16002) );
  OAI211_X1 U19213 ( .C1(n16093), .C2(n20155), .A(n16003), .B(n16002), .ZN(
        P1_U2984) );
  INV_X1 U19214 ( .A(n16004), .ZN(n16007) );
  OAI21_X1 U19215 ( .B1(n16007), .B2(n16006), .A(n16005), .ZN(n16011) );
  AOI22_X1 U19216 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16104), .B2(n16008), .ZN(n16010) );
  XNOR2_X1 U19217 ( .A(n16011), .B(n16010), .ZN(n16107) );
  AOI22_X1 U19218 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16015) );
  AOI22_X1 U19219 ( .A1(n16013), .A2(n20178), .B1(n16043), .B2(n16012), .ZN(
        n16014) );
  OAI211_X1 U19220 ( .C1(n16107), .C2(n20155), .A(n16015), .B(n16014), .ZN(
        P1_U2985) );
  OAI21_X1 U19221 ( .B1(n16026), .B2(n16018), .A(n16017), .ZN(n16019) );
  XOR2_X1 U19222 ( .A(n16020), .B(n16019), .Z(n16131) );
  AOI22_X1 U19223 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16024) );
  AOI22_X1 U19224 ( .A1(n16022), .A2(n20178), .B1(n16043), .B2(n16021), .ZN(
        n16023) );
  OAI211_X1 U19225 ( .C1(n16131), .C2(n20155), .A(n16024), .B(n16023), .ZN(
        P1_U2987) );
  AOI22_X1 U19226 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16032) );
  NOR2_X1 U19227 ( .A1(n16025), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16028) );
  NOR2_X1 U19228 ( .A1(n16026), .A2(n12685), .ZN(n16027) );
  MUX2_X1 U19229 ( .A(n16028), .B(n16027), .S(n10154), .Z(n16029) );
  XNOR2_X1 U19230 ( .A(n16029), .B(n12742), .ZN(n16133) );
  AOI22_X1 U19231 ( .A1(n16133), .A2(n16045), .B1(n16030), .B2(n20178), .ZN(
        n16031) );
  OAI211_X1 U19232 ( .C1(n20141), .C2(n16033), .A(n16032), .B(n16031), .ZN(
        P1_U2988) );
  AOI22_X1 U19233 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20149), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U19234 ( .A1(n16035), .A2(n16034), .ZN(n16036) );
  XNOR2_X1 U19235 ( .A(n16037), .B(n16036), .ZN(n16165) );
  INV_X1 U19236 ( .A(n16038), .ZN(n20082) );
  AOI22_X1 U19237 ( .A1(n16165), .A2(n16045), .B1(n20178), .B2(n20082), .ZN(
        n16039) );
  OAI211_X1 U19238 ( .C1(n20141), .C2(n20033), .A(n16040), .B(n16039), .ZN(
        P1_U2992) );
  XOR2_X1 U19239 ( .A(n16042), .B(n16041), .Z(n16183) );
  INV_X1 U19240 ( .A(n20058), .ZN(n16044) );
  AOI222_X1 U19241 ( .A1(n16183), .A2(n16045), .B1(n20178), .B2(n20085), .C1(
        n16044), .C2(n16043), .ZN(n16046) );
  NAND2_X1 U19242 ( .A1(n20149), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16174) );
  OAI211_X1 U19243 ( .C1(n20056), .C2(n16047), .A(n16046), .B(n16174), .ZN(
        P1_U2994) );
  AOI211_X1 U19244 ( .C1(n16049), .C2(n12408), .A(n16048), .B(n16064), .ZN(
        n16054) );
  INV_X1 U19245 ( .A(n16050), .ZN(n16051) );
  OAI21_X1 U19246 ( .B1(n16052), .B2(n16151), .A(n16051), .ZN(n16053) );
  AOI211_X1 U19247 ( .C1(n16057), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16054), .B(n16053), .ZN(n16055) );
  OAI21_X1 U19248 ( .B1(n20176), .B2(n16056), .A(n16055), .ZN(P1_U3005) );
  AOI22_X1 U19249 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16057), .B1(
        n20149), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n16063) );
  INV_X1 U19250 ( .A(n16058), .ZN(n16061) );
  INV_X1 U19251 ( .A(n16059), .ZN(n16060) );
  AOI22_X1 U19252 ( .A1(n16061), .A2(n16182), .B1(n20169), .B2(n16060), .ZN(
        n16062) );
  OAI211_X1 U19253 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n16064), .A(
        n16063), .B(n16062), .ZN(P1_U3006) );
  AOI22_X1 U19254 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16065), .B1(
        n20149), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16071) );
  INV_X1 U19255 ( .A(n16066), .ZN(n16069) );
  INV_X1 U19256 ( .A(n16067), .ZN(n16068) );
  AOI22_X1 U19257 ( .A1(n16069), .A2(n16182), .B1(n20169), .B2(n16068), .ZN(
        n16070) );
  OAI211_X1 U19258 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16072), .A(
        n16071), .B(n16070), .ZN(P1_U3008) );
  AOI22_X1 U19259 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16073), .B1(
        n20149), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16083) );
  INV_X1 U19260 ( .A(n16074), .ZN(n16076) );
  AOI22_X1 U19261 ( .A1(n16076), .A2(n16182), .B1(n20169), .B2(n16075), .ZN(
        n16082) );
  INV_X1 U19262 ( .A(n16077), .ZN(n16079) );
  OAI21_X1 U19263 ( .B1(n16080), .B2(n16079), .A(n16078), .ZN(n16081) );
  NAND3_X1 U19264 ( .A1(n16083), .A2(n16082), .A3(n16081), .ZN(P1_U3012) );
  NOR2_X1 U19265 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16084), .ZN(
        n16089) );
  AOI22_X1 U19266 ( .A1(n16086), .A2(n16182), .B1(n20169), .B2(n16085), .ZN(
        n16088) );
  NAND2_X1 U19267 ( .A1(n20149), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16087) );
  OAI211_X1 U19268 ( .C1(n16090), .C2(n16089), .A(n16088), .B(n16087), .ZN(
        P1_U3014) );
  INV_X1 U19269 ( .A(n16091), .ZN(n16096) );
  INV_X1 U19270 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20800) );
  OAI22_X1 U19271 ( .A1(n16092), .A2(n16151), .B1(n20800), .B2(n20140), .ZN(
        n16095) );
  NOR2_X1 U19272 ( .A1(n16093), .A2(n20176), .ZN(n16094) );
  AOI211_X1 U19273 ( .C1(n16098), .C2(n16096), .A(n16095), .B(n16094), .ZN(
        n16097) );
  OAI21_X1 U19274 ( .B1(n16099), .B2(n16098), .A(n16097), .ZN(P1_U3016) );
  AND2_X1 U19275 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16100), .ZN(
        n16105) );
  INV_X1 U19276 ( .A(n16101), .ZN(n16102) );
  OAI22_X1 U19277 ( .A1(n16102), .A2(n16151), .B1(n21232), .B2(n20140), .ZN(
        n16103) );
  AOI221_X1 U19278 ( .B1(n16105), .B2(n16104), .C1(n16112), .C2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n16103), .ZN(n16106) );
  OAI21_X1 U19279 ( .B1(n16107), .B2(n20176), .A(n16106), .ZN(P1_U3017) );
  INV_X1 U19280 ( .A(n16108), .ZN(n16109) );
  AOI21_X1 U19281 ( .B1(n16110), .B2(n20169), .A(n16109), .ZN(n16114) );
  AOI22_X1 U19282 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16112), .B1(
        n16182), .B2(n16111), .ZN(n16113) );
  OAI211_X1 U19283 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16115), .A(
        n16114), .B(n16113), .ZN(P1_U3018) );
  OR2_X1 U19284 ( .A1(n16119), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16137) );
  NOR2_X1 U19285 ( .A1(n16116), .A2(n16137), .ZN(n16125) );
  OAI21_X1 U19286 ( .B1(n16119), .B2(n16118), .A(n16117), .ZN(n16120) );
  OAI211_X1 U19287 ( .C1(n16127), .C2(n20162), .A(n16121), .B(n16120), .ZN(
        n16134) );
  OAI22_X1 U19288 ( .A1(n16123), .A2(n16151), .B1(n16122), .B2(n20140), .ZN(
        n16124) );
  AOI221_X1 U19289 ( .B1(n16125), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C1(n16134), .C2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16124), .ZN(
        n16130) );
  INV_X1 U19290 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16126) );
  NAND3_X1 U19291 ( .A1(n16128), .A2(n16127), .A3(n16126), .ZN(n16129) );
  OAI211_X1 U19292 ( .C1(n16131), .C2(n20176), .A(n16130), .B(n16129), .ZN(
        P1_U3019) );
  AOI22_X1 U19293 ( .A1(n16132), .A2(n20169), .B1(n20149), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16136) );
  AOI22_X1 U19294 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16134), .B1(
        n16182), .B2(n16133), .ZN(n16135) );
  OAI211_X1 U19295 ( .C1(n16138), .C2(n16137), .A(n16136), .B(n16135), .ZN(
        P1_U3020) );
  OAI211_X1 U19296 ( .C1(n16140), .C2(n16139), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16143), .ZN(n16142) );
  AOI21_X1 U19297 ( .B1(n20157), .B2(n16142), .A(n16141), .ZN(n16158) );
  NAND2_X1 U19298 ( .A1(n16143), .A2(n16164), .ZN(n16150) );
  AOI221_X1 U19299 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12685), .C2(n16157), .A(
        n16150), .ZN(n16146) );
  OAI22_X1 U19300 ( .A1(n16144), .A2(n16151), .B1(n21007), .B2(n20140), .ZN(
        n16145) );
  AOI211_X1 U19301 ( .C1(n16147), .C2(n16182), .A(n16146), .B(n16145), .ZN(
        n16148) );
  OAI21_X1 U19302 ( .B1(n16158), .B2(n12685), .A(n16148), .ZN(P1_U3021) );
  INV_X1 U19303 ( .A(n16149), .ZN(n16155) );
  NOR2_X1 U19304 ( .A1(n16150), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16154) );
  OAI22_X1 U19305 ( .A1(n16152), .A2(n16151), .B1(n21251), .B2(n20140), .ZN(
        n16153) );
  AOI211_X1 U19306 ( .C1(n16155), .C2(n16182), .A(n16154), .B(n16153), .ZN(
        n16156) );
  OAI21_X1 U19307 ( .B1(n16158), .B2(n16157), .A(n16156), .ZN(P1_U3022) );
  INV_X1 U19308 ( .A(n16173), .ZN(n16161) );
  AOI21_X1 U19309 ( .B1(n16161), .B2(n16160), .A(n16159), .ZN(n16163) );
  AOI22_X1 U19310 ( .A1(n10462), .A2(n20169), .B1(n20149), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16167) );
  AOI22_X1 U19311 ( .A1(n16165), .A2(n16182), .B1(n16164), .B2(n16168), .ZN(
        n16166) );
  OAI211_X1 U19312 ( .C1(n16169), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        P1_U3024) );
  NAND2_X1 U19313 ( .A1(n16171), .A2(n16170), .ZN(n16172) );
  AND2_X1 U19314 ( .A1(n16173), .A2(n16172), .ZN(n20084) );
  OAI21_X1 U19315 ( .B1(n16176), .B2(n16175), .A(n16174), .ZN(n16177) );
  AOI21_X1 U19316 ( .B1(n20169), .B2(n20084), .A(n16177), .ZN(n16178) );
  OAI21_X1 U19317 ( .B1(n16180), .B2(n16179), .A(n16178), .ZN(n16181) );
  AOI21_X1 U19318 ( .B1(n16183), .B2(n16182), .A(n16181), .ZN(n16185) );
  NAND2_X1 U19319 ( .A1(n16185), .A2(n16184), .ZN(P1_U3026) );
  INV_X1 U19320 ( .A(n20842), .ZN(n20844) );
  NAND4_X1 U19321 ( .A1(n16189), .A2(n16188), .A3(n16187), .A4(n16186), .ZN(
        n16190) );
  OAI21_X1 U19322 ( .B1(n20844), .B2(n11821), .A(n16190), .ZN(P1_U3468) );
  OAI221_X1 U19323 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n16196), .C2(n20880), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20768) );
  AOI21_X1 U19324 ( .B1(n16192), .B2(n20768), .A(n16191), .ZN(n16193) );
  AOI21_X1 U19325 ( .B1(n16195), .B2(n16194), .A(n16193), .ZN(P1_U3162) );
  NOR2_X1 U19326 ( .A1(n16197), .A2(n16196), .ZN(n20767) );
  OAI21_X1 U19327 ( .B1(n20767), .B2(n20466), .A(n16198), .ZN(P1_U3466) );
  INV_X1 U19328 ( .A(n16199), .ZN(n16202) );
  OAI21_X1 U19329 ( .B1(n16202), .B2(n16201), .A(n16200), .ZN(n16203) );
  AOI22_X1 U19330 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19167), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n16203), .ZN(n16209) );
  INV_X1 U19331 ( .A(n16204), .ZN(n19216) );
  NAND2_X1 U19332 ( .A1(n19108), .A2(n19152), .ZN(n16207) );
  INV_X1 U19333 ( .A(n16205), .ZN(n16206) );
  AOI22_X1 U19334 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19197), .ZN(n16219) );
  AOI22_X1 U19335 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19183), .B1(n16210), 
        .B2(n19205), .ZN(n16218) );
  AOI22_X1 U19336 ( .A1(n16212), .A2(n19199), .B1(n16211), .B2(n19185), .ZN(
        n16217) );
  OAI211_X1 U19337 ( .C1(n16215), .C2(n16214), .A(n19108), .B(n16213), .ZN(
        n16216) );
  NAND4_X1 U19338 ( .A1(n16219), .A2(n16218), .A3(n16217), .A4(n16216), .ZN(
        P2_U2826) );
  INV_X1 U19339 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n16221) );
  AOI22_X1 U19340 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19197), .ZN(n16220) );
  OAI21_X1 U19341 ( .B1(n16221), .B2(n19202), .A(n16220), .ZN(n16224) );
  NOR2_X1 U19342 ( .A1(n16222), .A2(n19158), .ZN(n16223) );
  AOI211_X1 U19343 ( .C1(n19205), .C2(n16225), .A(n16224), .B(n16223), .ZN(
        n16230) );
  OAI211_X1 U19344 ( .C1(n16228), .C2(n16227), .A(n19108), .B(n16226), .ZN(
        n16229) );
  OAI211_X1 U19345 ( .C1(n19207), .C2(n16231), .A(n16230), .B(n16229), .ZN(
        P2_U2827) );
  AOI22_X1 U19346 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19197), .ZN(n16241) );
  AOI22_X1 U19347 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19183), .B1(n16232), 
        .B2(n19205), .ZN(n16240) );
  AOI22_X1 U19348 ( .A1(n16234), .A2(n19199), .B1(n19185), .B2(n16233), .ZN(
        n16239) );
  OAI211_X1 U19349 ( .C1(n16237), .C2(n16236), .A(n19108), .B(n16235), .ZN(
        n16238) );
  NAND4_X1 U19350 ( .A1(n16241), .A2(n16240), .A3(n16239), .A4(n16238), .ZN(
        P2_U2828) );
  AOI22_X1 U19351 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19197), .ZN(n16252) );
  AOI22_X1 U19352 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19183), .B1(n16242), 
        .B2(n19205), .ZN(n16251) );
  NOR2_X1 U19353 ( .A1(n16243), .A2(n19207), .ZN(n16244) );
  AOI21_X1 U19354 ( .B1(n16245), .B2(n19199), .A(n16244), .ZN(n16250) );
  OAI211_X1 U19355 ( .C1(n16248), .C2(n16247), .A(n19108), .B(n16246), .ZN(
        n16249) );
  NAND4_X1 U19356 ( .A1(n16252), .A2(n16251), .A3(n16250), .A4(n16249), .ZN(
        P2_U2829) );
  AOI22_X1 U19357 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19197), .ZN(n16264) );
  INV_X1 U19358 ( .A(n16253), .ZN(n16254) );
  AOI22_X1 U19359 ( .A1(n16254), .A2(n19205), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19183), .ZN(n16263) );
  NOR2_X1 U19360 ( .A1(n16255), .A2(n19207), .ZN(n16256) );
  AOI21_X1 U19361 ( .B1(n16257), .B2(n19199), .A(n16256), .ZN(n16262) );
  OAI211_X1 U19362 ( .C1(n16260), .C2(n16259), .A(n19108), .B(n16258), .ZN(
        n16261) );
  NAND4_X1 U19363 ( .A1(n16264), .A2(n16263), .A3(n16262), .A4(n16261), .ZN(
        P2_U2830) );
  NOR2_X1 U19364 ( .A1(n16265), .A2(n19141), .ZN(n16269) );
  AOI22_X1 U19365 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19197), .ZN(n16266) );
  OAI21_X1 U19366 ( .B1(n16267), .B2(n19202), .A(n16266), .ZN(n16268) );
  AOI211_X1 U19367 ( .C1(n16288), .C2(n19199), .A(n16269), .B(n16268), .ZN(
        n16274) );
  OAI211_X1 U19368 ( .C1(n16272), .C2(n16271), .A(n19108), .B(n16270), .ZN(
        n16273) );
  OAI211_X1 U19369 ( .C1(n19207), .C2(n16275), .A(n16274), .B(n16273), .ZN(
        P2_U2831) );
  AOI22_X1 U19370 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19197), .ZN(n16285) );
  AOI22_X1 U19371 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19183), .B1(n16276), 
        .B2(n19205), .ZN(n16284) );
  AOI22_X1 U19372 ( .A1(n16278), .A2(n19199), .B1(n19185), .B2(n16277), .ZN(
        n16283) );
  OAI211_X1 U19373 ( .C1(n16281), .C2(n16280), .A(n19108), .B(n16279), .ZN(
        n16282) );
  NAND4_X1 U19374 ( .A1(n16285), .A2(n16284), .A3(n16283), .A4(n16282), .ZN(
        P2_U2832) );
  AOI22_X1 U19375 ( .A1(n16286), .A2(n19228), .B1(n19231), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16291) );
  AOI22_X1 U19376 ( .A1(n19217), .A2(BUF1_REG_24__SCAN_IN), .B1(n19215), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16290) );
  AOI22_X1 U19377 ( .A1(n16288), .A2(n19245), .B1(n19246), .B2(n16287), .ZN(
        n16289) );
  NAND3_X1 U19378 ( .A1(n16291), .A2(n16290), .A3(n16289), .ZN(P2_U2895) );
  AOI22_X1 U19379 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19286), .ZN(n16303) );
  NAND2_X1 U19380 ( .A1(n16293), .A2(n16292), .ZN(n16294) );
  NAND2_X1 U19381 ( .A1(n9852), .A2(n16294), .ZN(n16374) );
  AND2_X1 U19382 ( .A1(n16296), .A2(n16295), .ZN(n16297) );
  XNOR2_X1 U19383 ( .A(n16298), .B(n16297), .ZN(n16370) );
  NAND2_X1 U19384 ( .A1(n16370), .A2(n19291), .ZN(n16300) );
  NAND2_X1 U19385 ( .A1(n19290), .A2(n16371), .ZN(n16299) );
  OAI211_X1 U19386 ( .C1(n16374), .C2(n16358), .A(n16300), .B(n16299), .ZN(
        n16301) );
  INV_X1 U19387 ( .A(n16301), .ZN(n16302) );
  OAI211_X1 U19388 ( .C1(n19296), .C2(n19106), .A(n16303), .B(n16302), .ZN(
        P2_U3000) );
  AOI22_X1 U19389 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19286), .B1(n16355), 
        .B2(n16304), .ZN(n16310) );
  OAI22_X1 U19390 ( .A1(n16306), .A2(n16358), .B1(n16356), .B2(n16305), .ZN(
        n16307) );
  AOI21_X1 U19391 ( .B1(n19290), .B2(n16308), .A(n16307), .ZN(n16309) );
  OAI211_X1 U19392 ( .C1(n16365), .C2(n16311), .A(n16310), .B(n16309), .ZN(
        P2_U3001) );
  AOI22_X1 U19393 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19286), .ZN(n16315) );
  AOI222_X1 U19394 ( .A1(n16313), .A2(n10925), .B1(n19291), .B2(n16312), .C1(
        n19290), .C2(n19117), .ZN(n16314) );
  OAI211_X1 U19395 ( .C1(n19296), .C2(n19116), .A(n16315), .B(n16314), .ZN(
        P2_U3002) );
  AOI22_X1 U19396 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19286), .B1(n16355), 
        .B2(n19136), .ZN(n16321) );
  OAI22_X1 U19397 ( .A1(n16317), .A2(n16358), .B1(n16316), .B2(n16356), .ZN(
        n16318) );
  AOI21_X1 U19398 ( .B1(n19290), .B2(n16319), .A(n16318), .ZN(n16320) );
  OAI211_X1 U19399 ( .C1(n16365), .C2(n19126), .A(n16321), .B(n16320), .ZN(
        P2_U3003) );
  AOI22_X1 U19400 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19286), .ZN(n16326) );
  AOI222_X1 U19401 ( .A1(n16324), .A2(n19291), .B1(n19290), .B2(n16323), .C1(
        n10925), .C2(n16322), .ZN(n16325) );
  OAI211_X1 U19402 ( .C1(n19296), .C2(n16327), .A(n16326), .B(n16325), .ZN(
        P2_U3004) );
  AOI22_X1 U19403 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19286), .B1(n16355), 
        .B2(n16328), .ZN(n16334) );
  OAI22_X1 U19404 ( .A1(n16330), .A2(n16358), .B1(n16356), .B2(n16329), .ZN(
        n16331) );
  AOI21_X1 U19405 ( .B1(n19290), .B2(n16332), .A(n16331), .ZN(n16333) );
  OAI211_X1 U19406 ( .C1(n16365), .C2(n16335), .A(n16334), .B(n16333), .ZN(
        P2_U3005) );
  AOI22_X1 U19407 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19286), .ZN(n16346) );
  NAND2_X1 U19408 ( .A1(n16337), .A2(n16336), .ZN(n16342) );
  INV_X1 U19409 ( .A(n16338), .ZN(n16339) );
  AOI21_X1 U19410 ( .B1(n13982), .B2(n16340), .A(n16339), .ZN(n16341) );
  XOR2_X1 U19411 ( .A(n16342), .B(n16341), .Z(n16392) );
  XOR2_X1 U19412 ( .A(n16344), .B(n16343), .Z(n16387) );
  AOI222_X1 U19413 ( .A1(n16392), .A2(n19291), .B1(n19290), .B2(n16389), .C1(
        n10925), .C2(n16387), .ZN(n16345) );
  OAI211_X1 U19414 ( .C1(n19296), .C2(n19145), .A(n16346), .B(n16345), .ZN(
        P2_U3006) );
  AOI22_X1 U19415 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19286), .ZN(n16352) );
  INV_X1 U19416 ( .A(n16347), .ZN(n16350) );
  AOI222_X1 U19417 ( .A1(n10925), .A2(n16350), .B1(n16349), .B2(n19291), .C1(
        n19290), .C2(n16348), .ZN(n16351) );
  OAI211_X1 U19418 ( .C1(n19296), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        P2_U3008) );
  AOI22_X1 U19419 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19286), .B1(n16355), 
        .B2(n16354), .ZN(n16363) );
  OAI22_X1 U19420 ( .A1(n16359), .A2(n16358), .B1(n16357), .B2(n16356), .ZN(
        n16360) );
  AOI21_X1 U19421 ( .B1(n19290), .B2(n16361), .A(n16360), .ZN(n16362) );
  OAI211_X1 U19422 ( .C1(n16365), .C2(n16364), .A(n16363), .B(n16362), .ZN(
        P2_U3009) );
  AOI21_X1 U19423 ( .B1(n16368), .B2(n16367), .A(n16366), .ZN(n19220) );
  AOI22_X1 U19424 ( .A1(n16369), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19308), .B2(n19220), .ZN(n16382) );
  NAND2_X1 U19425 ( .A1(n16370), .A2(n16391), .ZN(n16373) );
  NAND2_X1 U19426 ( .A1(n16390), .A2(n16371), .ZN(n16372) );
  OAI211_X1 U19427 ( .C1(n16374), .C2(n19311), .A(n16373), .B(n16372), .ZN(
        n16375) );
  INV_X1 U19428 ( .A(n16375), .ZN(n16381) );
  NAND2_X1 U19429 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19286), .ZN(n16380) );
  OAI211_X1 U19430 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16378), .A(
        n16377), .B(n16376), .ZN(n16379) );
  NAND4_X1 U19431 ( .A1(n16382), .A2(n16381), .A3(n16380), .A4(n16379), .ZN(
        P2_U3032) );
  AOI21_X1 U19432 ( .B1(n16385), .B2(n16384), .A(n16383), .ZN(n19227) );
  AOI22_X1 U19433 ( .A1(n16386), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19308), .B2(n19227), .ZN(n16398) );
  AOI222_X1 U19434 ( .A1(n16392), .A2(n16391), .B1(n16390), .B2(n16389), .C1(
        n16388), .C2(n16387), .ZN(n16397) );
  NAND2_X1 U19435 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19286), .ZN(n16396) );
  OAI211_X1 U19436 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16394), .B(n16393), .ZN(n16395) );
  NAND4_X1 U19437 ( .A1(n16398), .A2(n16397), .A3(n16396), .A4(n16395), .ZN(
        P2_U3038) );
  INV_X1 U19438 ( .A(n19198), .ZN(n16399) );
  OR2_X1 U19439 ( .A1(n16400), .A2(n16399), .ZN(n16401) );
  OAI21_X1 U19440 ( .B1(n19311), .B2(n16402), .A(n16401), .ZN(n16403) );
  INV_X1 U19441 ( .A(n16403), .ZN(n16409) );
  INV_X1 U19442 ( .A(n19297), .ZN(n16407) );
  OAI22_X1 U19443 ( .A1(n19208), .A2(n19305), .B1(n19300), .B2(n16404), .ZN(
        n16405) );
  AOI211_X1 U19444 ( .C1(n16407), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16406), .B(n16405), .ZN(n16408) );
  OAI211_X1 U19445 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16410), .A(
        n16409), .B(n16408), .ZN(P2_U3046) );
  MUX2_X1 U19446 ( .A(n16414), .B(n16411), .S(n16427), .Z(n16429) );
  MUX2_X1 U19447 ( .A(n16413), .B(n16412), .S(n16427), .Z(n16428) );
  NOR2_X1 U19448 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16428), .ZN(
        n16423) );
  INV_X1 U19449 ( .A(n16414), .ZN(n16419) );
  AOI211_X1 U19450 ( .C1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16416), .A(
        n19994), .B(n16415), .ZN(n16417) );
  OAI21_X1 U19451 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16421), .A(
        n16417), .ZN(n16418) );
  OAI21_X1 U19452 ( .B1(n16419), .B2(n19966), .A(n16418), .ZN(n16420) );
  AOI211_X1 U19453 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16421), .A(
        n16427), .B(n16420), .ZN(n16422) );
  AOI222_X1 U19454 ( .A1(n16423), .A2(n16422), .B1(n16423), .B2(n19973), .C1(
        n16422), .C2(n19973), .ZN(n16424) );
  OAI21_X1 U19455 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16429), .A(
        n16424), .ZN(n16425) );
  AOI22_X1 U19456 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16427), .B1(
        n16426), .B2(n16425), .ZN(n16447) );
  INV_X1 U19457 ( .A(n16428), .ZN(n16445) );
  INV_X1 U19458 ( .A(n16429), .ZN(n16444) );
  NAND2_X1 U19459 ( .A1(n16434), .A2(n16433), .ZN(n16435) );
  AND2_X1 U19460 ( .A1(n16436), .A2(n16435), .ZN(n20002) );
  NAND2_X1 U19461 ( .A1(n16438), .A2(n16437), .ZN(n16442) );
  OAI21_X1 U19462 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16439), .ZN(n16441) );
  NAND4_X1 U19463 ( .A1(n20002), .A2(n16442), .A3(n16441), .A4(n16440), .ZN(
        n16443) );
  AOI21_X1 U19464 ( .B1(n16445), .B2(n16444), .A(n16443), .ZN(n16446) );
  NAND2_X1 U19465 ( .A1(n16447), .A2(n16446), .ZN(n16459) );
  INV_X1 U19466 ( .A(n19998), .ZN(n16448) );
  AOI22_X1 U19467 ( .A1(n19866), .A2(n16459), .B1(n16449), .B2(n16448), .ZN(
        n16467) );
  OR2_X1 U19468 ( .A1(n16451), .A2(n16450), .ZN(n16454) );
  NOR2_X1 U19469 ( .A1(n16452), .A2(n19798), .ZN(n16453) );
  NAND2_X1 U19470 ( .A1(n16454), .A2(n16453), .ZN(n16460) );
  OAI22_X1 U19471 ( .A1(n16457), .A2(n16456), .B1(n16455), .B2(n16460), .ZN(
        n16458) );
  INV_X1 U19472 ( .A(n16458), .ZN(n16463) );
  OAI21_X1 U19473 ( .B1(n16459), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16462) );
  INV_X1 U19474 ( .A(n16460), .ZN(n16461) );
  AND2_X1 U19475 ( .A1(n16462), .A2(n16461), .ZN(n19861) );
  INV_X1 U19476 ( .A(n19861), .ZN(n19864) );
  NAND2_X1 U19477 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19864), .ZN(n16468) );
  OAI21_X1 U19478 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16463), .A(n16468), 
        .ZN(n16465) );
  NAND4_X1 U19479 ( .A1(n16467), .A2(n16466), .A3(n16465), .A4(n16464), .ZN(
        P2_U3176) );
  INV_X1 U19480 ( .A(n16468), .ZN(n16470) );
  OAI21_X1 U19481 ( .B1(n16470), .B2(n19809), .A(n16469), .ZN(P2_U3593) );
  INV_X1 U19482 ( .A(n16471), .ZN(n18807) );
  NOR2_X1 U19483 ( .A1(n17793), .A2(n16474), .ZN(n16482) );
  OAI21_X1 U19484 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17793), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16475) );
  OAI221_X1 U19485 ( .B1(n16517), .B2(n16476), .C1(n17793), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16475), .ZN(n16481) );
  OAI21_X1 U19486 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16517), .A(
        n16476), .ZN(n16479) );
  NAND2_X1 U19487 ( .A1(n17793), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16477) );
  OAI22_X1 U19488 ( .A1(n17793), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n16477), .B2(n16517), .ZN(n16478) );
  OAI21_X1 U19489 ( .B1(n16482), .B2(n16479), .A(n16478), .ZN(n16480) );
  OAI21_X1 U19490 ( .B1(n16482), .B2(n16481), .A(n16480), .ZN(n16526) );
  INV_X1 U19491 ( .A(n17955), .ZN(n17830) );
  INV_X1 U19492 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18961) );
  NOR2_X1 U19493 ( .A1(n18216), .A2(n18961), .ZN(n16520) );
  NAND2_X1 U19494 ( .A1(n18877), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17748) );
  OR2_X1 U19495 ( .A1(n16483), .A2(n17833), .ZN(n16497) );
  XNOR2_X1 U19496 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16485) );
  INV_X1 U19497 ( .A(n17773), .ZN(n17658) );
  NOR2_X1 U19498 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17658), .ZN(
        n16508) );
  INV_X1 U19499 ( .A(n17748), .ZN(n17828) );
  NOR2_X1 U19500 ( .A1(n17987), .A2(n17670), .ZN(n17669) );
  INV_X1 U19501 ( .A(n17669), .ZN(n16674) );
  NOR2_X1 U19502 ( .A1(n16674), .A2(n17671), .ZN(n17631) );
  NAND2_X1 U19503 ( .A1(n17631), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16670) );
  INV_X1 U19504 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17649) );
  NOR2_X1 U19505 ( .A1(n16670), .A2(n17649), .ZN(n16669) );
  NAND2_X1 U19506 ( .A1(n16669), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16668) );
  AOI22_X1 U19507 ( .A1(n17828), .A2(n16668), .B1(n18752), .B2(n16483), .ZN(
        n16484) );
  NAND2_X1 U19508 ( .A1(n16484), .A2(n17995), .ZN(n16509) );
  NOR2_X1 U19509 ( .A1(n16508), .A2(n16509), .ZN(n16496) );
  OAI22_X1 U19510 ( .A1(n16497), .A2(n16485), .B1(n16496), .B2(n16688), .ZN(
        n16486) );
  AOI211_X1 U19511 ( .C1(n17808), .C2(n17001), .A(n16520), .B(n16486), .ZN(
        n16490) );
  NAND2_X1 U19512 ( .A1(n17494), .A2(n17978), .ZN(n17861) );
  INV_X1 U19513 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18986) );
  NOR2_X1 U19514 ( .A1(n16491), .A2(n16517), .ZN(n16487) );
  XNOR2_X1 U19515 ( .A(n18986), .B(n16487), .ZN(n16523) );
  OR2_X1 U19516 ( .A1(n16492), .A2(n16517), .ZN(n16488) );
  XOR2_X1 U19517 ( .A(n16488), .B(n18986), .Z(n16522) );
  AOI22_X1 U19518 ( .A1(n17905), .A2(n16523), .B1(n17986), .B2(n16522), .ZN(
        n16489) );
  OAI211_X1 U19519 ( .C1(n17903), .C2(n16526), .A(n16490), .B(n16489), .ZN(
        P3_U2799) );
  NAND2_X1 U19520 ( .A1(n17905), .A2(n16491), .ZN(n16501) );
  NAND2_X1 U19521 ( .A1(n17986), .A2(n16492), .ZN(n16502) );
  AND2_X1 U19522 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17665), .ZN(
        n17652) );
  INV_X1 U19523 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16692) );
  XNOR2_X1 U19524 ( .A(n16692), .B(n16507), .ZN(n16691) );
  AOI21_X1 U19525 ( .B1(n17808), .B2(n16691), .A(n16494), .ZN(n16495) );
  OAI221_X1 U19526 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16497), .C1(
        n16692), .C2(n16496), .A(n16495), .ZN(n16498) );
  OAI221_X1 U19527 ( .B1(n16517), .B2(n16501), .C1(n16517), .C2(n16502), .A(
        n16500), .ZN(P3_U2800) );
  AOI21_X1 U19528 ( .B1(n16528), .B2(n16518), .A(n16501), .ZN(n16505) );
  INV_X1 U19529 ( .A(n16535), .ZN(n16503) );
  AOI21_X1 U19530 ( .B1(n16503), .B2(n16518), .A(n16502), .ZN(n16504) );
  AOI211_X1 U19531 ( .C1(n17859), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        n16514) );
  INV_X1 U19532 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16702) );
  AOI21_X1 U19533 ( .B1(n16702), .B2(n16668), .A(n16507), .ZN(n16701) );
  OAI21_X1 U19534 ( .B1(n16508), .B2(n17808), .A(n16701), .ZN(n16512) );
  OAI221_X1 U19535 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18752), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16510), .A(n16509), .ZN(
        n16511) );
  NAND4_X1 U19536 ( .A1(n16514), .A2(n16513), .A3(n16512), .A4(n16511), .ZN(
        P3_U2801) );
  OAI21_X1 U19537 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18312), .A(
        n16515), .ZN(n16521) );
  NOR4_X1 U19538 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16518), .A3(
        n16517), .A4(n16516), .ZN(n16519) );
  AOI211_X1 U19539 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16521), .A(
        n16520), .B(n16519), .ZN(n16525) );
  AOI22_X1 U19540 ( .A1(n16523), .A2(n18242), .B1(n16522), .B2(n18322), .ZN(
        n16524) );
  OAI211_X1 U19541 ( .C1(n18229), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        P3_U2831) );
  NAND2_X1 U19542 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18330), .ZN(n17637) );
  NAND2_X1 U19543 ( .A1(n18809), .A2(n17494), .ZN(n18179) );
  INV_X1 U19544 ( .A(n18179), .ZN(n18199) );
  AOI211_X1 U19545 ( .C1(n18199), .C2(n16528), .A(n18056), .B(n16527), .ZN(
        n16534) );
  AOI21_X1 U19546 ( .B1(n17793), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16529), .ZN(n17630) );
  INV_X1 U19547 ( .A(n16530), .ZN(n16541) );
  NAND3_X1 U19548 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18216), .A3(
        n16536), .ZN(n16544) );
  INV_X1 U19549 ( .A(n17628), .ZN(n16537) );
  OAI22_X1 U19550 ( .A1(n18196), .A2(n18811), .B1(n18179), .B2(n18198), .ZN(
        n18113) );
  AOI21_X1 U19551 ( .B1(n18115), .B2(n18113), .A(n18025), .ZN(n18057) );
  OAI211_X1 U19552 ( .C1(n16540), .C2(n18064), .A(n16539), .B(n16538), .ZN(
        n16543) );
  OR3_X1 U19553 ( .A1(n16541), .A2(n18229), .A3(n17630), .ZN(n16542) );
  NAND4_X1 U19554 ( .A1(n17637), .A2(n16544), .A3(n16543), .A4(n16542), .ZN(
        P3_U2834) );
  NOR3_X1 U19555 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16546) );
  NOR4_X1 U19556 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16545) );
  INV_X2 U19557 ( .A(n16637), .ZN(U215) );
  NAND4_X1 U19558 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16546), .A3(n16545), .A4(
        U215), .ZN(U213) );
  INV_X1 U19559 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16639) );
  INV_X2 U19560 ( .A(U214), .ZN(n16600) );
  INV_X1 U19561 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16640) );
  OAI222_X1 U19562 ( .A1(U212), .A2(n16639), .B1(n16602), .B2(n16548), .C1(
        U214), .C2(n16640), .ZN(U216) );
  INV_X1 U19563 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16550) );
  AOI22_X1 U19564 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16585), .ZN(n16549) );
  OAI21_X1 U19565 ( .B1(n16550), .B2(n16602), .A(n16549), .ZN(U217) );
  INV_X1 U19566 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16552) );
  AOI22_X1 U19567 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16585), .ZN(n16551) );
  OAI21_X1 U19568 ( .B1(n16552), .B2(n16602), .A(n16551), .ZN(U218) );
  INV_X1 U19569 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16554) );
  AOI22_X1 U19570 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16585), .ZN(n16553) );
  OAI21_X1 U19571 ( .B1(n16554), .B2(n16602), .A(n16553), .ZN(U219) );
  INV_X1 U19572 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16556) );
  AOI22_X1 U19573 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16585), .ZN(n16555) );
  OAI21_X1 U19574 ( .B1(n16556), .B2(n16602), .A(n16555), .ZN(U220) );
  AOI22_X1 U19575 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16585), .ZN(n16557) );
  OAI21_X1 U19576 ( .B1(n16558), .B2(n16602), .A(n16557), .ZN(U221) );
  INV_X1 U19577 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16560) );
  AOI22_X1 U19578 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16585), .ZN(n16559) );
  OAI21_X1 U19579 ( .B1(n16560), .B2(n16602), .A(n16559), .ZN(U222) );
  AOI22_X1 U19580 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16585), .ZN(n16561) );
  OAI21_X1 U19581 ( .B1(n14564), .B2(n16602), .A(n16561), .ZN(U223) );
  AOI22_X1 U19582 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16585), .ZN(n16562) );
  OAI21_X1 U19583 ( .B1(n15056), .B2(n16602), .A(n16562), .ZN(U224) );
  AOI22_X1 U19584 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16585), .ZN(n16563) );
  OAI21_X1 U19585 ( .B1(n15067), .B2(n16602), .A(n16563), .ZN(U225) );
  AOI22_X1 U19586 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16585), .ZN(n16564) );
  OAI21_X1 U19587 ( .B1(n15074), .B2(n16602), .A(n16564), .ZN(U226) );
  AOI22_X1 U19588 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16585), .ZN(n16565) );
  OAI21_X1 U19589 ( .B1(n15086), .B2(n16602), .A(n16565), .ZN(U227) );
  AOI22_X1 U19590 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16585), .ZN(n16566) );
  OAI21_X1 U19591 ( .B1(n15093), .B2(n16602), .A(n16566), .ZN(U228) );
  INV_X1 U19592 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20199) );
  AOI22_X1 U19593 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16585), .ZN(n16567) );
  OAI21_X1 U19594 ( .B1(n20199), .B2(n16602), .A(n16567), .ZN(U229) );
  AOI22_X1 U19595 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16585), .ZN(n16568) );
  OAI21_X1 U19596 ( .B1(n15111), .B2(n16602), .A(n16568), .ZN(U230) );
  AOI22_X1 U19597 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16585), .ZN(n16569) );
  OAI21_X1 U19598 ( .B1(n13932), .B2(n16602), .A(n16569), .ZN(U231) );
  AOI22_X1 U19599 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16585), .ZN(n16570) );
  OAI21_X1 U19600 ( .B1(n13585), .B2(n16602), .A(n16570), .ZN(U232) );
  AOI22_X1 U19601 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16585), .ZN(n16571) );
  OAI21_X1 U19602 ( .B1(n16572), .B2(n16602), .A(n16571), .ZN(U233) );
  INV_X1 U19603 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16574) );
  AOI22_X1 U19604 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16585), .ZN(n16573) );
  OAI21_X1 U19605 ( .B1(n16574), .B2(n16602), .A(n16573), .ZN(U234) );
  AOI22_X1 U19606 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16585), .ZN(n16575) );
  OAI21_X1 U19607 ( .B1(n16576), .B2(n16602), .A(n16575), .ZN(U235) );
  INV_X1 U19608 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16578) );
  AOI22_X1 U19609 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16585), .ZN(n16577) );
  OAI21_X1 U19610 ( .B1(n16578), .B2(n16602), .A(n16577), .ZN(U236) );
  AOI22_X1 U19611 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16585), .ZN(n16579) );
  OAI21_X1 U19612 ( .B1(n16580), .B2(n16602), .A(n16579), .ZN(U237) );
  INV_X1 U19613 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16582) );
  AOI22_X1 U19614 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16585), .ZN(n16581) );
  OAI21_X1 U19615 ( .B1(n16582), .B2(n16602), .A(n16581), .ZN(U238) );
  AOI22_X1 U19616 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16585), .ZN(n16583) );
  OAI21_X1 U19617 ( .B1(n16584), .B2(n16602), .A(n16583), .ZN(U239) );
  INV_X1 U19618 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16587) );
  AOI22_X1 U19619 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16585), .ZN(n16586) );
  OAI21_X1 U19620 ( .B1(n16587), .B2(n16602), .A(n16586), .ZN(U240) );
  INV_X1 U19621 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16589) );
  AOI22_X1 U19622 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16585), .ZN(n16588) );
  OAI21_X1 U19623 ( .B1(n16589), .B2(n16602), .A(n16588), .ZN(U241) );
  INV_X1 U19624 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16591) );
  AOI22_X1 U19625 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16585), .ZN(n16590) );
  OAI21_X1 U19626 ( .B1(n16591), .B2(n16602), .A(n16590), .ZN(U242) );
  INV_X1 U19627 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U19628 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16585), .ZN(n16592) );
  OAI21_X1 U19629 ( .B1(n16593), .B2(n16602), .A(n16592), .ZN(U243) );
  INV_X1 U19630 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19631 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16585), .ZN(n16594) );
  OAI21_X1 U19632 ( .B1(n16595), .B2(n16602), .A(n16594), .ZN(U244) );
  INV_X1 U19633 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U19634 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16585), .ZN(n16596) );
  OAI21_X1 U19635 ( .B1(n16597), .B2(n16602), .A(n16596), .ZN(U245) );
  INV_X1 U19636 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16599) );
  AOI22_X1 U19637 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16585), .ZN(n16598) );
  OAI21_X1 U19638 ( .B1(n16599), .B2(n16602), .A(n16598), .ZN(U246) );
  INV_X1 U19639 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16603) );
  AOI22_X1 U19640 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16600), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16585), .ZN(n16601) );
  OAI21_X1 U19641 ( .B1(n16603), .B2(n16602), .A(n16601), .ZN(U247) );
  OAI22_X1 U19642 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16637), .ZN(n16604) );
  INV_X1 U19643 ( .A(n16604), .ZN(U251) );
  OAI22_X1 U19644 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16637), .ZN(n16605) );
  INV_X1 U19645 ( .A(n16605), .ZN(U252) );
  OAI22_X1 U19646 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16637), .ZN(n16606) );
  INV_X1 U19647 ( .A(n16606), .ZN(U253) );
  OAI22_X1 U19648 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16637), .ZN(n16607) );
  INV_X1 U19649 ( .A(n16607), .ZN(U254) );
  OAI22_X1 U19650 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16637), .ZN(n16608) );
  INV_X1 U19651 ( .A(n16608), .ZN(U255) );
  OAI22_X1 U19652 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16637), .ZN(n16609) );
  INV_X1 U19653 ( .A(n16609), .ZN(U256) );
  OAI22_X1 U19654 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16637), .ZN(n16610) );
  INV_X1 U19655 ( .A(n16610), .ZN(U257) );
  OAI22_X1 U19656 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16637), .ZN(n16611) );
  INV_X1 U19657 ( .A(n16611), .ZN(U258) );
  OAI22_X1 U19658 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16637), .ZN(n16612) );
  INV_X1 U19659 ( .A(n16612), .ZN(U259) );
  OAI22_X1 U19660 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16631), .ZN(n16613) );
  INV_X1 U19661 ( .A(n16613), .ZN(U260) );
  OAI22_X1 U19662 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16631), .ZN(n16614) );
  INV_X1 U19663 ( .A(n16614), .ZN(U261) );
  OAI22_X1 U19664 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16637), .ZN(n16615) );
  INV_X1 U19665 ( .A(n16615), .ZN(U262) );
  OAI22_X1 U19666 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16637), .ZN(n16616) );
  INV_X1 U19667 ( .A(n16616), .ZN(U263) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16637), .ZN(n16617) );
  INV_X1 U19669 ( .A(n16617), .ZN(U264) );
  OAI22_X1 U19670 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16637), .ZN(n16618) );
  INV_X1 U19671 ( .A(n16618), .ZN(U265) );
  OAI22_X1 U19672 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16631), .ZN(n16619) );
  INV_X1 U19673 ( .A(n16619), .ZN(U266) );
  OAI22_X1 U19674 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16631), .ZN(n16620) );
  INV_X1 U19675 ( .A(n16620), .ZN(U267) );
  OAI22_X1 U19676 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16631), .ZN(n16621) );
  INV_X1 U19677 ( .A(n16621), .ZN(U268) );
  OAI22_X1 U19678 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16631), .ZN(n16622) );
  INV_X1 U19679 ( .A(n16622), .ZN(U269) );
  OAI22_X1 U19680 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16631), .ZN(n16623) );
  INV_X1 U19681 ( .A(n16623), .ZN(U270) );
  OAI22_X1 U19682 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16631), .ZN(n16624) );
  INV_X1 U19683 ( .A(n16624), .ZN(U271) );
  OAI22_X1 U19684 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16637), .ZN(n16625) );
  INV_X1 U19685 ( .A(n16625), .ZN(U272) );
  OAI22_X1 U19686 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16637), .ZN(n16626) );
  INV_X1 U19687 ( .A(n16626), .ZN(U273) );
  OAI22_X1 U19688 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16631), .ZN(n16627) );
  INV_X1 U19689 ( .A(n16627), .ZN(U274) );
  OAI22_X1 U19690 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16637), .ZN(n16628) );
  INV_X1 U19691 ( .A(n16628), .ZN(U275) );
  OAI22_X1 U19692 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16637), .ZN(n16629) );
  INV_X1 U19693 ( .A(n16629), .ZN(U276) );
  OAI22_X1 U19694 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16637), .ZN(n16630) );
  INV_X1 U19695 ( .A(n16630), .ZN(U277) );
  OAI22_X1 U19696 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16631), .ZN(n16632) );
  INV_X1 U19697 ( .A(n16632), .ZN(U278) );
  OAI22_X1 U19698 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16637), .ZN(n16633) );
  INV_X1 U19699 ( .A(n16633), .ZN(U279) );
  OAI22_X1 U19700 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16637), .ZN(n16634) );
  INV_X1 U19701 ( .A(n16634), .ZN(U280) );
  OAI22_X1 U19702 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16637), .ZN(n16636) );
  INV_X1 U19703 ( .A(n16636), .ZN(U281) );
  INV_X1 U19704 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18380) );
  AOI22_X1 U19705 ( .A1(n16637), .A2(n16639), .B1(n18380), .B2(U215), .ZN(U282) );
  INV_X1 U19706 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16638) );
  AOI222_X1 U19707 ( .A1(n16640), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16639), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16638), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16641) );
  INV_X2 U19708 ( .A(n16643), .ZN(n16642) );
  INV_X1 U19709 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18919) );
  INV_X1 U19710 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U19711 ( .A1(n16642), .A2(n18919), .B1(n19909), .B2(n16643), .ZN(
        U347) );
  INV_X1 U19712 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18917) );
  INV_X1 U19713 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U19714 ( .A1(n16642), .A2(n18917), .B1(n19907), .B2(n16643), .ZN(
        U348) );
  INV_X1 U19715 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18914) );
  INV_X1 U19716 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19717 ( .A1(n16642), .A2(n18914), .B1(n19905), .B2(n16643), .ZN(
        U349) );
  INV_X1 U19718 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18913) );
  INV_X1 U19719 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U19720 ( .A1(n16642), .A2(n18913), .B1(n19903), .B2(n16643), .ZN(
        U350) );
  INV_X1 U19721 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18911) );
  INV_X1 U19722 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U19723 ( .A1(n16642), .A2(n18911), .B1(n19901), .B2(n16643), .ZN(
        U351) );
  INV_X1 U19724 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18909) );
  INV_X1 U19725 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U19726 ( .A1(n16642), .A2(n18909), .B1(n19899), .B2(n16643), .ZN(
        U352) );
  INV_X1 U19727 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18907) );
  INV_X1 U19728 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19729 ( .A1(n16642), .A2(n18907), .B1(n19897), .B2(n16643), .ZN(
        U353) );
  INV_X1 U19730 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18905) );
  AOI22_X1 U19731 ( .A1(n16642), .A2(n18905), .B1(n19895), .B2(n16643), .ZN(
        U354) );
  INV_X1 U19732 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18958) );
  INV_X1 U19733 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19945) );
  AOI22_X1 U19734 ( .A1(n16642), .A2(n18958), .B1(n19945), .B2(n16643), .ZN(
        U356) );
  INV_X1 U19735 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18955) );
  INV_X1 U19736 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19943) );
  AOI22_X1 U19737 ( .A1(n16642), .A2(n18955), .B1(n19943), .B2(n16643), .ZN(
        U357) );
  INV_X1 U19738 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18952) );
  INV_X1 U19739 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19940) );
  AOI22_X1 U19740 ( .A1(n16642), .A2(n18952), .B1(n19940), .B2(n16643), .ZN(
        U358) );
  INV_X1 U19741 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18951) );
  INV_X1 U19742 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19939) );
  AOI22_X1 U19743 ( .A1(n16642), .A2(n18951), .B1(n19939), .B2(n16643), .ZN(
        U359) );
  INV_X1 U19744 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18949) );
  INV_X1 U19745 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19937) );
  AOI22_X1 U19746 ( .A1(n16642), .A2(n18949), .B1(n19937), .B2(n16643), .ZN(
        U360) );
  INV_X1 U19747 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18947) );
  INV_X1 U19748 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19935) );
  AOI22_X1 U19749 ( .A1(n16642), .A2(n18947), .B1(n19935), .B2(n16643), .ZN(
        U361) );
  INV_X1 U19750 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18944) );
  INV_X1 U19751 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19933) );
  AOI22_X1 U19752 ( .A1(n16642), .A2(n18944), .B1(n19933), .B2(n16643), .ZN(
        U362) );
  INV_X1 U19753 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18943) );
  INV_X1 U19754 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U19755 ( .A1(n16642), .A2(n18943), .B1(n19931), .B2(n16643), .ZN(
        U363) );
  INV_X1 U19756 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18941) );
  INV_X1 U19757 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U19758 ( .A1(n16642), .A2(n18941), .B1(n19930), .B2(n16643), .ZN(
        U364) );
  INV_X1 U19759 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18902) );
  INV_X1 U19760 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U19761 ( .A1(n16642), .A2(n18902), .B1(n19893), .B2(n16643), .ZN(
        U365) );
  INV_X1 U19762 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18939) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19928) );
  AOI22_X1 U19764 ( .A1(n16642), .A2(n18939), .B1(n19928), .B2(n16643), .ZN(
        U366) );
  INV_X1 U19765 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18937) );
  INV_X1 U19766 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19926) );
  AOI22_X1 U19767 ( .A1(n16642), .A2(n18937), .B1(n19926), .B2(n16643), .ZN(
        U367) );
  INV_X1 U19768 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18935) );
  INV_X1 U19769 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19924) );
  AOI22_X1 U19770 ( .A1(n16642), .A2(n18935), .B1(n19924), .B2(n16643), .ZN(
        U368) );
  INV_X1 U19771 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18932) );
  INV_X1 U19772 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19922) );
  AOI22_X1 U19773 ( .A1(n16642), .A2(n18932), .B1(n19922), .B2(n16643), .ZN(
        U369) );
  INV_X1 U19774 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18931) );
  INV_X1 U19775 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19920) );
  AOI22_X1 U19776 ( .A1(n16642), .A2(n18931), .B1(n19920), .B2(n16643), .ZN(
        U370) );
  INV_X1 U19777 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18929) );
  INV_X1 U19778 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19918) );
  AOI22_X1 U19779 ( .A1(n16642), .A2(n18929), .B1(n19918), .B2(n16643), .ZN(
        U371) );
  INV_X1 U19780 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18926) );
  INV_X1 U19781 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19916) );
  AOI22_X1 U19782 ( .A1(n16642), .A2(n18926), .B1(n19916), .B2(n16643), .ZN(
        U372) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18925) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19785 ( .A1(n16642), .A2(n18925), .B1(n19914), .B2(n16643), .ZN(
        U373) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18923) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U19788 ( .A1(n16642), .A2(n18923), .B1(n19913), .B2(n16643), .ZN(
        U374) );
  INV_X1 U19789 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18921) );
  INV_X1 U19790 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19911) );
  AOI22_X1 U19791 ( .A1(n16642), .A2(n18921), .B1(n19911), .B2(n16643), .ZN(
        U375) );
  INV_X1 U19792 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18900) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19794 ( .A1(n16642), .A2(n18900), .B1(n19891), .B2(n16643), .ZN(
        U376) );
  INV_X1 U19795 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18899) );
  NAND2_X1 U19796 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18899), .ZN(n18890) );
  AOI22_X1 U19797 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18890), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18897), .ZN(n18971) );
  AOI21_X1 U19798 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18971), .ZN(n16644) );
  INV_X1 U19799 ( .A(n16644), .ZN(P3_U2633) );
  OAI21_X1 U19800 ( .B1(n16645), .B2(n17560), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16646) );
  OAI21_X1 U19801 ( .B1(n16647), .B2(n17994), .A(n16646), .ZN(P3_U2634) );
  AOI21_X1 U19802 ( .B1(n18897), .B2(n18899), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16648) );
  AOI22_X1 U19803 ( .A1(n18966), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16648), 
        .B2(n19033), .ZN(P3_U2635) );
  OAI21_X1 U19804 ( .B1(n18885), .B2(BS16), .A(n18971), .ZN(n18969) );
  OAI21_X1 U19805 ( .B1(n18971), .B2(n19024), .A(n18969), .ZN(P3_U2636) );
  AND3_X1 U19806 ( .A1(n18806), .A2(n16650), .A3(n16649), .ZN(n18813) );
  NOR2_X1 U19807 ( .A1(n18813), .A2(n18874), .ZN(n19017) );
  INV_X1 U19808 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18337) );
  OAI21_X1 U19809 ( .B1(n19017), .B2(n18337), .A(n16651), .ZN(P3_U2637) );
  NOR4_X1 U19810 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16655) );
  NOR4_X1 U19811 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16654) );
  NOR4_X1 U19812 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16653) );
  NOR4_X1 U19813 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16652) );
  NAND4_X1 U19814 ( .A1(n16655), .A2(n16654), .A3(n16653), .A4(n16652), .ZN(
        n16661) );
  NOR4_X1 U19815 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16659) );
  AOI211_X1 U19816 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16658) );
  NOR4_X1 U19817 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16657) );
  NOR4_X1 U19818 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16656) );
  NAND4_X1 U19819 ( .A1(n16659), .A2(n16658), .A3(n16657), .A4(n16656), .ZN(
        n16660) );
  NOR2_X1 U19820 ( .A1(n16661), .A2(n16660), .ZN(n19015) );
  INV_X1 U19821 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16663) );
  NOR3_X1 U19822 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16664) );
  OAI21_X1 U19823 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16664), .A(n19015), .ZN(
        n16662) );
  OAI21_X1 U19824 ( .B1(n19015), .B2(n16663), .A(n16662), .ZN(P3_U2638) );
  INV_X1 U19825 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18970) );
  AOI21_X1 U19826 ( .B1(n19008), .B2(n18970), .A(n16664), .ZN(n16666) );
  INV_X1 U19827 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16665) );
  INV_X1 U19828 ( .A(n19015), .ZN(n19010) );
  AOI22_X1 U19829 ( .A1(n19015), .A2(n16666), .B1(n16665), .B2(n19010), .ZN(
        P3_U2639) );
  INV_X1 U19830 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18948) );
  INV_X1 U19831 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18945) );
  INV_X1 U19832 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18924) );
  INV_X1 U19833 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18920) );
  INV_X1 U19834 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18910) );
  INV_X1 U19835 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18906) );
  NAND3_X1 U19836 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16990) );
  NOR2_X1 U19837 ( .A1(n18906), .A2(n16990), .ZN(n16973) );
  NAND2_X1 U19838 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16973), .ZN(n16967) );
  NOR2_X1 U19839 ( .A1(n18910), .A2(n16967), .ZN(n16939) );
  NAND3_X1 U19840 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(n16939), .ZN(n16911) );
  INV_X1 U19841 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18918) );
  INV_X1 U19842 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18916) );
  NOR2_X1 U19843 ( .A1(n18918), .A2(n18916), .ZN(n16901) );
  INV_X1 U19844 ( .A(n16901), .ZN(n16912) );
  NOR3_X1 U19845 ( .A1(n18920), .A2(n16911), .A3(n16912), .ZN(n16875) );
  NAND2_X1 U19846 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16875), .ZN(n16876) );
  NOR2_X1 U19847 ( .A1(n18924), .A2(n16876), .ZN(n16868) );
  NAND2_X1 U19848 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16868), .ZN(n16774) );
  INV_X1 U19849 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18940) );
  INV_X1 U19850 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18933) );
  NAND2_X1 U19851 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16830) );
  NOR2_X1 U19852 ( .A1(n18933), .A2(n16830), .ZN(n16776) );
  NAND4_X1 U19853 ( .A1(n16776), .A2(P3_REIP_REG_20__SCAN_IN), .A3(
        P3_REIP_REG_19__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16775) );
  NOR2_X1 U19854 ( .A1(n18940), .A2(n16775), .ZN(n16778) );
  NAND2_X1 U19855 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16778), .ZN(n16763) );
  NOR3_X1 U19856 ( .A1(n18945), .A2(n16774), .A3(n16763), .ZN(n16755) );
  NAND2_X1 U19857 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16755), .ZN(n16746) );
  NOR2_X1 U19858 ( .A1(n18948), .A2(n16746), .ZN(n16732) );
  NAND2_X1 U19859 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16732), .ZN(n16680) );
  NOR2_X1 U19860 ( .A1(n17026), .A2(n16680), .ZN(n16727) );
  NAND4_X1 U19861 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16727), .ZN(n16682) );
  NOR3_X1 U19862 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18959), .A3(n16682), 
        .ZN(n16667) );
  AOI21_X1 U19863 ( .B1(n17014), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16667), .ZN(
        n16687) );
  NOR3_X1 U19864 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17024) );
  NAND2_X1 U19865 ( .A1(n17024), .A2(n17008), .ZN(n17006) );
  NOR2_X1 U19866 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17006), .ZN(n16989) );
  NAND2_X1 U19867 ( .A1(n16989), .A2(n16985), .ZN(n16982) );
  NAND2_X1 U19868 ( .A1(n16965), .A2(n17344), .ZN(n16956) );
  NAND2_X1 U19869 ( .A1(n16938), .A2(n16933), .ZN(n16932) );
  NAND2_X1 U19870 ( .A1(n16910), .A2(n17277), .ZN(n16906) );
  INV_X1 U19871 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16882) );
  NAND2_X1 U19872 ( .A1(n16889), .A2(n16882), .ZN(n16881) );
  INV_X1 U19873 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16860) );
  NAND2_X1 U19874 ( .A1(n16865), .A2(n16860), .ZN(n16859) );
  INV_X1 U19875 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16839) );
  NAND2_X1 U19876 ( .A1(n16845), .A2(n16839), .ZN(n16838) );
  INV_X1 U19877 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16816) );
  NAND2_X1 U19878 ( .A1(n16823), .A2(n16816), .ZN(n16815) );
  NAND2_X1 U19879 ( .A1(n16796), .A2(n16791), .ZN(n16789) );
  INV_X1 U19880 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17099) );
  NAND2_X1 U19881 ( .A1(n16782), .A2(n17099), .ZN(n16770) );
  NAND2_X1 U19882 ( .A1(n16756), .A2(n16750), .ZN(n16749) );
  NOR2_X1 U19883 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16749), .ZN(n16733) );
  NAND2_X1 U19884 ( .A1(n16733), .A2(n16729), .ZN(n16728) );
  NOR2_X1 U19885 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16728), .ZN(n16712) );
  INV_X1 U19886 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16708) );
  NAND2_X1 U19887 ( .A1(n16712), .A2(n16708), .ZN(n16689) );
  NOR2_X1 U19888 ( .A1(n17036), .A2(n16689), .ZN(n16696) );
  INV_X1 U19889 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17049) );
  OAI21_X1 U19890 ( .B1(n16669), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16668), .ZN(n17638) );
  INV_X1 U19891 ( .A(n17638), .ZN(n16715) );
  AOI21_X1 U19892 ( .B1(n16670), .B2(n17649), .A(n16669), .ZN(n17645) );
  OAI21_X1 U19893 ( .B1(n17631), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16670), .ZN(n16671) );
  INV_X1 U19894 ( .A(n16671), .ZN(n17659) );
  INV_X1 U19895 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17683) );
  NOR2_X1 U19896 ( .A1(n16674), .A2(n17683), .ZN(n16673) );
  INV_X1 U19897 ( .A(n17631), .ZN(n16672) );
  OAI21_X1 U19898 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16673), .A(
        n16672), .ZN(n17673) );
  INV_X1 U19899 ( .A(n17673), .ZN(n16744) );
  AOI21_X1 U19900 ( .B1(n16674), .B2(n17683), .A(n16673), .ZN(n17681) );
  INV_X1 U19901 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17713) );
  NAND3_X1 U19902 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17710), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16675) );
  NOR2_X1 U19903 ( .A1(n17713), .A2(n16675), .ZN(n17695) );
  OAI21_X1 U19904 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17695), .A(
        n16674), .ZN(n17707) );
  INV_X1 U19905 ( .A(n17707), .ZN(n16766) );
  AOI21_X1 U19906 ( .B1(n17713), .B2(n16675), .A(n17695), .ZN(n17716) );
  INV_X1 U19907 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17724) );
  NAND2_X1 U19908 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17710), .ZN(
        n16677) );
  INV_X1 U19909 ( .A(n16675), .ZN(n16676) );
  AOI21_X1 U19910 ( .B1(n17724), .B2(n16677), .A(n16676), .ZN(n17727) );
  INV_X1 U19911 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17766) );
  INV_X1 U19912 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17750) );
  INV_X1 U19913 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17800) );
  INV_X1 U19914 ( .A(n16678), .ZN(n17814) );
  NAND2_X1 U19915 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17814), .ZN(
        n16974) );
  NOR2_X1 U19916 ( .A1(n17929), .A2(n16974), .ZN(n16959) );
  NAND2_X1 U19917 ( .A1(n17831), .A2(n16959), .ZN(n17827) );
  INV_X1 U19918 ( .A(n17827), .ZN(n16899) );
  NAND2_X1 U19919 ( .A1(n16863), .A2(n16899), .ZN(n16877) );
  INV_X1 U19920 ( .A(n16877), .ZN(n16864) );
  NAND2_X1 U19921 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16864), .ZN(
        n17785) );
  NOR2_X1 U19922 ( .A1(n17800), .A2(n17785), .ZN(n16852) );
  NAND2_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16852), .ZN(
        n16843) );
  NOR2_X1 U19924 ( .A1(n17775), .A2(n16843), .ZN(n17749) );
  INV_X1 U19925 ( .A(n17749), .ZN(n16819) );
  NOR3_X1 U19926 ( .A1(n17766), .A2(n17750), .A3(n16819), .ZN(n16679) );
  INV_X1 U19927 ( .A(n16679), .ZN(n17708) );
  AOI22_X1 U19928 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17710), .B1(
        n17736), .B2(n17708), .ZN(n17738) );
  INV_X1 U19929 ( .A(n16852), .ZN(n16834) );
  OAI21_X1 U19930 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16834), .A(
        n17001), .ZN(n16853) );
  OAI21_X1 U19931 ( .B1(n16679), .B2(n16975), .A(n16853), .ZN(n16800) );
  NOR2_X1 U19932 ( .A1(n17716), .A2(n16781), .ZN(n16780) );
  NOR2_X1 U19933 ( .A1(n16780), .A2(n16975), .ZN(n16765) );
  NOR2_X1 U19934 ( .A1(n16766), .A2(n16765), .ZN(n16764) );
  NOR2_X1 U19935 ( .A1(n16764), .A2(n16975), .ZN(n16758) );
  NOR2_X1 U19936 ( .A1(n17681), .A2(n16758), .ZN(n16757) );
  NOR2_X1 U19937 ( .A1(n16757), .A2(n16975), .ZN(n16743) );
  NOR2_X1 U19938 ( .A1(n16744), .A2(n16743), .ZN(n16742) );
  NOR2_X1 U19939 ( .A1(n16742), .A2(n16975), .ZN(n16735) );
  NOR2_X1 U19940 ( .A1(n17659), .A2(n16735), .ZN(n16734) );
  NOR2_X1 U19941 ( .A1(n16734), .A2(n16975), .ZN(n16724) );
  NOR2_X1 U19942 ( .A1(n17645), .A2(n16724), .ZN(n16723) );
  NOR2_X1 U19943 ( .A1(n16699), .A2(n16975), .ZN(n16690) );
  NAND2_X1 U19944 ( .A1(n17001), .A2(n18878), .ZN(n16961) );
  NOR3_X1 U19945 ( .A1(n16691), .A2(n16690), .A3(n16961), .ZN(n16685) );
  NAND3_X1 U19946 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16681) );
  AOI21_X1 U19947 ( .B1(n16680), .B2(n16998), .A(n17035), .ZN(n16741) );
  INV_X1 U19948 ( .A(n16741), .ZN(n16718) );
  AOI21_X1 U19949 ( .B1(n16998), .B2(n16681), .A(n16718), .ZN(n16711) );
  NOR2_X1 U19950 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16682), .ZN(n16694) );
  INV_X1 U19951 ( .A(n16694), .ZN(n16683) );
  AOI21_X1 U19952 ( .B1(n16711), .B2(n16683), .A(n18961), .ZN(n16684) );
  AOI211_X1 U19953 ( .C1(n16696), .C2(n17049), .A(n16685), .B(n16684), .ZN(
        n16686) );
  OAI211_X1 U19954 ( .C1(n16688), .C2(n17003), .A(n16687), .B(n16686), .ZN(
        P3_U2640) );
  NAND2_X1 U19955 ( .A1(n17007), .A2(n16689), .ZN(n16706) );
  XOR2_X1 U19956 ( .A(n16691), .B(n16690), .Z(n16695) );
  OAI22_X1 U19957 ( .A1(n16711), .A2(n18959), .B1(n16692), .B2(n17003), .ZN(
        n16693) );
  AOI211_X1 U19958 ( .C1(n16695), .C2(n18878), .A(n16694), .B(n16693), .ZN(
        n16698) );
  OAI21_X1 U19959 ( .B1(n17014), .B2(n16696), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16697) );
  INV_X1 U19960 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18957) );
  AOI211_X1 U19961 ( .C1(n16701), .C2(n16700), .A(n16699), .B(n17019), .ZN(
        n16705) );
  NAND3_X1 U19962 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16727), .ZN(n16703) );
  OAI22_X1 U19963 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16703), .B1(n16702), 
        .B2(n17003), .ZN(n16704) );
  AOI211_X1 U19964 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17014), .A(n16705), .B(
        n16704), .ZN(n16710) );
  INV_X1 U19965 ( .A(n16706), .ZN(n16707) );
  OAI21_X1 U19966 ( .B1(n16712), .B2(n16708), .A(n16707), .ZN(n16709) );
  OAI211_X1 U19967 ( .C1(n16711), .C2(n18957), .A(n16710), .B(n16709), .ZN(
        P3_U2642) );
  AOI22_X1 U19968 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17030), .B1(
        n17014), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16722) );
  AOI211_X1 U19969 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16728), .A(n16712), .B(
        n17036), .ZN(n16717) );
  AOI211_X1 U19970 ( .C1(n16715), .C2(n16714), .A(n16713), .B(n17019), .ZN(
        n16716) );
  AOI211_X1 U19971 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16718), .A(n16717), 
        .B(n16716), .ZN(n16721) );
  NAND2_X1 U19972 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16719) );
  OAI211_X1 U19973 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16727), .B(n16719), .ZN(n16720) );
  NAND3_X1 U19974 ( .A1(n16722), .A2(n16721), .A3(n16720), .ZN(P3_U2643) );
  INV_X1 U19975 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18953) );
  AOI211_X1 U19976 ( .C1(n17645), .C2(n16724), .A(n16723), .B(n17019), .ZN(
        n16726) );
  OAI22_X1 U19977 ( .A1(n17649), .A2(n17003), .B1(n17037), .B2(n16729), .ZN(
        n16725) );
  AOI211_X1 U19978 ( .C1(n16727), .C2(n18953), .A(n16726), .B(n16725), .ZN(
        n16731) );
  OAI211_X1 U19979 ( .C1(n16733), .C2(n16729), .A(n17007), .B(n16728), .ZN(
        n16730) );
  OAI211_X1 U19980 ( .C1(n16741), .C2(n18953), .A(n16731), .B(n16730), .ZN(
        P3_U2644) );
  AOI21_X1 U19981 ( .B1(n16998), .B2(n16732), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16740) );
  AOI22_X1 U19982 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17030), .B1(
        n17014), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16739) );
  AOI211_X1 U19983 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16749), .A(n16733), .B(
        n17036), .ZN(n16737) );
  AOI211_X1 U19984 ( .C1(n17659), .C2(n16735), .A(n16734), .B(n17019), .ZN(
        n16736) );
  NOR2_X1 U19985 ( .A1(n16737), .A2(n16736), .ZN(n16738) );
  OAI211_X1 U19986 ( .C1(n16741), .C2(n16740), .A(n16739), .B(n16738), .ZN(
        P3_U2645) );
  INV_X1 U19987 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18946) );
  OAI21_X1 U19988 ( .B1(n16755), .B2(n17026), .A(n17017), .ZN(n16768) );
  AOI21_X1 U19989 ( .B1(n16998), .B2(n18946), .A(n16768), .ZN(n16753) );
  AOI211_X1 U19990 ( .C1(n16744), .C2(n16743), .A(n16742), .B(n17019), .ZN(
        n16748) );
  NAND2_X1 U19991 ( .A1(n16998), .A2(n18948), .ZN(n16745) );
  OAI22_X1 U19992 ( .A1(n17037), .A2(n16750), .B1(n16746), .B2(n16745), .ZN(
        n16747) );
  AOI211_X1 U19993 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16748), .B(n16747), .ZN(n16752) );
  OAI211_X1 U19994 ( .C1(n16756), .C2(n16750), .A(n17007), .B(n16749), .ZN(
        n16751) );
  OAI211_X1 U19995 ( .C1(n16753), .C2(n18948), .A(n16752), .B(n16751), .ZN(
        P3_U2646) );
  NOR2_X1 U19996 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17026), .ZN(n16754) );
  AOI22_X1 U19997 ( .A1(n17014), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16755), 
        .B2(n16754), .ZN(n16762) );
  AOI211_X1 U19998 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16770), .A(n16756), .B(
        n17036), .ZN(n16760) );
  AOI211_X1 U19999 ( .C1(n17681), .C2(n16758), .A(n16757), .B(n17019), .ZN(
        n16759) );
  AOI211_X1 U20000 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16768), .A(n16760), 
        .B(n16759), .ZN(n16761) );
  OAI211_X1 U20001 ( .C1(n17683), .C2(n17003), .A(n16762), .B(n16761), .ZN(
        P3_U2647) );
  AOI22_X1 U20002 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17030), .B1(
        n17014), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16773) );
  NAND3_X1 U20003 ( .A1(n16998), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16868), 
        .ZN(n16848) );
  NOR2_X1 U20004 ( .A1(n16763), .A2(n16848), .ZN(n16769) );
  AOI211_X1 U20005 ( .C1(n16766), .C2(n16765), .A(n16764), .B(n17019), .ZN(
        n16767) );
  AOI221_X1 U20006 ( .B1(n16769), .B2(n18945), .C1(n16768), .C2(
        P3_REIP_REG_23__SCAN_IN), .A(n16767), .ZN(n16772) );
  OAI211_X1 U20007 ( .C1(n16782), .C2(n17099), .A(n17007), .B(n16770), .ZN(
        n16771) );
  NAND3_X1 U20008 ( .A1(n16773), .A2(n16772), .A3(n16771), .ZN(P3_U2648) );
  INV_X1 U20009 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18942) );
  OR2_X1 U20010 ( .A1(n16774), .A2(n17035), .ZN(n16869) );
  NAND2_X1 U20011 ( .A1(n17017), .A2(n17026), .ZN(n17040) );
  OAI21_X1 U20012 ( .B1(n16775), .B2(n16869), .A(n17040), .ZN(n16805) );
  INV_X1 U20013 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18938) );
  NAND2_X1 U20014 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16807) );
  NOR2_X1 U20015 ( .A1(n18938), .A2(n16807), .ZN(n16777) );
  INV_X1 U20016 ( .A(n16776), .ZN(n16806) );
  NOR2_X1 U20017 ( .A1(n16806), .A2(n16848), .ZN(n16798) );
  NAND3_X1 U20018 ( .A1(n16777), .A2(n16798), .A3(n18940), .ZN(n16794) );
  INV_X1 U20019 ( .A(n16778), .ZN(n16779) );
  NOR3_X1 U20020 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16779), .A3(n16848), 
        .ZN(n16786) );
  AOI211_X1 U20021 ( .C1(n17716), .C2(n16781), .A(n16780), .B(n17019), .ZN(
        n16785) );
  AOI211_X1 U20022 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16789), .A(n16782), .B(
        n17036), .ZN(n16784) );
  INV_X1 U20023 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17098) );
  OAI22_X1 U20024 ( .A1(n17713), .A2(n17003), .B1(n17037), .B2(n17098), .ZN(
        n16783) );
  NOR4_X1 U20025 ( .A1(n16786), .A2(n16785), .A3(n16784), .A4(n16783), .ZN(
        n16787) );
  OAI221_X1 U20026 ( .B1(n18942), .B2(n16805), .C1(n18942), .C2(n16794), .A(
        n16787), .ZN(P3_U2649) );
  AOI211_X1 U20027 ( .C1(n17727), .C2(n16788), .A(n9912), .B(n17019), .ZN(
        n16793) );
  OAI211_X1 U20028 ( .C1(n16796), .C2(n16791), .A(n17007), .B(n16789), .ZN(
        n16790) );
  OAI21_X1 U20029 ( .B1(n16791), .B2(n17037), .A(n16790), .ZN(n16792) );
  AOI211_X1 U20030 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16793), .B(n16792), .ZN(n16795) );
  OAI211_X1 U20031 ( .C1(n16805), .C2(n18940), .A(n16795), .B(n16794), .ZN(
        P3_U2650) );
  AOI211_X1 U20032 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16815), .A(n16796), .B(
        n17036), .ZN(n16797) );
  AOI21_X1 U20033 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17014), .A(n16797), .ZN(
        n16804) );
  INV_X1 U20034 ( .A(n16798), .ZN(n16829) );
  NOR3_X1 U20035 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16807), .A3(n16829), 
        .ZN(n16802) );
  AOI211_X1 U20036 ( .C1(n17738), .C2(n16800), .A(n16799), .B(n17019), .ZN(
        n16801) );
  AOI211_X1 U20037 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16802), .B(n16801), .ZN(n16803) );
  OAI211_X1 U20038 ( .C1(n18938), .C2(n16805), .A(n16804), .B(n16803), .ZN(
        P3_U2651) );
  OAI21_X1 U20039 ( .B1(n16806), .B2(n16869), .A(n17040), .ZN(n16828) );
  INV_X1 U20040 ( .A(n16828), .ZN(n16833) );
  INV_X1 U20041 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18936) );
  INV_X1 U20042 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18934) );
  INV_X1 U20043 ( .A(n16807), .ZN(n16808) );
  AOI211_X1 U20044 ( .C1(n18936), .C2(n18934), .A(n16808), .B(n16829), .ZN(
        n16814) );
  NOR2_X1 U20045 ( .A1(n17766), .A2(n16819), .ZN(n16809) );
  OAI21_X1 U20046 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16809), .A(
        n17708), .ZN(n17752) );
  INV_X1 U20047 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17034) );
  NAND2_X1 U20048 ( .A1(n17749), .A2(n17034), .ZN(n16820) );
  OAI21_X1 U20049 ( .B1(n17766), .B2(n16820), .A(n17001), .ZN(n16811) );
  AOI21_X1 U20050 ( .B1(n17752), .B2(n16811), .A(n17019), .ZN(n16810) );
  OAI21_X1 U20051 ( .B1(n17752), .B2(n16811), .A(n16810), .ZN(n16812) );
  OAI211_X1 U20052 ( .C1(n17037), .C2(n16816), .A(n18216), .B(n16812), .ZN(
        n16813) );
  AOI211_X1 U20053 ( .C1(n16833), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16814), 
        .B(n16813), .ZN(n16818) );
  OAI211_X1 U20054 ( .C1(n16823), .C2(n16816), .A(n17007), .B(n16815), .ZN(
        n16817) );
  OAI211_X1 U20055 ( .C1(n17003), .C2(n17750), .A(n16818), .B(n16817), .ZN(
        P3_U2652) );
  AOI22_X1 U20056 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16819), .B1(
        n17749), .B2(n17766), .ZN(n17763) );
  NAND2_X1 U20057 ( .A1(n17001), .A2(n16820), .ZN(n16822) );
  OAI21_X1 U20058 ( .B1(n17763), .B2(n16822), .A(n18878), .ZN(n16821) );
  AOI21_X1 U20059 ( .B1(n17763), .B2(n16822), .A(n16821), .ZN(n16826) );
  AOI211_X1 U20060 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16838), .A(n16823), .B(
        n17036), .ZN(n16825) );
  OAI22_X1 U20061 ( .A1(n17766), .A2(n17003), .B1(n17037), .B2(n17170), .ZN(
        n16824) );
  NOR4_X1 U20062 ( .A1(n18330), .A2(n16826), .A3(n16825), .A4(n16824), .ZN(
        n16827) );
  OAI221_X1 U20063 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16829), .C1(n18934), 
        .C2(n16828), .A(n16827), .ZN(P3_U2653) );
  NOR2_X1 U20064 ( .A1(n16830), .A2(n16848), .ZN(n16832) );
  OAI22_X1 U20065 ( .A1(n17775), .A2(n17003), .B1(n17037), .B2(n16839), .ZN(
        n16831) );
  AOI221_X1 U20066 ( .B1(n16833), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16832), 
        .C2(n18933), .A(n16831), .ZN(n16842) );
  AOI21_X1 U20067 ( .B1(n17775), .B2(n16843), .A(n17749), .ZN(n17778) );
  NOR2_X1 U20068 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16834), .ZN(
        n16835) );
  AOI21_X1 U20069 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16835), .A(
        n16975), .ZN(n16837) );
  AOI21_X1 U20070 ( .B1(n17778), .B2(n16837), .A(n17019), .ZN(n16836) );
  OAI21_X1 U20071 ( .B1(n17778), .B2(n16837), .A(n16836), .ZN(n16841) );
  OAI211_X1 U20072 ( .C1(n16845), .C2(n16839), .A(n17007), .B(n16838), .ZN(
        n16840) );
  NAND4_X1 U20073 ( .A1(n16842), .A2(n18216), .A3(n16841), .A4(n16840), .ZN(
        P3_U2654) );
  OAI21_X1 U20074 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16852), .A(
        n16843), .ZN(n17786) );
  XOR2_X1 U20075 ( .A(n16853), .B(n17786), .Z(n16844) );
  AOI22_X1 U20076 ( .A1(n17014), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n18878), 
        .B2(n16844), .ZN(n16851) );
  INV_X1 U20077 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18928) );
  NOR3_X1 U20078 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18928), .A3(n16848), 
        .ZN(n16847) );
  AOI211_X1 U20079 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16859), .A(n16845), .B(
        n17036), .ZN(n16846) );
  AOI211_X1 U20080 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16847), .B(n16846), .ZN(n16850) );
  AND2_X1 U20081 ( .A1(n17040), .A2(n16869), .ZN(n16871) );
  NOR2_X1 U20082 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16848), .ZN(n16858) );
  OAI21_X1 U20083 ( .B1(n16871), .B2(n16858), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16849) );
  NAND4_X1 U20084 ( .A1(n16851), .A2(n16850), .A3(n18216), .A4(n16849), .ZN(
        P3_U2655) );
  AOI21_X1 U20085 ( .B1(n17800), .B2(n17785), .A(n16852), .ZN(n17807) );
  AOI21_X1 U20086 ( .B1(n17001), .B2(n17785), .A(n16960), .ZN(n16855) );
  NOR3_X1 U20087 ( .A1(n17807), .A2(n16853), .A3(n17019), .ZN(n16854) );
  AOI211_X1 U20088 ( .C1(n17807), .C2(n16855), .A(n18330), .B(n16854), .ZN(
        n16856) );
  OAI21_X1 U20089 ( .B1(n17037), .B2(n16860), .A(n16856), .ZN(n16857) );
  AOI211_X1 U20090 ( .C1(n16871), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16858), 
        .B(n16857), .ZN(n16862) );
  OAI211_X1 U20091 ( .C1(n16865), .C2(n16860), .A(n17007), .B(n16859), .ZN(
        n16861) );
  OAI211_X1 U20092 ( .C1(n17003), .C2(n17800), .A(n16862), .B(n16861), .ZN(
        P3_U2656) );
  AOI22_X1 U20093 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17030), .B1(
        n17014), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16874) );
  NOR2_X1 U20094 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17827), .ZN(
        n16890) );
  AOI21_X1 U20095 ( .B1(n16863), .B2(n16890), .A(n16961), .ZN(n16880) );
  OAI21_X1 U20096 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16864), .A(
        n17785), .ZN(n17816) );
  AOI211_X1 U20097 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16881), .A(n16865), .B(
        n17036), .ZN(n16867) );
  AOI211_X1 U20098 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17001), .A(
        n17816), .B(n16960), .ZN(n16866) );
  AOI211_X1 U20099 ( .C1(n16880), .C2(n17816), .A(n16867), .B(n16866), .ZN(
        n16873) );
  AND2_X1 U20100 ( .A1(n16998), .A2(n16868), .ZN(n16870) );
  AOI22_X1 U20101 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16871), .B1(n16870), 
        .B2(n16869), .ZN(n16872) );
  NAND4_X1 U20102 ( .A1(n16874), .A2(n16873), .A3(n16872), .A4(n18216), .ZN(
        P3_U2657) );
  INV_X1 U20103 ( .A(n16875), .ZN(n16898) );
  AOI21_X1 U20104 ( .B1(n16998), .B2(n16898), .A(n17035), .ZN(n16903) );
  INV_X1 U20105 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18922) );
  NAND2_X1 U20106 ( .A1(n16998), .A2(n18922), .ZN(n16897) );
  NOR3_X1 U20107 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17026), .A3(n16876), 
        .ZN(n16887) );
  NOR2_X1 U20108 ( .A1(n17848), .A2(n17827), .ZN(n16878) );
  OAI21_X1 U20109 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16878), .A(
        n16877), .ZN(n17837) );
  AOI211_X1 U20110 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17001), .A(
        n17837), .B(n16960), .ZN(n16879) );
  AOI211_X1 U20111 ( .C1(n16880), .C2(n17837), .A(n18330), .B(n16879), .ZN(
        n16884) );
  OAI211_X1 U20112 ( .C1(n16889), .C2(n16882), .A(n17007), .B(n16881), .ZN(
        n16883) );
  OAI211_X1 U20113 ( .C1(n17003), .C2(n16885), .A(n16884), .B(n16883), .ZN(
        n16886) );
  AOI211_X1 U20114 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n17014), .A(n16887), .B(
        n16886), .ZN(n16888) );
  OAI221_X1 U20115 ( .B1(n18924), .B2(n16903), .C1(n18924), .C2(n16897), .A(
        n16888), .ZN(P3_U2658) );
  AOI211_X1 U20116 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16906), .A(n16889), .B(
        n17036), .ZN(n16895) );
  NOR2_X1 U20117 ( .A1(n16890), .A2(n16975), .ZN(n16891) );
  AOI22_X1 U20118 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17827), .B1(
        n16899), .B2(n17848), .ZN(n17844) );
  XNOR2_X1 U20119 ( .A(n16891), .B(n17844), .ZN(n16892) );
  AOI22_X1 U20120 ( .A1(n17014), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n18878), 
        .B2(n16892), .ZN(n16893) );
  OAI211_X1 U20121 ( .C1(n16903), .C2(n18922), .A(n16893), .B(n18216), .ZN(
        n16894) );
  AOI211_X1 U20122 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16895), .B(n16894), .ZN(n16896) );
  OAI21_X1 U20123 ( .B1(n16898), .B2(n16897), .A(n16896), .ZN(P3_U2659) );
  INV_X1 U20124 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16923) );
  AND3_X1 U20125 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17894), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16947) );
  NAND2_X1 U20126 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16947), .ZN(
        n16937) );
  NOR2_X1 U20127 ( .A1(n16923), .A2(n16937), .ZN(n16922) );
  NAND2_X1 U20128 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16922), .ZN(
        n16913) );
  AOI21_X1 U20129 ( .B1(n16909), .B2(n16913), .A(n16899), .ZN(n17856) );
  OAI21_X1 U20130 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16913), .A(
        n17001), .ZN(n16900) );
  XNOR2_X1 U20131 ( .A(n17856), .B(n16900), .ZN(n16905) );
  NOR2_X1 U20132 ( .A1(n17026), .A2(n16911), .ZN(n16931) );
  AOI21_X1 U20133 ( .B1(n16901), .B2(n16931), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16902) );
  OAI22_X1 U20134 ( .A1(n16903), .A2(n16902), .B1(n17037), .B2(n17277), .ZN(
        n16904) );
  AOI211_X1 U20135 ( .C1(n18878), .C2(n16905), .A(n18330), .B(n16904), .ZN(
        n16908) );
  OAI211_X1 U20136 ( .C1(n16910), .C2(n17277), .A(n17007), .B(n16906), .ZN(
        n16907) );
  OAI211_X1 U20137 ( .C1(n17003), .C2(n16909), .A(n16908), .B(n16907), .ZN(
        P3_U2660) );
  INV_X1 U20138 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16921) );
  AOI211_X1 U20139 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16932), .A(n16910), .B(
        n17036), .ZN(n16919) );
  AOI21_X1 U20140 ( .B1(n16998), .B2(n16911), .A(n17035), .ZN(n16942) );
  OAI211_X1 U20141 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16931), .B(n16912), .ZN(n16917) );
  OAI21_X1 U20142 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16922), .A(
        n16913), .ZN(n16914) );
  INV_X1 U20143 ( .A(n16914), .ZN(n17878) );
  AOI21_X1 U20144 ( .B1(n16922), .B2(n17034), .A(n16975), .ZN(n16926) );
  AOI21_X1 U20145 ( .B1(n17878), .B2(n16926), .A(n17019), .ZN(n16915) );
  OAI21_X1 U20146 ( .B1(n17878), .B2(n16926), .A(n16915), .ZN(n16916) );
  OAI211_X1 U20147 ( .C1(n16942), .C2(n18918), .A(n16917), .B(n16916), .ZN(
        n16918) );
  AOI211_X1 U20148 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17014), .A(n16919), .B(
        n16918), .ZN(n16920) );
  OAI211_X1 U20149 ( .C1(n16921), .C2(n17003), .A(n16920), .B(n18216), .ZN(
        P3_U2661) );
  AOI22_X1 U20150 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17030), .B1(
        n17014), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16936) );
  INV_X1 U20151 ( .A(n16942), .ZN(n16930) );
  AOI21_X1 U20152 ( .B1(n16923), .B2(n16937), .A(n16922), .ZN(n17886) );
  INV_X1 U20153 ( .A(n17886), .ZN(n16927) );
  NAND2_X1 U20154 ( .A1(n16959), .A2(n17034), .ZN(n16949) );
  NOR3_X1 U20155 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16924), .A3(
        n16949), .ZN(n16925) );
  AOI221_X1 U20156 ( .B1(n17886), .B2(n16975), .C1(n16927), .C2(n16926), .A(
        n16925), .ZN(n16928) );
  NOR2_X1 U20157 ( .A1(n16928), .A2(n17019), .ZN(n16929) );
  AOI221_X1 U20158 ( .B1(n16931), .B2(n18916), .C1(n16930), .C2(
        P3_REIP_REG_9__SCAN_IN), .A(n16929), .ZN(n16935) );
  OAI211_X1 U20159 ( .C1(n16938), .C2(n16933), .A(n17007), .B(n16932), .ZN(
        n16934) );
  NAND4_X1 U20160 ( .A1(n16936), .A2(n16935), .A3(n18216), .A4(n16934), .ZN(
        P3_U2662) );
  OAI21_X1 U20161 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16947), .A(
        n16937), .ZN(n17908) );
  INV_X1 U20162 ( .A(n16949), .ZN(n16962) );
  AOI21_X1 U20163 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16962), .A(
        n16975), .ZN(n16951) );
  XOR2_X1 U20164 ( .A(n17908), .B(n16951), .Z(n16946) );
  AOI211_X1 U20165 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16956), .A(n16938), .B(
        n17036), .ZN(n16944) );
  AND2_X1 U20166 ( .A1(n16998), .A2(n16939), .ZN(n16955) );
  AOI21_X1 U20167 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16955), .A(
        P3_REIP_REG_8__SCAN_IN), .ZN(n16941) );
  OAI22_X1 U20168 ( .A1(n16942), .A2(n16941), .B1(n17037), .B2(n16940), .ZN(
        n16943) );
  AOI211_X1 U20169 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16944), .B(n16943), .ZN(n16945) );
  OAI211_X1 U20170 ( .C1(n17019), .C2(n16946), .A(n16945), .B(n18216), .ZN(
        P3_U2663) );
  INV_X1 U20171 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18912) );
  AOI21_X1 U20172 ( .B1(n16998), .B2(n16967), .A(n17035), .ZN(n16979) );
  OAI21_X1 U20173 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17026), .A(n16979), .ZN(
        n16954) );
  INV_X1 U20174 ( .A(n16959), .ZN(n16948) );
  AOI21_X1 U20175 ( .B1(n17912), .B2(n16948), .A(n16947), .ZN(n17917) );
  NOR2_X1 U20176 ( .A1(n17001), .A2(n17019), .ZN(n17023) );
  AOI21_X1 U20177 ( .B1(n17917), .B2(n16949), .A(n17019), .ZN(n16950) );
  OAI22_X1 U20178 ( .A1(n17917), .A2(n16951), .B1(n17023), .B2(n16950), .ZN(
        n16952) );
  OAI211_X1 U20179 ( .C1(n17037), .C2(n17344), .A(n18216), .B(n16952), .ZN(
        n16953) );
  AOI221_X1 U20180 ( .B1(n16955), .B2(n18912), .C1(n16954), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n16953), .ZN(n16958) );
  OAI211_X1 U20181 ( .C1(n16965), .C2(n17344), .A(n17007), .B(n16956), .ZN(
        n16957) );
  OAI211_X1 U20182 ( .C1(n17003), .C2(n17912), .A(n16958), .B(n16957), .ZN(
        P3_U2664) );
  AOI21_X1 U20183 ( .B1(n17929), .B2(n16974), .A(n16959), .ZN(n17932) );
  AOI21_X1 U20184 ( .B1(n17001), .B2(n16974), .A(n16960), .ZN(n16964) );
  NOR3_X1 U20185 ( .A1(n17932), .A2(n16962), .A3(n16961), .ZN(n16963) );
  AOI211_X1 U20186 ( .C1(n17932), .C2(n16964), .A(n18330), .B(n16963), .ZN(
        n16971) );
  AOI211_X1 U20187 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16982), .A(n16965), .B(
        n17036), .ZN(n16969) );
  NAND2_X1 U20188 ( .A1(n16998), .A2(n18910), .ZN(n16966) );
  OAI22_X1 U20189 ( .A1(n18910), .A2(n16979), .B1(n16967), .B2(n16966), .ZN(
        n16968) );
  AOI211_X1 U20190 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16969), .B(n16968), .ZN(n16970) );
  OAI211_X1 U20191 ( .C1(n17037), .C2(n16972), .A(n16971), .B(n16970), .ZN(
        P3_U2665) );
  AOI21_X1 U20192 ( .B1(n16998), .B2(n16973), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16980) );
  AND2_X1 U20193 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17939), .ZN(
        n16986) );
  OAI21_X1 U20194 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16986), .A(
        n16974), .ZN(n17942) );
  INV_X1 U20195 ( .A(n17942), .ZN(n16977) );
  AOI21_X1 U20196 ( .B1(n17034), .B2(n16986), .A(n16975), .ZN(n16976) );
  INV_X1 U20197 ( .A(n16976), .ZN(n16988) );
  OAI221_X1 U20198 ( .B1(n16977), .B2(n16976), .C1(n17942), .C2(n16988), .A(
        n18878), .ZN(n16978) );
  OAI211_X1 U20199 ( .C1(n16980), .C2(n16979), .A(n18216), .B(n16978), .ZN(
        n16981) );
  AOI21_X1 U20200 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17030), .A(
        n16981), .ZN(n16984) );
  OAI211_X1 U20201 ( .C1(n16989), .C2(n16985), .A(n17007), .B(n16982), .ZN(
        n16983) );
  OAI211_X1 U20202 ( .C1(n16985), .C2(n17037), .A(n16984), .B(n16983), .ZN(
        P3_U2666) );
  AOI21_X1 U20203 ( .B1(n16998), .B2(n16990), .A(n17035), .ZN(n17012) );
  AOI22_X1 U20204 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17030), .B1(
        n17014), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16997) );
  NAND2_X1 U20205 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16987), .ZN(
        n17000) );
  AOI21_X1 U20206 ( .B1(n17956), .B2(n17000), .A(n16986), .ZN(n17958) );
  NAND2_X1 U20207 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17034), .ZN(
        n17020) );
  NAND2_X1 U20208 ( .A1(n17956), .A2(n16987), .ZN(n17948) );
  OAI22_X1 U20209 ( .A1(n17958), .A2(n16988), .B1(n17020), .B2(n17948), .ZN(
        n16995) );
  AOI211_X1 U20210 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17006), .A(n16989), .B(
        n17036), .ZN(n16994) );
  NOR3_X1 U20211 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17026), .A3(n16990), .ZN(
        n16991) );
  AOI211_X1 U20212 ( .C1(n17958), .C2(n17023), .A(n18330), .B(n16991), .ZN(
        n16992) );
  OAI221_X1 U20213 ( .B1(n17042), .B2(n15691), .C1(n17042), .C2(n18863), .A(
        n16992), .ZN(n16993) );
  AOI211_X1 U20214 ( .C1(n18878), .C2(n16995), .A(n16994), .B(n16993), .ZN(
        n16996) );
  OAI211_X1 U20215 ( .C1(n17012), .C2(n18906), .A(n16997), .B(n16996), .ZN(
        P3_U2667) );
  INV_X1 U20216 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18901) );
  NOR2_X1 U20217 ( .A1(n19008), .A2(n18901), .ZN(n17027) );
  AOI21_X1 U20218 ( .B1(n16998), .B2(n17027), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n17011) );
  INV_X1 U20219 ( .A(n18824), .ZN(n16999) );
  AOI21_X1 U20220 ( .B1(n18981), .B2(n16999), .A(n15554), .ZN(n18976) );
  NOR2_X1 U20221 ( .A1(n17987), .A2(n17016), .ZN(n17015) );
  OAI21_X1 U20222 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17015), .A(
        n17000), .ZN(n17967) );
  OAI21_X1 U20223 ( .B1(n17016), .B2(n17020), .A(n17001), .ZN(n17018) );
  OAI21_X1 U20224 ( .B1(n17967), .B2(n17018), .A(n18878), .ZN(n17002) );
  AOI21_X1 U20225 ( .B1(n17967), .B2(n17018), .A(n17002), .ZN(n17005) );
  OAI22_X1 U20226 ( .A1(n17971), .A2(n17003), .B1(n17037), .B2(n17008), .ZN(
        n17004) );
  AOI211_X1 U20227 ( .C1(n17013), .C2(n18976), .A(n17005), .B(n17004), .ZN(
        n17010) );
  OAI211_X1 U20228 ( .C1(n17024), .C2(n17008), .A(n17007), .B(n17006), .ZN(
        n17009) );
  OAI211_X1 U20229 ( .C1(n17012), .C2(n17011), .A(n17010), .B(n17009), .ZN(
        P3_U2668) );
  AOI21_X1 U20230 ( .B1(n18992), .B2(n18828), .A(n18824), .ZN(n18988) );
  AOI22_X1 U20231 ( .A1(n17014), .A2(P3_EBX_REG_2__SCAN_IN), .B1(n18988), .B2(
        n17013), .ZN(n17033) );
  AOI21_X1 U20232 ( .B1(n17987), .B2(n17016), .A(n17015), .ZN(n17976) );
  NOR2_X1 U20233 ( .A1(n17017), .A2(n18901), .ZN(n17022) );
  AOI211_X1 U20234 ( .C1(n17976), .C2(n17020), .A(n17019), .B(n17018), .ZN(
        n17021) );
  AOI211_X1 U20235 ( .C1(n17023), .C2(n17976), .A(n17022), .B(n17021), .ZN(
        n17032) );
  AOI211_X1 U20236 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17025), .A(n17024), .B(
        n17036), .ZN(n17029) );
  AOI211_X1 U20237 ( .C1(n19008), .C2(n18901), .A(n17027), .B(n17026), .ZN(
        n17028) );
  AOI211_X1 U20238 ( .C1(n17030), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17029), .B(n17028), .ZN(n17031) );
  NAND3_X1 U20239 ( .A1(n17033), .A2(n17032), .A3(n17031), .ZN(P3_U2669) );
  INV_X1 U20240 ( .A(n18979), .ZN(n19002) );
  NOR3_X1 U20241 ( .A1(n19002), .A2(n17035), .A3(n17034), .ZN(n17039) );
  AOI21_X1 U20242 ( .B1(n17037), .B2(n17036), .A(n17367), .ZN(n17038) );
  AOI211_X1 U20243 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n17040), .A(n17039), .B(
        n17038), .ZN(n17041) );
  OAI21_X1 U20244 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n17042), .A(
        n17041), .ZN(P3_U2671) );
  NAND3_X1 U20245 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .ZN(n17044) );
  NAND4_X1 U20246 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17043)
         );
  NOR2_X1 U20247 ( .A1(n17044), .A2(n17043), .ZN(n17045) );
  NAND4_X1 U20248 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(n17125), .A4(n17045), .ZN(n17048) );
  NOR2_X1 U20249 ( .A1(n17049), .A2(n17048), .ZN(n17075) );
  NAND2_X1 U20250 ( .A1(n17360), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U20251 ( .A1(n17075), .A2(n17371), .ZN(n17046) );
  OAI22_X1 U20252 ( .A1(n17075), .A2(n17047), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17046), .ZN(P3_U2672) );
  NAND2_X1 U20253 ( .A1(n17049), .A2(n17048), .ZN(n17050) );
  NAND2_X1 U20254 ( .A1(n17050), .A2(n17360), .ZN(n17074) );
  AOI22_X1 U20255 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17062) );
  OAI22_X1 U20256 ( .A1(n17306), .A2(n18507), .B1(n17283), .B2(n17051), .ZN(
        n17059) );
  AOI22_X1 U20257 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20258 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20259 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17308), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17052) );
  OAI211_X1 U20260 ( .C1(n17161), .C2(n18716), .A(n17053), .B(n17052), .ZN(
        n17054) );
  AOI21_X1 U20261 ( .B1(n15554), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17054), .ZN(n17055) );
  OAI211_X1 U20262 ( .C1(n17186), .C2(n17057), .A(n17056), .B(n17055), .ZN(
        n17058) );
  AOI211_X1 U20263 ( .C1(n9813), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17061) );
  AOI22_X1 U20264 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17060) );
  NAND3_X1 U20265 ( .A1(n17062), .A2(n17061), .A3(n17060), .ZN(n17073) );
  OAI22_X1 U20266 ( .A1(n17111), .A2(n17186), .B1(n17121), .B2(n9846), .ZN(
        n17072) );
  AOI22_X1 U20267 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12915), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20268 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n17330), .ZN(n17069) );
  AOI22_X1 U20269 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17063) );
  OAI21_X1 U20270 ( .B1(n17235), .B2(n15691), .A(n17063), .ZN(n17067) );
  AOI22_X1 U20271 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17325), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20272 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17064) );
  OAI211_X1 U20273 ( .C1(n18709), .C2(n17161), .A(n17065), .B(n17064), .ZN(
        n17066) );
  AOI211_X1 U20274 ( .C1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .C2(n15686), .A(
        n17067), .B(n17066), .ZN(n17068) );
  NAND3_X1 U20275 ( .A1(n17070), .A2(n17069), .A3(n17068), .ZN(n17071) );
  AOI211_X1 U20276 ( .C1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .C2(n17331), .A(
        n17072), .B(n17071), .ZN(n17078) );
  NOR2_X1 U20277 ( .A1(n17078), .A2(n17077), .ZN(n17076) );
  XNOR2_X1 U20278 ( .A(n17073), .B(n17076), .ZN(n17379) );
  OAI22_X1 U20279 ( .A1(n17075), .A2(n17074), .B1(n17379), .B2(n17360), .ZN(
        P3_U2673) );
  AOI21_X1 U20280 ( .B1(n17078), .B2(n17077), .A(n17076), .ZN(n17380) );
  INV_X1 U20281 ( .A(n17380), .ZN(n17080) );
  NAND3_X1 U20282 ( .A1(n17081), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17360), 
        .ZN(n17079) );
  OAI221_X1 U20283 ( .B1(n17081), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17360), 
        .C2(n17080), .A(n17079), .ZN(P3_U2674) );
  INV_X1 U20284 ( .A(n17082), .ZN(n17091) );
  AOI21_X1 U20285 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17360), .A(n17091), .ZN(
        n17086) );
  AOI21_X1 U20286 ( .B1(n17084), .B2(n17088), .A(n17083), .ZN(n17389) );
  INV_X1 U20287 ( .A(n17389), .ZN(n17085) );
  OAI22_X1 U20288 ( .A1(n17087), .A2(n17086), .B1(n17360), .B2(n17085), .ZN(
        P3_U2676) );
  AOI21_X1 U20289 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17360), .A(n17097), .ZN(
        n17090) );
  OAI21_X1 U20290 ( .B1(n17093), .B2(n17089), .A(n17088), .ZN(n17396) );
  OAI22_X1 U20291 ( .A1(n17091), .A2(n17090), .B1(n17360), .B2(n17396), .ZN(
        P3_U2677) );
  INV_X1 U20292 ( .A(n17092), .ZN(n17104) );
  AOI21_X1 U20293 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17360), .A(n17104), .ZN(
        n17096) );
  AOI21_X1 U20294 ( .B1(n17094), .B2(n17100), .A(n17093), .ZN(n17397) );
  INV_X1 U20295 ( .A(n17397), .ZN(n17095) );
  OAI22_X1 U20296 ( .A1(n17097), .A2(n17096), .B1(n17360), .B2(n17095), .ZN(
        P3_U2678) );
  INV_X1 U20297 ( .A(n17105), .ZN(n17124) );
  NOR3_X1 U20298 ( .A1(n17099), .A2(n17098), .A3(n17124), .ZN(n17109) );
  AOI21_X1 U20299 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17360), .A(n17109), .ZN(
        n17103) );
  OAI21_X1 U20300 ( .B1(n17102), .B2(n17101), .A(n17100), .ZN(n17407) );
  OAI22_X1 U20301 ( .A1(n17104), .A2(n17103), .B1(n17360), .B2(n17407), .ZN(
        P3_U2679) );
  AOI22_X1 U20302 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17360), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n17105), .ZN(n17108) );
  XNOR2_X1 U20303 ( .A(n17107), .B(n17106), .ZN(n17412) );
  OAI22_X1 U20304 ( .A1(n17109), .A2(n17108), .B1(n17360), .B2(n17412), .ZN(
        P3_U2680) );
  AOI22_X1 U20305 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n15676), .B1(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n17330), .ZN(n17120) );
  AOI22_X1 U20306 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17110) );
  OAI21_X1 U20307 ( .B1(n9850), .B2(n17111), .A(n17110), .ZN(n17118) );
  AOI22_X1 U20308 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20309 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n9811), .ZN(n17113) );
  AOI22_X1 U20310 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17326), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17112) );
  OAI211_X1 U20311 ( .C1(n15691), .C2(n17230), .A(n17113), .B(n17112), .ZN(
        n17114) );
  AOI21_X1 U20312 ( .B1(n15694), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17114), .ZN(n17115) );
  OAI211_X1 U20313 ( .C1(n17287), .C2(n18379), .A(n17116), .B(n17115), .ZN(
        n17117) );
  AOI211_X1 U20314 ( .C1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .C2(n15715), .A(
        n17118), .B(n17117), .ZN(n17119) );
  OAI211_X1 U20315 ( .C1(n17186), .C2(n17121), .A(n17120), .B(n17119), .ZN(
        n17413) );
  INV_X1 U20316 ( .A(n17413), .ZN(n17123) );
  NAND3_X1 U20317 ( .A1(n17124), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17360), 
        .ZN(n17122) );
  OAI221_X1 U20318 ( .B1(n17124), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17360), 
        .C2(n17123), .A(n17122), .ZN(P3_U2681) );
  NOR2_X1 U20319 ( .A1(n17365), .A2(n17125), .ZN(n17151) );
  AOI22_X1 U20320 ( .A1(n15607), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20321 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20322 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17126) );
  OAI211_X1 U20323 ( .C1(n17306), .C2(n17128), .A(n17127), .B(n17126), .ZN(
        n17134) );
  AOI22_X1 U20324 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20325 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20326 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17130) );
  NAND2_X1 U20327 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n17129) );
  NAND4_X1 U20328 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17133) );
  AOI211_X1 U20329 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17134), .B(n17133), .ZN(n17135) );
  OAI211_X1 U20330 ( .C1(n10447), .C2(n17137), .A(n17136), .B(n17135), .ZN(
        n17420) );
  AOI22_X1 U20331 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17151), .B1(n17365), 
        .B2(n17420), .ZN(n17138) );
  OAI21_X1 U20332 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17139), .A(n17138), .ZN(
        P3_U2682) );
  AOI22_X1 U20333 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20334 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17149) );
  OAI22_X1 U20335 ( .A1(n9844), .A2(n18701), .B1(n17287), .B2(n18368), .ZN(
        n17147) );
  OAI22_X1 U20336 ( .A1(n9850), .A2(n17140), .B1(n17186), .B2(n17259), .ZN(
        n17141) );
  AOI21_X1 U20337 ( .B1(n15694), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17141), .ZN(n17145) );
  AOI22_X1 U20338 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15714), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20339 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20340 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17142) );
  NAND4_X1 U20341 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17146) );
  AOI211_X1 U20342 ( .C1(n9811), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n17147), .B(n17146), .ZN(n17148) );
  NAND3_X1 U20343 ( .A1(n17150), .A2(n17149), .A3(n17148), .ZN(n17424) );
  INV_X1 U20344 ( .A(n17424), .ZN(n17154) );
  OAI21_X1 U20345 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17152), .A(n17151), .ZN(
        n17153) );
  OAI21_X1 U20346 ( .B1(n17154), .B2(n17360), .A(n17153), .ZN(P3_U2683) );
  AOI22_X1 U20347 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20348 ( .B1(n17317), .B2(n17156), .A(n17155), .ZN(n17167) );
  AOI22_X1 U20349 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20350 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20351 ( .B1(n17158), .B2(n18613), .A(n17157), .ZN(n17163) );
  AOI22_X1 U20352 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20353 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17159) );
  OAI211_X1 U20354 ( .C1(n17161), .C2(n17273), .A(n17160), .B(n17159), .ZN(
        n17162) );
  AOI211_X1 U20355 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17163), .B(n17162), .ZN(n17164) );
  OAI211_X1 U20356 ( .C1(n17287), .C2(n18363), .A(n17165), .B(n17164), .ZN(
        n17166) );
  AOI211_X1 U20357 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17167), .B(n17166), .ZN(n17433) );
  OAI21_X1 U20358 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17183), .A(n17168), .ZN(
        n17169) );
  AOI22_X1 U20359 ( .A1(n17365), .A2(n17433), .B1(n17169), .B2(n17360), .ZN(
        P3_U2684) );
  AOI21_X1 U20360 ( .B1(n17170), .B2(n17196), .A(n17365), .ZN(n17171) );
  INV_X1 U20361 ( .A(n17171), .ZN(n17182) );
  INV_X1 U20362 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20363 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20364 ( .B1(n17317), .B2(n17286), .A(n17172), .ZN(n17181) );
  AOI22_X1 U20365 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17179) );
  INV_X1 U20366 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U20367 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20368 ( .B1(n17306), .B2(n17284), .A(n17173), .ZN(n17177) );
  AOI22_X1 U20369 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20370 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17174) );
  OAI211_X1 U20371 ( .C1(n15691), .C2(n17282), .A(n17175), .B(n17174), .ZN(
        n17176) );
  AOI211_X1 U20372 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17177), .B(n17176), .ZN(n17178) );
  OAI211_X1 U20373 ( .C1(n17287), .C2(n18358), .A(n17179), .B(n17178), .ZN(
        n17180) );
  AOI211_X1 U20374 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n17181), .B(n17180), .ZN(n17437) );
  OAI22_X1 U20375 ( .A1(n17183), .A2(n17182), .B1(n17437), .B2(n17360), .ZN(
        P3_U2685) );
  AOI22_X1 U20376 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20377 ( .B1(n17304), .B2(n17185), .A(n17184), .ZN(n17195) );
  AOI22_X1 U20378 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17193) );
  OAI22_X1 U20379 ( .A1(n17186), .A2(n17307), .B1(n17283), .B2(n17305), .ZN(
        n17191) );
  AOI22_X1 U20380 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20381 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20382 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17187) );
  NAND3_X1 U20383 ( .A1(n17189), .A2(n17188), .A3(n17187), .ZN(n17190) );
  AOI211_X1 U20384 ( .C1(n15714), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n17191), .B(n17190), .ZN(n17192) );
  OAI211_X1 U20385 ( .C1(n17287), .C2(n18354), .A(n17193), .B(n17192), .ZN(
        n17194) );
  AOI211_X1 U20386 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17195), .B(n17194), .ZN(n17443) );
  OAI21_X1 U20387 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17197), .A(n17196), .ZN(
        n17198) );
  AOI22_X1 U20388 ( .A1(n17365), .A2(n17443), .B1(n17198), .B2(n17360), .ZN(
        P3_U2686) );
  AOI22_X1 U20389 ( .A1(n15735), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17199) );
  OAI21_X1 U20390 ( .B1(n9844), .B2(n18685), .A(n17199), .ZN(n17209) );
  AOI22_X1 U20391 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17207) );
  OAI22_X1 U20392 ( .A1(n17287), .A2(n18349), .B1(n17306), .B2(n17200), .ZN(
        n17205) );
  AOI22_X1 U20393 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20394 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20395 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17201) );
  NAND3_X1 U20396 ( .A1(n17203), .A2(n17202), .A3(n17201), .ZN(n17204) );
  AOI211_X1 U20397 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17205), .B(n17204), .ZN(n17206) );
  OAI211_X1 U20398 ( .C1(n9827), .C2(n18487), .A(n17207), .B(n17206), .ZN(
        n17208) );
  AOI211_X1 U20399 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17209), .B(n17208), .ZN(n17449) );
  INV_X1 U20400 ( .A(n17225), .ZN(n17210) );
  OAI33_X1 U20401 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18384), .A3(n17225), 
        .B1(n17211), .B2(n17365), .B3(n17210), .ZN(n17212) );
  INV_X1 U20402 ( .A(n17212), .ZN(n17213) );
  OAI21_X1 U20403 ( .B1(n17449), .B2(n17360), .A(n17213), .ZN(P3_U2687) );
  AOI22_X1 U20404 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17214) );
  OAI21_X1 U20405 ( .B1(n17304), .B2(n18627), .A(n17214), .ZN(n17224) );
  AOI22_X1 U20406 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17222) );
  OAI22_X1 U20407 ( .A1(n17287), .A2(n17215), .B1(n15691), .B2(n18415), .ZN(
        n17220) );
  AOI22_X1 U20408 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20409 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20410 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15686), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17216) );
  NAND3_X1 U20411 ( .A1(n17218), .A2(n17217), .A3(n17216), .ZN(n17219) );
  AOI211_X1 U20412 ( .C1(n17280), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n17220), .B(n17219), .ZN(n17221) );
  OAI211_X1 U20413 ( .C1(n10447), .C2(n18716), .A(n17222), .B(n17221), .ZN(
        n17223) );
  AOI211_X1 U20414 ( .C1(n15714), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n17224), .B(n17223), .ZN(n17453) );
  OAI211_X1 U20415 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17226), .A(n17225), .B(
        n17360), .ZN(n17227) );
  OAI21_X1 U20416 ( .B1(n17453), .B2(n17360), .A(n17227), .ZN(P3_U2688) );
  AOI22_X1 U20417 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17229) );
  OAI21_X1 U20418 ( .B1(n17230), .B2(n17283), .A(n17229), .ZN(n17241) );
  INV_X1 U20419 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18622) );
  AOI22_X1 U20420 ( .A1(n15607), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n17326), .ZN(n17239) );
  INV_X1 U20421 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18410) );
  AOI22_X1 U20422 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17231), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17232) );
  OAI21_X1 U20423 ( .B1(n15691), .B2(n18410), .A(n17232), .ZN(n17237) );
  AOI22_X1 U20424 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20425 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n9811), .ZN(n17233) );
  OAI211_X1 U20426 ( .C1(n17235), .C2(n17306), .A(n17234), .B(n17233), .ZN(
        n17236) );
  AOI211_X1 U20427 ( .C1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .C2(n15694), .A(
        n17237), .B(n17236), .ZN(n17238) );
  OAI211_X1 U20428 ( .C1(n18622), .C2(n17304), .A(n17239), .B(n17238), .ZN(
        n17240) );
  AOI211_X1 U20429 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n17241), .B(n17240), .ZN(n17461) );
  INV_X1 U20430 ( .A(n17461), .ZN(n17245) );
  NOR2_X1 U20431 ( .A1(n17243), .A2(n17242), .ZN(n17244) );
  AOI22_X1 U20432 ( .A1(n17365), .A2(n17245), .B1(n17244), .B2(n17248), .ZN(
        n17246) );
  OAI21_X1 U20433 ( .B1(n17248), .B2(n17247), .A(n17246), .ZN(P3_U2689) );
  AOI22_X1 U20434 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17249) );
  OAI21_X1 U20435 ( .B1(n9844), .B2(n17250), .A(n17249), .ZN(n17261) );
  AOI22_X1 U20436 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17258) );
  INV_X1 U20437 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20438 ( .A1(n15607), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20439 ( .B1(n17306), .B2(n17252), .A(n17251), .ZN(n17256) );
  AOI22_X1 U20440 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20441 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17280), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17253) );
  OAI211_X1 U20442 ( .C1(n15691), .C2(n18404), .A(n17254), .B(n17253), .ZN(
        n17255) );
  AOI211_X1 U20443 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17256), .B(n17255), .ZN(n17257) );
  OAI211_X1 U20444 ( .C1(n9850), .C2(n17259), .A(n17258), .B(n17257), .ZN(
        n17260) );
  AOI211_X1 U20445 ( .C1(n15714), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17261), .B(n17260), .ZN(n17467) );
  OAI21_X1 U20446 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17276), .A(n17360), .ZN(
        n17262) );
  OAI22_X1 U20447 ( .A1(n17467), .A2(n17360), .B1(n17263), .B2(n17262), .ZN(
        P3_U2691) );
  AOI22_X1 U20448 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U20449 ( .B1(n10447), .B2(n18696), .A(n17264), .ZN(n17275) );
  AOI22_X1 U20450 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17272) );
  INV_X1 U20451 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18401) );
  AOI22_X1 U20452 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17265) );
  OAI21_X1 U20453 ( .B1(n15691), .B2(n18401), .A(n17265), .ZN(n17270) );
  AOI22_X1 U20454 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20455 ( .A1(n15676), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17266) );
  OAI211_X1 U20456 ( .C1(n17306), .C2(n17268), .A(n17267), .B(n17266), .ZN(
        n17269) );
  AOI211_X1 U20457 ( .C1(n15694), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17270), .B(n17269), .ZN(n17271) );
  OAI211_X1 U20458 ( .C1(n9844), .C2(n17273), .A(n17272), .B(n17271), .ZN(
        n17274) );
  AOI211_X1 U20459 ( .C1(n15714), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n17275), .B(n17274), .ZN(n17471) );
  OR2_X1 U20460 ( .A1(n17299), .A2(n17320), .ZN(n17301) );
  AOI21_X1 U20461 ( .B1(n17277), .B2(n17301), .A(n17276), .ZN(n17278) );
  INV_X1 U20462 ( .A(n17278), .ZN(n17279) );
  AOI22_X1 U20463 ( .A1(n17365), .A2(n17471), .B1(n17279), .B2(n17360), .ZN(
        P3_U2692) );
  AOI22_X1 U20464 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17280), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20465 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17297) );
  OAI22_X1 U20466 ( .A1(n9827), .A2(n17284), .B1(n17283), .B2(n17282), .ZN(
        n17295) );
  OAI22_X1 U20467 ( .A1(n17287), .A2(n17286), .B1(n17306), .B2(n17285), .ZN(
        n17288) );
  AOI21_X1 U20468 ( .B1(n17331), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n17288), .ZN(n17293) );
  AOI22_X1 U20469 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15654), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20470 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20471 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17290) );
  NAND4_X1 U20472 ( .A1(n17293), .A2(n17292), .A3(n17291), .A4(n17290), .ZN(
        n17294) );
  AOI211_X1 U20473 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n17295), .B(n17294), .ZN(n17296) );
  NAND3_X1 U20474 ( .A1(n17298), .A2(n17297), .A3(n17296), .ZN(n17476) );
  AOI21_X1 U20475 ( .B1(n17299), .B2(n17320), .A(n17365), .ZN(n17300) );
  AOI22_X1 U20476 ( .A1(n17476), .A2(n17365), .B1(n17301), .B2(n17300), .ZN(
        n17302) );
  INV_X1 U20477 ( .A(n17302), .ZN(P3_U2693) );
  AOI22_X1 U20478 ( .A1(n15714), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17303) );
  OAI21_X1 U20479 ( .B1(n17304), .B2(n18608), .A(n17303), .ZN(n17319) );
  AOI22_X1 U20480 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17315) );
  OAI22_X1 U20481 ( .A1(n9850), .A2(n17307), .B1(n17306), .B2(n17305), .ZN(
        n17313) );
  AOI22_X1 U20482 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U20483 ( .A1(n17308), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20484 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17309) );
  NAND3_X1 U20485 ( .A1(n17311), .A2(n17310), .A3(n17309), .ZN(n17312) );
  AOI211_X1 U20486 ( .C1(n9813), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n17313), .B(n17312), .ZN(n17314) );
  OAI211_X1 U20487 ( .C1(n17317), .C2(n17316), .A(n17315), .B(n17314), .ZN(
        n17318) );
  AOI211_X1 U20488 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n17319), .B(n17318), .ZN(n17480) );
  OAI21_X1 U20489 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17321), .A(n17320), .ZN(
        n17322) );
  AOI22_X1 U20490 ( .A1(n17365), .A2(n17480), .B1(n17322), .B2(n17360), .ZN(
        P3_U2694) );
  NAND2_X1 U20491 ( .A1(n17323), .A2(n17352), .ZN(n17342) );
  AOI21_X1 U20492 ( .B1(n17349), .B2(n17323), .A(n17365), .ZN(n17343) );
  AOI22_X1 U20493 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17340) );
  AOI22_X1 U20494 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20495 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17328) );
  OAI211_X1 U20496 ( .C1(n15691), .C2(n18392), .A(n17329), .B(n17328), .ZN(
        n17338) );
  AOI22_X1 U20497 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20498 ( .A1(n12915), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17335) );
  AOI22_X1 U20499 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17334) );
  NAND2_X1 U20500 ( .A1(n15694), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n17333) );
  NAND4_X1 U20501 ( .A1(n17336), .A2(n17335), .A3(n17334), .A4(n17333), .ZN(
        n17337) );
  AOI211_X1 U20502 ( .C1(n15686), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17338), .B(n17337), .ZN(n17339) );
  OAI211_X1 U20503 ( .C1(n15688), .C2(n18487), .A(n17340), .B(n17339), .ZN(
        n17488) );
  AOI22_X1 U20504 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17343), .B1(n17365), .B2(
        n17488), .ZN(n17341) );
  OAI21_X1 U20505 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17342), .A(n17341), .ZN(
        P3_U2695) );
  AOI22_X1 U20506 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17365), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17343), .ZN(n17346) );
  NAND4_X1 U20507 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17352), .A4(n17344), .ZN(n17345) );
  NAND2_X1 U20508 ( .A1(n17346), .A2(n17345), .ZN(P3_U2696) );
  NAND2_X1 U20509 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17352), .ZN(n17348) );
  NAND3_X1 U20510 ( .A1(n17348), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17360), .ZN(
        n17347) );
  OAI221_X1 U20511 ( .B1(n17348), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17360), 
        .C2(n18379), .A(n17347), .ZN(P3_U2697) );
  OAI211_X1 U20512 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17349), .A(n17348), .B(
        n17360), .ZN(n17350) );
  OAI21_X1 U20513 ( .B1(n17360), .B2(n18374), .A(n17350), .ZN(P3_U2698) );
  NAND2_X1 U20514 ( .A1(n17371), .A2(n17368), .ZN(n17363) );
  INV_X1 U20515 ( .A(n17363), .ZN(n17364) );
  AOI22_X1 U20516 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17360), .B1(n17353), .B2(
        n17364), .ZN(n17351) );
  OAI22_X1 U20517 ( .A1(n17352), .A2(n17351), .B1(n18368), .B2(n17360), .ZN(
        P3_U2699) );
  AND2_X1 U20518 ( .A1(n17353), .A2(n17364), .ZN(n17356) );
  NOR2_X1 U20519 ( .A1(n17354), .A2(n17363), .ZN(n17358) );
  AOI21_X1 U20520 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17360), .A(n17358), .ZN(
        n17355) );
  OAI22_X1 U20521 ( .A1(n17356), .A2(n17355), .B1(n18363), .B2(n17360), .ZN(
        P3_U2700) );
  AOI21_X1 U20522 ( .B1(n17368), .B2(n17357), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17359) );
  AOI221_X1 U20523 ( .B1(n17359), .B2(n17360), .C1(n18358), .C2(n17365), .A(
        n17358), .ZN(P3_U2701) );
  OAI222_X1 U20524 ( .A1(n17363), .A2(n17362), .B1(n17361), .B2(n17368), .C1(
        n18354), .C2(n17360), .ZN(P3_U2702) );
  AOI22_X1 U20525 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17365), .B1(
        n17364), .B2(n17367), .ZN(n17366) );
  OAI21_X1 U20526 ( .B1(n17368), .B2(n17367), .A(n17366), .ZN(P3_U2703) );
  INV_X1 U20527 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17586) );
  INV_X1 U20528 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17583) );
  INV_X1 U20529 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17576) );
  INV_X1 U20530 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17566) );
  INV_X1 U20531 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17627) );
  INV_X1 U20532 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17602) );
  NAND3_X1 U20533 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17492) );
  NAND4_X1 U20534 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_7__SCAN_IN), .A4(P3_EAX_REG_6__SCAN_IN), .ZN(n17369) );
  NOR3_X1 U20535 ( .A1(n17602), .A2(n17492), .A3(n17369), .ZN(n17454) );
  NAND2_X1 U20536 ( .A1(n17513), .A2(n17454), .ZN(n17486) );
  NAND3_X1 U20537 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .ZN(n17456) );
  NAND2_X1 U20538 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17457) );
  NOR3_X1 U20539 ( .A1(n17486), .A2(n17456), .A3(n17457), .ZN(n17370) );
  NAND3_X1 U20540 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(n17370), .ZN(n17458) );
  NAND4_X1 U20541 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n17419)
         );
  NAND2_X1 U20542 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17404), .ZN(n17403) );
  NAND2_X1 U20543 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17384), .ZN(n17381) );
  NAND2_X1 U20544 ( .A1(n17376), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17375) );
  NAND2_X1 U20545 ( .A1(n18376), .A2(n17485), .ZN(n17402) );
  OAI22_X1 U20546 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17491), .B1(n17485), 
        .B2(n17376), .ZN(n17373) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17444), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17373), .ZN(n17374) );
  OAI21_X1 U20548 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17375), .A(n17374), .ZN(
        P3_U2704) );
  NOR2_X2 U20549 ( .A1(n18371), .A2(n17520), .ZN(n17445) );
  AOI22_X1 U20550 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17444), .ZN(n17378) );
  OAI211_X1 U20551 ( .C1(n17376), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17520), .B(
        n17375), .ZN(n17377) );
  OAI211_X1 U20552 ( .C1(n17379), .C2(n17506), .A(n17378), .B(n17377), .ZN(
        P3_U2705) );
  INV_X1 U20553 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U20554 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17445), .B1(n17517), .B2(
        n17380), .ZN(n17383) );
  OAI211_X1 U20555 ( .C1(n17384), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17520), .B(
        n17381), .ZN(n17382) );
  OAI211_X1 U20556 ( .C1(n17402), .C2(n18369), .A(n17383), .B(n17382), .ZN(
        P3_U2706) );
  AOI22_X1 U20557 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17444), .ZN(n17387) );
  AOI211_X1 U20558 ( .C1(n17586), .C2(n17390), .A(n17384), .B(n17485), .ZN(
        n17385) );
  INV_X1 U20559 ( .A(n17385), .ZN(n17386) );
  OAI211_X1 U20560 ( .C1(n17388), .C2(n17506), .A(n17387), .B(n17386), .ZN(
        P3_U2707) );
  INV_X1 U20561 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U20562 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17445), .B1(n17517), .B2(
        n17389), .ZN(n17392) );
  OAI211_X1 U20563 ( .C1(n9857), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17520), .B(
        n17390), .ZN(n17391) );
  OAI211_X1 U20564 ( .C1(n17402), .C2(n18359), .A(n17392), .B(n17391), .ZN(
        P3_U2708) );
  AOI22_X1 U20565 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17444), .ZN(n17395) );
  AOI211_X1 U20566 ( .C1(n17583), .C2(n17398), .A(n9857), .B(n17485), .ZN(
        n17393) );
  INV_X1 U20567 ( .A(n17393), .ZN(n17394) );
  OAI211_X1 U20568 ( .C1(n17396), .C2(n17506), .A(n17395), .B(n17394), .ZN(
        P3_U2709) );
  INV_X1 U20569 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U20570 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17445), .B1(n17517), .B2(
        n17397), .ZN(n17401) );
  OAI211_X1 U20571 ( .C1(n17399), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17520), .B(
        n17398), .ZN(n17400) );
  OAI211_X1 U20572 ( .C1(n17402), .C2(n18351), .A(n17401), .B(n17400), .ZN(
        P3_U2710) );
  AOI22_X1 U20573 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17444), .ZN(n17406) );
  OAI211_X1 U20574 ( .C1(n17404), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17520), .B(
        n17403), .ZN(n17405) );
  OAI211_X1 U20575 ( .C1(n17407), .C2(n17506), .A(n17406), .B(n17405), .ZN(
        P3_U2711) );
  AOI22_X1 U20576 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17444), .ZN(n17411) );
  OAI211_X1 U20577 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17409), .A(n17520), .B(
        n17408), .ZN(n17410) );
  OAI211_X1 U20578 ( .C1(n17412), .C2(n17506), .A(n17411), .B(n17410), .ZN(
        P3_U2712) );
  NAND2_X1 U20579 ( .A1(n17438), .A2(n17576), .ZN(n17418) );
  AOI22_X1 U20580 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17444), .B1(n17517), .B2(
        n17413), .ZN(n17417) );
  INV_X1 U20581 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17572) );
  INV_X1 U20582 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17570) );
  NAND2_X1 U20583 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17438), .ZN(n17434) );
  NOR3_X1 U20584 ( .A1(n17572), .A2(n17570), .A3(n17434), .ZN(n17428) );
  NOR2_X1 U20585 ( .A1(n17485), .A2(n17428), .ZN(n17425) );
  INV_X1 U20586 ( .A(n17425), .ZN(n17414) );
  OAI21_X1 U20587 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17491), .A(n17414), .ZN(
        n17415) );
  AOI22_X1 U20588 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17445), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17415), .ZN(n17416) );
  OAI211_X1 U20589 ( .C1(n17419), .C2(n17418), .A(n17417), .B(n17416), .ZN(
        P3_U2713) );
  INV_X1 U20590 ( .A(n17428), .ZN(n17423) );
  AOI22_X1 U20591 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17444), .B1(n17517), .B2(
        n17420), .ZN(n17422) );
  AOI22_X1 U20592 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17445), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17425), .ZN(n17421) );
  OAI211_X1 U20593 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17423), .A(n17422), .B(
        n17421), .ZN(P3_U2714) );
  INV_X1 U20594 ( .A(n17434), .ZN(n17430) );
  NAND2_X1 U20595 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17430), .ZN(n17429) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17444), .B1(n17517), .B2(
        n17424), .ZN(n17427) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17445), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n17425), .ZN(n17426) );
  OAI211_X1 U20598 ( .C1(n17428), .C2(n17429), .A(n17427), .B(n17426), .ZN(
        P3_U2715) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17444), .ZN(n17432) );
  OAI211_X1 U20600 ( .C1(n17430), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17520), .B(
        n17429), .ZN(n17431) );
  OAI211_X1 U20601 ( .C1(n17433), .C2(n17506), .A(n17432), .B(n17431), .ZN(
        P3_U2716) );
  AOI22_X1 U20602 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17444), .ZN(n17436) );
  OAI211_X1 U20603 ( .C1(n17438), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17520), .B(
        n17434), .ZN(n17435) );
  OAI211_X1 U20604 ( .C1(n17437), .C2(n17506), .A(n17436), .B(n17435), .ZN(
        P3_U2717) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17444), .ZN(n17442) );
  INV_X1 U20606 ( .A(n17446), .ZN(n17440) );
  INV_X1 U20607 ( .A(n17438), .ZN(n17439) );
  OAI211_X1 U20608 ( .C1(n17440), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17520), .B(
        n17439), .ZN(n17441) );
  OAI211_X1 U20609 ( .C1(n17443), .C2(n17506), .A(n17442), .B(n17441), .ZN(
        P3_U2718) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17445), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17444), .ZN(n17448) );
  OAI211_X1 U20611 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17450), .A(n17520), .B(
        n17446), .ZN(n17447) );
  OAI211_X1 U20612 ( .C1(n17449), .C2(n17506), .A(n17448), .B(n17447), .ZN(
        P3_U2719) );
  AOI211_X1 U20613 ( .C1(n17627), .C2(n17458), .A(n17485), .B(n17450), .ZN(
        n17451) );
  AOI21_X1 U20614 ( .B1(n17518), .B2(BUF2_REG_15__SCAN_IN), .A(n17451), .ZN(
        n17452) );
  OAI21_X1 U20615 ( .B1(n17453), .B2(n17506), .A(n17452), .ZN(P3_U2720) );
  INV_X1 U20616 ( .A(n17454), .ZN(n17455) );
  NOR2_X1 U20617 ( .A1(n17455), .A2(n17491), .ZN(n17496) );
  INV_X1 U20618 ( .A(n17496), .ZN(n17475) );
  NAND2_X1 U20619 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17479), .ZN(n17466) );
  NOR2_X1 U20620 ( .A1(n17457), .A2(n17466), .ZN(n17463) );
  INV_X1 U20621 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U20622 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17518), .B1(n17463), .B2(
        n17622), .ZN(n17460) );
  NAND3_X1 U20623 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17520), .A3(n17458), 
        .ZN(n17459) );
  OAI211_X1 U20624 ( .C1(n17461), .C2(n17506), .A(n17460), .B(n17459), .ZN(
        P3_U2721) );
  INV_X1 U20625 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17465) );
  INV_X1 U20626 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17618) );
  NOR2_X1 U20627 ( .A1(n17618), .A2(n17466), .ZN(n17469) );
  AOI21_X1 U20628 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17520), .A(n17469), .ZN(
        n17464) );
  OAI222_X1 U20629 ( .A1(n17509), .A2(n17465), .B1(n17464), .B2(n17463), .C1(
        n17506), .C2(n17462), .ZN(P3_U2722) );
  INV_X1 U20630 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17470) );
  INV_X1 U20631 ( .A(n17466), .ZN(n17473) );
  AOI21_X1 U20632 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17520), .A(n17473), .ZN(
        n17468) );
  OAI222_X1 U20633 ( .A1(n17509), .A2(n17470), .B1(n17469), .B2(n17468), .C1(
        n17506), .C2(n17467), .ZN(P3_U2723) );
  INV_X1 U20634 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17474) );
  AOI21_X1 U20635 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17520), .A(n17479), .ZN(
        n17472) );
  OAI222_X1 U20636 ( .A1(n17509), .A2(n17474), .B1(n17473), .B2(n17472), .C1(
        n17506), .C2(n17471), .ZN(P3_U2724) );
  INV_X1 U20637 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17608) );
  NOR2_X1 U20638 ( .A1(n17608), .A2(n17475), .ZN(n17484) );
  AND2_X1 U20639 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17484), .ZN(n17482) );
  OAI21_X1 U20640 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17482), .A(n17520), .ZN(
        n17478) );
  AOI22_X1 U20641 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17518), .B1(n17517), .B2(
        n17476), .ZN(n17477) );
  OAI21_X1 U20642 ( .B1(n17479), .B2(n17478), .A(n17477), .ZN(P3_U2725) );
  INV_X1 U20643 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17483) );
  AOI21_X1 U20644 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17520), .A(n17484), .ZN(
        n17481) );
  OAI222_X1 U20645 ( .A1(n17509), .A2(n17483), .B1(n17482), .B2(n17481), .C1(
        n17506), .C2(n17480), .ZN(P3_U2726) );
  AOI211_X1 U20646 ( .C1(n17486), .C2(n17608), .A(n17485), .B(n17484), .ZN(
        n17487) );
  AOI21_X1 U20647 ( .B1(n17517), .B2(n17488), .A(n17487), .ZN(n17489) );
  OAI21_X1 U20648 ( .B1(n17490), .B2(n17509), .A(n17489), .ZN(P3_U2727) );
  INV_X1 U20649 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18381) );
  INV_X1 U20650 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17604) );
  NAND2_X1 U20651 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n17493) );
  NOR2_X1 U20652 ( .A1(n17492), .A2(n17491), .ZN(n17504) );
  INV_X1 U20653 ( .A(n17504), .ZN(n17512) );
  NOR2_X1 U20654 ( .A1(n17493), .A2(n17512), .ZN(n17508) );
  NAND2_X1 U20655 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17508), .ZN(n17497) );
  NOR2_X1 U20656 ( .A1(n17604), .A2(n17497), .ZN(n17499) );
  AOI21_X1 U20657 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17520), .A(n17499), .ZN(
        n17495) );
  OAI222_X1 U20658 ( .A1(n17509), .A2(n18381), .B1(n17496), .B2(n17495), .C1(
        n17506), .C2(n17494), .ZN(P3_U2728) );
  INV_X1 U20659 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18375) );
  INV_X1 U20660 ( .A(n17497), .ZN(n17502) );
  AOI21_X1 U20661 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17520), .A(n17502), .ZN(
        n17500) );
  OAI222_X1 U20662 ( .A1(n17509), .A2(n18375), .B1(n17500), .B2(n17499), .C1(
        n17506), .C2(n17498), .ZN(P3_U2729) );
  INV_X1 U20663 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18370) );
  AOI21_X1 U20664 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17520), .A(n17508), .ZN(
        n17503) );
  OAI222_X1 U20665 ( .A1(n17509), .A2(n18370), .B1(n17503), .B2(n17502), .C1(
        n17506), .C2(n17501), .ZN(P3_U2730) );
  INV_X1 U20666 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18364) );
  AOI22_X1 U20667 ( .A1(n17504), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17520), .ZN(n17507) );
  OAI222_X1 U20668 ( .A1(n18364), .A2(n17509), .B1(n17508), .B2(n17507), .C1(
        n17506), .C2(n17505), .ZN(P3_U2731) );
  INV_X1 U20669 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17598) );
  NAND2_X1 U20670 ( .A1(n17520), .A2(n17512), .ZN(n17516) );
  AOI22_X1 U20671 ( .A1(n17518), .A2(BUF2_REG_3__SCAN_IN), .B1(n17517), .B2(
        n17510), .ZN(n17511) );
  OAI221_X1 U20672 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17512), .C1(n17598), 
        .C2(n17516), .A(n17511), .ZN(P3_U2732) );
  INV_X1 U20673 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17596) );
  NAND3_X1 U20674 ( .A1(n17513), .A2(P3_EAX_REG_1__SCAN_IN), .A3(
        P3_EAX_REG_0__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20675 ( .A1(n17518), .A2(BUF2_REG_2__SCAN_IN), .B1(n17517), .B2(
        n17514), .ZN(n17515) );
  OAI221_X1 U20676 ( .B1(n17516), .B2(n17596), .C1(n17516), .C2(n17519), .A(
        n17515), .ZN(P3_U2733) );
  AOI22_X1 U20677 ( .A1(n17518), .A2(BUF2_REG_1__SCAN_IN), .B1(n17517), .B2(
        n10112), .ZN(n17523) );
  OAI211_X1 U20678 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17521), .A(n17520), .B(
        n17519), .ZN(n17522) );
  NAND2_X1 U20679 ( .A1(n17523), .A2(n17522), .ZN(P3_U2734) );
  NOR2_X2 U20680 ( .A1(n18985), .A2(n17748), .ZN(n19022) );
  NOR2_X4 U20681 ( .A1(n19022), .A2(n17542), .ZN(n17539) );
  AND2_X1 U20682 ( .A1(n17539), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20683 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17590) );
  AOI22_X1 U20684 ( .A1(n19022), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17539), .ZN(n17525) );
  OAI21_X1 U20685 ( .B1(n17590), .B2(n17541), .A(n17525), .ZN(P3_U2737) );
  INV_X1 U20686 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20687 ( .A1(n19022), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U20688 ( .B1(n17588), .B2(n17541), .A(n17526), .ZN(P3_U2738) );
  AOI22_X1 U20689 ( .A1(n19022), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U20690 ( .B1(n17586), .B2(n17541), .A(n17527), .ZN(P3_U2739) );
  AOI22_X1 U20691 ( .A1(n19022), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20692 ( .B1(n10099), .B2(n17541), .A(n17528), .ZN(P3_U2740) );
  AOI22_X1 U20693 ( .A1(n19022), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17529) );
  OAI21_X1 U20694 ( .B1(n17583), .B2(n17541), .A(n17529), .ZN(P3_U2741) );
  AOI22_X1 U20695 ( .A1(n19022), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17530) );
  OAI21_X1 U20696 ( .B1(n10098), .B2(n17541), .A(n17530), .ZN(P3_U2742) );
  INV_X1 U20697 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17580) );
  AOI22_X1 U20698 ( .A1(n19022), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20699 ( .B1(n17580), .B2(n17541), .A(n17531), .ZN(P3_U2743) );
  INV_X1 U20700 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17578) );
  AOI22_X1 U20701 ( .A1(n19022), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17532) );
  OAI21_X1 U20702 ( .B1(n17578), .B2(n17541), .A(n17532), .ZN(P3_U2744) );
  CLKBUF_X1 U20703 ( .A(n19022), .Z(n18865) );
  AOI22_X1 U20704 ( .A1(n18865), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20705 ( .B1(n17576), .B2(n17541), .A(n17533), .ZN(P3_U2745) );
  INV_X1 U20706 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U20707 ( .A1(n18865), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17534) );
  OAI21_X1 U20708 ( .B1(n17574), .B2(n17541), .A(n17534), .ZN(P3_U2746) );
  AOI22_X1 U20709 ( .A1(n18865), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20710 ( .B1(n17572), .B2(n17541), .A(n17535), .ZN(P3_U2747) );
  AOI22_X1 U20711 ( .A1(n18865), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U20712 ( .B1(n17570), .B2(n17541), .A(n17536), .ZN(P3_U2748) );
  INV_X1 U20713 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U20714 ( .A1(n18865), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U20715 ( .B1(n17568), .B2(n17541), .A(n17537), .ZN(P3_U2749) );
  AOI22_X1 U20716 ( .A1(n18865), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17538) );
  OAI21_X1 U20717 ( .B1(n17566), .B2(n17541), .A(n17538), .ZN(P3_U2750) );
  INV_X1 U20718 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17564) );
  AOI22_X1 U20719 ( .A1(n18865), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17540) );
  OAI21_X1 U20720 ( .B1(n17564), .B2(n17541), .A(n17540), .ZN(P3_U2751) );
  AOI22_X1 U20721 ( .A1(n18865), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17543) );
  OAI21_X1 U20722 ( .B1(n17627), .B2(n17559), .A(n17543), .ZN(P3_U2752) );
  AOI22_X1 U20723 ( .A1(n18865), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17544) );
  OAI21_X1 U20724 ( .B1(n17622), .B2(n17559), .A(n17544), .ZN(P3_U2753) );
  INV_X1 U20725 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U20726 ( .A1(n18865), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17545) );
  OAI21_X1 U20727 ( .B1(n17620), .B2(n17559), .A(n17545), .ZN(P3_U2754) );
  AOI22_X1 U20728 ( .A1(n18865), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17546) );
  OAI21_X1 U20729 ( .B1(n17618), .B2(n17559), .A(n17546), .ZN(P3_U2755) );
  INV_X1 U20730 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U20731 ( .A1(n18865), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17547) );
  OAI21_X1 U20732 ( .B1(n17614), .B2(n17559), .A(n17547), .ZN(P3_U2756) );
  INV_X1 U20733 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U20734 ( .A1(n18865), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17548) );
  OAI21_X1 U20735 ( .B1(n17612), .B2(n17559), .A(n17548), .ZN(P3_U2757) );
  INV_X1 U20736 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17610) );
  AOI22_X1 U20737 ( .A1(n18865), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17549) );
  OAI21_X1 U20738 ( .B1(n17610), .B2(n17559), .A(n17549), .ZN(P3_U2758) );
  AOI22_X1 U20739 ( .A1(n18865), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17550) );
  OAI21_X1 U20740 ( .B1(n17608), .B2(n17559), .A(n17550), .ZN(P3_U2759) );
  INV_X1 U20741 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U20742 ( .A1(n18865), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17551) );
  OAI21_X1 U20743 ( .B1(n17606), .B2(n17559), .A(n17551), .ZN(P3_U2760) );
  AOI22_X1 U20744 ( .A1(n18865), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17552) );
  OAI21_X1 U20745 ( .B1(n17604), .B2(n17559), .A(n17552), .ZN(P3_U2761) );
  AOI22_X1 U20746 ( .A1(n18865), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17553) );
  OAI21_X1 U20747 ( .B1(n17602), .B2(n17559), .A(n17553), .ZN(P3_U2762) );
  INV_X1 U20748 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17600) );
  AOI22_X1 U20749 ( .A1(n18865), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17554) );
  OAI21_X1 U20750 ( .B1(n17600), .B2(n17559), .A(n17554), .ZN(P3_U2763) );
  AOI22_X1 U20751 ( .A1(n18865), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17555) );
  OAI21_X1 U20752 ( .B1(n17598), .B2(n17559), .A(n17555), .ZN(P3_U2764) );
  AOI22_X1 U20753 ( .A1(n18865), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17556) );
  OAI21_X1 U20754 ( .B1(n17596), .B2(n17559), .A(n17556), .ZN(P3_U2765) );
  INV_X1 U20755 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U20756 ( .A1(n18865), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17557) );
  OAI21_X1 U20757 ( .B1(n17594), .B2(n17559), .A(n17557), .ZN(P3_U2766) );
  AOI22_X1 U20758 ( .A1(n18865), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17539), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17558) );
  OAI21_X1 U20759 ( .B1(n17592), .B2(n17559), .A(n17558), .ZN(P3_U2767) );
  NAND2_X2 U20760 ( .A1(n19025), .A2(n17562), .ZN(n17626) );
  AOI22_X1 U20761 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17615), .ZN(n17563) );
  OAI21_X1 U20762 ( .B1(n17564), .B2(n17626), .A(n17563), .ZN(P3_U2768) );
  AOI22_X1 U20763 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17615), .ZN(n17565) );
  OAI21_X1 U20764 ( .B1(n17566), .B2(n17626), .A(n17565), .ZN(P3_U2769) );
  AOI22_X1 U20765 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17615), .ZN(n17567) );
  OAI21_X1 U20766 ( .B1(n17568), .B2(n17626), .A(n17567), .ZN(P3_U2770) );
  AOI22_X1 U20767 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17615), .ZN(n17569) );
  OAI21_X1 U20768 ( .B1(n17570), .B2(n17626), .A(n17569), .ZN(P3_U2771) );
  AOI22_X1 U20769 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17615), .ZN(n17571) );
  OAI21_X1 U20770 ( .B1(n17572), .B2(n17626), .A(n17571), .ZN(P3_U2772) );
  AOI22_X1 U20771 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17615), .ZN(n17573) );
  OAI21_X1 U20772 ( .B1(n17574), .B2(n17626), .A(n17573), .ZN(P3_U2773) );
  AOI22_X1 U20773 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17615), .ZN(n17575) );
  OAI21_X1 U20774 ( .B1(n17576), .B2(n17626), .A(n17575), .ZN(P3_U2774) );
  AOI22_X1 U20775 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17615), .ZN(n17577) );
  OAI21_X1 U20776 ( .B1(n17578), .B2(n17626), .A(n17577), .ZN(P3_U2775) );
  AOI22_X1 U20777 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17615), .ZN(n17579) );
  OAI21_X1 U20778 ( .B1(n17580), .B2(n17626), .A(n17579), .ZN(P3_U2776) );
  AOI22_X1 U20779 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17615), .ZN(n17581) );
  OAI21_X1 U20780 ( .B1(n10098), .B2(n17626), .A(n17581), .ZN(P3_U2777) );
  AOI22_X1 U20781 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17615), .ZN(n17582) );
  OAI21_X1 U20782 ( .B1(n17583), .B2(n17626), .A(n17582), .ZN(P3_U2778) );
  AOI22_X1 U20783 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17616), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17615), .ZN(n17584) );
  OAI21_X1 U20784 ( .B1(n10099), .B2(n17626), .A(n17584), .ZN(P3_U2779) );
  AOI22_X1 U20785 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17615), .ZN(n17585) );
  OAI21_X1 U20786 ( .B1(n17586), .B2(n17626), .A(n17585), .ZN(P3_U2780) );
  AOI22_X1 U20787 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17615), .ZN(n17587) );
  OAI21_X1 U20788 ( .B1(n17588), .B2(n17626), .A(n17587), .ZN(P3_U2781) );
  AOI22_X1 U20789 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17615), .ZN(n17589) );
  OAI21_X1 U20790 ( .B1(n17590), .B2(n17626), .A(n17589), .ZN(P3_U2782) );
  AOI22_X1 U20791 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17615), .ZN(n17591) );
  OAI21_X1 U20792 ( .B1(n17592), .B2(n17626), .A(n17591), .ZN(P3_U2783) );
  AOI22_X1 U20793 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17615), .ZN(n17593) );
  OAI21_X1 U20794 ( .B1(n17594), .B2(n17626), .A(n17593), .ZN(P3_U2784) );
  AOI22_X1 U20795 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17615), .ZN(n17595) );
  OAI21_X1 U20796 ( .B1(n17596), .B2(n17626), .A(n17595), .ZN(P3_U2785) );
  AOI22_X1 U20797 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17615), .ZN(n17597) );
  OAI21_X1 U20798 ( .B1(n17598), .B2(n17626), .A(n17597), .ZN(P3_U2786) );
  AOI22_X1 U20799 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17623), .ZN(n17599) );
  OAI21_X1 U20800 ( .B1(n17600), .B2(n17626), .A(n17599), .ZN(P3_U2787) );
  AOI22_X1 U20801 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17623), .ZN(n17601) );
  OAI21_X1 U20802 ( .B1(n17602), .B2(n17626), .A(n17601), .ZN(P3_U2788) );
  AOI22_X1 U20803 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17623), .ZN(n17603) );
  OAI21_X1 U20804 ( .B1(n17604), .B2(n17626), .A(n17603), .ZN(P3_U2789) );
  AOI22_X1 U20805 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17623), .ZN(n17605) );
  OAI21_X1 U20806 ( .B1(n17606), .B2(n17626), .A(n17605), .ZN(P3_U2790) );
  AOI22_X1 U20807 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17623), .ZN(n17607) );
  OAI21_X1 U20808 ( .B1(n17608), .B2(n17626), .A(n17607), .ZN(P3_U2791) );
  AOI22_X1 U20809 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17623), .ZN(n17609) );
  OAI21_X1 U20810 ( .B1(n17610), .B2(n17626), .A(n17609), .ZN(P3_U2792) );
  AOI22_X1 U20811 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17616), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17615), .ZN(n17611) );
  OAI21_X1 U20812 ( .B1(n17612), .B2(n17626), .A(n17611), .ZN(P3_U2793) );
  AOI22_X1 U20813 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17623), .ZN(n17613) );
  OAI21_X1 U20814 ( .B1(n17614), .B2(n17626), .A(n17613), .ZN(P3_U2794) );
  AOI22_X1 U20815 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17616), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17615), .ZN(n17617) );
  OAI21_X1 U20816 ( .B1(n17618), .B2(n17626), .A(n17617), .ZN(P3_U2795) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17623), .ZN(n17619) );
  OAI21_X1 U20818 ( .B1(n17620), .B2(n17626), .A(n17619), .ZN(P3_U2796) );
  AOI22_X1 U20819 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17623), .ZN(n17621) );
  OAI21_X1 U20820 ( .B1(n17622), .B2(n17626), .A(n17621), .ZN(P3_U2797) );
  AOI22_X1 U20821 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17623), .ZN(n17625) );
  OAI21_X1 U20822 ( .B1(n17627), .B2(n17626), .A(n17625), .ZN(P3_U2798) );
  OAI21_X1 U20823 ( .B1(n17630), .B2(n17629), .A(n17628), .ZN(n17644) );
  OAI21_X1 U20824 ( .B1(n17631), .B2(n17748), .A(n17995), .ZN(n17632) );
  AOI21_X1 U20825 ( .B1(n17955), .B2(n17634), .A(n17632), .ZN(n17662) );
  OAI21_X1 U20826 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17658), .A(
        n17662), .ZN(n17646) );
  NOR3_X1 U20827 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17633), .A3(
        n17783), .ZN(n17640) );
  NOR2_X1 U20828 ( .A1(n17833), .A2(n17634), .ZN(n17650) );
  OAI211_X1 U20829 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17650), .B(n17635), .ZN(n17636) );
  OAI211_X1 U20830 ( .C1(n17845), .C2(n17638), .A(n17637), .B(n17636), .ZN(
        n17639) );
  AOI211_X1 U20831 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17646), .A(
        n17640), .B(n17639), .ZN(n17643) );
  OAI22_X1 U20832 ( .A1(n18000), .A2(n17641), .B1(n17861), .B2(n18009), .ZN(
        n17664) );
  OR2_X1 U20833 ( .A1(n18016), .A2(n17664), .ZN(n17651) );
  OAI211_X1 U20834 ( .C1(n17905), .C2(n17986), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17651), .ZN(n17642) );
  OAI211_X1 U20835 ( .C1(n17903), .C2(n17644), .A(n17643), .B(n17642), .ZN(
        P3_U2802) );
  AOI22_X1 U20836 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17646), .B1(
        n17808), .B2(n17645), .ZN(n17655) );
  OAI21_X1 U20837 ( .B1(n17793), .B2(n17648), .A(n17647), .ZN(n18013) );
  AOI22_X1 U20838 ( .A1(n17859), .A2(n18013), .B1(n17650), .B2(n17649), .ZN(
        n17654) );
  OAI21_X1 U20839 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17652), .A(
        n17651), .ZN(n17653) );
  NAND2_X1 U20840 ( .A1(n18330), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18014) );
  NAND4_X1 U20841 ( .A1(n17655), .A2(n17654), .A3(n17653), .A4(n18014), .ZN(
        P3_U2803) );
  AOI21_X1 U20842 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17657), .A(
        n17656), .ZN(n18018) );
  INV_X1 U20843 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18019) );
  AOI21_X1 U20844 ( .B1(n18752), .B2(n9918), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17661) );
  OAI21_X1 U20845 ( .B1(n17808), .B2(n17773), .A(n17659), .ZN(n17660) );
  NAND2_X1 U20846 ( .A1(n18330), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18021) );
  OAI211_X1 U20847 ( .C1(n17662), .C2(n17661), .A(n17660), .B(n18021), .ZN(
        n17663) );
  AOI221_X1 U20848 ( .B1(n17665), .B2(n18019), .C1(n17664), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17663), .ZN(n17666) );
  OAI21_X1 U20849 ( .B1(n18018), .B2(n17903), .A(n17666), .ZN(P3_U2804) );
  NOR2_X1 U20850 ( .A1(n18034), .A2(n18029), .ZN(n18017) );
  AOI22_X1 U20851 ( .A1(n18034), .A2(n17667), .B1(n18017), .B2(n18068), .ZN(
        n17668) );
  INV_X1 U20852 ( .A(n17668), .ZN(n18035) );
  AOI21_X1 U20853 ( .B1(n18752), .B2(n17670), .A(n17953), .ZN(n17694) );
  OAI21_X1 U20854 ( .B1(n17669), .B2(n17748), .A(n17694), .ZN(n17682) );
  NOR2_X1 U20855 ( .A1(n17833), .A2(n17670), .ZN(n17684) );
  OAI211_X1 U20856 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17684), .B(n17671), .ZN(n17672) );
  NAND2_X1 U20857 ( .A1(n18330), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18033) );
  OAI211_X1 U20858 ( .C1(n17845), .C2(n17673), .A(n17672), .B(n18033), .ZN(
        n17679) );
  XOR2_X1 U20859 ( .A(n17674), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18041) );
  OAI21_X1 U20860 ( .B1(n17902), .B2(n17676), .A(n17675), .ZN(n17677) );
  XOR2_X1 U20861 ( .A(n17677), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18036) );
  OAI22_X1 U20862 ( .A1(n17861), .A2(n18041), .B1(n17903), .B2(n18036), .ZN(
        n17678) );
  AOI211_X1 U20863 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17682), .A(
        n17679), .B(n17678), .ZN(n17680) );
  OAI21_X1 U20864 ( .B1(n18000), .B2(n18035), .A(n17680), .ZN(P3_U2805) );
  INV_X1 U20865 ( .A(n17681), .ZN(n17693) );
  NOR2_X1 U20866 ( .A1(n18216), .A2(n18946), .ZN(n18052) );
  AOI221_X1 U20867 ( .B1(n17684), .B2(n17683), .C1(n17682), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18052), .ZN(n17692) );
  NOR2_X1 U20868 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17685), .ZN(
        n18053) );
  NAND2_X1 U20869 ( .A1(n17686), .A2(n18068), .ZN(n18046) );
  INV_X1 U20870 ( .A(n18044), .ZN(n17687) );
  AOI22_X1 U20871 ( .A1(n17986), .A2(n18046), .B1(n17905), .B2(n17687), .ZN(
        n17701) );
  INV_X1 U20872 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18049) );
  AOI21_X1 U20873 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17689), .A(
        n17688), .ZN(n18055) );
  OAI22_X1 U20874 ( .A1(n17701), .A2(n18049), .B1(n18055), .B2(n17903), .ZN(
        n17690) );
  AOI21_X1 U20875 ( .B1(n17795), .B2(n18053), .A(n17690), .ZN(n17691) );
  OAI211_X1 U20876 ( .C1(n17845), .C2(n17693), .A(n17692), .B(n17691), .ZN(
        P3_U2806) );
  OAI21_X1 U20877 ( .B1(n17695), .B2(n17748), .A(n17694), .ZN(n17697) );
  NOR2_X1 U20878 ( .A1(n18216), .A2(n18945), .ZN(n18059) );
  NAND2_X1 U20879 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17711) );
  INV_X1 U20880 ( .A(n17833), .ZN(n17784) );
  NAND2_X1 U20881 ( .A1(n17710), .A2(n17784), .ZN(n17725) );
  NOR3_X1 U20882 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17711), .A3(
        n17725), .ZN(n17696) );
  AOI211_X1 U20883 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n17697), .A(
        n18059), .B(n17696), .ZN(n17706) );
  AOI22_X1 U20884 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17902), .B1(
        n17698), .B2(n17717), .ZN(n17699) );
  NAND2_X1 U20885 ( .A1(n17744), .A2(n17699), .ZN(n17700) );
  XOR2_X1 U20886 ( .A(n17700), .B(n18002), .Z(n18060) );
  NOR2_X1 U20887 ( .A1(n18073), .A2(n17783), .ZN(n17703) );
  INV_X1 U20888 ( .A(n17701), .ZN(n17702) );
  MUX2_X1 U20889 ( .A(n17703), .B(n17702), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17704) );
  AOI21_X1 U20890 ( .B1(n17859), .B2(n18060), .A(n17704), .ZN(n17705) );
  OAI211_X1 U20891 ( .C1(n17845), .C2(n17707), .A(n17706), .B(n17705), .ZN(
        P3_U2807) );
  NAND2_X1 U20892 ( .A1(n18071), .A2(n17795), .ZN(n17722) );
  NAND2_X1 U20893 ( .A1(n18330), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18080) );
  INV_X1 U20894 ( .A(n18080), .ZN(n17715) );
  NAND2_X1 U20895 ( .A1(n17828), .A2(n17708), .ZN(n17709) );
  OAI211_X1 U20896 ( .C1(n17710), .C2(n17830), .A(n17995), .B(n17709), .ZN(
        n17742) );
  AOI21_X1 U20897 ( .B1(n17773), .B2(n17736), .A(n17742), .ZN(n17723) );
  OAI21_X1 U20898 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17711), .ZN(n17712) );
  OAI22_X1 U20899 ( .A1(n17723), .A2(n17713), .B1(n17725), .B2(n17712), .ZN(
        n17714) );
  AOI211_X1 U20900 ( .C1(n17716), .C2(n17808), .A(n17715), .B(n17714), .ZN(
        n17721) );
  NOR2_X1 U20901 ( .A1(n17905), .A2(n17986), .ZN(n17743) );
  AOI22_X1 U20902 ( .A1(n17986), .A2(n18150), .B1(n17905), .B2(n18067), .ZN(
        n17798) );
  OAI21_X1 U20903 ( .B1(n18071), .B2(n17743), .A(n17798), .ZN(n17733) );
  INV_X1 U20904 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18082) );
  INV_X1 U20905 ( .A(n17717), .ZN(n17718) );
  OAI221_X1 U20906 ( .B1(n17718), .B2(n18071), .C1(n17718), .C2(n17792), .A(
        n17744), .ZN(n17719) );
  XOR2_X1 U20907 ( .A(n18082), .B(n17719), .Z(n18079) );
  AOI22_X1 U20908 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17733), .B1(
        n17859), .B2(n18079), .ZN(n17720) );
  OAI211_X1 U20909 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17722), .A(
        n17721), .B(n17720), .ZN(P3_U2808) );
  INV_X1 U20910 ( .A(n18087), .ZN(n17731) );
  NAND2_X1 U20911 ( .A1(n17731), .A2(n18088), .ZN(n18094) );
  NAND2_X1 U20912 ( .A1(n18065), .A2(n17795), .ZN(n17761) );
  NAND2_X1 U20913 ( .A1(n18330), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18092) );
  OAI221_X1 U20914 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17725), .C1(
        n17724), .C2(n17723), .A(n18092), .ZN(n17726) );
  AOI21_X1 U20915 ( .B1(n17808), .B2(n17727), .A(n17726), .ZN(n17735) );
  INV_X1 U20916 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18123) );
  NOR3_X1 U20917 ( .A1(n17902), .A2(n18123), .A3(n17728), .ZN(n17756) );
  INV_X1 U20918 ( .A(n17729), .ZN(n17769) );
  AOI22_X1 U20919 ( .A1(n17731), .A2(n17756), .B1(n17769), .B2(n17730), .ZN(
        n17732) );
  XOR2_X1 U20920 ( .A(n18088), .B(n17732), .Z(n18091) );
  AOI22_X1 U20921 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17733), .B1(
        n17859), .B2(n18091), .ZN(n17734) );
  OAI211_X1 U20922 ( .C1(n18094), .C2(n17761), .A(n17735), .B(n17734), .ZN(
        P3_U2809) );
  INV_X1 U20923 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18098) );
  NAND2_X1 U20924 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18098), .ZN(
        n18104) );
  OAI21_X1 U20925 ( .B1(n17737), .B2(n18680), .A(n17736), .ZN(n17741) );
  INV_X1 U20926 ( .A(n17738), .ZN(n17739) );
  AOI21_X1 U20927 ( .B1(n17845), .B2(n17658), .A(n17739), .ZN(n17740) );
  NOR2_X1 U20928 ( .A1(n18216), .A2(n18938), .ZN(n18101) );
  AOI211_X1 U20929 ( .C1(n17742), .C2(n17741), .A(n17740), .B(n18101), .ZN(
        n17747) );
  NOR2_X1 U20930 ( .A1(n18083), .A2(n18109), .ZN(n18095) );
  OAI21_X1 U20931 ( .B1(n17743), .B2(n18095), .A(n17798), .ZN(n17758) );
  OAI221_X1 U20932 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17768), 
        .C1(n18109), .C2(n17756), .A(n17744), .ZN(n17745) );
  XOR2_X1 U20933 ( .A(n18098), .B(n17745), .Z(n18102) );
  AOI22_X1 U20934 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17758), .B1(
        n17859), .B2(n18102), .ZN(n17746) );
  OAI211_X1 U20935 ( .C1(n17761), .C2(n18104), .A(n17747), .B(n17746), .ZN(
        P3_U2810) );
  INV_X1 U20936 ( .A(n17751), .ZN(n17762) );
  AOI21_X1 U20937 ( .B1(n17955), .B2(n17762), .A(n17953), .ZN(n17774) );
  OAI21_X1 U20938 ( .B1(n17749), .B2(n17748), .A(n17774), .ZN(n17765) );
  NOR2_X1 U20939 ( .A1(n18216), .A2(n18936), .ZN(n18105) );
  NOR2_X1 U20940 ( .A1(n17766), .A2(n17750), .ZN(n17754) );
  OAI211_X1 U20941 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17751), .B(n17784), .ZN(n17753) );
  OAI22_X1 U20942 ( .A1(n17754), .A2(n17753), .B1(n17752), .B2(n17845), .ZN(
        n17755) );
  AOI211_X1 U20943 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17765), .A(
        n18105), .B(n17755), .ZN(n17760) );
  AOI21_X1 U20944 ( .B1(n17768), .B2(n17769), .A(n17756), .ZN(n17757) );
  XOR2_X1 U20945 ( .A(n18109), .B(n17757), .Z(n18106) );
  AOI22_X1 U20946 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17758), .B1(
        n17859), .B2(n18106), .ZN(n17759) );
  OAI211_X1 U20947 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17761), .A(
        n17760), .B(n17759), .ZN(P3_U2811) );
  NAND2_X1 U20948 ( .A1(n18120), .A2(n18123), .ZN(n18128) );
  NOR2_X1 U20949 ( .A1(n17833), .A2(n17762), .ZN(n17767) );
  OAI22_X1 U20950 ( .A1(n18216), .A2(n18934), .B1(n17845), .B2(n17763), .ZN(
        n17764) );
  AOI221_X1 U20951 ( .B1(n17767), .B2(n17766), .C1(n17765), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17764), .ZN(n17772) );
  OAI21_X1 U20952 ( .B1(n18120), .B2(n17783), .A(n17798), .ZN(n17780) );
  AOI21_X1 U20953 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17793), .A(
        n17768), .ZN(n17770) );
  XOR2_X1 U20954 ( .A(n17770), .B(n17769), .Z(n18125) );
  AOI22_X1 U20955 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17780), .B1(
        n17859), .B2(n18125), .ZN(n17771) );
  OAI211_X1 U20956 ( .C1(n17783), .C2(n18128), .A(n17772), .B(n17771), .ZN(
        P3_U2812) );
  NAND2_X1 U20957 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18129), .ZN(
        n18135) );
  NOR2_X1 U20958 ( .A1(n18216), .A2(n18933), .ZN(n18132) );
  AOI221_X1 U20959 ( .B1(n17776), .B2(n17775), .C1(n18680), .C2(n17775), .A(
        n17774), .ZN(n17777) );
  AOI211_X1 U20960 ( .C1(n17778), .C2(n17988), .A(n18132), .B(n17777), .ZN(
        n17782) );
  OAI21_X1 U20961 ( .B1(n10446), .B2(n18129), .A(n17779), .ZN(n18133) );
  AOI22_X1 U20962 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17780), .B1(
        n17859), .B2(n18133), .ZN(n17781) );
  OAI211_X1 U20963 ( .C1(n17783), .C2(n18135), .A(n17782), .B(n17781), .ZN(
        P3_U2813) );
  INV_X1 U20964 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17787) );
  NAND2_X1 U20965 ( .A1(n9923), .A2(n17784), .ZN(n17801) );
  AOI221_X1 U20966 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17800), .C2(n17787), .A(
        n17801), .ZN(n17789) );
  OAI21_X1 U20967 ( .B1(n9923), .B2(n17830), .A(n17995), .ZN(n17819) );
  AOI21_X1 U20968 ( .B1(n17828), .B2(n17785), .A(n17819), .ZN(n17799) );
  OAI22_X1 U20969 ( .A1(n17799), .A2(n17787), .B1(n17845), .B2(n17786), .ZN(
        n17788) );
  AOI211_X1 U20970 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n18330), .A(n17789), 
        .B(n17788), .ZN(n17797) );
  NAND4_X1 U20971 ( .A1(n17793), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n17790), .ZN(n17884) );
  OAI22_X1 U20972 ( .A1(n17793), .A2(n17792), .B1(n17884), .B2(n17791), .ZN(
        n17794) );
  XOR2_X1 U20973 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17794), .Z(
        n18146) );
  AOI22_X1 U20974 ( .A1(n17859), .A2(n18146), .B1(n17795), .B2(n18142), .ZN(
        n17796) );
  OAI211_X1 U20975 ( .C1(n17798), .C2(n18142), .A(n17797), .B(n17796), .ZN(
        P3_U2814) );
  NOR3_X1 U20976 ( .A1(n18198), .A2(n18170), .A3(n17820), .ZN(n17821) );
  NOR2_X1 U20977 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17821), .ZN(
        n18154) );
  NAND2_X1 U20978 ( .A1(n17905), .A2(n18067), .ZN(n17810) );
  NAND2_X1 U20979 ( .A1(n18330), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18160) );
  OAI221_X1 U20980 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17801), .C1(
        n17800), .C2(n17799), .A(n18160), .ZN(n17806) );
  NOR3_X1 U20981 ( .A1(n18196), .A2(n17820), .A3(n18170), .ZN(n17823) );
  NOR2_X1 U20982 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17823), .ZN(
        n18156) );
  NAND2_X1 U20983 ( .A1(n17986), .A2(n18150), .ZN(n17804) );
  NOR2_X1 U20984 ( .A1(n17839), .A2(n17884), .ZN(n17811) );
  NAND2_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n10398), .ZN(
        n18187) );
  OAI221_X1 U20986 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17812), 
        .C1(n18170), .C2(n17811), .A(n18187), .ZN(n17802) );
  XOR2_X1 U20987 ( .A(n15817), .B(n17802), .Z(n18158) );
  INV_X1 U20988 ( .A(n18158), .ZN(n17803) );
  OAI22_X1 U20989 ( .A1(n18156), .A2(n17804), .B1(n17903), .B2(n17803), .ZN(
        n17805) );
  AOI211_X1 U20990 ( .C1(n17808), .C2(n17807), .A(n17806), .B(n17805), .ZN(
        n17809) );
  OAI21_X1 U20991 ( .B1(n18154), .B2(n17810), .A(n17809), .ZN(P3_U2815) );
  OAI21_X1 U20992 ( .B1(n17812), .B2(n17811), .A(n18187), .ZN(n17813) );
  XOR2_X1 U20993 ( .A(n17813), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18176) );
  NAND2_X1 U20994 ( .A1(n17814), .A2(n18752), .ZN(n17930) );
  NOR2_X1 U20995 ( .A1(n17929), .A2(n17930), .ZN(n17913) );
  NAND2_X1 U20996 ( .A1(n17831), .A2(n17913), .ZN(n17865) );
  OAI21_X1 U20997 ( .B1(n17834), .B2(n17865), .A(n17815), .ZN(n17818) );
  INV_X1 U20998 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18927) );
  OAI22_X1 U20999 ( .A1(n17968), .A2(n17816), .B1(n18216), .B2(n18927), .ZN(
        n17817) );
  AOI21_X1 U21000 ( .B1(n17819), .B2(n17818), .A(n17817), .ZN(n17826) );
  INV_X1 U21001 ( .A(n17820), .ZN(n18167) );
  NAND2_X1 U21002 ( .A1(n17862), .A2(n18167), .ZN(n17822) );
  AOI21_X1 U21003 ( .B1(n18170), .B2(n17822), .A(n17821), .ZN(n18173) );
  NAND2_X1 U21004 ( .A1(n18167), .A2(n17860), .ZN(n17824) );
  AOI21_X1 U21005 ( .B1(n18170), .B2(n17824), .A(n17823), .ZN(n18172) );
  AOI22_X1 U21006 ( .A1(n17905), .A2(n18173), .B1(n17986), .B2(n18172), .ZN(
        n17825) );
  OAI211_X1 U21007 ( .C1(n17903), .C2(n18176), .A(n17826), .B(n17825), .ZN(
        P3_U2816) );
  NAND2_X1 U21008 ( .A1(n18178), .A2(n17891), .ZN(n17855) );
  OAI21_X1 U21009 ( .B1(n17894), .B2(n17830), .A(n17995), .ZN(n17911) );
  AOI21_X1 U21010 ( .B1(n17828), .B2(n17827), .A(n17911), .ZN(n17829) );
  OAI21_X1 U21011 ( .B1(n17831), .B2(n17830), .A(n17829), .ZN(n17847) );
  NOR2_X1 U21012 ( .A1(n17833), .A2(n17832), .ZN(n17849) );
  OAI211_X1 U21013 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17849), .B(n17834), .ZN(n17836) );
  NAND2_X1 U21014 ( .A1(n18330), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17835) );
  OAI211_X1 U21015 ( .C1(n17845), .C2(n17837), .A(n17836), .B(n17835), .ZN(
        n17838) );
  AOI21_X1 U21016 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17847), .A(
        n17838), .ZN(n17843) );
  NOR2_X1 U21017 ( .A1(n18196), .A2(n17839), .ZN(n18181) );
  NOR2_X1 U21018 ( .A1(n18198), .A2(n17839), .ZN(n18180) );
  OAI22_X1 U21019 ( .A1(n18181), .A2(n18000), .B1(n18180), .B2(n17861), .ZN(
        n17852) );
  AOI22_X1 U21020 ( .A1(n18162), .A2(n17874), .B1(n17902), .B2(n18195), .ZN(
        n17840) );
  AOI21_X1 U21021 ( .B1(n17850), .B2(n17902), .A(n17840), .ZN(n17841) );
  XOR2_X1 U21022 ( .A(n17841), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18177) );
  AOI22_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17852), .B1(
        n17859), .B2(n18177), .ZN(n17842) );
  OAI211_X1 U21024 ( .C1(n18187), .C2(n17855), .A(n17843), .B(n17842), .ZN(
        P3_U2817) );
  NAND2_X1 U21025 ( .A1(n18330), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18193) );
  OAI21_X1 U21026 ( .B1(n17845), .B2(n17844), .A(n18193), .ZN(n17846) );
  AOI221_X1 U21027 ( .B1(n17849), .B2(n17848), .C1(n17847), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17846), .ZN(n17854) );
  OAI21_X1 U21028 ( .B1(n17857), .B2(n9893), .A(n17850), .ZN(n17851) );
  XOR2_X1 U21029 ( .A(n17851), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18192) );
  AOI22_X1 U21030 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17852), .B1(
        n17859), .B2(n18192), .ZN(n17853) );
  OAI211_X1 U21031 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17855), .A(
        n17854), .B(n17853), .ZN(P3_U2818) );
  AOI22_X1 U21032 ( .A1(n18330), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17856), 
        .B2(n17988), .ZN(n17869) );
  XOR2_X1 U21033 ( .A(n17858), .B(n17857), .Z(n18208) );
  NOR2_X1 U21034 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18204), .ZN(
        n18207) );
  AOI22_X1 U21035 ( .A1(n17859), .A2(n18208), .B1(n18207), .B2(n17891), .ZN(
        n17868) );
  AND2_X1 U21036 ( .A1(n18204), .A2(n17891), .ZN(n17863) );
  OAI22_X1 U21037 ( .A1(n17862), .A2(n17861), .B1(n18000), .B2(n17860), .ZN(
        n17892) );
  OAI21_X1 U21038 ( .B1(n17863), .B2(n17892), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17867) );
  NAND2_X1 U21039 ( .A1(n17895), .A2(n17913), .ZN(n17889) );
  NOR2_X1 U21040 ( .A1(n17864), .A2(n17889), .ZN(n17882) );
  OAI211_X1 U21041 ( .C1(n17882), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17989), .B(n17865), .ZN(n17866) );
  NAND4_X1 U21042 ( .A1(n17869), .A2(n17868), .A3(n17867), .A4(n17866), .ZN(
        P3_U2819) );
  INV_X1 U21043 ( .A(n17889), .ZN(n17870) );
  AOI22_X1 U21044 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17870), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17989), .ZN(n17881) );
  NOR2_X1 U21045 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17876) );
  AOI22_X1 U21046 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17892), .B1(
        n18204), .B2(n17891), .ZN(n17875) );
  INV_X1 U21047 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18220) );
  NAND3_X1 U21048 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17902), .A3(
        n18220), .ZN(n17873) );
  INV_X1 U21049 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17871) );
  OAI221_X1 U21050 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17883), .C1(
        n18220), .C2(n17884), .A(n17871), .ZN(n17872) );
  OAI211_X1 U21051 ( .C1(n17874), .C2(n17873), .A(n17872), .B(n9893), .ZN(
        n18219) );
  OAI22_X1 U21052 ( .A1(n17876), .A2(n17875), .B1(n18219), .B2(n17903), .ZN(
        n17877) );
  AOI21_X1 U21053 ( .B1(n17878), .B2(n17988), .A(n17877), .ZN(n17880) );
  NAND2_X1 U21054 ( .A1(n18330), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17879) );
  OAI211_X1 U21055 ( .C1(n17882), .C2(n17881), .A(n17880), .B(n17879), .ZN(
        P3_U2820) );
  NAND2_X1 U21056 ( .A1(n17884), .A2(n17883), .ZN(n17885) );
  XOR2_X1 U21057 ( .A(n17885), .B(n18220), .Z(n18230) );
  NAND3_X1 U21058 ( .A1(n17989), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17889), .ZN(n17888) );
  AOI22_X1 U21059 ( .A1(n18330), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17886), 
        .B2(n17988), .ZN(n17887) );
  OAI211_X1 U21060 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17889), .A(
        n17888), .B(n17887), .ZN(n17890) );
  AOI221_X1 U21061 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17892), .C1(
        n18220), .C2(n17891), .A(n17890), .ZN(n17893) );
  OAI21_X1 U21062 ( .B1(n18230), .B2(n17903), .A(n17893), .ZN(P3_U2821) );
  INV_X1 U21063 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18915) );
  NOR2_X1 U21064 ( .A1(n18216), .A2(n18915), .ZN(n18235) );
  NAND2_X1 U21065 ( .A1(n17894), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17896) );
  AOI211_X1 U21066 ( .C1(n17897), .C2(n17896), .A(n17895), .B(n18680), .ZN(
        n17898) );
  AOI211_X1 U21067 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17911), .A(
        n18235), .B(n17898), .ZN(n17907) );
  OAI21_X1 U21068 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17900), .A(
        n17899), .ZN(n18246) );
  OAI21_X1 U21069 ( .B1(n18243), .B2(n17902), .A(n17901), .ZN(n18239) );
  OAI22_X1 U21070 ( .A1(n18000), .A2(n18246), .B1(n17903), .B2(n18239), .ZN(
        n17904) );
  AOI21_X1 U21071 ( .B1(n18243), .B2(n17905), .A(n17904), .ZN(n17906) );
  OAI211_X1 U21072 ( .C1(n17968), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        P3_U2822) );
  OAI21_X1 U21073 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17910), .A(
        n17909), .ZN(n18257) );
  NOR2_X1 U21074 ( .A1(n18216), .A2(n18912), .ZN(n18247) );
  AOI221_X1 U21075 ( .B1(n17913), .B2(n17912), .C1(n17911), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18247), .ZN(n17919) );
  NOR2_X1 U21076 ( .A1(n17915), .A2(n17914), .ZN(n17916) );
  XOR2_X1 U21077 ( .A(n17916), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18248) );
  AOI22_X1 U21078 ( .A1(n17986), .A2(n18248), .B1(n17917), .B2(n17988), .ZN(
        n17918) );
  OAI211_X1 U21079 ( .C1(n17999), .C2(n18257), .A(n17919), .B(n17918), .ZN(
        P3_U2823) );
  OAI21_X1 U21080 ( .B1(n17922), .B2(n17921), .A(n17920), .ZN(n18264) );
  NAND2_X1 U21081 ( .A1(n17989), .A2(n17930), .ZN(n17940) );
  AOI22_X1 U21082 ( .A1(n17925), .A2(n17936), .B1(n17924), .B2(n17923), .ZN(
        n17927) );
  XOR2_X1 U21083 ( .A(n17927), .B(n17926), .Z(n18261) );
  AOI22_X1 U21084 ( .A1(n18330), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17986), 
        .B2(n18261), .ZN(n17928) );
  OAI221_X1 U21085 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17930), .C1(
        n17929), .C2(n17940), .A(n17928), .ZN(n17931) );
  AOI21_X1 U21086 ( .B1(n17932), .B2(n17988), .A(n17931), .ZN(n17933) );
  OAI21_X1 U21087 ( .B1(n17999), .B2(n18264), .A(n17933), .ZN(P3_U2824) );
  OAI21_X1 U21088 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17935), .A(
        n17934), .ZN(n18273) );
  AOI21_X1 U21089 ( .B1(n17938), .B2(n17937), .A(n17936), .ZN(n18265) );
  AOI21_X1 U21090 ( .B1(n17939), .B2(n17995), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17941) );
  OAI22_X1 U21091 ( .A1(n17968), .A2(n17942), .B1(n17941), .B2(n17940), .ZN(
        n17943) );
  AOI21_X1 U21092 ( .B1(n17986), .B2(n18265), .A(n17943), .ZN(n17944) );
  NAND2_X1 U21093 ( .A1(n18330), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18266) );
  OAI211_X1 U21094 ( .C1(n17999), .C2(n18273), .A(n17944), .B(n18266), .ZN(
        P3_U2825) );
  AOI21_X1 U21095 ( .B1(n17947), .B2(n17946), .A(n17945), .ZN(n18279) );
  INV_X1 U21096 ( .A(n17948), .ZN(n17949) );
  AOI22_X1 U21097 ( .A1(n17986), .A2(n18279), .B1(n18752), .B2(n17949), .ZN(
        n17960) );
  OAI21_X1 U21098 ( .B1(n17952), .B2(n17951), .A(n17950), .ZN(n18282) );
  AOI21_X1 U21099 ( .B1(n17955), .B2(n17954), .A(n17953), .ZN(n17972) );
  OAI22_X1 U21100 ( .A1(n17999), .A2(n18282), .B1(n17956), .B2(n17972), .ZN(
        n17957) );
  AOI21_X1 U21101 ( .B1(n17958), .B2(n17988), .A(n17957), .ZN(n17959) );
  OAI211_X1 U21102 ( .C1(n18216), .C2(n18906), .A(n17960), .B(n17959), .ZN(
        P3_U2826) );
  NAND2_X1 U21103 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17995), .ZN(
        n17977) );
  AOI21_X1 U21104 ( .B1(n17963), .B2(n17962), .A(n17961), .ZN(n18286) );
  INV_X1 U21105 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18904) );
  NOR2_X1 U21106 ( .A1(n18216), .A2(n18904), .ZN(n18285) );
  OAI21_X1 U21107 ( .B1(n17966), .B2(n17965), .A(n17964), .ZN(n18283) );
  OAI22_X1 U21108 ( .A1(n17968), .A2(n17967), .B1(n17999), .B2(n18283), .ZN(
        n17969) );
  AOI211_X1 U21109 ( .C1(n17986), .C2(n18286), .A(n18285), .B(n17969), .ZN(
        n17970) );
  OAI221_X1 U21110 ( .B1(n17972), .B2(n17971), .C1(n17972), .C2(n17977), .A(
        n17970), .ZN(P3_U2827) );
  AOI21_X1 U21111 ( .B1(n17975), .B2(n17974), .A(n17973), .ZN(n18308) );
  AOI22_X1 U21112 ( .A1(n17986), .A2(n18308), .B1(n17976), .B2(n17988), .ZN(
        n17981) );
  OAI21_X1 U21113 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18752), .A(
        n17977), .ZN(n17980) );
  NAND2_X1 U21114 ( .A1(n18330), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18309) );
  OAI211_X1 U21115 ( .C1(n18294), .C2(n18293), .A(n17978), .B(n18292), .ZN(
        n17979) );
  NAND4_X1 U21116 ( .A1(n17981), .A2(n17980), .A3(n18309), .A4(n17979), .ZN(
        P3_U2828) );
  OAI21_X1 U21117 ( .B1(n17993), .B2(n17983), .A(n17982), .ZN(n18319) );
  OAI21_X1 U21118 ( .B1(n17992), .B2(n17985), .A(n17984), .ZN(n18321) );
  AOI22_X1 U21119 ( .A1(n18330), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17986), 
        .B2(n18321), .ZN(n17991) );
  AOI22_X1 U21120 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17989), .B1(
        n17988), .B2(n17987), .ZN(n17990) );
  OAI211_X1 U21121 ( .C1(n17999), .C2(n18319), .A(n17991), .B(n17990), .ZN(
        P3_U2829) );
  NOR2_X1 U21122 ( .A1(n17993), .A2(n17992), .ZN(n18335) );
  INV_X1 U21123 ( .A(n18335), .ZN(n18333) );
  INV_X1 U21124 ( .A(n17994), .ZN(n17996) );
  NOR2_X1 U21125 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19028) );
  OAI21_X1 U21126 ( .B1(n17996), .B2(n19028), .A(n17995), .ZN(n17997) );
  AOI22_X1 U21127 ( .A1(n18330), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17997), .ZN(n17998) );
  OAI221_X1 U21128 ( .B1(n18335), .B2(n18000), .C1(n18333), .C2(n17999), .A(
        n17998), .ZN(P3_U2830) );
  NOR2_X1 U21129 ( .A1(n18057), .A2(n18001), .ZN(n18012) );
  NOR2_X1 U21130 ( .A1(n18002), .A2(n18049), .ZN(n18005) );
  INV_X1 U21131 ( .A(n18137), .ZN(n18003) );
  OAI211_X1 U21132 ( .C1(n18224), .C2(n18003), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18071), .ZN(n18004) );
  OAI21_X1 U21133 ( .B1(n18117), .B2(n18004), .A(n18231), .ZN(n18043) );
  OAI21_X1 U21134 ( .B1(n18005), .B2(n18296), .A(n18043), .ZN(n18027) );
  NAND2_X1 U21135 ( .A1(n18006), .A2(n18231), .ZN(n18007) );
  OAI211_X1 U21136 ( .C1(n18009), .C2(n18179), .A(n18008), .B(n18007), .ZN(
        n18010) );
  OAI211_X1 U21137 ( .C1(n18317), .C2(n18016), .A(n18015), .B(n18014), .ZN(
        P3_U2835) );
  AOI22_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18315), .B1(
        n18064), .B2(n18017), .ZN(n18023) );
  OAI22_X1 U21139 ( .A1(n18019), .A2(n18317), .B1(n18229), .B2(n18018), .ZN(
        n18020) );
  INV_X1 U21140 ( .A(n18020), .ZN(n18022) );
  OAI211_X1 U21141 ( .C1(n18024), .C2(n18023), .A(n18022), .B(n18021), .ZN(
        P3_U2836) );
  INV_X1 U21142 ( .A(n18025), .ZN(n18026) );
  NOR2_X1 U21143 ( .A1(n18026), .A2(n18029), .ZN(n18032) );
  AOI221_X1 U21144 ( .B1(n18029), .B2(n10244), .C1(n18028), .C2(n10244), .A(
        n18027), .ZN(n18030) );
  INV_X1 U21145 ( .A(n18030), .ZN(n18031) );
  MUX2_X1 U21146 ( .A(n18032), .B(n18031), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n18039) );
  OAI21_X1 U21147 ( .B1(n18317), .B2(n18034), .A(n18033), .ZN(n18038) );
  OAI22_X1 U21148 ( .A1(n18229), .A2(n18036), .B1(n18334), .B2(n18035), .ZN(
        n18037) );
  AOI211_X1 U21149 ( .C1(n18325), .C2(n18039), .A(n18038), .B(n18037), .ZN(
        n18040) );
  OAI21_X1 U21150 ( .B1(n18042), .B2(n18041), .A(n18040), .ZN(P3_U2837) );
  OAI211_X1 U21151 ( .C1(n18044), .C2(n18179), .A(n18317), .B(n18043), .ZN(
        n18045) );
  AOI21_X1 U21152 ( .B1(n18197), .B2(n18046), .A(n18045), .ZN(n18050) );
  OAI211_X1 U21153 ( .C1(n18047), .C2(n18835), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18050), .ZN(n18048) );
  NAND2_X1 U21154 ( .A1(n18216), .A2(n18048), .ZN(n18062) );
  AOI211_X1 U21155 ( .C1(n18050), .C2(n18144), .A(n18049), .B(n18062), .ZN(
        n18051) );
  AOI211_X1 U21156 ( .C1(n18053), .C2(n18064), .A(n18052), .B(n18051), .ZN(
        n18054) );
  OAI21_X1 U21157 ( .B1(n18055), .B2(n18229), .A(n18054), .ZN(P3_U2838) );
  NOR3_X1 U21158 ( .A1(n18057), .A2(n18073), .A3(n18056), .ZN(n18058) );
  NOR2_X1 U21159 ( .A1(n18058), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18063) );
  AOI21_X1 U21160 ( .B1(n18060), .B2(n18241), .A(n18059), .ZN(n18061) );
  OAI21_X1 U21161 ( .B1(n18063), .B2(n18062), .A(n18061), .ZN(P3_U2839) );
  NAND2_X1 U21162 ( .A1(n18065), .A2(n18064), .ZN(n18110) );
  OAI22_X1 U21163 ( .A1(n18072), .A2(n18110), .B1(n18082), .B2(n18305), .ZN(
        n18078) );
  AOI21_X1 U21164 ( .B1(n18066), .B2(n18095), .A(n10247), .ZN(n18069) );
  NAND2_X1 U21165 ( .A1(n18199), .A2(n18067), .ZN(n18155) );
  OAI21_X1 U21166 ( .B1(n18068), .B2(n18811), .A(n18155), .ZN(n18136) );
  AOI211_X1 U21167 ( .C1(n10244), .C2(n18070), .A(n18069), .B(n18136), .ZN(
        n18085) );
  NAND2_X1 U21168 ( .A1(n18179), .A2(n18811), .ZN(n18203) );
  INV_X1 U21169 ( .A(n18203), .ZN(n18119) );
  OAI22_X1 U21170 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10247), .B1(
        n18071), .B2(n18119), .ZN(n18086) );
  INV_X1 U21171 ( .A(n18086), .ZN(n18076) );
  AOI22_X1 U21172 ( .A1(n10244), .A2(n18072), .B1(n18088), .B2(n18826), .ZN(
        n18075) );
  OAI22_X1 U21173 ( .A1(n18082), .A2(n18841), .B1(n18073), .B2(n18137), .ZN(
        n18074) );
  NAND4_X1 U21174 ( .A1(n18085), .A2(n18076), .A3(n18075), .A4(n18074), .ZN(
        n18077) );
  AOI22_X1 U21175 ( .A1(n18241), .A2(n18079), .B1(n18078), .B2(n18077), .ZN(
        n18081) );
  OAI211_X1 U21176 ( .C1(n18317), .C2(n18082), .A(n18081), .B(n18080), .ZN(
        P3_U2840) );
  OAI21_X1 U21177 ( .B1(n18083), .B2(n18137), .A(n18841), .ZN(n18084) );
  NAND3_X1 U21178 ( .A1(n18085), .A2(n18315), .A3(n18084), .ZN(n18097) );
  AOI211_X1 U21179 ( .C1(n18087), .C2(n18316), .A(n18097), .B(n18086), .ZN(
        n18089) );
  NOR3_X1 U21180 ( .A1(n18330), .A2(n18089), .A3(n18088), .ZN(n18090) );
  AOI21_X1 U21181 ( .B1(n18241), .B2(n18091), .A(n18090), .ZN(n18093) );
  OAI211_X1 U21182 ( .C1(n18094), .C2(n18110), .A(n18093), .B(n18092), .ZN(
        P3_U2841) );
  NOR2_X1 U21183 ( .A1(n18095), .A2(n18119), .ZN(n18096) );
  OAI21_X1 U21184 ( .B1(n18097), .B2(n18096), .A(n18216), .ZN(n18108) );
  NAND3_X1 U21185 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18109), .A3(n18316), 
        .ZN(n18099) );
  AOI21_X1 U21186 ( .B1(n18108), .B2(n18099), .A(n18098), .ZN(n18100) );
  AOI211_X1 U21187 ( .C1(n18102), .C2(n18241), .A(n18101), .B(n18100), .ZN(
        n18103) );
  OAI21_X1 U21188 ( .B1(n18104), .B2(n18110), .A(n18103), .ZN(P3_U2842) );
  AOI21_X1 U21189 ( .B1(n18241), .B2(n18106), .A(n18105), .ZN(n18107) );
  OAI221_X1 U21190 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18110), 
        .C1(n18109), .C2(n18108), .A(n18107), .ZN(P3_U2843) );
  OAI22_X1 U21191 ( .A1(n18111), .A2(n18835), .B1(n18232), .B2(n18298), .ZN(
        n18288) );
  OAI21_X1 U21192 ( .B1(n18113), .B2(n18166), .A(n18325), .ZN(n18114) );
  NAND2_X1 U21193 ( .A1(n18115), .A2(n18221), .ZN(n18149) );
  AOI21_X1 U21194 ( .B1(n18120), .B2(n18116), .A(n18835), .ZN(n18122) );
  NOR2_X1 U21195 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18224), .ZN(
        n18295) );
  NOR3_X1 U21196 ( .A1(n18295), .A2(n18117), .A3(n18142), .ZN(n18118) );
  OAI22_X1 U21197 ( .A1(n18120), .A2(n18119), .B1(n18296), .B2(n18118), .ZN(
        n18121) );
  NOR4_X1 U21198 ( .A1(n18122), .A2(n18136), .A3(n18305), .A4(n18121), .ZN(
        n18130) );
  AOI221_X1 U21199 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18130), 
        .C1(n18296), .C2(n18130), .A(n18123), .ZN(n18124) );
  AOI22_X1 U21200 ( .A1(n18125), .A2(n18241), .B1(n18124), .B2(n18216), .ZN(
        n18127) );
  NAND2_X1 U21201 ( .A1(n18330), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18126) );
  OAI211_X1 U21202 ( .C1(n18128), .C2(n18149), .A(n18127), .B(n18126), .ZN(
        P3_U2844) );
  NOR3_X1 U21203 ( .A1(n18330), .A2(n18130), .A3(n18129), .ZN(n18131) );
  AOI211_X1 U21204 ( .C1(n18241), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        n18134) );
  OAI21_X1 U21205 ( .B1(n18149), .B2(n18135), .A(n18134), .ZN(P3_U2845) );
  NOR2_X1 U21206 ( .A1(n18305), .A2(n18136), .ZN(n18143) );
  OAI21_X1 U21207 ( .B1(n18841), .B2(n15817), .A(n18137), .ZN(n18140) );
  NAND2_X1 U21208 ( .A1(n10244), .A2(n18138), .ZN(n18201) );
  NAND2_X1 U21209 ( .A1(n18826), .A2(n18139), .ZN(n18212) );
  AND2_X1 U21210 ( .A1(n18201), .A2(n18212), .ZN(n18223) );
  OAI211_X1 U21211 ( .C1(n18151), .C2(n18214), .A(n18140), .B(n18223), .ZN(
        n18141) );
  INV_X1 U21212 ( .A(n18141), .ZN(n18152) );
  AOI221_X1 U21213 ( .B1(n18144), .B2(n18143), .C1(n18152), .C2(n18143), .A(
        n18142), .ZN(n18145) );
  AOI22_X1 U21214 ( .A1(n18241), .A2(n18146), .B1(n18145), .B2(n18216), .ZN(
        n18148) );
  NAND2_X1 U21215 ( .A1(n18330), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18147) );
  OAI211_X1 U21216 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18149), .A(
        n18148), .B(n18147), .ZN(P3_U2846) );
  NAND2_X1 U21217 ( .A1(n18197), .A2(n18150), .ZN(n18157) );
  AOI21_X1 U21218 ( .B1(n18151), .B2(n18166), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18153) );
  OAI222_X1 U21219 ( .A1(n18157), .A2(n18156), .B1(n18155), .B2(n18154), .C1(
        n18153), .C2(n18152), .ZN(n18159) );
  AOI22_X1 U21220 ( .A1(n18325), .A2(n18159), .B1(n18241), .B2(n18158), .ZN(
        n18161) );
  OAI211_X1 U21221 ( .C1(n18317), .C2(n15817), .A(n18161), .B(n18160), .ZN(
        P3_U2847) );
  OAI221_X1 U21222 ( .B1(n18224), .B2(n18162), .C1(n18224), .C2(n18222), .A(
        n18201), .ZN(n18183) );
  AOI21_X1 U21223 ( .B1(n18212), .B2(n18167), .A(n18214), .ZN(n18163) );
  AOI211_X1 U21224 ( .C1(n10398), .C2(n18316), .A(n18170), .B(n18163), .ZN(
        n18164) );
  INV_X1 U21225 ( .A(n18164), .ZN(n18165) );
  OAI21_X1 U21226 ( .B1(n18183), .B2(n18165), .A(n18325), .ZN(n18169) );
  NAND2_X1 U21227 ( .A1(n18167), .A2(n18166), .ZN(n18168) );
  AOI222_X1 U21228 ( .A1(n18170), .A2(n18169), .B1(n18170), .B2(n18168), .C1(
        n18169), .C2(n18317), .ZN(n18171) );
  AOI21_X1 U21229 ( .B1(n18330), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18171), 
        .ZN(n18175) );
  AOI22_X1 U21230 ( .A1(n18242), .A2(n18173), .B1(n18322), .B2(n18172), .ZN(
        n18174) );
  OAI211_X1 U21231 ( .C1(n18229), .C2(n18176), .A(n18175), .B(n18174), .ZN(
        P3_U2848) );
  NAND2_X1 U21232 ( .A1(n18178), .A2(n18221), .ZN(n18189) );
  AOI22_X1 U21233 ( .A1(n18330), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18241), 
        .B2(n18177), .ZN(n18186) );
  AOI21_X1 U21234 ( .B1(n18178), .B2(n18212), .A(n18214), .ZN(n18206) );
  OAI22_X1 U21235 ( .A1(n18181), .A2(n18811), .B1(n18180), .B2(n18179), .ZN(
        n18182) );
  NOR3_X1 U21236 ( .A1(n18206), .A2(n18183), .A3(n18182), .ZN(n18190) );
  OAI211_X1 U21237 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18214), .A(
        n18325), .B(n18190), .ZN(n18184) );
  NAND3_X1 U21238 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18216), .A3(
        n18184), .ZN(n18185) );
  OAI211_X1 U21239 ( .C1(n18187), .C2(n18189), .A(n18186), .B(n18185), .ZN(
        P3_U2849) );
  NAND2_X1 U21240 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18325), .ZN(
        n18188) );
  AOI22_X1 U21241 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18190), .B1(
        n18189), .B2(n18188), .ZN(n18191) );
  AOI21_X1 U21242 ( .B1(n18241), .B2(n18192), .A(n18191), .ZN(n18194) );
  OAI211_X1 U21243 ( .C1(n18317), .C2(n18195), .A(n18194), .B(n18193), .ZN(
        P3_U2850) );
  AOI22_X1 U21244 ( .A1(n18199), .A2(n18198), .B1(n18197), .B2(n18196), .ZN(
        n18200) );
  NAND2_X1 U21245 ( .A1(n18315), .A2(n18200), .ZN(n18225) );
  OAI221_X1 U21246 ( .B1(n18224), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18224), .C2(n18222), .A(n18201), .ZN(n18202) );
  AOI211_X1 U21247 ( .C1(n18204), .C2(n18203), .A(n18225), .B(n18202), .ZN(
        n18213) );
  OAI21_X1 U21248 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18224), .A(
        n18213), .ZN(n18205) );
  OAI21_X1 U21249 ( .B1(n18206), .B2(n18205), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U21250 ( .A1(n18241), .A2(n18208), .B1(n18221), .B2(n18207), .ZN(
        n18209) );
  OAI221_X1 U21251 ( .B1(n18330), .B2(n18210), .C1(n18216), .C2(n18920), .A(
        n18209), .ZN(P3_U2851) );
  NOR2_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18220), .ZN(
        n18211) );
  AOI22_X1 U21253 ( .A1(n18330), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18221), 
        .B2(n18211), .ZN(n18218) );
  OAI211_X1 U21254 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18214), .A(
        n18213), .B(n18212), .ZN(n18215) );
  NAND3_X1 U21255 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18216), .A3(
        n18215), .ZN(n18217) );
  OAI211_X1 U21256 ( .C1(n18219), .C2(n18229), .A(n18218), .B(n18217), .ZN(
        P3_U2852) );
  AOI22_X1 U21257 ( .A1(n18330), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18221), 
        .B2(n18220), .ZN(n18228) );
  AOI21_X1 U21258 ( .B1(n18224), .B2(n18223), .A(n18222), .ZN(n18226) );
  OAI211_X1 U21259 ( .C1(n18226), .C2(n18225), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18216), .ZN(n18227) );
  OAI211_X1 U21260 ( .C1(n18230), .C2(n18229), .A(n18228), .B(n18227), .ZN(
        P3_U2853) );
  NAND2_X1 U21261 ( .A1(n18315), .A2(n18288), .ZN(n18276) );
  NOR2_X1 U21262 ( .A1(n18234), .A2(n18276), .ZN(n18238) );
  OAI21_X1 U21263 ( .B1(n18295), .B2(n18232), .A(n18231), .ZN(n18233) );
  OAI21_X1 U21264 ( .B1(n18300), .B2(n18835), .A(n18233), .ZN(n18287) );
  NOR2_X1 U21265 ( .A1(n18234), .A2(n18287), .ZN(n18252) );
  OAI21_X1 U21266 ( .B1(n18312), .B2(n18252), .A(n18317), .ZN(n18236) );
  AOI221_X1 U21267 ( .B1(n18238), .B2(n18237), .C1(n18236), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18235), .ZN(n18245) );
  INV_X1 U21268 ( .A(n18239), .ZN(n18240) );
  AOI22_X1 U21269 ( .A1(n18243), .A2(n18242), .B1(n18241), .B2(n18240), .ZN(
        n18244) );
  OAI211_X1 U21270 ( .C1(n18334), .C2(n18246), .A(n18245), .B(n18244), .ZN(
        P3_U2854) );
  AOI21_X1 U21271 ( .B1(n18248), .B2(n18322), .A(n18247), .ZN(n18256) );
  NAND2_X1 U21272 ( .A1(n18315), .A2(n18249), .ZN(n18251) );
  OAI22_X1 U21273 ( .A1(n18252), .A2(n18251), .B1(n18250), .B2(n18317), .ZN(
        n18253) );
  OAI221_X1 U21274 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18254), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18288), .A(n18253), .ZN(
        n18255) );
  OAI211_X1 U21275 ( .C1(n18257), .C2(n18332), .A(n18256), .B(n18255), .ZN(
        P3_U2855) );
  NOR3_X1 U21276 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18259), .A3(
        n18276), .ZN(n18258) );
  AOI21_X1 U21277 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n18330), .A(n18258), .ZN(
        n18263) );
  NOR2_X1 U21278 ( .A1(n18287), .A2(n18259), .ZN(n18260) );
  OAI21_X1 U21279 ( .B1(n18260), .B2(n18312), .A(n18317), .ZN(n18269) );
  AOI22_X1 U21280 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18269), .B1(
        n18322), .B2(n18261), .ZN(n18262) );
  OAI211_X1 U21281 ( .C1(n18332), .C2(n18264), .A(n18263), .B(n18262), .ZN(
        P3_U2856) );
  NOR3_X1 U21282 ( .A1(n18274), .A2(n18291), .A3(n18276), .ZN(n18271) );
  INV_X1 U21283 ( .A(n18265), .ZN(n18267) );
  OAI21_X1 U21284 ( .B1(n18267), .B2(n18334), .A(n18266), .ZN(n18268) );
  AOI221_X1 U21285 ( .B1(n18271), .B2(n18270), .C1(n18269), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18268), .ZN(n18272) );
  OAI21_X1 U21286 ( .B1(n18332), .B2(n18273), .A(n18272), .ZN(P3_U2857) );
  NOR2_X1 U21287 ( .A1(n18291), .A2(n18287), .ZN(n18275) );
  AOI221_X1 U21288 ( .B1(n18312), .B2(n18317), .C1(n18275), .C2(n18317), .A(
        n18274), .ZN(n18278) );
  NOR3_X1 U21289 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18291), .A3(
        n18276), .ZN(n18277) );
  AOI211_X1 U21290 ( .C1(n18279), .C2(n18322), .A(n18278), .B(n18277), .ZN(
        n18281) );
  NAND2_X1 U21291 ( .A1(n18330), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18280) );
  OAI211_X1 U21292 ( .C1(n18282), .C2(n18332), .A(n18281), .B(n18280), .ZN(
        P3_U2858) );
  NOR2_X1 U21293 ( .A1(n18332), .A2(n18283), .ZN(n18284) );
  AOI211_X1 U21294 ( .C1(n18322), .C2(n18286), .A(n18285), .B(n18284), .ZN(
        n18290) );
  OAI221_X1 U21295 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18288), .C1(
        n18291), .C2(n18287), .A(n18325), .ZN(n18289) );
  OAI211_X1 U21296 ( .C1(n18317), .C2(n18291), .A(n18290), .B(n18289), .ZN(
        P3_U2859) );
  OAI21_X1 U21297 ( .B1(n18294), .B2(n18293), .A(n18292), .ZN(n18311) );
  INV_X1 U21298 ( .A(n18295), .ZN(n18297) );
  AOI211_X1 U21299 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18297), .A(
        n18296), .B(n18304), .ZN(n18303) );
  NOR3_X1 U21300 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18987), .A3(
        n18298), .ZN(n18302) );
  AOI21_X1 U21301 ( .B1(n18300), .B2(n18299), .A(n18835), .ZN(n18301) );
  NOR3_X1 U21302 ( .A1(n18303), .A2(n18302), .A3(n18301), .ZN(n18306) );
  OAI22_X1 U21303 ( .A1(n18306), .A2(n18305), .B1(n18304), .B2(n18317), .ZN(
        n18307) );
  AOI21_X1 U21304 ( .B1(n18322), .B2(n18308), .A(n18307), .ZN(n18310) );
  OAI211_X1 U21305 ( .C1(n18332), .C2(n18311), .A(n18310), .B(n18309), .ZN(
        P3_U2860) );
  INV_X1 U21306 ( .A(n18312), .ZN(n18313) );
  NAND2_X1 U21307 ( .A1(n18314), .A2(n18313), .ZN(n18324) );
  NAND2_X1 U21308 ( .A1(n18316), .A2(n18315), .ZN(n18326) );
  OAI21_X1 U21309 ( .B1(n18326), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18317), .ZN(n18318) );
  INV_X1 U21310 ( .A(n18318), .ZN(n18328) );
  OAI22_X1 U21311 ( .A1(n18216), .A2(n19008), .B1(n18332), .B2(n18319), .ZN(
        n18320) );
  AOI21_X1 U21312 ( .B1(n18322), .B2(n18321), .A(n18320), .ZN(n18323) );
  OAI221_X1 U21313 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18324), .C1(
        n18987), .C2(n18328), .A(n18323), .ZN(P3_U2861) );
  NAND2_X1 U21314 ( .A1(n18325), .A2(n18826), .ZN(n18327) );
  AOI22_X1 U21315 ( .A1(n18328), .A2(n18327), .B1(n19003), .B2(n18326), .ZN(
        n18329) );
  AOI21_X1 U21316 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18330), .A(n18329), .ZN(
        n18331) );
  OAI221_X1 U21317 ( .B1(n18335), .B2(n18334), .C1(n18333), .C2(n18332), .A(
        n18331), .ZN(P3_U2862) );
  AOI211_X1 U21318 ( .C1(n18337), .C2(n18336), .A(n18985), .B(n18869), .ZN(
        n18871) );
  OAI21_X1 U21319 ( .B1(n18871), .B2(n18389), .A(n18342), .ZN(n18338) );
  OAI221_X1 U21320 ( .B1(n18845), .B2(n19019), .C1(n18845), .C2(n18342), .A(
        n18338), .ZN(P3_U2863) );
  INV_X1 U21321 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18855) );
  NAND2_X1 U21322 ( .A1(n18852), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18652) );
  INV_X1 U21323 ( .A(n18652), .ZN(n18629) );
  NAND2_X1 U21324 ( .A1(n18855), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18508) );
  INV_X1 U21325 ( .A(n18508), .ZN(n18534) );
  NOR2_X1 U21326 ( .A1(n18629), .A2(n18534), .ZN(n18340) );
  OAI22_X1 U21327 ( .A1(n18341), .A2(n18855), .B1(n18340), .B2(n18339), .ZN(
        P3_U2866) );
  NOR2_X1 U21328 ( .A1(n18856), .A2(n18342), .ZN(P3_U2867) );
  NAND2_X1 U21329 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18532), .ZN(
        n18748) );
  NOR2_X2 U21330 ( .A1(n18845), .A2(n18748), .ZN(n18744) );
  NAND2_X1 U21331 ( .A1(n18847), .A2(n18845), .ZN(n18848) );
  NOR2_X1 U21332 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18439) );
  INV_X1 U21333 ( .A(n18439), .ZN(n18416) );
  NOR2_X1 U21334 ( .A1(n18848), .A2(n18416), .ZN(n18421) );
  NOR2_X1 U21335 ( .A1(n18744), .A2(n18455), .ZN(n18417) );
  OAI21_X1 U21336 ( .B1(n18975), .B2(n18845), .A(n18511), .ZN(n18718) );
  NAND2_X1 U21337 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18678) );
  INV_X1 U21338 ( .A(n18678), .ZN(n18346) );
  NAND2_X1 U21339 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18845), .ZN(
        n18599) );
  NOR2_X1 U21340 ( .A1(n18845), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18484) );
  INV_X1 U21341 ( .A(n18484), .ZN(n18577) );
  NAND2_X1 U21342 ( .A1(n18599), .A2(n18577), .ZN(n18655) );
  NAND2_X1 U21343 ( .A1(n18346), .A2(n18655), .ZN(n18721) );
  OAI22_X1 U21344 ( .A1(n18417), .A2(n18718), .B1(n18680), .B2(n18721), .ZN(
        n18387) );
  AND2_X1 U21345 ( .A1(n18752), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18747) );
  NOR2_X2 U21346 ( .A1(n18678), .A2(n18599), .ZN(n18717) );
  AND2_X1 U21347 ( .A1(n18511), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18746) );
  NOR2_X1 U21348 ( .A1(n18745), .A2(n18417), .ZN(n18382) );
  AOI22_X1 U21349 ( .A1(n18747), .A2(n18717), .B1(n18746), .B2(n18382), .ZN(
        n18348) );
  NOR2_X1 U21350 ( .A1(n18344), .A2(n18343), .ZN(n18383) );
  NAND2_X1 U21351 ( .A1(n18345), .A2(n18383), .ZN(n18756) );
  INV_X1 U21352 ( .A(n18756), .ZN(n18682) );
  NAND2_X1 U21353 ( .A1(n18346), .A2(n18847), .ZN(n18681) );
  NOR2_X1 U21354 ( .A1(n18845), .A2(n18681), .ZN(n18789) );
  CLKBUF_X1 U21355 ( .A(n18789), .Z(n18797) );
  AND2_X1 U21356 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18752), .ZN(n18753) );
  AOI22_X1 U21357 ( .A1(n18455), .A2(n18682), .B1(n18797), .B2(n18753), .ZN(
        n18347) );
  OAI211_X1 U21358 ( .C1(n18349), .C2(n18387), .A(n18348), .B(n18347), .ZN(
        P3_U2868) );
  AND2_X1 U21359 ( .A1(n18752), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18759) );
  AND2_X1 U21360 ( .A1(n18511), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18757) );
  AOI22_X1 U21361 ( .A1(n18717), .A2(n18759), .B1(n18382), .B2(n18757), .ZN(
        n18353) );
  NAND2_X1 U21362 ( .A1(n18350), .A2(n18383), .ZN(n18762) );
  INV_X1 U21363 ( .A(n18762), .ZN(n18686) );
  NOR2_X2 U21364 ( .A1(n18351), .A2(n18680), .ZN(n18758) );
  AOI22_X1 U21365 ( .A1(n18421), .A2(n18686), .B1(n18797), .B2(n18758), .ZN(
        n18352) );
  OAI211_X1 U21366 ( .C1(n18354), .C2(n18387), .A(n18353), .B(n18352), .ZN(
        P3_U2869) );
  AND2_X1 U21367 ( .A1(n18511), .A2(BUF2_REG_2__SCAN_IN), .ZN(n18763) );
  AOI22_X1 U21368 ( .A1(n18797), .A2(n18764), .B1(n18382), .B2(n18763), .ZN(
        n18357) );
  NAND2_X1 U21369 ( .A1(n18355), .A2(n18383), .ZN(n18768) );
  INV_X1 U21370 ( .A(n18768), .ZN(n18690) );
  AND2_X1 U21371 ( .A1(n18752), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18765) );
  AOI22_X1 U21372 ( .A1(n18421), .A2(n18690), .B1(n18717), .B2(n18765), .ZN(
        n18356) );
  OAI211_X1 U21373 ( .C1(n18358), .C2(n18387), .A(n18357), .B(n18356), .ZN(
        P3_U2870) );
  NOR2_X2 U21374 ( .A1(n18359), .A2(n18680), .ZN(n18770) );
  AND2_X1 U21375 ( .A1(n18511), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18769) );
  AOI22_X1 U21376 ( .A1(n18797), .A2(n18770), .B1(n18382), .B2(n18769), .ZN(
        n18362) );
  NAND2_X1 U21377 ( .A1(n18360), .A2(n18383), .ZN(n18774) );
  INV_X1 U21378 ( .A(n18774), .ZN(n18693) );
  AND2_X1 U21379 ( .A1(n18752), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18771) );
  AOI22_X1 U21380 ( .A1(n18421), .A2(n18693), .B1(n18717), .B2(n18771), .ZN(
        n18361) );
  OAI211_X1 U21381 ( .C1(n18363), .C2(n18387), .A(n18362), .B(n18361), .ZN(
        P3_U2871) );
  AND2_X1 U21382 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18752), .ZN(n18777) );
  NOR2_X2 U21383 ( .A1(n18364), .A2(n18653), .ZN(n18775) );
  AOI22_X1 U21384 ( .A1(n18717), .A2(n18777), .B1(n18382), .B2(n18775), .ZN(
        n18367) );
  NAND2_X1 U21385 ( .A1(n18365), .A2(n18383), .ZN(n18780) );
  INV_X1 U21386 ( .A(n18780), .ZN(n18698) );
  AND2_X1 U21387 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18752), .ZN(n18776) );
  AOI22_X1 U21388 ( .A1(n18421), .A2(n18698), .B1(n18797), .B2(n18776), .ZN(
        n18366) );
  OAI211_X1 U21389 ( .C1(n18368), .C2(n18387), .A(n18367), .B(n18366), .ZN(
        P3_U2872) );
  NOR2_X2 U21390 ( .A1(n18369), .A2(n18680), .ZN(n18783) );
  NOR2_X2 U21391 ( .A1(n18370), .A2(n18653), .ZN(n18781) );
  AOI22_X1 U21392 ( .A1(n18797), .A2(n18783), .B1(n18382), .B2(n18781), .ZN(
        n18373) );
  NAND2_X1 U21393 ( .A1(n18371), .A2(n18383), .ZN(n18786) );
  INV_X1 U21394 ( .A(n18786), .ZN(n18702) );
  AND2_X1 U21395 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18752), .ZN(n18782) );
  AOI22_X1 U21396 ( .A1(n18421), .A2(n18702), .B1(n18717), .B2(n18782), .ZN(
        n18372) );
  OAI211_X1 U21397 ( .C1(n18374), .C2(n18387), .A(n18373), .B(n18372), .ZN(
        P3_U2873) );
  AND2_X1 U21398 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18752), .ZN(n18790) );
  NOR2_X2 U21399 ( .A1(n18375), .A2(n18653), .ZN(n18787) );
  AOI22_X1 U21400 ( .A1(n18789), .A2(n18790), .B1(n18382), .B2(n18787), .ZN(
        n18378) );
  NAND2_X1 U21401 ( .A1(n18376), .A2(n18383), .ZN(n18793) );
  INV_X1 U21402 ( .A(n18793), .ZN(n18706) );
  AND2_X1 U21403 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18752), .ZN(n18788) );
  AOI22_X1 U21404 ( .A1(n18421), .A2(n18706), .B1(n18717), .B2(n18788), .ZN(
        n18377) );
  OAI211_X1 U21405 ( .C1(n18379), .C2(n18387), .A(n18378), .B(n18377), .ZN(
        P3_U2874) );
  NOR2_X2 U21406 ( .A1(n18680), .A2(n18380), .ZN(n18799) );
  NOR2_X2 U21407 ( .A1(n18381), .A2(n18653), .ZN(n18795) );
  AOI22_X1 U21408 ( .A1(n18797), .A2(n18799), .B1(n18382), .B2(n18795), .ZN(
        n18386) );
  NAND2_X1 U21409 ( .A1(n18384), .A2(n18383), .ZN(n18803) );
  INV_X1 U21410 ( .A(n18803), .ZN(n18712) );
  AOI22_X1 U21411 ( .A1(n18421), .A2(n18712), .B1(n18717), .B2(n18796), .ZN(
        n18385) );
  OAI211_X1 U21412 ( .C1(n18388), .C2(n18387), .A(n18386), .B(n18385), .ZN(
        P3_U2875) );
  NOR2_X1 U21413 ( .A1(n18389), .A2(n18653), .ZN(n18749) );
  NAND2_X1 U21414 ( .A1(n18749), .A2(n18847), .ZN(n18677) );
  OAI22_X1 U21415 ( .A1(n18680), .A2(n18748), .B1(n18416), .B2(n18677), .ZN(
        n18414) );
  AOI22_X1 U21416 ( .A1(n18744), .A2(n18747), .B1(n18746), .B2(n18411), .ZN(
        n18391) );
  NOR2_X1 U21417 ( .A1(n18577), .A2(n18416), .ZN(n18462) );
  AOI22_X1 U21418 ( .A1(n18753), .A2(n18717), .B1(n18682), .B2(n18478), .ZN(
        n18390) );
  OAI211_X1 U21419 ( .C1(n18392), .C2(n18414), .A(n18391), .B(n18390), .ZN(
        P3_U2876) );
  INV_X1 U21420 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18395) );
  AOI22_X1 U21421 ( .A1(n18717), .A2(n18758), .B1(n18757), .B2(n18411), .ZN(
        n18394) );
  AOI22_X1 U21422 ( .A1(n18744), .A2(n18759), .B1(n18686), .B2(n18478), .ZN(
        n18393) );
  OAI211_X1 U21423 ( .C1(n18395), .C2(n18414), .A(n18394), .B(n18393), .ZN(
        P3_U2877) );
  INV_X1 U21424 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18398) );
  AOI22_X1 U21425 ( .A1(n18744), .A2(n18765), .B1(n18763), .B2(n18411), .ZN(
        n18397) );
  AOI22_X1 U21426 ( .A1(n18717), .A2(n18764), .B1(n18690), .B2(n18478), .ZN(
        n18396) );
  OAI211_X1 U21427 ( .C1(n18398), .C2(n18414), .A(n18397), .B(n18396), .ZN(
        P3_U2878) );
  AOI22_X1 U21428 ( .A1(n18744), .A2(n18771), .B1(n18769), .B2(n18411), .ZN(
        n18400) );
  AOI22_X1 U21429 ( .A1(n18717), .A2(n18770), .B1(n18693), .B2(n18462), .ZN(
        n18399) );
  OAI211_X1 U21430 ( .C1(n18401), .C2(n18414), .A(n18400), .B(n18399), .ZN(
        P3_U2879) );
  AOI22_X1 U21431 ( .A1(n18717), .A2(n18776), .B1(n18775), .B2(n18411), .ZN(
        n18403) );
  AOI22_X1 U21432 ( .A1(n18744), .A2(n18777), .B1(n18698), .B2(n18462), .ZN(
        n18402) );
  OAI211_X1 U21433 ( .C1(n18404), .C2(n18414), .A(n18403), .B(n18402), .ZN(
        P3_U2880) );
  AOI22_X1 U21434 ( .A1(n18744), .A2(n18782), .B1(n18781), .B2(n18411), .ZN(
        n18406) );
  AOI22_X1 U21435 ( .A1(n18717), .A2(n18783), .B1(n18702), .B2(n18462), .ZN(
        n18405) );
  OAI211_X1 U21436 ( .C1(n18407), .C2(n18414), .A(n18406), .B(n18405), .ZN(
        P3_U2881) );
  AOI22_X1 U21437 ( .A1(n18717), .A2(n18790), .B1(n18787), .B2(n18411), .ZN(
        n18409) );
  AOI22_X1 U21438 ( .A1(n18744), .A2(n18788), .B1(n18706), .B2(n18462), .ZN(
        n18408) );
  OAI211_X1 U21439 ( .C1(n18410), .C2(n18414), .A(n18409), .B(n18408), .ZN(
        P3_U2882) );
  AOI22_X1 U21440 ( .A1(n18744), .A2(n18796), .B1(n18795), .B2(n18411), .ZN(
        n18413) );
  AOI22_X1 U21441 ( .A1(n18717), .A2(n18799), .B1(n18712), .B2(n18462), .ZN(
        n18412) );
  OAI211_X1 U21442 ( .C1(n18415), .C2(n18414), .A(n18413), .B(n18412), .ZN(
        P3_U2883) );
  NOR2_X2 U21443 ( .A1(n18599), .A2(n18416), .ZN(n18503) );
  INV_X1 U21444 ( .A(n18503), .ZN(n18438) );
  NOR2_X1 U21445 ( .A1(n18478), .A2(n18503), .ZN(n18460) );
  NOR2_X1 U21446 ( .A1(n18745), .A2(n18460), .ZN(n18434) );
  AOI22_X1 U21447 ( .A1(n18421), .A2(n18747), .B1(n18746), .B2(n18434), .ZN(
        n18420) );
  OAI21_X1 U21448 ( .B1(n18417), .B2(n18720), .A(n18460), .ZN(n18418) );
  OAI211_X1 U21449 ( .C1(n18503), .C2(n18975), .A(n18511), .B(n18418), .ZN(
        n18435) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18435), .B1(
        n18744), .B2(n18753), .ZN(n18419) );
  OAI211_X1 U21451 ( .C1(n18756), .C2(n18438), .A(n18420), .B(n18419), .ZN(
        P3_U2884) );
  AOI22_X1 U21452 ( .A1(n18744), .A2(n18758), .B1(n18757), .B2(n18434), .ZN(
        n18423) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18435), .B1(
        n18421), .B2(n18759), .ZN(n18422) );
  OAI211_X1 U21454 ( .C1(n18762), .C2(n18438), .A(n18423), .B(n18422), .ZN(
        P3_U2885) );
  AOI22_X1 U21455 ( .A1(n18455), .A2(n18765), .B1(n18763), .B2(n18434), .ZN(
        n18425) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18435), .B1(
        n18744), .B2(n18764), .ZN(n18424) );
  OAI211_X1 U21457 ( .C1(n18768), .C2(n18438), .A(n18425), .B(n18424), .ZN(
        P3_U2886) );
  AOI22_X1 U21458 ( .A1(n18744), .A2(n18770), .B1(n18769), .B2(n18434), .ZN(
        n18427) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18435), .B1(
        n18455), .B2(n18771), .ZN(n18426) );
  OAI211_X1 U21460 ( .C1(n18774), .C2(n18438), .A(n18427), .B(n18426), .ZN(
        P3_U2887) );
  AOI22_X1 U21461 ( .A1(n18455), .A2(n18777), .B1(n18775), .B2(n18434), .ZN(
        n18429) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18435), .B1(
        n18744), .B2(n18776), .ZN(n18428) );
  OAI211_X1 U21463 ( .C1(n18780), .C2(n18438), .A(n18429), .B(n18428), .ZN(
        P3_U2888) );
  AOI22_X1 U21464 ( .A1(n18455), .A2(n18782), .B1(n18781), .B2(n18434), .ZN(
        n18431) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18435), .B1(
        n18744), .B2(n18783), .ZN(n18430) );
  OAI211_X1 U21466 ( .C1(n18786), .C2(n18438), .A(n18431), .B(n18430), .ZN(
        P3_U2889) );
  AOI22_X1 U21467 ( .A1(n18455), .A2(n18788), .B1(n18787), .B2(n18434), .ZN(
        n18433) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18435), .B1(
        n18744), .B2(n18790), .ZN(n18432) );
  OAI211_X1 U21469 ( .C1(n18793), .C2(n18438), .A(n18433), .B(n18432), .ZN(
        P3_U2890) );
  AOI22_X1 U21470 ( .A1(n18744), .A2(n18799), .B1(n18795), .B2(n18434), .ZN(
        n18437) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18435), .B1(
        n18455), .B2(n18796), .ZN(n18436) );
  OAI211_X1 U21472 ( .C1(n18803), .C2(n18438), .A(n18437), .B(n18436), .ZN(
        P3_U2891) );
  NAND2_X1 U21473 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18439), .ZN(
        n18483) );
  NOR2_X2 U21474 ( .A1(n18845), .A2(n18483), .ZN(n18527) );
  NOR2_X1 U21475 ( .A1(n18745), .A2(n18483), .ZN(n18454) );
  AOI22_X1 U21476 ( .A1(n18455), .A2(n18753), .B1(n18746), .B2(n18454), .ZN(
        n18441) );
  AOI21_X1 U21477 ( .B1(n18847), .B2(n18720), .A(n18653), .ZN(n18533) );
  OAI211_X1 U21478 ( .C1(n18527), .C2(n18975), .A(n18439), .B(n18533), .ZN(
        n18456) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18456), .B1(
        n18747), .B2(n18478), .ZN(n18440) );
  OAI211_X1 U21480 ( .C1(n18756), .C2(n18459), .A(n18441), .B(n18440), .ZN(
        P3_U2892) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18456), .B1(
        n18757), .B2(n18454), .ZN(n18443) );
  AOI22_X1 U21482 ( .A1(n18455), .A2(n18758), .B1(n18759), .B2(n18462), .ZN(
        n18442) );
  OAI211_X1 U21483 ( .C1(n18762), .C2(n18459), .A(n18443), .B(n18442), .ZN(
        P3_U2893) );
  AOI22_X1 U21484 ( .A1(n18455), .A2(n18764), .B1(n18763), .B2(n18454), .ZN(
        n18445) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18456), .B1(
        n18765), .B2(n18462), .ZN(n18444) );
  OAI211_X1 U21486 ( .C1(n18768), .C2(n18459), .A(n18445), .B(n18444), .ZN(
        P3_U2894) );
  AOI22_X1 U21487 ( .A1(n18771), .A2(n18478), .B1(n18769), .B2(n18454), .ZN(
        n18447) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18456), .B1(
        n18455), .B2(n18770), .ZN(n18446) );
  OAI211_X1 U21489 ( .C1(n18774), .C2(n18459), .A(n18447), .B(n18446), .ZN(
        P3_U2895) );
  AOI22_X1 U21490 ( .A1(n18455), .A2(n18776), .B1(n18775), .B2(n18454), .ZN(
        n18449) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18456), .B1(
        n18777), .B2(n18462), .ZN(n18448) );
  OAI211_X1 U21492 ( .C1(n18780), .C2(n18459), .A(n18449), .B(n18448), .ZN(
        P3_U2896) );
  AOI22_X1 U21493 ( .A1(n18782), .A2(n18478), .B1(n18781), .B2(n18454), .ZN(
        n18451) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18456), .B1(
        n18455), .B2(n18783), .ZN(n18450) );
  OAI211_X1 U21495 ( .C1(n18786), .C2(n18459), .A(n18451), .B(n18450), .ZN(
        P3_U2897) );
  AOI22_X1 U21496 ( .A1(n18455), .A2(n18790), .B1(n18787), .B2(n18454), .ZN(
        n18453) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18456), .B1(
        n18788), .B2(n18462), .ZN(n18452) );
  OAI211_X1 U21498 ( .C1(n18793), .C2(n18459), .A(n18453), .B(n18452), .ZN(
        P3_U2898) );
  AOI22_X1 U21499 ( .A1(n18455), .A2(n18799), .B1(n18795), .B2(n18454), .ZN(
        n18458) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18456), .B1(
        n18796), .B2(n18478), .ZN(n18457) );
  OAI211_X1 U21501 ( .C1(n18803), .C2(n18459), .A(n18458), .B(n18457), .ZN(
        P3_U2899) );
  NOR2_X2 U21502 ( .A1(n18848), .A2(n18508), .ZN(n18550) );
  AOI21_X1 U21503 ( .B1(n18459), .B2(n18482), .A(n18745), .ZN(n18477) );
  AOI22_X1 U21504 ( .A1(n18747), .A2(n18503), .B1(n18746), .B2(n18477), .ZN(
        n18464) );
  AOI221_X1 U21505 ( .B1(n18460), .B2(n18459), .C1(n18720), .C2(n18459), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18461) );
  OAI21_X1 U21506 ( .B1(n18550), .B2(n18461), .A(n18511), .ZN(n18479) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18479), .B1(
        n18753), .B2(n18462), .ZN(n18463) );
  OAI211_X1 U21508 ( .C1(n18756), .C2(n18482), .A(n18464), .B(n18463), .ZN(
        P3_U2900) );
  AOI22_X1 U21509 ( .A1(n18758), .A2(n18478), .B1(n18757), .B2(n18477), .ZN(
        n18466) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18479), .B1(
        n18759), .B2(n18503), .ZN(n18465) );
  OAI211_X1 U21511 ( .C1(n18762), .C2(n18482), .A(n18466), .B(n18465), .ZN(
        P3_U2901) );
  AOI22_X1 U21512 ( .A1(n18765), .A2(n18503), .B1(n18763), .B2(n18477), .ZN(
        n18468) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18479), .B1(
        n18764), .B2(n18478), .ZN(n18467) );
  OAI211_X1 U21514 ( .C1(n18768), .C2(n18482), .A(n18468), .B(n18467), .ZN(
        P3_U2902) );
  AOI22_X1 U21515 ( .A1(n18771), .A2(n18503), .B1(n18769), .B2(n18477), .ZN(
        n18470) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18479), .B1(
        n18770), .B2(n18478), .ZN(n18469) );
  OAI211_X1 U21517 ( .C1(n18774), .C2(n18482), .A(n18470), .B(n18469), .ZN(
        P3_U2903) );
  AOI22_X1 U21518 ( .A1(n18776), .A2(n18478), .B1(n18775), .B2(n18477), .ZN(
        n18472) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18479), .B1(
        n18777), .B2(n18503), .ZN(n18471) );
  OAI211_X1 U21520 ( .C1(n18780), .C2(n18482), .A(n18472), .B(n18471), .ZN(
        P3_U2904) );
  AOI22_X1 U21521 ( .A1(n18783), .A2(n18478), .B1(n18781), .B2(n18477), .ZN(
        n18474) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18479), .B1(
        n18782), .B2(n18503), .ZN(n18473) );
  OAI211_X1 U21523 ( .C1(n18786), .C2(n18482), .A(n18474), .B(n18473), .ZN(
        P3_U2905) );
  AOI22_X1 U21524 ( .A1(n18790), .A2(n18478), .B1(n18787), .B2(n18477), .ZN(
        n18476) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18479), .B1(
        n18788), .B2(n18503), .ZN(n18475) );
  OAI211_X1 U21526 ( .C1(n18793), .C2(n18482), .A(n18476), .B(n18475), .ZN(
        P3_U2906) );
  AOI22_X1 U21527 ( .A1(n18799), .A2(n18478), .B1(n18795), .B2(n18477), .ZN(
        n18481) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18479), .B1(
        n18796), .B2(n18503), .ZN(n18480) );
  OAI211_X1 U21529 ( .C1(n18803), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2907) );
  OAI22_X1 U21530 ( .A1(n18680), .A2(n18483), .B1(n18508), .B2(n18677), .ZN(
        n18506) );
  AOI22_X1 U21531 ( .A1(n18747), .A2(n18527), .B1(n18746), .B2(n18502), .ZN(
        n18486) );
  NAND2_X1 U21532 ( .A1(n18534), .A2(n18484), .ZN(n18501) );
  AOI22_X1 U21533 ( .A1(n18753), .A2(n18503), .B1(n18682), .B2(n18572), .ZN(
        n18485) );
  OAI211_X1 U21534 ( .C1(n18487), .C2(n18506), .A(n18486), .B(n18485), .ZN(
        P3_U2908) );
  AOI22_X1 U21535 ( .A1(n18757), .A2(n18502), .B1(n18759), .B2(n18527), .ZN(
        n18489) );
  INV_X1 U21536 ( .A(n18506), .ZN(n18498) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18498), .B1(
        n18758), .B2(n18503), .ZN(n18488) );
  OAI211_X1 U21538 ( .C1(n18762), .C2(n18501), .A(n18489), .B(n18488), .ZN(
        P3_U2909) );
  AOI22_X1 U21539 ( .A1(n18764), .A2(n18503), .B1(n18763), .B2(n18502), .ZN(
        n18491) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18498), .B1(
        n18765), .B2(n18527), .ZN(n18490) );
  OAI211_X1 U21541 ( .C1(n18768), .C2(n18501), .A(n18491), .B(n18490), .ZN(
        P3_U2910) );
  AOI22_X1 U21542 ( .A1(n18771), .A2(n18527), .B1(n18769), .B2(n18502), .ZN(
        n18493) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18498), .B1(
        n18770), .B2(n18503), .ZN(n18492) );
  OAI211_X1 U21544 ( .C1(n18774), .C2(n18501), .A(n18493), .B(n18492), .ZN(
        P3_U2911) );
  AOI22_X1 U21545 ( .A1(n18777), .A2(n18527), .B1(n18775), .B2(n18502), .ZN(
        n18495) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18498), .B1(
        n18776), .B2(n18503), .ZN(n18494) );
  OAI211_X1 U21547 ( .C1(n18780), .C2(n18501), .A(n18495), .B(n18494), .ZN(
        P3_U2912) );
  AOI22_X1 U21548 ( .A1(n18782), .A2(n18527), .B1(n18781), .B2(n18502), .ZN(
        n18497) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18498), .B1(
        n18783), .B2(n18503), .ZN(n18496) );
  OAI211_X1 U21550 ( .C1(n18786), .C2(n18501), .A(n18497), .B(n18496), .ZN(
        P3_U2913) );
  AOI22_X1 U21551 ( .A1(n18788), .A2(n18527), .B1(n18787), .B2(n18502), .ZN(
        n18500) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18498), .B1(
        n18790), .B2(n18503), .ZN(n18499) );
  OAI211_X1 U21553 ( .C1(n18793), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        P3_U2914) );
  AOI22_X1 U21554 ( .A1(n18799), .A2(n18503), .B1(n18795), .B2(n18502), .ZN(
        n18505) );
  AOI22_X1 U21555 ( .A1(n18796), .A2(n18527), .B1(n18712), .B2(n18572), .ZN(
        n18504) );
  OAI211_X1 U21556 ( .C1(n18507), .C2(n18506), .A(n18505), .B(n18504), .ZN(
        P3_U2915) );
  NOR2_X2 U21557 ( .A1(n18508), .A2(n18599), .ZN(n18595) );
  INV_X1 U21558 ( .A(n18595), .ZN(n18531) );
  NOR2_X1 U21559 ( .A1(n18572), .A2(n18595), .ZN(n18555) );
  NOR2_X1 U21560 ( .A1(n18745), .A2(n18555), .ZN(n18526) );
  AOI22_X1 U21561 ( .A1(n18753), .A2(n18527), .B1(n18746), .B2(n18526), .ZN(
        n18513) );
  NOR2_X1 U21562 ( .A1(n18527), .A2(n18550), .ZN(n18509) );
  OAI21_X1 U21563 ( .B1(n18509), .B2(n18720), .A(n18555), .ZN(n18510) );
  OAI211_X1 U21564 ( .C1(n18595), .C2(n18975), .A(n18511), .B(n18510), .ZN(
        n18528) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18528), .B1(
        n18747), .B2(n18550), .ZN(n18512) );
  OAI211_X1 U21566 ( .C1(n18756), .C2(n18531), .A(n18513), .B(n18512), .ZN(
        P3_U2916) );
  AOI22_X1 U21567 ( .A1(n18758), .A2(n18527), .B1(n18757), .B2(n18526), .ZN(
        n18515) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18528), .B1(
        n18759), .B2(n18550), .ZN(n18514) );
  OAI211_X1 U21569 ( .C1(n18762), .C2(n18531), .A(n18515), .B(n18514), .ZN(
        P3_U2917) );
  AOI22_X1 U21570 ( .A1(n18765), .A2(n18550), .B1(n18763), .B2(n18526), .ZN(
        n18517) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18528), .B1(
        n18764), .B2(n18527), .ZN(n18516) );
  OAI211_X1 U21572 ( .C1(n18768), .C2(n18531), .A(n18517), .B(n18516), .ZN(
        P3_U2918) );
  AOI22_X1 U21573 ( .A1(n18770), .A2(n18527), .B1(n18769), .B2(n18526), .ZN(
        n18519) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18528), .B1(
        n18771), .B2(n18550), .ZN(n18518) );
  OAI211_X1 U21575 ( .C1(n18774), .C2(n18531), .A(n18519), .B(n18518), .ZN(
        P3_U2919) );
  AOI22_X1 U21576 ( .A1(n18776), .A2(n18527), .B1(n18775), .B2(n18526), .ZN(
        n18521) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18528), .B1(
        n18777), .B2(n18550), .ZN(n18520) );
  OAI211_X1 U21578 ( .C1(n18780), .C2(n18531), .A(n18521), .B(n18520), .ZN(
        P3_U2920) );
  AOI22_X1 U21579 ( .A1(n18782), .A2(n18550), .B1(n18781), .B2(n18526), .ZN(
        n18523) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18528), .B1(
        n18783), .B2(n18527), .ZN(n18522) );
  OAI211_X1 U21581 ( .C1(n18786), .C2(n18531), .A(n18523), .B(n18522), .ZN(
        P3_U2921) );
  AOI22_X1 U21582 ( .A1(n18790), .A2(n18527), .B1(n18787), .B2(n18526), .ZN(
        n18525) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18528), .B1(
        n18788), .B2(n18550), .ZN(n18524) );
  OAI211_X1 U21584 ( .C1(n18793), .C2(n18531), .A(n18525), .B(n18524), .ZN(
        P3_U2922) );
  AOI22_X1 U21585 ( .A1(n18796), .A2(n18550), .B1(n18795), .B2(n18526), .ZN(
        n18530) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18528), .B1(
        n18799), .B2(n18527), .ZN(n18529) );
  OAI211_X1 U21587 ( .C1(n18803), .C2(n18531), .A(n18530), .B(n18529), .ZN(
        P3_U2923) );
  NAND2_X1 U21588 ( .A1(n18855), .A2(n18532), .ZN(n18578) );
  NOR2_X2 U21589 ( .A1(n18845), .A2(n18578), .ZN(n18624) );
  INV_X1 U21590 ( .A(n18624), .ZN(n18554) );
  OAI211_X1 U21591 ( .C1(n18624), .C2(n18975), .A(n18534), .B(n18533), .ZN(
        n18551) );
  NOR2_X1 U21592 ( .A1(n18745), .A2(n18578), .ZN(n18549) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18551), .B1(
        n18746), .B2(n18549), .ZN(n18536) );
  AOI22_X1 U21594 ( .A1(n18753), .A2(n18550), .B1(n18747), .B2(n18572), .ZN(
        n18535) );
  OAI211_X1 U21595 ( .C1(n18756), .C2(n18554), .A(n18536), .B(n18535), .ZN(
        P3_U2924) );
  AOI22_X1 U21596 ( .A1(n18758), .A2(n18550), .B1(n18757), .B2(n18549), .ZN(
        n18538) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18551), .B1(
        n18759), .B2(n18572), .ZN(n18537) );
  OAI211_X1 U21598 ( .C1(n18762), .C2(n18554), .A(n18538), .B(n18537), .ZN(
        P3_U2925) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18551), .B1(
        n18763), .B2(n18549), .ZN(n18540) );
  AOI22_X1 U21600 ( .A1(n18765), .A2(n18572), .B1(n18764), .B2(n18550), .ZN(
        n18539) );
  OAI211_X1 U21601 ( .C1(n18768), .C2(n18554), .A(n18540), .B(n18539), .ZN(
        P3_U2926) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18551), .B1(
        n18769), .B2(n18549), .ZN(n18542) );
  AOI22_X1 U21603 ( .A1(n18771), .A2(n18572), .B1(n18770), .B2(n18550), .ZN(
        n18541) );
  OAI211_X1 U21604 ( .C1(n18774), .C2(n18554), .A(n18542), .B(n18541), .ZN(
        P3_U2927) );
  AOI22_X1 U21605 ( .A1(n18776), .A2(n18550), .B1(n18775), .B2(n18549), .ZN(
        n18544) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18551), .B1(
        n18777), .B2(n18572), .ZN(n18543) );
  OAI211_X1 U21607 ( .C1(n18780), .C2(n18554), .A(n18544), .B(n18543), .ZN(
        P3_U2928) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18551), .B1(
        n18781), .B2(n18549), .ZN(n18546) );
  AOI22_X1 U21609 ( .A1(n18782), .A2(n18572), .B1(n18783), .B2(n18550), .ZN(
        n18545) );
  OAI211_X1 U21610 ( .C1(n18786), .C2(n18554), .A(n18546), .B(n18545), .ZN(
        P3_U2929) );
  AOI22_X1 U21611 ( .A1(n18788), .A2(n18572), .B1(n18787), .B2(n18549), .ZN(
        n18548) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18551), .B1(
        n18790), .B2(n18550), .ZN(n18547) );
  OAI211_X1 U21613 ( .C1(n18793), .C2(n18554), .A(n18548), .B(n18547), .ZN(
        P3_U2930) );
  AOI22_X1 U21614 ( .A1(n18796), .A2(n18572), .B1(n18795), .B2(n18549), .ZN(
        n18553) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18551), .B1(
        n18799), .B2(n18550), .ZN(n18552) );
  OAI211_X1 U21616 ( .C1(n18803), .C2(n18554), .A(n18553), .B(n18552), .ZN(
        P3_U2931) );
  NOR2_X2 U21617 ( .A1(n18848), .A2(n18652), .ZN(n18647) );
  INV_X1 U21618 ( .A(n18647), .ZN(n18576) );
  NOR2_X1 U21619 ( .A1(n18624), .A2(n18647), .ZN(n18601) );
  NOR2_X1 U21620 ( .A1(n18745), .A2(n18601), .ZN(n18571) );
  AOI22_X1 U21621 ( .A1(n18747), .A2(n18595), .B1(n18746), .B2(n18571), .ZN(
        n18558) );
  OAI22_X1 U21622 ( .A1(n18555), .A2(n18680), .B1(n18601), .B2(n18653), .ZN(
        n18556) );
  OAI21_X1 U21623 ( .B1(n18647), .B2(n18975), .A(n18556), .ZN(n18573) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18573), .B1(
        n18753), .B2(n18572), .ZN(n18557) );
  OAI211_X1 U21625 ( .C1(n18756), .C2(n18576), .A(n18558), .B(n18557), .ZN(
        P3_U2932) );
  AOI22_X1 U21626 ( .A1(n18757), .A2(n18571), .B1(n18759), .B2(n18595), .ZN(
        n18560) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18573), .B1(
        n18758), .B2(n18572), .ZN(n18559) );
  OAI211_X1 U21628 ( .C1(n18762), .C2(n18576), .A(n18560), .B(n18559), .ZN(
        P3_U2933) );
  AOI22_X1 U21629 ( .A1(n18765), .A2(n18595), .B1(n18763), .B2(n18571), .ZN(
        n18562) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18573), .B1(
        n18764), .B2(n18572), .ZN(n18561) );
  OAI211_X1 U21631 ( .C1(n18768), .C2(n18576), .A(n18562), .B(n18561), .ZN(
        P3_U2934) );
  AOI22_X1 U21632 ( .A1(n18770), .A2(n18572), .B1(n18769), .B2(n18571), .ZN(
        n18564) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18573), .B1(
        n18771), .B2(n18595), .ZN(n18563) );
  OAI211_X1 U21634 ( .C1(n18774), .C2(n18576), .A(n18564), .B(n18563), .ZN(
        P3_U2935) );
  AOI22_X1 U21635 ( .A1(n18777), .A2(n18595), .B1(n18775), .B2(n18571), .ZN(
        n18566) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18573), .B1(
        n18776), .B2(n18572), .ZN(n18565) );
  OAI211_X1 U21637 ( .C1(n18780), .C2(n18576), .A(n18566), .B(n18565), .ZN(
        P3_U2936) );
  AOI22_X1 U21638 ( .A1(n18782), .A2(n18595), .B1(n18781), .B2(n18571), .ZN(
        n18568) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18573), .B1(
        n18783), .B2(n18572), .ZN(n18567) );
  OAI211_X1 U21640 ( .C1(n18786), .C2(n18576), .A(n18568), .B(n18567), .ZN(
        P3_U2937) );
  AOI22_X1 U21641 ( .A1(n18788), .A2(n18595), .B1(n18787), .B2(n18571), .ZN(
        n18570) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18573), .B1(
        n18790), .B2(n18572), .ZN(n18569) );
  OAI211_X1 U21643 ( .C1(n18793), .C2(n18576), .A(n18570), .B(n18569), .ZN(
        P3_U2938) );
  AOI22_X1 U21644 ( .A1(n18799), .A2(n18572), .B1(n18795), .B2(n18571), .ZN(
        n18575) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18573), .B1(
        n18796), .B2(n18595), .ZN(n18574) );
  OAI211_X1 U21646 ( .C1(n18803), .C2(n18576), .A(n18575), .B(n18574), .ZN(
        P3_U2939) );
  NOR2_X2 U21647 ( .A1(n18652), .A2(n18577), .ZN(n18673) );
  AOI22_X1 U21648 ( .A1(n18747), .A2(n18624), .B1(n18746), .B2(n18594), .ZN(
        n18581) );
  INV_X1 U21649 ( .A(n18578), .ZN(n18579) );
  NOR2_X1 U21650 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18652), .ZN(
        n18631) );
  AOI22_X1 U21651 ( .A1(n18752), .A2(n18579), .B1(n18749), .B2(n18631), .ZN(
        n18596) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18596), .B1(
        n18753), .B2(n18595), .ZN(n18580) );
  OAI211_X1 U21653 ( .C1(n18756), .C2(n18602), .A(n18581), .B(n18580), .ZN(
        P3_U2940) );
  AOI22_X1 U21654 ( .A1(n18758), .A2(n18595), .B1(n18757), .B2(n18594), .ZN(
        n18583) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18596), .B1(
        n18759), .B2(n18624), .ZN(n18582) );
  OAI211_X1 U21656 ( .C1(n18762), .C2(n18602), .A(n18583), .B(n18582), .ZN(
        P3_U2941) );
  AOI22_X1 U21657 ( .A1(n18764), .A2(n18595), .B1(n18763), .B2(n18594), .ZN(
        n18585) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18596), .B1(
        n18765), .B2(n18624), .ZN(n18584) );
  OAI211_X1 U21659 ( .C1(n18768), .C2(n18602), .A(n18585), .B(n18584), .ZN(
        P3_U2942) );
  AOI22_X1 U21660 ( .A1(n18770), .A2(n18595), .B1(n18769), .B2(n18594), .ZN(
        n18587) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18596), .B1(
        n18771), .B2(n18624), .ZN(n18586) );
  OAI211_X1 U21662 ( .C1(n18774), .C2(n18602), .A(n18587), .B(n18586), .ZN(
        P3_U2943) );
  AOI22_X1 U21663 ( .A1(n18777), .A2(n18624), .B1(n18775), .B2(n18594), .ZN(
        n18589) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18596), .B1(
        n18776), .B2(n18595), .ZN(n18588) );
  OAI211_X1 U21665 ( .C1(n18780), .C2(n18602), .A(n18589), .B(n18588), .ZN(
        P3_U2944) );
  AOI22_X1 U21666 ( .A1(n18783), .A2(n18595), .B1(n18781), .B2(n18594), .ZN(
        n18591) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18596), .B1(
        n18782), .B2(n18624), .ZN(n18590) );
  OAI211_X1 U21668 ( .C1(n18786), .C2(n18602), .A(n18591), .B(n18590), .ZN(
        P3_U2945) );
  AOI22_X1 U21669 ( .A1(n18790), .A2(n18595), .B1(n18787), .B2(n18594), .ZN(
        n18593) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18596), .B1(
        n18788), .B2(n18624), .ZN(n18592) );
  OAI211_X1 U21671 ( .C1(n18793), .C2(n18602), .A(n18593), .B(n18592), .ZN(
        P3_U2946) );
  AOI22_X1 U21672 ( .A1(n18799), .A2(n18595), .B1(n18795), .B2(n18594), .ZN(
        n18598) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18596), .B1(
        n18796), .B2(n18624), .ZN(n18597) );
  OAI211_X1 U21674 ( .C1(n18803), .C2(n18602), .A(n18598), .B(n18597), .ZN(
        P3_U2947) );
  NOR2_X1 U21675 ( .A1(n18652), .A2(n18599), .ZN(n18711) );
  NOR2_X1 U21676 ( .A1(n18673), .A2(n18697), .ZN(n18600) );
  AOI221_X1 U21677 ( .B1(n18601), .B2(n18600), .C1(n18720), .C2(n18600), .A(
        n18718), .ZN(n18628) );
  INV_X1 U21678 ( .A(n18711), .ZN(n18619) );
  AOI21_X1 U21679 ( .B1(n18602), .B2(n18619), .A(n18745), .ZN(n18623) );
  AOI22_X1 U21680 ( .A1(n18753), .A2(n18624), .B1(n18746), .B2(n18623), .ZN(
        n18604) );
  AOI22_X1 U21681 ( .A1(n18682), .A2(n18697), .B1(n18747), .B2(n18647), .ZN(
        n18603) );
  OAI211_X1 U21682 ( .C1(n18628), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2948) );
  AOI22_X1 U21683 ( .A1(n18758), .A2(n18624), .B1(n18757), .B2(n18623), .ZN(
        n18607) );
  AOI22_X1 U21684 ( .A1(n18686), .A2(n18697), .B1(n18759), .B2(n18647), .ZN(
        n18606) );
  OAI211_X1 U21685 ( .C1(n18628), .C2(n18608), .A(n18607), .B(n18606), .ZN(
        P3_U2949) );
  AOI22_X1 U21686 ( .A1(n18764), .A2(n18624), .B1(n18763), .B2(n18623), .ZN(
        n18610) );
  INV_X1 U21687 ( .A(n18628), .ZN(n18616) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18616), .B1(
        n18765), .B2(n18647), .ZN(n18609) );
  OAI211_X1 U21689 ( .C1(n18768), .C2(n18619), .A(n18610), .B(n18609), .ZN(
        P3_U2950) );
  AOI22_X1 U21690 ( .A1(n18770), .A2(n18624), .B1(n18769), .B2(n18623), .ZN(
        n18612) );
  AOI22_X1 U21691 ( .A1(n18771), .A2(n18647), .B1(n18693), .B2(n18697), .ZN(
        n18611) );
  OAI211_X1 U21692 ( .C1(n18628), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P3_U2951) );
  AOI22_X1 U21693 ( .A1(n18777), .A2(n18647), .B1(n18775), .B2(n18623), .ZN(
        n18615) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18616), .B1(
        n18776), .B2(n18624), .ZN(n18614) );
  OAI211_X1 U21695 ( .C1(n18780), .C2(n18619), .A(n18615), .B(n18614), .ZN(
        P3_U2952) );
  AOI22_X1 U21696 ( .A1(n18782), .A2(n18647), .B1(n18781), .B2(n18623), .ZN(
        n18618) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18616), .B1(
        n18783), .B2(n18624), .ZN(n18617) );
  OAI211_X1 U21698 ( .C1(n18786), .C2(n18619), .A(n18618), .B(n18617), .ZN(
        P3_U2953) );
  AOI22_X1 U21699 ( .A1(n18790), .A2(n18624), .B1(n18787), .B2(n18623), .ZN(
        n18621) );
  AOI22_X1 U21700 ( .A1(n18788), .A2(n18647), .B1(n18706), .B2(n18711), .ZN(
        n18620) );
  OAI211_X1 U21701 ( .C1(n18628), .C2(n18622), .A(n18621), .B(n18620), .ZN(
        P3_U2954) );
  AOI22_X1 U21702 ( .A1(n18799), .A2(n18624), .B1(n18795), .B2(n18623), .ZN(
        n18626) );
  AOI22_X1 U21703 ( .A1(n18796), .A2(n18647), .B1(n18712), .B2(n18711), .ZN(
        n18625) );
  OAI211_X1 U21704 ( .C1(n18628), .C2(n18627), .A(n18626), .B(n18625), .ZN(
        P3_U2955) );
  NAND2_X1 U21705 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18629), .ZN(
        n18679) );
  NOR2_X2 U21706 ( .A1(n18845), .A2(n18679), .ZN(n18739) );
  NOR2_X1 U21707 ( .A1(n18745), .A2(n18679), .ZN(n18646) );
  AOI22_X1 U21708 ( .A1(n18753), .A2(n18647), .B1(n18746), .B2(n18646), .ZN(
        n18633) );
  INV_X1 U21709 ( .A(n18679), .ZN(n18630) );
  AOI22_X1 U21710 ( .A1(n18752), .A2(n18631), .B1(n18749), .B2(n18630), .ZN(
        n18648) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18648), .B1(
        n18747), .B2(n18673), .ZN(n18632) );
  OAI211_X1 U21712 ( .C1(n18756), .C2(n18651), .A(n18633), .B(n18632), .ZN(
        P3_U2956) );
  AOI22_X1 U21713 ( .A1(n18757), .A2(n18646), .B1(n18759), .B2(n18673), .ZN(
        n18635) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18648), .B1(
        n18758), .B2(n18647), .ZN(n18634) );
  OAI211_X1 U21715 ( .C1(n18762), .C2(n18651), .A(n18635), .B(n18634), .ZN(
        P3_U2957) );
  AOI22_X1 U21716 ( .A1(n18764), .A2(n18647), .B1(n18763), .B2(n18646), .ZN(
        n18637) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18648), .B1(
        n18765), .B2(n18673), .ZN(n18636) );
  OAI211_X1 U21718 ( .C1(n18768), .C2(n18651), .A(n18637), .B(n18636), .ZN(
        P3_U2958) );
  AOI22_X1 U21719 ( .A1(n18770), .A2(n18647), .B1(n18769), .B2(n18646), .ZN(
        n18639) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18648), .B1(
        n18771), .B2(n18673), .ZN(n18638) );
  OAI211_X1 U21721 ( .C1(n18774), .C2(n18651), .A(n18639), .B(n18638), .ZN(
        P3_U2959) );
  AOI22_X1 U21722 ( .A1(n18777), .A2(n18673), .B1(n18775), .B2(n18646), .ZN(
        n18641) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18648), .B1(
        n18776), .B2(n18647), .ZN(n18640) );
  OAI211_X1 U21724 ( .C1(n18780), .C2(n18651), .A(n18641), .B(n18640), .ZN(
        P3_U2960) );
  AOI22_X1 U21725 ( .A1(n18783), .A2(n18647), .B1(n18781), .B2(n18646), .ZN(
        n18643) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18648), .B1(
        n18782), .B2(n18673), .ZN(n18642) );
  OAI211_X1 U21727 ( .C1(n18786), .C2(n18651), .A(n18643), .B(n18642), .ZN(
        P3_U2961) );
  AOI22_X1 U21728 ( .A1(n18788), .A2(n18673), .B1(n18787), .B2(n18646), .ZN(
        n18645) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18648), .B1(
        n18790), .B2(n18647), .ZN(n18644) );
  OAI211_X1 U21730 ( .C1(n18793), .C2(n18651), .A(n18645), .B(n18644), .ZN(
        P3_U2962) );
  AOI22_X1 U21731 ( .A1(n18796), .A2(n18673), .B1(n18795), .B2(n18646), .ZN(
        n18650) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18648), .B1(
        n18799), .B2(n18647), .ZN(n18649) );
  OAI211_X1 U21733 ( .C1(n18803), .C2(n18651), .A(n18650), .B(n18649), .ZN(
        P3_U2963) );
  INV_X1 U21734 ( .A(n18681), .ZN(n18751) );
  NAND2_X1 U21735 ( .A1(n18751), .A2(n18845), .ZN(n18723) );
  NAND2_X1 U21736 ( .A1(n18651), .A2(n18723), .ZN(n18657) );
  INV_X1 U21737 ( .A(n18657), .ZN(n18719) );
  NOR2_X1 U21738 ( .A1(n18745), .A2(n18719), .ZN(n18672) );
  AOI22_X1 U21739 ( .A1(n18747), .A2(n18711), .B1(n18746), .B2(n18672), .ZN(
        n18659) );
  NOR2_X1 U21740 ( .A1(n18720), .A2(n18652), .ZN(n18656) );
  AOI21_X1 U21741 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18723), .A(n18653), 
        .ZN(n18654) );
  OAI221_X1 U21742 ( .B1(n18657), .B2(n18656), .C1(n18657), .C2(n18655), .A(
        n18654), .ZN(n18674) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18674), .B1(
        n18753), .B2(n18673), .ZN(n18658) );
  OAI211_X1 U21744 ( .C1(n18756), .C2(n18723), .A(n18659), .B(n18658), .ZN(
        P3_U2964) );
  AOI22_X1 U21745 ( .A1(n18758), .A2(n18673), .B1(n18757), .B2(n18672), .ZN(
        n18661) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18674), .B1(
        n18759), .B2(n18697), .ZN(n18660) );
  OAI211_X1 U21747 ( .C1(n18762), .C2(n18723), .A(n18661), .B(n18660), .ZN(
        P3_U2965) );
  AOI22_X1 U21748 ( .A1(n18764), .A2(n18673), .B1(n18763), .B2(n18672), .ZN(
        n18663) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18674), .B1(
        n18765), .B2(n18711), .ZN(n18662) );
  OAI211_X1 U21750 ( .C1(n18768), .C2(n18723), .A(n18663), .B(n18662), .ZN(
        P3_U2966) );
  AOI22_X1 U21751 ( .A1(n18770), .A2(n18673), .B1(n18769), .B2(n18672), .ZN(
        n18665) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18674), .B1(
        n18771), .B2(n18697), .ZN(n18664) );
  OAI211_X1 U21753 ( .C1(n18774), .C2(n18723), .A(n18665), .B(n18664), .ZN(
        P3_U2967) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18674), .B1(
        n18775), .B2(n18672), .ZN(n18667) );
  AOI22_X1 U21755 ( .A1(n18776), .A2(n18673), .B1(n18777), .B2(n18697), .ZN(
        n18666) );
  OAI211_X1 U21756 ( .C1(n18780), .C2(n18723), .A(n18667), .B(n18666), .ZN(
        P3_U2968) );
  AOI22_X1 U21757 ( .A1(n18782), .A2(n18697), .B1(n18781), .B2(n18672), .ZN(
        n18669) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18674), .B1(
        n18783), .B2(n18673), .ZN(n18668) );
  OAI211_X1 U21759 ( .C1(n18786), .C2(n18723), .A(n18669), .B(n18668), .ZN(
        P3_U2969) );
  AOI22_X1 U21760 ( .A1(n18790), .A2(n18673), .B1(n18787), .B2(n18672), .ZN(
        n18671) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18674), .B1(
        n18788), .B2(n18711), .ZN(n18670) );
  OAI211_X1 U21762 ( .C1(n18793), .C2(n18723), .A(n18671), .B(n18670), .ZN(
        P3_U2970) );
  AOI22_X1 U21763 ( .A1(n18799), .A2(n18673), .B1(n18795), .B2(n18672), .ZN(
        n18676) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18674), .B1(
        n18796), .B2(n18697), .ZN(n18675) );
  OAI211_X1 U21765 ( .C1(n18803), .C2(n18723), .A(n18676), .B(n18675), .ZN(
        P3_U2971) );
  OAI22_X1 U21766 ( .A1(n18680), .A2(n18679), .B1(n18678), .B2(n18677), .ZN(
        n18715) );
  NOR2_X1 U21767 ( .A1(n18745), .A2(n18681), .ZN(n18710) );
  AOI22_X1 U21768 ( .A1(n18753), .A2(n18697), .B1(n18746), .B2(n18710), .ZN(
        n18684) );
  AOI22_X1 U21769 ( .A1(n18789), .A2(n18682), .B1(n18747), .B2(n18739), .ZN(
        n18683) );
  OAI211_X1 U21770 ( .C1(n18685), .C2(n18715), .A(n18684), .B(n18683), .ZN(
        P3_U2972) );
  INV_X1 U21771 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18689) );
  AOI22_X1 U21772 ( .A1(n18758), .A2(n18697), .B1(n18757), .B2(n18710), .ZN(
        n18688) );
  AOI22_X1 U21773 ( .A1(n18789), .A2(n18686), .B1(n18759), .B2(n18739), .ZN(
        n18687) );
  OAI211_X1 U21774 ( .C1(n18689), .C2(n18715), .A(n18688), .B(n18687), .ZN(
        P3_U2973) );
  AOI22_X1 U21775 ( .A1(n18765), .A2(n18739), .B1(n18763), .B2(n18710), .ZN(
        n18692) );
  AOI22_X1 U21776 ( .A1(n18789), .A2(n18690), .B1(n18764), .B2(n18711), .ZN(
        n18691) );
  OAI211_X1 U21777 ( .C1(n10402), .C2(n18715), .A(n18692), .B(n18691), .ZN(
        P3_U2974) );
  AOI22_X1 U21778 ( .A1(n18771), .A2(n18739), .B1(n18769), .B2(n18710), .ZN(
        n18695) );
  AOI22_X1 U21779 ( .A1(n18789), .A2(n18693), .B1(n18770), .B2(n18711), .ZN(
        n18694) );
  OAI211_X1 U21780 ( .C1(n18696), .C2(n18715), .A(n18695), .B(n18694), .ZN(
        P3_U2975) );
  AOI22_X1 U21781 ( .A1(n18776), .A2(n18697), .B1(n18775), .B2(n18710), .ZN(
        n18700) );
  AOI22_X1 U21782 ( .A1(n18789), .A2(n18698), .B1(n18777), .B2(n18739), .ZN(
        n18699) );
  OAI211_X1 U21783 ( .C1(n18701), .C2(n18715), .A(n18700), .B(n18699), .ZN(
        P3_U2976) );
  INV_X1 U21784 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18705) );
  AOI22_X1 U21785 ( .A1(n18783), .A2(n18711), .B1(n18781), .B2(n18710), .ZN(
        n18704) );
  AOI22_X1 U21786 ( .A1(n18789), .A2(n18702), .B1(n18782), .B2(n18739), .ZN(
        n18703) );
  OAI211_X1 U21787 ( .C1(n18705), .C2(n18715), .A(n18704), .B(n18703), .ZN(
        P3_U2977) );
  AOI22_X1 U21788 ( .A1(n18788), .A2(n18739), .B1(n18787), .B2(n18710), .ZN(
        n18708) );
  AOI22_X1 U21789 ( .A1(n18789), .A2(n18706), .B1(n18790), .B2(n18711), .ZN(
        n18707) );
  OAI211_X1 U21790 ( .C1(n18709), .C2(n18715), .A(n18708), .B(n18707), .ZN(
        P3_U2978) );
  AOI22_X1 U21791 ( .A1(n18796), .A2(n18739), .B1(n18795), .B2(n18710), .ZN(
        n18714) );
  AOI22_X1 U21792 ( .A1(n18789), .A2(n18712), .B1(n18799), .B2(n18711), .ZN(
        n18713) );
  OAI211_X1 U21793 ( .C1(n18716), .C2(n18715), .A(n18714), .B(n18713), .ZN(
        P3_U2979) );
  INV_X1 U21794 ( .A(n18717), .ZN(n18743) );
  NOR2_X1 U21795 ( .A1(n18745), .A2(n18721), .ZN(n18738) );
  AOI22_X1 U21796 ( .A1(n18753), .A2(n18739), .B1(n18746), .B2(n18738), .ZN(
        n18725) );
  AOI221_X1 U21797 ( .B1(n18721), .B2(n18720), .C1(n18721), .C2(n18719), .A(
        n18718), .ZN(n18722) );
  INV_X1 U21798 ( .A(n18722), .ZN(n18740) );
  INV_X1 U21799 ( .A(n18723), .ZN(n18798) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18740), .B1(
        n18747), .B2(n18798), .ZN(n18724) );
  OAI211_X1 U21801 ( .C1(n18756), .C2(n18743), .A(n18725), .B(n18724), .ZN(
        P3_U2980) );
  AOI22_X1 U21802 ( .A1(n18757), .A2(n18738), .B1(n18759), .B2(n18798), .ZN(
        n18727) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18740), .B1(
        n18758), .B2(n18739), .ZN(n18726) );
  OAI211_X1 U21804 ( .C1(n18743), .C2(n18762), .A(n18727), .B(n18726), .ZN(
        P3_U2981) );
  AOI22_X1 U21805 ( .A1(n18764), .A2(n18739), .B1(n18763), .B2(n18738), .ZN(
        n18729) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18740), .B1(
        n18765), .B2(n18798), .ZN(n18728) );
  OAI211_X1 U21807 ( .C1(n18743), .C2(n18768), .A(n18729), .B(n18728), .ZN(
        P3_U2982) );
  AOI22_X1 U21808 ( .A1(n18771), .A2(n18798), .B1(n18769), .B2(n18738), .ZN(
        n18731) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18740), .B1(
        n18770), .B2(n18739), .ZN(n18730) );
  OAI211_X1 U21810 ( .C1(n18743), .C2(n18774), .A(n18731), .B(n18730), .ZN(
        P3_U2983) );
  AOI22_X1 U21811 ( .A1(n18776), .A2(n18739), .B1(n18775), .B2(n18738), .ZN(
        n18733) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18740), .B1(
        n18777), .B2(n18798), .ZN(n18732) );
  OAI211_X1 U21813 ( .C1(n18743), .C2(n18780), .A(n18733), .B(n18732), .ZN(
        P3_U2984) );
  AOI22_X1 U21814 ( .A1(n18783), .A2(n18739), .B1(n18781), .B2(n18738), .ZN(
        n18735) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18740), .B1(
        n18782), .B2(n18798), .ZN(n18734) );
  OAI211_X1 U21816 ( .C1(n18743), .C2(n18786), .A(n18735), .B(n18734), .ZN(
        P3_U2985) );
  AOI22_X1 U21817 ( .A1(n18790), .A2(n18739), .B1(n18787), .B2(n18738), .ZN(
        n18737) );
  AOI22_X1 U21818 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18740), .B1(
        n18788), .B2(n18798), .ZN(n18736) );
  OAI211_X1 U21819 ( .C1(n18743), .C2(n18793), .A(n18737), .B(n18736), .ZN(
        P3_U2986) );
  AOI22_X1 U21820 ( .A1(n18796), .A2(n18798), .B1(n18795), .B2(n18738), .ZN(
        n18742) );
  AOI22_X1 U21821 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18740), .B1(
        n18799), .B2(n18739), .ZN(n18741) );
  OAI211_X1 U21822 ( .C1(n18743), .C2(n18803), .A(n18742), .B(n18741), .ZN(
        P3_U2987) );
  INV_X1 U21823 ( .A(n18744), .ZN(n18804) );
  NOR2_X1 U21824 ( .A1(n18745), .A2(n18748), .ZN(n18794) );
  AOI22_X1 U21825 ( .A1(n18797), .A2(n18747), .B1(n18746), .B2(n18794), .ZN(
        n18755) );
  INV_X1 U21826 ( .A(n18748), .ZN(n18750) );
  AOI22_X1 U21827 ( .A1(n18752), .A2(n18751), .B1(n18750), .B2(n18749), .ZN(
        n18800) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18800), .B1(
        n18753), .B2(n18798), .ZN(n18754) );
  OAI211_X1 U21829 ( .C1(n18804), .C2(n18756), .A(n18755), .B(n18754), .ZN(
        P3_U2988) );
  AOI22_X1 U21830 ( .A1(n18758), .A2(n18798), .B1(n18757), .B2(n18794), .ZN(
        n18761) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18800), .B1(
        n18797), .B2(n18759), .ZN(n18760) );
  OAI211_X1 U21832 ( .C1(n18804), .C2(n18762), .A(n18761), .B(n18760), .ZN(
        P3_U2989) );
  AOI22_X1 U21833 ( .A1(n18764), .A2(n18798), .B1(n18763), .B2(n18794), .ZN(
        n18767) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18800), .B1(
        n18797), .B2(n18765), .ZN(n18766) );
  OAI211_X1 U21835 ( .C1(n18804), .C2(n18768), .A(n18767), .B(n18766), .ZN(
        P3_U2990) );
  AOI22_X1 U21836 ( .A1(n18770), .A2(n18798), .B1(n18769), .B2(n18794), .ZN(
        n18773) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18800), .B1(
        n18797), .B2(n18771), .ZN(n18772) );
  OAI211_X1 U21838 ( .C1(n18804), .C2(n18774), .A(n18773), .B(n18772), .ZN(
        P3_U2991) );
  AOI22_X1 U21839 ( .A1(n18776), .A2(n18798), .B1(n18775), .B2(n18794), .ZN(
        n18779) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18800), .B1(
        n18797), .B2(n18777), .ZN(n18778) );
  OAI211_X1 U21841 ( .C1(n18804), .C2(n18780), .A(n18779), .B(n18778), .ZN(
        P3_U2992) );
  AOI22_X1 U21842 ( .A1(n18789), .A2(n18782), .B1(n18781), .B2(n18794), .ZN(
        n18785) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18800), .B1(
        n18783), .B2(n18798), .ZN(n18784) );
  OAI211_X1 U21844 ( .C1(n18804), .C2(n18786), .A(n18785), .B(n18784), .ZN(
        P3_U2993) );
  AOI22_X1 U21845 ( .A1(n18789), .A2(n18788), .B1(n18787), .B2(n18794), .ZN(
        n18792) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18800), .B1(
        n18790), .B2(n18798), .ZN(n18791) );
  OAI211_X1 U21847 ( .C1(n18804), .C2(n18793), .A(n18792), .B(n18791), .ZN(
        P3_U2994) );
  AOI22_X1 U21848 ( .A1(n18797), .A2(n18796), .B1(n18795), .B2(n18794), .ZN(
        n18802) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18800), .B1(
        n18799), .B2(n18798), .ZN(n18801) );
  OAI211_X1 U21850 ( .C1(n18804), .C2(n18803), .A(n18802), .B(n18801), .ZN(
        P3_U2995) );
  NOR2_X1 U21851 ( .A1(n18806), .A2(n18805), .ZN(n18808) );
  OAI21_X1 U21852 ( .B1(n18809), .B2(n18808), .A(n18807), .ZN(n18810) );
  OAI221_X1 U21853 ( .B1(n18812), .B2(n18835), .C1(n18812), .C2(n18811), .A(
        n18810), .ZN(n19018) );
  OAI21_X1 U21854 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18813), .ZN(n18815) );
  OAI211_X1 U21855 ( .C1(n18840), .C2(n18863), .A(n18815), .B(n18814), .ZN(
        n18861) );
  NOR2_X1 U21856 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18826), .ZN(
        n18843) );
  INV_X1 U21857 ( .A(n18843), .ZN(n18816) );
  NAND2_X1 U21858 ( .A1(n18992), .A2(n18828), .ZN(n18823) );
  AOI22_X1 U21859 ( .A1(n18817), .A2(n18816), .B1(n10244), .B2(n18823), .ZN(
        n18818) );
  NOR2_X1 U21860 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18818), .ZN(
        n18977) );
  INV_X1 U21861 ( .A(n18819), .ZN(n18822) );
  AOI21_X1 U21862 ( .B1(n18822), .B2(n18821), .A(n18820), .ZN(n18829) );
  OAI21_X1 U21863 ( .B1(n18824), .B2(n18829), .A(n18823), .ZN(n18825) );
  AOI21_X1 U21864 ( .B1(n18832), .B2(n18826), .A(n18825), .ZN(n18978) );
  NAND2_X1 U21865 ( .A1(n18840), .A2(n18978), .ZN(n18827) );
  AOI22_X1 U21866 ( .A1(n18840), .A2(n18977), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18827), .ZN(n18859) );
  INV_X1 U21867 ( .A(n18840), .ZN(n18850) );
  AND2_X1 U21868 ( .A1(n18828), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18839) );
  OAI21_X1 U21869 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18831), .A(
        n18829), .ZN(n18838) );
  NAND2_X1 U21870 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18841), .ZN(
        n18830) );
  AOI211_X1 U21871 ( .C1(n18831), .C2(n18830), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18999), .ZN(n18837) );
  OAI21_X1 U21872 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18832), .ZN(n18833) );
  OAI22_X1 U21873 ( .A1(n18988), .A2(n18835), .B1(n18834), .B2(n18833), .ZN(
        n18836) );
  AOI211_X1 U21874 ( .C1(n18839), .C2(n18838), .A(n18837), .B(n18836), .ZN(
        n18984) );
  AOI22_X1 U21875 ( .A1(n18850), .A2(n18992), .B1(n18984), .B2(n18840), .ZN(
        n18854) );
  NOR2_X1 U21876 ( .A1(n18842), .A2(n18841), .ZN(n18844) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10247), .B1(
        n18844), .B2(n19006), .ZN(n19001) );
  OAI22_X1 U21878 ( .A1(n18844), .A2(n18993), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18843), .ZN(n18997) );
  OR3_X1 U21879 ( .A1(n19001), .A2(n18847), .A3(n18845), .ZN(n18846) );
  AOI22_X1 U21880 ( .A1(n19001), .A2(n18847), .B1(n18997), .B2(n18846), .ZN(
        n18849) );
  OAI21_X1 U21881 ( .B1(n18850), .B2(n18849), .A(n18848), .ZN(n18853) );
  AND2_X1 U21882 ( .A1(n18854), .A2(n18853), .ZN(n18851) );
  OAI221_X1 U21883 ( .B1(n18854), .B2(n18853), .C1(n18852), .C2(n18851), .A(
        n18856), .ZN(n18858) );
  AOI21_X1 U21884 ( .B1(n18856), .B2(n18855), .A(n18854), .ZN(n18857) );
  AOI222_X1 U21885 ( .A1(n18859), .A2(n18858), .B1(n18859), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18858), .C2(n18857), .ZN(
        n18860) );
  NOR4_X1 U21886 ( .A1(n18862), .A2(n19018), .A3(n18861), .A4(n18860), .ZN(
        n18875) );
  INV_X1 U21887 ( .A(n18870), .ZN(n18864) );
  AOI22_X1 U21888 ( .A1(n18865), .A2(n18884), .B1(n18864), .B2(n18863), .ZN(
        n18872) );
  NAND3_X1 U21889 ( .A1(n19025), .A2(n18867), .A3(n18866), .ZN(n18868) );
  NAND3_X1 U21890 ( .A1(n18875), .A2(n19020), .A3(n18868), .ZN(n18974) );
  NAND2_X1 U21891 ( .A1(n18884), .A2(n18869), .ZN(n18876) );
  NAND4_X1 U21892 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18974), .A3(n18870), 
        .A4(n18876), .ZN(n18880) );
  OAI22_X1 U21893 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18872), .B1(n18871), 
        .B2(n18880), .ZN(n18873) );
  OAI21_X1 U21894 ( .B1(n18875), .B2(n18874), .A(n18873), .ZN(P3_U2996) );
  NOR3_X1 U21895 ( .A1(n18877), .A2(n18985), .A3(n18876), .ZN(n18881) );
  AOI211_X1 U21896 ( .C1(n18884), .C2(n19022), .A(n18878), .B(n18881), .ZN(
        n18879) );
  OAI21_X1 U21897 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18880), .A(n18879), 
        .ZN(P3_U2997) );
  NOR4_X1 U21898 ( .A1(n19028), .A2(n18882), .A3(n18881), .A4(n18972), .ZN(
        P3_U2998) );
  AND2_X1 U21899 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18883), .ZN(
        P3_U2999) );
  AND2_X1 U21900 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18883), .ZN(
        P3_U3000) );
  AND2_X1 U21901 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18883), .ZN(
        P3_U3001) );
  AND2_X1 U21902 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18883), .ZN(
        P3_U3002) );
  AND2_X1 U21903 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18883), .ZN(
        P3_U3003) );
  AND2_X1 U21904 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18883), .ZN(
        P3_U3004) );
  AND2_X1 U21905 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18883), .ZN(
        P3_U3005) );
  AND2_X1 U21906 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18883), .ZN(
        P3_U3006) );
  AND2_X1 U21907 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18883), .ZN(
        P3_U3007) );
  AND2_X1 U21908 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18883), .ZN(
        P3_U3008) );
  AND2_X1 U21909 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18883), .ZN(
        P3_U3009) );
  AND2_X1 U21910 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18883), .ZN(
        P3_U3010) );
  AND2_X1 U21911 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18883), .ZN(
        P3_U3011) );
  AND2_X1 U21912 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18883), .ZN(
        P3_U3012) );
  AND2_X1 U21913 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18883), .ZN(
        P3_U3013) );
  AND2_X1 U21914 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18883), .ZN(
        P3_U3014) );
  AND2_X1 U21915 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18883), .ZN(
        P3_U3015) );
  AND2_X1 U21916 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18883), .ZN(
        P3_U3016) );
  AND2_X1 U21917 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18883), .ZN(
        P3_U3017) );
  AND2_X1 U21918 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18883), .ZN(
        P3_U3018) );
  AND2_X1 U21919 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18883), .ZN(
        P3_U3019) );
  AND2_X1 U21920 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18883), .ZN(
        P3_U3020) );
  AND2_X1 U21921 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18883), .ZN(P3_U3021) );
  AND2_X1 U21922 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18883), .ZN(P3_U3022) );
  AND2_X1 U21923 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18883), .ZN(P3_U3023) );
  AND2_X1 U21924 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18883), .ZN(P3_U3024) );
  AND2_X1 U21925 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18883), .ZN(P3_U3025) );
  AND2_X1 U21926 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18883), .ZN(P3_U3026) );
  AND2_X1 U21927 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18883), .ZN(P3_U3027) );
  AND2_X1 U21928 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18883), .ZN(P3_U3028) );
  NAND2_X1 U21929 ( .A1(n18884), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18893) );
  INV_X1 U21930 ( .A(n18893), .ZN(n18891) );
  OAI21_X1 U21931 ( .B1(n18885), .B2(n21001), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18886) );
  AOI22_X1 U21932 ( .A1(n18891), .A2(n18899), .B1(n19033), .B2(n18886), .ZN(
        n18887) );
  INV_X1 U21933 ( .A(NA), .ZN(n19871) );
  OR3_X1 U21934 ( .A1(n19871), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18892) );
  OAI211_X1 U21935 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18887), .B(n18892), .ZN(P3_U3029) );
  NOR2_X1 U21936 ( .A1(n18899), .A2(n21001), .ZN(n18895) );
  NOR2_X1 U21937 ( .A1(n18897), .A2(n18895), .ZN(n18888) );
  AOI21_X1 U21938 ( .B1(n18888), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n18891), .ZN(n18889) );
  OAI211_X1 U21939 ( .C1(n21001), .C2(n18890), .A(n18889), .B(n19023), .ZN(
        P3_U3030) );
  AOI21_X1 U21940 ( .B1(n18897), .B2(n18892), .A(n18891), .ZN(n18898) );
  OAI22_X1 U21941 ( .A1(NA), .A2(n18893), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18894) );
  OAI22_X1 U21942 ( .A1(n18895), .A2(n18894), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18896) );
  OAI22_X1 U21943 ( .A1(n18898), .A2(n18899), .B1(n18897), .B2(n18896), .ZN(
        P3_U3031) );
  INV_X2 U21944 ( .A(n18903), .ZN(n18956) );
  OAI222_X1 U21945 ( .A1(n19008), .A2(n18956), .B1(n18900), .B2(n18966), .C1(
        n18901), .C2(n18962), .ZN(P3_U3032) );
  OAI222_X1 U21946 ( .A1(n18962), .A2(n18904), .B1(n18902), .B2(n18966), .C1(
        n18901), .C2(n18956), .ZN(P3_U3033) );
  OAI222_X1 U21947 ( .A1(n18962), .A2(n18906), .B1(n18905), .B2(n18966), .C1(
        n18904), .C2(n18956), .ZN(P3_U3034) );
  INV_X1 U21948 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18908) );
  OAI222_X1 U21949 ( .A1(n18962), .A2(n18908), .B1(n18907), .B2(n18966), .C1(
        n18906), .C2(n18956), .ZN(P3_U3035) );
  OAI222_X1 U21950 ( .A1(n18962), .A2(n18910), .B1(n18909), .B2(n18966), .C1(
        n18908), .C2(n18956), .ZN(P3_U3036) );
  OAI222_X1 U21951 ( .A1(n18962), .A2(n18912), .B1(n18911), .B2(n18966), .C1(
        n18910), .C2(n18956), .ZN(P3_U3037) );
  OAI222_X1 U21952 ( .A1(n18962), .A2(n18915), .B1(n18913), .B2(n18966), .C1(
        n18912), .C2(n18956), .ZN(P3_U3038) );
  OAI222_X1 U21953 ( .A1(n18915), .A2(n18956), .B1(n18914), .B2(n18966), .C1(
        n18916), .C2(n18962), .ZN(P3_U3039) );
  OAI222_X1 U21954 ( .A1(n18962), .A2(n18918), .B1(n18917), .B2(n18966), .C1(
        n18916), .C2(n18956), .ZN(P3_U3040) );
  OAI222_X1 U21955 ( .A1(n18962), .A2(n18920), .B1(n18919), .B2(n18966), .C1(
        n18918), .C2(n18956), .ZN(P3_U3041) );
  OAI222_X1 U21956 ( .A1(n18962), .A2(n18922), .B1(n18921), .B2(n18966), .C1(
        n18920), .C2(n18956), .ZN(P3_U3042) );
  OAI222_X1 U21957 ( .A1(n18962), .A2(n18924), .B1(n18923), .B2(n18966), .C1(
        n18922), .C2(n18956), .ZN(P3_U3043) );
  OAI222_X1 U21958 ( .A1(n18962), .A2(n18927), .B1(n18925), .B2(n18966), .C1(
        n18924), .C2(n18956), .ZN(P3_U3044) );
  OAI222_X1 U21959 ( .A1(n18927), .A2(n18956), .B1(n18926), .B2(n18966), .C1(
        n18928), .C2(n18962), .ZN(P3_U3045) );
  INV_X1 U21960 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18930) );
  OAI222_X1 U21961 ( .A1(n18962), .A2(n18930), .B1(n18929), .B2(n18966), .C1(
        n18928), .C2(n18956), .ZN(P3_U3046) );
  OAI222_X1 U21962 ( .A1(n18962), .A2(n18933), .B1(n18931), .B2(n18966), .C1(
        n18930), .C2(n18956), .ZN(P3_U3047) );
  OAI222_X1 U21963 ( .A1(n18933), .A2(n18956), .B1(n18932), .B2(n18966), .C1(
        n18934), .C2(n18962), .ZN(P3_U3048) );
  OAI222_X1 U21964 ( .A1(n18962), .A2(n18936), .B1(n18935), .B2(n18966), .C1(
        n18934), .C2(n18956), .ZN(P3_U3049) );
  OAI222_X1 U21965 ( .A1(n18962), .A2(n18938), .B1(n18937), .B2(n18966), .C1(
        n18936), .C2(n18956), .ZN(P3_U3050) );
  OAI222_X1 U21966 ( .A1(n18962), .A2(n18940), .B1(n18939), .B2(n18966), .C1(
        n18938), .C2(n18956), .ZN(P3_U3051) );
  OAI222_X1 U21967 ( .A1(n18962), .A2(n18942), .B1(n18941), .B2(n18966), .C1(
        n18940), .C2(n18956), .ZN(P3_U3052) );
  OAI222_X1 U21968 ( .A1(n18962), .A2(n18945), .B1(n18943), .B2(n18966), .C1(
        n18942), .C2(n18956), .ZN(P3_U3053) );
  OAI222_X1 U21969 ( .A1(n18945), .A2(n18956), .B1(n18944), .B2(n18966), .C1(
        n18946), .C2(n18962), .ZN(P3_U3054) );
  OAI222_X1 U21970 ( .A1(n18962), .A2(n18948), .B1(n18947), .B2(n18966), .C1(
        n18946), .C2(n18956), .ZN(P3_U3055) );
  INV_X1 U21971 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18950) );
  OAI222_X1 U21972 ( .A1(n18962), .A2(n18950), .B1(n18949), .B2(n18966), .C1(
        n18948), .C2(n18956), .ZN(P3_U3056) );
  OAI222_X1 U21973 ( .A1(n18962), .A2(n18953), .B1(n18951), .B2(n18966), .C1(
        n18950), .C2(n18956), .ZN(P3_U3057) );
  INV_X1 U21974 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18954) );
  OAI222_X1 U21975 ( .A1(n18956), .A2(n18953), .B1(n18952), .B2(n18966), .C1(
        n18954), .C2(n18962), .ZN(P3_U3058) );
  OAI222_X1 U21976 ( .A1(n18962), .A2(n18957), .B1(n18955), .B2(n18966), .C1(
        n18954), .C2(n18956), .ZN(P3_U3059) );
  OAI222_X1 U21977 ( .A1(n18962), .A2(n18959), .B1(n18958), .B2(n18966), .C1(
        n18957), .C2(n18956), .ZN(P3_U3060) );
  INV_X1 U21978 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18960) );
  OAI222_X1 U21979 ( .A1(n18962), .A2(n18961), .B1(n18960), .B2(n18966), .C1(
        n18959), .C2(n18956), .ZN(P3_U3061) );
  OAI22_X1 U21980 ( .A1(n19033), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18966), .ZN(n18963) );
  INV_X1 U21981 ( .A(n18963), .ZN(P3_U3274) );
  OAI22_X1 U21982 ( .A1(n19033), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18966), .ZN(n18964) );
  INV_X1 U21983 ( .A(n18964), .ZN(P3_U3275) );
  OAI22_X1 U21984 ( .A1(n19033), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18966), .ZN(n18965) );
  INV_X1 U21985 ( .A(n18965), .ZN(P3_U3276) );
  OAI22_X1 U21986 ( .A1(n19033), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18966), .ZN(n18967) );
  INV_X1 U21987 ( .A(n18967), .ZN(P3_U3277) );
  OAI21_X1 U21988 ( .B1(n18971), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18969), 
        .ZN(n18968) );
  INV_X1 U21989 ( .A(n18968), .ZN(P3_U3280) );
  OAI21_X1 U21990 ( .B1(n18971), .B2(n18970), .A(n18969), .ZN(P3_U3281) );
  INV_X1 U21991 ( .A(n18972), .ZN(n18973) );
  OAI221_X1 U21992 ( .B1(n18975), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18975), 
        .C2(n18974), .A(n18973), .ZN(P3_U3282) );
  AOI22_X1 U21993 ( .A1(n19002), .A2(n18977), .B1(n19000), .B2(n18976), .ZN(
        n18983) );
  OAI21_X1 U21994 ( .B1(n18979), .B2(n18978), .A(n19004), .ZN(n18980) );
  INV_X1 U21995 ( .A(n18980), .ZN(n18982) );
  OAI22_X1 U21996 ( .A1(n19007), .A2(n18983), .B1(n18982), .B2(n18981), .ZN(
        P3_U3285) );
  INV_X1 U21997 ( .A(n18984), .ZN(n18990) );
  NOR2_X1 U21998 ( .A1(n18985), .A2(n19003), .ZN(n18994) );
  OAI22_X1 U21999 ( .A1(n18987), .A2(n18986), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18995) );
  INV_X1 U22000 ( .A(n18995), .ZN(n18989) );
  AOI222_X1 U22001 ( .A1(n18990), .A2(n19002), .B1(n18994), .B2(n18989), .C1(
        n19000), .C2(n18988), .ZN(n18991) );
  AOI22_X1 U22002 ( .A1(n19007), .A2(n18992), .B1(n18991), .B2(n19004), .ZN(
        P3_U3288) );
  INV_X1 U22003 ( .A(n18993), .ZN(n18996) );
  AOI222_X1 U22004 ( .A1(n18997), .A2(n19002), .B1(n19000), .B2(n18996), .C1(
        n18995), .C2(n18994), .ZN(n18998) );
  AOI22_X1 U22005 ( .A1(n19007), .A2(n18999), .B1(n18998), .B2(n19004), .ZN(
        P3_U3289) );
  AOI222_X1 U22006 ( .A1(n19003), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19002), 
        .B2(n19001), .C1(n19006), .C2(n19000), .ZN(n19005) );
  AOI22_X1 U22007 ( .A1(n19007), .A2(n19006), .B1(n19005), .B2(n19004), .ZN(
        P3_U3290) );
  AOI21_X1 U22008 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19009) );
  AOI22_X1 U22009 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19009), .B2(n19008), .ZN(n19012) );
  INV_X1 U22010 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19011) );
  AOI22_X1 U22011 ( .A1(n19015), .A2(n19012), .B1(n19011), .B2(n19010), .ZN(
        P3_U3292) );
  INV_X1 U22012 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19014) );
  OAI21_X1 U22013 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19015), .ZN(n19013) );
  OAI21_X1 U22014 ( .B1(n19015), .B2(n19014), .A(n19013), .ZN(P3_U3293) );
  INV_X1 U22015 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19016) );
  AOI22_X1 U22016 ( .A1(n18966), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19016), 
        .B2(n19033), .ZN(P3_U3294) );
  MUX2_X1 U22017 ( .A(P3_MORE_REG_SCAN_IN), .B(n19018), .S(n19017), .Z(
        P3_U3295) );
  OAI21_X1 U22018 ( .B1(n19020), .B2(n19019), .A(n19036), .ZN(n19021) );
  AOI21_X1 U22019 ( .B1(n19022), .B2(n19026), .A(n19021), .ZN(n19032) );
  AOI21_X1 U22020 ( .B1(n19025), .B2(n19024), .A(n19023), .ZN(n19027) );
  OAI211_X1 U22021 ( .C1(n19027), .C2(n19034), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19026), .ZN(n19029) );
  AOI21_X1 U22022 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19029), .A(n19028), 
        .ZN(n19031) );
  NAND2_X1 U22023 ( .A1(n19032), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19030) );
  OAI21_X1 U22024 ( .B1(n19032), .B2(n19031), .A(n19030), .ZN(P3_U3296) );
  MUX2_X1 U22025 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19033), .Z(P3_U3297) );
  OAI21_X1 U22026 ( .B1(n19037), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19036), 
        .ZN(n19035) );
  OAI21_X1 U22027 ( .B1(n10241), .B2(n19036), .A(n19035), .ZN(P3_U3298) );
  NOR2_X1 U22028 ( .A1(n19037), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19039)
         );
  OAI21_X1 U22029 ( .B1(n19040), .B2(n19039), .A(n19038), .ZN(P3_U3299) );
  NAND2_X1 U22030 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19889), .ZN(n19882) );
  OR2_X1 U22031 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19879) );
  OAI21_X1 U22032 ( .B1(n19878), .B2(n19882), .A(n19879), .ZN(n19956) );
  AOI21_X1 U22033 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19956), .ZN(n19041) );
  INV_X1 U22034 ( .A(n19041), .ZN(P2_U2815) );
  AOI22_X1 U22035 ( .A1(n19043), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_0__SCAN_IN), .B2(n19042), .ZN(n19044) );
  INV_X1 U22036 ( .A(n19044), .ZN(P2_U2816) );
  INV_X1 U22037 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19045) );
  AOI22_X1 U22038 ( .A1(n20005), .A2(n19045), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20006), .ZN(n19046) );
  OAI21_X1 U22039 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19883), .A(n19046), 
        .ZN(P2_U2817) );
  OAI21_X1 U22040 ( .B1(n19873), .B2(BS16), .A(n19956), .ZN(n19954) );
  OAI21_X1 U22041 ( .B1(n19956), .B2(n19633), .A(n19954), .ZN(P2_U2818) );
  NOR4_X1 U22042 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19050) );
  NOR4_X1 U22043 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19049) );
  NOR4_X1 U22044 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19048) );
  NOR4_X1 U22045 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19047) );
  NAND4_X1 U22046 ( .A1(n19050), .A2(n19049), .A3(n19048), .A4(n19047), .ZN(
        n19056) );
  NOR4_X1 U22047 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19054) );
  AOI211_X1 U22048 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19053) );
  NOR4_X1 U22049 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19052) );
  NOR4_X1 U22050 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19051) );
  NAND4_X1 U22051 ( .A1(n19054), .A2(n19053), .A3(n19052), .A4(n19051), .ZN(
        n19055) );
  NOR2_X1 U22052 ( .A1(n19056), .A2(n19055), .ZN(n19067) );
  INV_X1 U22053 ( .A(n19067), .ZN(n19065) );
  NOR2_X1 U22054 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19065), .ZN(n19059) );
  INV_X1 U22055 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19057) );
  AOI22_X1 U22056 ( .A1(n19059), .A2(n19060), .B1(n19065), .B2(n19057), .ZN(
        P2_U2820) );
  OR3_X1 U22057 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19064) );
  INV_X1 U22058 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19058) );
  AOI22_X1 U22059 ( .A1(n19059), .A2(n19064), .B1(n19065), .B2(n19058), .ZN(
        P2_U2821) );
  INV_X1 U22060 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19955) );
  NAND2_X1 U22061 ( .A1(n19059), .A2(n19955), .ZN(n19063) );
  INV_X1 U22062 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19890) );
  OAI21_X1 U22063 ( .B1(n19890), .B2(n19060), .A(n19067), .ZN(n19061) );
  OAI21_X1 U22064 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19067), .A(n19061), 
        .ZN(n19062) );
  OAI221_X1 U22065 ( .B1(n19063), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19063), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19062), .ZN(P2_U2822) );
  INV_X1 U22066 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19066) );
  OAI221_X1 U22067 ( .B1(n19067), .B2(n19066), .C1(n19065), .C2(n19064), .A(
        n19063), .ZN(P2_U2823) );
  NOR2_X1 U22068 ( .A1(n19068), .A2(n19141), .ZN(n19071) );
  AOI22_X1 U22069 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19197), .ZN(n19069) );
  OAI21_X1 U22070 ( .B1(n19202), .B2(n11156), .A(n19069), .ZN(n19070) );
  AOI211_X1 U22071 ( .C1(n19072), .C2(n19199), .A(n19071), .B(n19070), .ZN(
        n19077) );
  OAI211_X1 U22072 ( .C1(n19075), .C2(n19074), .A(n19108), .B(n19073), .ZN(
        n19076) );
  OAI211_X1 U22073 ( .C1(n19207), .C2(n19078), .A(n19077), .B(n19076), .ZN(
        P2_U2835) );
  XOR2_X1 U22074 ( .A(n19080), .B(n19079), .Z(n19089) );
  INV_X1 U22075 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U22076 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19183), .B1(n19081), 
        .B2(n19205), .ZN(n19082) );
  OAI211_X1 U22077 ( .C1(n19923), .C2(n19179), .A(n19082), .B(n19170), .ZN(
        n19083) );
  AOI21_X1 U22078 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19167), .A(
        n19083), .ZN(n19088) );
  INV_X1 U22079 ( .A(n19084), .ZN(n19085) );
  AOI22_X1 U22080 ( .A1(n19086), .A2(n19199), .B1(n19085), .B2(n19185), .ZN(
        n19087) );
  OAI211_X1 U22081 ( .C1(n19869), .C2(n19089), .A(n19088), .B(n19087), .ZN(
        P2_U2837) );
  NOR2_X1 U22082 ( .A1(n19165), .A2(n19090), .ZN(n19092) );
  XOR2_X1 U22083 ( .A(n19092), .B(n19091), .Z(n19101) );
  OAI21_X1 U22084 ( .B1(n19919), .B2(n19179), .A(n19170), .ZN(n19096) );
  OAI22_X1 U22085 ( .A1(n19094), .A2(n19141), .B1(n19093), .B2(n19210), .ZN(
        n19095) );
  AOI211_X1 U22086 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19183), .A(n19096), .B(
        n19095), .ZN(n19100) );
  AOI22_X1 U22087 ( .A1(n19098), .A2(n19199), .B1(n19097), .B2(n19185), .ZN(
        n19099) );
  OAI211_X1 U22088 ( .C1(n19869), .C2(n19101), .A(n19100), .B(n19099), .ZN(
        P2_U2839) );
  AOI22_X1 U22089 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n19183), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19167), .ZN(n19102) );
  OAI21_X1 U22090 ( .B1(n19103), .B2(n19141), .A(n19102), .ZN(n19104) );
  AOI211_X1 U22091 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19197), .A(n19286), 
        .B(n19104), .ZN(n19111) );
  NOR2_X1 U22092 ( .A1(n19165), .A2(n19105), .ZN(n19107) );
  XNOR2_X1 U22093 ( .A(n19107), .B(n19106), .ZN(n19109) );
  AOI22_X1 U22094 ( .A1(n19109), .A2(n19108), .B1(n19199), .B2(n19220), .ZN(
        n19110) );
  OAI211_X1 U22095 ( .C1(n19112), .C2(n19207), .A(n19111), .B(n19110), .ZN(
        P2_U2841) );
  OAI22_X1 U22096 ( .A1(n19113), .A2(n19141), .B1(n10211), .B2(n19210), .ZN(
        n19114) );
  AOI211_X1 U22097 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19197), .A(n19286), 
        .B(n19114), .ZN(n19122) );
  NOR2_X1 U22098 ( .A1(n19165), .A2(n19115), .ZN(n19134) );
  XNOR2_X1 U22099 ( .A(n19116), .B(n19134), .ZN(n19120) );
  INV_X1 U22100 ( .A(n19117), .ZN(n19118) );
  OAI22_X1 U22101 ( .A1(n19226), .A2(n19158), .B1(n19207), .B2(n19118), .ZN(
        n19119) );
  AOI21_X1 U22102 ( .B1(n19120), .B2(n19108), .A(n19119), .ZN(n19121) );
  OAI211_X1 U22103 ( .C1(n19202), .C2(n11124), .A(n19122), .B(n19121), .ZN(
        P2_U2843) );
  INV_X1 U22104 ( .A(n19123), .ZN(n19125) );
  AOI211_X1 U22105 ( .C1(n19125), .C2(P2_EBX_REG_11__SCAN_IN), .A(n19124), .B(
        n19141), .ZN(n19128) );
  OAI22_X1 U22106 ( .A1(n19126), .A2(n19210), .B1(n19910), .B2(n19179), .ZN(
        n19127) );
  NOR3_X1 U22107 ( .A1(n19128), .A2(n19286), .A3(n19127), .ZN(n19129) );
  OAI21_X1 U22108 ( .B1(n19130), .B2(n19158), .A(n19129), .ZN(n19131) );
  AOI21_X1 U22109 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(n19183), .A(n19131), .ZN(
        n19138) );
  AOI21_X1 U22110 ( .B1(n19136), .B2(n19132), .A(n19869), .ZN(n19133) );
  AOI22_X1 U22111 ( .A1(n19136), .A2(n19135), .B1(n19134), .B2(n19133), .ZN(
        n19137) );
  OAI211_X1 U22112 ( .C1(n19139), .C2(n19207), .A(n19138), .B(n19137), .ZN(
        P2_U2844) );
  AOI22_X1 U22113 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19183), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19167), .ZN(n19140) );
  OAI21_X1 U22114 ( .B1(n19142), .B2(n19141), .A(n19140), .ZN(n19143) );
  AOI211_X1 U22115 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19197), .A(n19286), .B(
        n19143), .ZN(n19149) );
  NOR2_X1 U22116 ( .A1(n19165), .A2(n19144), .ZN(n19146) );
  XNOR2_X1 U22117 ( .A(n19146), .B(n19145), .ZN(n19147) );
  AOI22_X1 U22118 ( .A1(n19147), .A2(n19108), .B1(n19199), .B2(n19227), .ZN(
        n19148) );
  OAI211_X1 U22119 ( .C1(n19207), .C2(n19150), .A(n19149), .B(n19148), .ZN(
        P2_U2847) );
  NAND2_X1 U22120 ( .A1(n19152), .A2(n19151), .ZN(n19154) );
  XOR2_X1 U22121 ( .A(n19154), .B(n19153), .Z(n19163) );
  AOI22_X1 U22122 ( .A1(n19155), .A2(n19205), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19167), .ZN(n19156) );
  OAI211_X1 U22123 ( .C1(n19902), .C2(n19179), .A(n19156), .B(n19170), .ZN(
        n19161) );
  OAI22_X1 U22124 ( .A1(n19159), .A2(n19158), .B1(n19207), .B2(n19157), .ZN(
        n19160) );
  AOI211_X1 U22125 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19183), .A(n19161), .B(
        n19160), .ZN(n19162) );
  OAI21_X1 U22126 ( .B1(n19163), .B2(n19869), .A(n19162), .ZN(P2_U2848) );
  NOR2_X1 U22127 ( .A1(n19165), .A2(n19164), .ZN(n19166) );
  XOR2_X1 U22128 ( .A(n19295), .B(n19166), .Z(n19178) );
  AOI22_X1 U22129 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19167), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19197), .ZN(n19172) );
  AOI22_X1 U22130 ( .A1(n19205), .A2(n19169), .B1(n19168), .B2(n19199), .ZN(
        n19171) );
  NAND3_X1 U22131 ( .A1(n19172), .A2(n19171), .A3(n19170), .ZN(n19176) );
  INV_X1 U22132 ( .A(n19213), .ZN(n19174) );
  OAI22_X1 U22133 ( .A1(n19233), .A2(n19174), .B1(n19207), .B2(n19173), .ZN(
        n19175) );
  AOI211_X1 U22134 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n19183), .A(n19176), .B(
        n19175), .ZN(n19177) );
  OAI21_X1 U22135 ( .B1(n19869), .B2(n19178), .A(n19177), .ZN(P2_U2851) );
  OAI22_X1 U22136 ( .A1(n19180), .A2(n19210), .B1(n19890), .B2(n19179), .ZN(
        n19181) );
  INV_X1 U22137 ( .A(n19181), .ZN(n19189) );
  INV_X1 U22138 ( .A(n19182), .ZN(n19184) );
  AOI22_X1 U22139 ( .A1(n19205), .A2(n19184), .B1(n19183), .B2(
        P2_EBX_REG_1__SCAN_IN), .ZN(n19188) );
  NAND2_X1 U22140 ( .A1(n19185), .A2(n13222), .ZN(n19187) );
  NAND2_X1 U22141 ( .A1(n19977), .A2(n19199), .ZN(n19186) );
  NAND4_X1 U22142 ( .A1(n19189), .A2(n19188), .A3(n19187), .A4(n19186), .ZN(
        n19190) );
  AOI21_X1 U22143 ( .B1(n19981), .B2(n19213), .A(n19190), .ZN(n19191) );
  OAI21_X1 U22144 ( .B1(n19192), .B2(n19869), .A(n19191), .ZN(n19193) );
  INV_X1 U22145 ( .A(n19193), .ZN(n19194) );
  OAI21_X1 U22146 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19195), .A(
        n19194), .ZN(P2_U2854) );
  AOI22_X1 U22147 ( .A1(n19199), .A2(n19198), .B1(n19197), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22148 ( .B1(n19202), .B2(n19201), .A(n19200), .ZN(n19203) );
  AOI21_X1 U22149 ( .B1(n19205), .B2(n19204), .A(n19203), .ZN(n19206) );
  OAI21_X1 U22150 ( .B1(n19208), .B2(n19207), .A(n19206), .ZN(n19212) );
  NOR2_X1 U22151 ( .A1(n19210), .A2(n19209), .ZN(n19211) );
  AOI211_X1 U22152 ( .C1(n19316), .C2(n19213), .A(n19212), .B(n19211), .ZN(
        n19214) );
  OAI21_X1 U22153 ( .B1(n19869), .B2(n15510), .A(n19214), .ZN(P2_U2855) );
  AOI22_X1 U22154 ( .A1(n19216), .A2(n19245), .B1(n19215), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U22155 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19231), .B1(n19217), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19218) );
  NAND2_X1 U22156 ( .A1(n19219), .A2(n19218), .ZN(P2_U2888) );
  INV_X1 U22157 ( .A(n19220), .ZN(n19223) );
  AOI22_X1 U22158 ( .A1(n19243), .A2(n19221), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19231), .ZN(n19222) );
  OAI21_X1 U22159 ( .B1(n19239), .B2(n19223), .A(n19222), .ZN(P2_U2905) );
  AOI22_X1 U22160 ( .A1(n19243), .A2(n19224), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19231), .ZN(n19225) );
  OAI21_X1 U22161 ( .B1(n19239), .B2(n19226), .A(n19225), .ZN(P2_U2907) );
  INV_X1 U22162 ( .A(n19227), .ZN(n19230) );
  AOI22_X1 U22163 ( .A1(n19243), .A2(n19228), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19231), .ZN(n19229) );
  OAI21_X1 U22164 ( .B1(n19239), .B2(n19230), .A(n19229), .ZN(P2_U2911) );
  AOI22_X1 U22165 ( .A1(n19243), .A2(n19232), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19231), .ZN(n19237) );
  INV_X1 U22166 ( .A(n19233), .ZN(n19234) );
  NAND3_X1 U22167 ( .A1(n19235), .A2(n19234), .A3(n19246), .ZN(n19236) );
  OAI211_X1 U22168 ( .C1(n19239), .C2(n19238), .A(n19237), .B(n19236), .ZN(
        P2_U2914) );
  INV_X1 U22169 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19279) );
  OAI21_X1 U22170 ( .B1(n19242), .B2(n19241), .A(n19240), .ZN(n19247) );
  AOI222_X1 U22171 ( .A1(n19247), .A2(n19246), .B1(n19971), .B2(n19245), .C1(
        n19244), .C2(n19243), .ZN(n19248) );
  OAI21_X1 U22172 ( .B1(n19249), .B2(n19279), .A(n19248), .ZN(P2_U2917) );
  AND2_X1 U22173 ( .A1(n19267), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22174 ( .A1(n19282), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22175 ( .B1(n19252), .B2(n19284), .A(n19251), .ZN(P2_U2936) );
  AOI22_X1 U22176 ( .A1(n19282), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19253) );
  OAI21_X1 U22177 ( .B1(n19254), .B2(n19284), .A(n19253), .ZN(P2_U2937) );
  AOI22_X1 U22178 ( .A1(n19282), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19255) );
  OAI21_X1 U22179 ( .B1(n19256), .B2(n19284), .A(n19255), .ZN(P2_U2938) );
  AOI22_X1 U22180 ( .A1(n19282), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19257) );
  OAI21_X1 U22181 ( .B1(n19258), .B2(n19284), .A(n19257), .ZN(P2_U2939) );
  AOI22_X1 U22182 ( .A1(n19282), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19259) );
  OAI21_X1 U22183 ( .B1(n19260), .B2(n19284), .A(n19259), .ZN(P2_U2940) );
  AOI22_X1 U22184 ( .A1(n19282), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19261) );
  OAI21_X1 U22185 ( .B1(n19262), .B2(n19284), .A(n19261), .ZN(P2_U2941) );
  AOI22_X1 U22186 ( .A1(n19282), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19263) );
  OAI21_X1 U22187 ( .B1(n19264), .B2(n19284), .A(n19263), .ZN(P2_U2942) );
  AOI22_X1 U22188 ( .A1(n19282), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19265) );
  OAI21_X1 U22189 ( .B1(n19266), .B2(n19284), .A(n19265), .ZN(P2_U2943) );
  AOI22_X1 U22190 ( .A1(n19282), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19268) );
  OAI21_X1 U22191 ( .B1(n19269), .B2(n19284), .A(n19268), .ZN(P2_U2944) );
  AOI22_X1 U22192 ( .A1(n19282), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19270) );
  OAI21_X1 U22193 ( .B1(n19271), .B2(n19284), .A(n19270), .ZN(P2_U2945) );
  INV_X1 U22194 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19273) );
  AOI22_X1 U22195 ( .A1(n19282), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19272) );
  OAI21_X1 U22196 ( .B1(n19273), .B2(n19284), .A(n19272), .ZN(P2_U2946) );
  INV_X1 U22197 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19275) );
  AOI22_X1 U22198 ( .A1(n19282), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19274) );
  OAI21_X1 U22199 ( .B1(n19275), .B2(n19284), .A(n19274), .ZN(P2_U2947) );
  INV_X1 U22200 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19277) );
  AOI22_X1 U22201 ( .A1(n19282), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19276) );
  OAI21_X1 U22202 ( .B1(n19277), .B2(n19284), .A(n19276), .ZN(P2_U2948) );
  AOI22_X1 U22203 ( .A1(n19282), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19278) );
  OAI21_X1 U22204 ( .B1(n19279), .B2(n19284), .A(n19278), .ZN(P2_U2949) );
  INV_X1 U22205 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19281) );
  AOI22_X1 U22206 ( .A1(n19282), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19280) );
  OAI21_X1 U22207 ( .B1(n19281), .B2(n19284), .A(n19280), .ZN(P2_U2950) );
  INV_X1 U22208 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19285) );
  AOI22_X1 U22209 ( .A1(n19282), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19267), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19283) );
  OAI21_X1 U22210 ( .B1(n19285), .B2(n19284), .A(n19283), .ZN(P2_U2951) );
  AOI22_X1 U22211 ( .A1(n19287), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19286), .ZN(n19294) );
  AOI222_X1 U22212 ( .A1(n19292), .A2(n19291), .B1(n19290), .B2(n19289), .C1(
        n10925), .C2(n19288), .ZN(n19293) );
  OAI211_X1 U22213 ( .C1(n19296), .C2(n19295), .A(n19294), .B(n19293), .ZN(
        P2_U3010) );
  OAI22_X1 U22214 ( .A1(n19300), .A2(n19299), .B1(n19298), .B2(n19297), .ZN(
        n19307) );
  OAI211_X1 U22215 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19302), .B(n19301), .ZN(n19303) );
  OAI21_X1 U22216 ( .B1(n19305), .B2(n19304), .A(n19303), .ZN(n19306) );
  AOI211_X1 U22217 ( .C1(n19308), .C2(n19977), .A(n19307), .B(n19306), .ZN(
        n19310) );
  OAI211_X1 U22218 ( .C1(n19312), .C2(n19311), .A(n19310), .B(n19309), .ZN(
        P2_U3045) );
  AOI22_X2 U22219 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19349), .ZN(n19766) );
  AOI22_X1 U22220 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19349), .ZN(n19813) );
  INV_X1 U22221 ( .A(n19802), .ZN(n19543) );
  NOR2_X2 U22222 ( .A1(n19317), .A2(n19351), .ZN(n19800) );
  NAND2_X1 U22223 ( .A1(n19966), .A2(n19973), .ZN(n19417) );
  INV_X1 U22224 ( .A(n19417), .ZN(n19388) );
  NAND2_X1 U22225 ( .A1(n19388), .A2(n19984), .ZN(n19361) );
  NOR2_X1 U22226 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19361), .ZN(
        n19353) );
  AOI22_X1 U22227 ( .A1(n19753), .A2(n19855), .B1(n19800), .B2(n19353), .ZN(
        n19328) );
  OAI21_X1 U22228 ( .B1(n19855), .B2(n19384), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19318) );
  NAND2_X1 U22229 ( .A1(n19318), .A2(n19961), .ZN(n19326) );
  NOR2_X1 U22230 ( .A1(n19326), .A2(n19851), .ZN(n19319) );
  AOI211_X1 U22231 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19320), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19319), .ZN(n19321) );
  OAI21_X1 U22232 ( .B1(n19321), .B2(n19353), .A(n19807), .ZN(n19356) );
  NOR2_X2 U22233 ( .A1(n19322), .A2(n19546), .ZN(n19801) );
  NOR2_X1 U22234 ( .A1(n19851), .A2(n19353), .ZN(n19325) );
  OAI21_X1 U22235 ( .B1(n19323), .B2(n19353), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19324) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19356), .B1(
        n19801), .B2(n19355), .ZN(n19327) );
  OAI211_X1 U22237 ( .C1(n19766), .C2(n19381), .A(n19328), .B(n19327), .ZN(
        P2_U3048) );
  AOI22_X1 U22238 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19349), .ZN(n19770) );
  AOI22_X1 U22239 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19349), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19350), .ZN(n19819) );
  NOR2_X2 U22240 ( .A1(n9992), .A2(n19351), .ZN(n19814) );
  AOI22_X1 U22241 ( .A1(n19767), .A2(n19855), .B1(n19814), .B2(n19353), .ZN(
        n19331) );
  NOR2_X2 U22242 ( .A1(n19329), .A2(n19546), .ZN(n19815) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19356), .B1(
        n19815), .B2(n19355), .ZN(n19330) );
  OAI211_X1 U22244 ( .C1(n19770), .C2(n19381), .A(n19331), .B(n19330), .ZN(
        P2_U3049) );
  AOI22_X1 U22245 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19349), .ZN(n19735) );
  AOI22_X1 U22246 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19349), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19350), .ZN(n19825) );
  NOR2_X2 U22247 ( .A1(n19332), .A2(n19351), .ZN(n19820) );
  AOI22_X1 U22248 ( .A1(n19732), .A2(n19855), .B1(n19820), .B2(n19353), .ZN(
        n19335) );
  NOR2_X2 U22249 ( .A1(n19333), .A2(n19546), .ZN(n19821) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19356), .B1(
        n19821), .B2(n19355), .ZN(n19334) );
  OAI211_X1 U22251 ( .C1(n19735), .C2(n19381), .A(n19335), .B(n19334), .ZN(
        P2_U3050) );
  AOI22_X1 U22252 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19349), .ZN(n19739) );
  AOI22_X1 U22253 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19349), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19350), .ZN(n19831) );
  NOR2_X2 U22254 ( .A1(n10591), .A2(n19351), .ZN(n19826) );
  AOI22_X1 U22255 ( .A1(n19736), .A2(n19855), .B1(n19826), .B2(n19353), .ZN(
        n19338) );
  NOR2_X2 U22256 ( .A1(n19336), .A2(n19546), .ZN(n19827) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19356), .B1(
        n19827), .B2(n19355), .ZN(n19337) );
  OAI211_X1 U22258 ( .C1(n19739), .C2(n19381), .A(n19338), .B(n19337), .ZN(
        P2_U3051) );
  AOI22_X1 U22259 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19349), .ZN(n19780) );
  AOI22_X1 U22260 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19349), .ZN(n19837) );
  INV_X1 U22261 ( .A(n19837), .ZN(n19777) );
  AOI22_X1 U22262 ( .A1(n19777), .A2(n19855), .B1(n19832), .B2(n19353), .ZN(
        n19342) );
  NOR2_X2 U22263 ( .A1(n19340), .A2(n19546), .ZN(n19833) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19356), .B1(
        n19833), .B2(n19355), .ZN(n19341) );
  OAI211_X1 U22265 ( .C1(n19780), .C2(n19381), .A(n19342), .B(n19341), .ZN(
        P2_U3052) );
  AOI22_X1 U22266 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19349), .ZN(n19784) );
  AOI22_X1 U22267 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19349), .ZN(n19843) );
  NOR2_X2 U22268 ( .A1(n11071), .A2(n19351), .ZN(n19838) );
  AOI22_X1 U22269 ( .A1(n19781), .A2(n19855), .B1(n19838), .B2(n19353), .ZN(
        n19345) );
  NOR2_X2 U22270 ( .A1(n19343), .A2(n19546), .ZN(n19839) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19356), .B1(
        n19839), .B2(n19355), .ZN(n19344) );
  OAI211_X1 U22272 ( .C1(n19784), .C2(n19381), .A(n19345), .B(n19344), .ZN(
        P2_U3053) );
  AOI22_X2 U22273 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19349), .ZN(n19788) );
  AOI22_X1 U22274 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19349), .ZN(n19849) );
  NOR2_X2 U22275 ( .A1(n13165), .A2(n19351), .ZN(n19844) );
  AOI22_X1 U22276 ( .A1(n19785), .A2(n19855), .B1(n19844), .B2(n19353), .ZN(
        n19348) );
  NOR2_X2 U22277 ( .A1(n19346), .A2(n19546), .ZN(n19845) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19356), .B1(
        n19845), .B2(n19355), .ZN(n19347) );
  OAI211_X1 U22279 ( .C1(n19788), .C2(n19381), .A(n19348), .B(n19347), .ZN(
        P2_U3054) );
  AOI22_X2 U22280 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19349), .ZN(n19796) );
  AOI22_X1 U22281 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19350), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19349), .ZN(n19860) );
  NOR2_X2 U22282 ( .A1(n19352), .A2(n19351), .ZN(n19850) );
  AOI22_X1 U22283 ( .A1(n19791), .A2(n19855), .B1(n19850), .B2(n19353), .ZN(
        n19358) );
  NOR2_X2 U22284 ( .A1(n19354), .A2(n19546), .ZN(n19852) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19356), .B1(
        n19852), .B2(n19355), .ZN(n19357) );
  OAI211_X1 U22286 ( .C1(n19796), .C2(n19381), .A(n19358), .B(n19357), .ZN(
        P2_U3055) );
  NAND2_X1 U22287 ( .A1(n19984), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19600) );
  NOR2_X1 U22288 ( .A1(n19600), .A2(n19417), .ZN(n19382) );
  OAI21_X1 U22289 ( .B1(n19362), .B2(n19382), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19359) );
  OAI21_X1 U22290 ( .B1(n19361), .B2(n19756), .A(n19359), .ZN(n19383) );
  AOI22_X1 U22291 ( .A1(n19383), .A2(n19801), .B1(n19800), .B2(n19382), .ZN(
        n19368) );
  NAND2_X1 U22292 ( .A1(n19360), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19544) );
  OAI21_X1 U22293 ( .B1(n19544), .B2(n19601), .A(n19361), .ZN(n19366) );
  INV_X1 U22294 ( .A(n19362), .ZN(n19364) );
  INV_X1 U22295 ( .A(n19382), .ZN(n19363) );
  OAI211_X1 U22296 ( .C1(n19364), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19363), 
        .B(n19756), .ZN(n19365) );
  NAND3_X1 U22297 ( .A1(n19366), .A2(n19807), .A3(n19365), .ZN(n19385) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19753), .ZN(n19367) );
  OAI211_X1 U22299 ( .C1(n19766), .C2(n19391), .A(n19368), .B(n19367), .ZN(
        P2_U3056) );
  AOI22_X1 U22300 ( .A1(n19383), .A2(n19815), .B1(n19814), .B2(n19382), .ZN(
        n19370) );
  INV_X1 U22301 ( .A(n19770), .ZN(n19816) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19385), .B1(
        n19413), .B2(n19816), .ZN(n19369) );
  OAI211_X1 U22303 ( .C1(n19819), .C2(n19381), .A(n19370), .B(n19369), .ZN(
        P2_U3057) );
  AOI22_X1 U22304 ( .A1(n19383), .A2(n19821), .B1(n19820), .B2(n19382), .ZN(
        n19372) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19732), .ZN(n19371) );
  OAI211_X1 U22306 ( .C1(n19735), .C2(n19391), .A(n19372), .B(n19371), .ZN(
        P2_U3058) );
  AOI22_X1 U22307 ( .A1(n19383), .A2(n19827), .B1(n19826), .B2(n19382), .ZN(
        n19374) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19736), .ZN(n19373) );
  OAI211_X1 U22309 ( .C1(n19739), .C2(n19391), .A(n19374), .B(n19373), .ZN(
        P2_U3059) );
  AOI22_X1 U22310 ( .A1(n19383), .A2(n19833), .B1(n19832), .B2(n19382), .ZN(
        n19376) );
  INV_X1 U22311 ( .A(n19780), .ZN(n19834) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19385), .B1(
        n19413), .B2(n19834), .ZN(n19375) );
  OAI211_X1 U22313 ( .C1(n19837), .C2(n19381), .A(n19376), .B(n19375), .ZN(
        P2_U3060) );
  AOI22_X1 U22314 ( .A1(n19383), .A2(n19839), .B1(n19838), .B2(n19382), .ZN(
        n19378) );
  INV_X1 U22315 ( .A(n19784), .ZN(n19840) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19385), .B1(
        n19413), .B2(n19840), .ZN(n19377) );
  OAI211_X1 U22317 ( .C1(n19843), .C2(n19381), .A(n19378), .B(n19377), .ZN(
        P2_U3061) );
  AOI22_X1 U22318 ( .A1(n19383), .A2(n19845), .B1(n19844), .B2(n19382), .ZN(
        n19380) );
  INV_X1 U22319 ( .A(n19788), .ZN(n19846) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19385), .B1(
        n19413), .B2(n19846), .ZN(n19379) );
  OAI211_X1 U22321 ( .C1(n19849), .C2(n19381), .A(n19380), .B(n19379), .ZN(
        P2_U3062) );
  AOI22_X1 U22322 ( .A1(n19383), .A2(n19852), .B1(n19850), .B2(n19382), .ZN(
        n19387) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19791), .ZN(n19386) );
  OAI211_X1 U22324 ( .C1(n19796), .C2(n19391), .A(n19387), .B(n19386), .ZN(
        P2_U3063) );
  NOR2_X1 U22325 ( .A1(n19984), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19630) );
  AND2_X1 U22326 ( .A1(n19630), .A2(n19388), .ZN(n19411) );
  OAI21_X1 U22327 ( .B1(n10802), .B2(n19411), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19390) );
  NOR2_X1 U22328 ( .A1(n19632), .A2(n19417), .ZN(n19392) );
  INV_X1 U22329 ( .A(n19392), .ZN(n19389) );
  NAND2_X1 U22330 ( .A1(n19390), .A2(n19389), .ZN(n19412) );
  AOI22_X1 U22331 ( .A1(n19412), .A2(n19801), .B1(n19800), .B2(n19411), .ZN(
        n19398) );
  AOI21_X1 U22332 ( .B1(n19446), .B2(n19391), .A(n19633), .ZN(n19393) );
  NOR2_X1 U22333 ( .A1(n19393), .A2(n19392), .ZN(n19395) );
  AOI21_X1 U22334 ( .B1(n10802), .B2(n19809), .A(n19411), .ZN(n19394) );
  MUX2_X1 U22335 ( .A(n19395), .B(n19394), .S(n19756), .Z(n19396) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19753), .ZN(n19397) );
  OAI211_X1 U22337 ( .C1(n19766), .C2(n19446), .A(n19398), .B(n19397), .ZN(
        P2_U3064) );
  AOI22_X1 U22338 ( .A1(n19412), .A2(n19815), .B1(n19814), .B2(n19411), .ZN(
        n19400) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19767), .ZN(n19399) );
  OAI211_X1 U22340 ( .C1(n19770), .C2(n19446), .A(n19400), .B(n19399), .ZN(
        P2_U3065) );
  AOI22_X1 U22341 ( .A1(n19412), .A2(n19821), .B1(n19820), .B2(n19411), .ZN(
        n19402) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19732), .ZN(n19401) );
  OAI211_X1 U22343 ( .C1(n19735), .C2(n19446), .A(n19402), .B(n19401), .ZN(
        P2_U3066) );
  AOI22_X1 U22344 ( .A1(n19412), .A2(n19827), .B1(n19826), .B2(n19411), .ZN(
        n19404) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19736), .ZN(n19403) );
  OAI211_X1 U22346 ( .C1(n19739), .C2(n19446), .A(n19404), .B(n19403), .ZN(
        P2_U3067) );
  AOI22_X1 U22347 ( .A1(n19412), .A2(n19833), .B1(n9927), .B2(n19411), .ZN(
        n19406) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19777), .ZN(n19405) );
  OAI211_X1 U22349 ( .C1(n19780), .C2(n19446), .A(n19406), .B(n19405), .ZN(
        P2_U3068) );
  AOI22_X1 U22350 ( .A1(n19412), .A2(n19839), .B1(n19838), .B2(n19411), .ZN(
        n19408) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19781), .ZN(n19407) );
  OAI211_X1 U22352 ( .C1(n19784), .C2(n19446), .A(n19408), .B(n19407), .ZN(
        P2_U3069) );
  AOI22_X1 U22353 ( .A1(n19412), .A2(n19845), .B1(n19844), .B2(n19411), .ZN(
        n19410) );
  AOI22_X1 U22354 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19785), .ZN(n19409) );
  OAI211_X1 U22355 ( .C1(n19788), .C2(n19446), .A(n19410), .B(n19409), .ZN(
        P2_U3070) );
  AOI22_X1 U22356 ( .A1(n19412), .A2(n19852), .B1(n19850), .B2(n19411), .ZN(
        n19416) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19414), .B1(
        n19413), .B2(n19791), .ZN(n19415) );
  OAI211_X1 U22358 ( .C1(n19796), .C2(n19446), .A(n19416), .B(n19415), .ZN(
        P2_U3071) );
  INV_X1 U22359 ( .A(n19766), .ZN(n19810) );
  NOR2_X1 U22360 ( .A1(n19662), .A2(n19417), .ZN(n19441) );
  AOI22_X1 U22361 ( .A1(n19810), .A2(n19476), .B1(n19441), .B2(n19800), .ZN(
        n19427) );
  OAI21_X1 U22362 ( .B1(n19544), .B2(n19669), .A(n19961), .ZN(n19425) );
  NOR2_X1 U22363 ( .A1(n19984), .A2(n19417), .ZN(n19421) );
  INV_X1 U22364 ( .A(n19441), .ZN(n19418) );
  OAI211_X1 U22365 ( .C1(n19419), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19418), 
        .B(n19756), .ZN(n19420) );
  OAI211_X1 U22366 ( .C1(n19425), .C2(n19421), .A(n19807), .B(n19420), .ZN(
        n19443) );
  INV_X1 U22367 ( .A(n19421), .ZN(n19424) );
  OAI21_X1 U22368 ( .B1(n19422), .B2(n19441), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19423) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19443), .B1(
        n19801), .B2(n19442), .ZN(n19426) );
  OAI211_X1 U22370 ( .C1(n19813), .C2(n19446), .A(n19427), .B(n19426), .ZN(
        P2_U3072) );
  AOI22_X1 U22371 ( .A1(n19816), .A2(n19476), .B1(n19441), .B2(n19814), .ZN(
        n19429) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19443), .B1(
        n19815), .B2(n19442), .ZN(n19428) );
  OAI211_X1 U22373 ( .C1(n19819), .C2(n19446), .A(n19429), .B(n19428), .ZN(
        P2_U3073) );
  INV_X1 U22374 ( .A(n19735), .ZN(n19822) );
  AOI22_X1 U22375 ( .A1(n19822), .A2(n19476), .B1(n19441), .B2(n19820), .ZN(
        n19431) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19443), .B1(
        n19821), .B2(n19442), .ZN(n19430) );
  OAI211_X1 U22377 ( .C1(n19825), .C2(n19446), .A(n19431), .B(n19430), .ZN(
        P2_U3074) );
  INV_X1 U22378 ( .A(n19739), .ZN(n19828) );
  AOI22_X1 U22379 ( .A1(n19828), .A2(n19476), .B1(n19441), .B2(n19826), .ZN(
        n19433) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19443), .B1(
        n19827), .B2(n19442), .ZN(n19432) );
  OAI211_X1 U22381 ( .C1(n19831), .C2(n19446), .A(n19433), .B(n19432), .ZN(
        P2_U3075) );
  AOI22_X1 U22382 ( .A1(n19834), .A2(n19476), .B1(n19441), .B2(n19832), .ZN(
        n19435) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19443), .B1(
        n19833), .B2(n19442), .ZN(n19434) );
  OAI211_X1 U22384 ( .C1(n19837), .C2(n19446), .A(n19435), .B(n19434), .ZN(
        P2_U3076) );
  INV_X1 U22385 ( .A(n19446), .ZN(n19438) );
  AOI22_X1 U22386 ( .A1(n19781), .A2(n19438), .B1(n19441), .B2(n19838), .ZN(
        n19437) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19443), .B1(
        n19839), .B2(n19442), .ZN(n19436) );
  OAI211_X1 U22388 ( .C1(n19784), .C2(n19454), .A(n19437), .B(n19436), .ZN(
        P2_U3077) );
  AOI22_X1 U22389 ( .A1(n19785), .A2(n19438), .B1(n19441), .B2(n19844), .ZN(
        n19440) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19443), .B1(
        n19845), .B2(n19442), .ZN(n19439) );
  OAI211_X1 U22391 ( .C1(n19788), .C2(n19454), .A(n19440), .B(n19439), .ZN(
        P2_U3078) );
  INV_X1 U22392 ( .A(n19796), .ZN(n19854) );
  AOI22_X1 U22393 ( .A1(n19854), .A2(n19476), .B1(n19441), .B2(n19850), .ZN(
        n19445) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19443), .B1(
        n19852), .B2(n19442), .ZN(n19444) );
  OAI211_X1 U22395 ( .C1(n19860), .C2(n19446), .A(n19445), .B(n19444), .ZN(
        P2_U3079) );
  OR2_X1 U22396 ( .A1(n19451), .A2(n19450), .ZN(n19695) );
  NOR2_X1 U22397 ( .A1(n19695), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19459) );
  INV_X1 U22398 ( .A(n19459), .ZN(n19453) );
  NOR3_X1 U22399 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n19973), .ZN(n19483) );
  INV_X1 U22400 ( .A(n19483), .ZN(n19485) );
  NOR2_X1 U22401 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19485), .ZN(
        n19474) );
  OAI21_X1 U22402 ( .B1(n10809), .B2(n19474), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19452) );
  OAI21_X1 U22403 ( .B1(n19756), .B2(n19453), .A(n19452), .ZN(n19475) );
  AOI22_X1 U22404 ( .A1(n19475), .A2(n19801), .B1(n19800), .B2(n19474), .ZN(
        n19461) );
  AOI21_X1 U22405 ( .B1(n19454), .B2(n19497), .A(n19633), .ZN(n19458) );
  INV_X1 U22406 ( .A(n19474), .ZN(n19455) );
  OAI211_X1 U22407 ( .C1(n19456), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19455), 
        .B(n19756), .ZN(n19457) );
  OAI211_X1 U22408 ( .C1(n19459), .C2(n19458), .A(n19457), .B(n19807), .ZN(
        n19477) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19753), .ZN(n19460) );
  OAI211_X1 U22410 ( .C1(n19766), .C2(n19497), .A(n19461), .B(n19460), .ZN(
        P2_U3080) );
  AOI22_X1 U22411 ( .A1(n19475), .A2(n19815), .B1(n19814), .B2(n19474), .ZN(
        n19463) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19767), .ZN(n19462) );
  OAI211_X1 U22413 ( .C1(n19770), .C2(n19497), .A(n19463), .B(n19462), .ZN(
        P2_U3081) );
  AOI22_X1 U22414 ( .A1(n19475), .A2(n19821), .B1(n19820), .B2(n19474), .ZN(
        n19465) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19732), .ZN(n19464) );
  OAI211_X1 U22416 ( .C1(n19735), .C2(n19497), .A(n19465), .B(n19464), .ZN(
        P2_U3082) );
  AOI22_X1 U22417 ( .A1(n19475), .A2(n19827), .B1(n19826), .B2(n19474), .ZN(
        n19467) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19736), .ZN(n19466) );
  OAI211_X1 U22419 ( .C1(n19739), .C2(n19497), .A(n19467), .B(n19466), .ZN(
        P2_U3083) );
  AOI22_X1 U22420 ( .A1(n19475), .A2(n19833), .B1(n9927), .B2(n19474), .ZN(
        n19469) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19777), .ZN(n19468) );
  OAI211_X1 U22422 ( .C1(n19780), .C2(n19497), .A(n19469), .B(n19468), .ZN(
        P2_U3084) );
  AOI22_X1 U22423 ( .A1(n19475), .A2(n19839), .B1(n19838), .B2(n19474), .ZN(
        n19471) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19781), .ZN(n19470) );
  OAI211_X1 U22425 ( .C1(n19784), .C2(n19497), .A(n19471), .B(n19470), .ZN(
        P2_U3085) );
  AOI22_X1 U22426 ( .A1(n19475), .A2(n19845), .B1(n19844), .B2(n19474), .ZN(
        n19473) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19785), .ZN(n19472) );
  OAI211_X1 U22428 ( .C1(n19788), .C2(n19497), .A(n19473), .B(n19472), .ZN(
        P2_U3086) );
  AOI22_X1 U22429 ( .A1(n19475), .A2(n19852), .B1(n19850), .B2(n19474), .ZN(
        n19479) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19791), .ZN(n19478) );
  OAI211_X1 U22431 ( .C1(n19796), .C2(n19497), .A(n19479), .B(n19478), .ZN(
        P2_U3087) );
  INV_X1 U22432 ( .A(n19497), .ZN(n19502) );
  NAND2_X1 U22433 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19483), .ZN(
        n19509) );
  INV_X1 U22434 ( .A(n19509), .ZN(n19514) );
  AOI22_X1 U22435 ( .A1(n19753), .A2(n19502), .B1(n19800), .B2(n19514), .ZN(
        n19488) );
  OAI21_X1 U22436 ( .B1(n19544), .B2(n19726), .A(n19961), .ZN(n19486) );
  OAI211_X1 U22437 ( .C1(n19481), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19509), 
        .B(n19756), .ZN(n19482) );
  OAI211_X1 U22438 ( .C1(n19486), .C2(n19483), .A(n19807), .B(n19482), .ZN(
        n19504) );
  OAI21_X1 U22439 ( .B1(n10808), .B2(n19514), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19484) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19504), .B1(
        n19801), .B2(n19503), .ZN(n19487) );
  OAI211_X1 U22441 ( .C1(n19766), .C2(n19507), .A(n19488), .B(n19487), .ZN(
        P2_U3088) );
  AOI22_X1 U22442 ( .A1(n19767), .A2(n19502), .B1(n19514), .B2(n19814), .ZN(
        n19490) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19504), .B1(
        n19815), .B2(n19503), .ZN(n19489) );
  OAI211_X1 U22444 ( .C1(n19770), .C2(n19507), .A(n19490), .B(n19489), .ZN(
        P2_U3089) );
  AOI22_X1 U22445 ( .A1(n19732), .A2(n19502), .B1(n19514), .B2(n19820), .ZN(
        n19492) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19504), .B1(
        n19821), .B2(n19503), .ZN(n19491) );
  OAI211_X1 U22447 ( .C1(n19735), .C2(n19507), .A(n19492), .B(n19491), .ZN(
        P2_U3090) );
  AOI22_X1 U22448 ( .A1(n19828), .A2(n19534), .B1(n19514), .B2(n19826), .ZN(
        n19494) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19504), .B1(
        n19827), .B2(n19503), .ZN(n19493) );
  OAI211_X1 U22450 ( .C1(n19831), .C2(n19497), .A(n19494), .B(n19493), .ZN(
        P2_U3091) );
  AOI22_X1 U22451 ( .A1(n19834), .A2(n19534), .B1(n19514), .B2(n19832), .ZN(
        n19496) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19504), .B1(
        n19833), .B2(n19503), .ZN(n19495) );
  OAI211_X1 U22453 ( .C1(n19837), .C2(n19497), .A(n19496), .B(n19495), .ZN(
        P2_U3092) );
  AOI22_X1 U22454 ( .A1(n19781), .A2(n19502), .B1(n19514), .B2(n19838), .ZN(
        n19499) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19504), .B1(
        n19839), .B2(n19503), .ZN(n19498) );
  OAI211_X1 U22456 ( .C1(n19784), .C2(n19507), .A(n19499), .B(n19498), .ZN(
        P2_U3093) );
  AOI22_X1 U22457 ( .A1(n19785), .A2(n19502), .B1(n19514), .B2(n19844), .ZN(
        n19501) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19504), .B1(
        n19845), .B2(n19503), .ZN(n19500) );
  OAI211_X1 U22459 ( .C1(n19788), .C2(n19507), .A(n19501), .B(n19500), .ZN(
        P2_U3094) );
  AOI22_X1 U22460 ( .A1(n19791), .A2(n19502), .B1(n19514), .B2(n19850), .ZN(
        n19506) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19504), .B1(
        n19852), .B2(n19503), .ZN(n19505) );
  OAI211_X1 U22462 ( .C1(n19796), .C2(n19507), .A(n19506), .B(n19505), .ZN(
        P2_U3095) );
  NAND2_X1 U22463 ( .A1(n19966), .A2(n19797), .ZN(n19541) );
  INV_X1 U22464 ( .A(n19541), .ZN(n19549) );
  NAND2_X1 U22465 ( .A1(n19549), .A2(n19994), .ZN(n19510) );
  AND2_X1 U22466 ( .A1(n19510), .A2(n19509), .ZN(n19513) );
  INV_X1 U22467 ( .A(n19510), .ZN(n19532) );
  OAI21_X1 U22468 ( .B1(n19511), .B2(n19532), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19512) );
  OAI21_X1 U22469 ( .B1(n19513), .B2(n19756), .A(n19512), .ZN(n19533) );
  AOI22_X1 U22470 ( .A1(n19533), .A2(n19801), .B1(n19800), .B2(n19532), .ZN(
        n19519) );
  AOI221_X1 U22471 ( .B1(n19534), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19565), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19514), .ZN(n19515) );
  AOI211_X1 U22472 ( .C1(n19516), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19515), .ZN(n19517) );
  OAI21_X1 U22473 ( .B1(n19517), .B2(n19532), .A(n19807), .ZN(n19535) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19753), .ZN(n19518) );
  OAI211_X1 U22475 ( .C1(n19766), .C2(n19538), .A(n19519), .B(n19518), .ZN(
        P2_U3096) );
  AOI22_X1 U22476 ( .A1(n19533), .A2(n19815), .B1(n19814), .B2(n19532), .ZN(
        n19521) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19767), .ZN(n19520) );
  OAI211_X1 U22478 ( .C1(n19770), .C2(n19538), .A(n19521), .B(n19520), .ZN(
        P2_U3097) );
  AOI22_X1 U22479 ( .A1(n19533), .A2(n19821), .B1(n19820), .B2(n19532), .ZN(
        n19523) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19732), .ZN(n19522) );
  OAI211_X1 U22481 ( .C1(n19735), .C2(n19538), .A(n19523), .B(n19522), .ZN(
        P2_U3098) );
  AOI22_X1 U22482 ( .A1(n19533), .A2(n19827), .B1(n19826), .B2(n19532), .ZN(
        n19525) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19736), .ZN(n19524) );
  OAI211_X1 U22484 ( .C1(n19739), .C2(n19538), .A(n19525), .B(n19524), .ZN(
        P2_U3099) );
  AOI22_X1 U22485 ( .A1(n19533), .A2(n19833), .B1(n9927), .B2(n19532), .ZN(
        n19527) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19777), .ZN(n19526) );
  OAI211_X1 U22487 ( .C1(n19780), .C2(n19538), .A(n19527), .B(n19526), .ZN(
        P2_U3100) );
  AOI22_X1 U22488 ( .A1(n19533), .A2(n19839), .B1(n19838), .B2(n19532), .ZN(
        n19529) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19781), .ZN(n19528) );
  OAI211_X1 U22490 ( .C1(n19784), .C2(n19538), .A(n19529), .B(n19528), .ZN(
        P2_U3101) );
  AOI22_X1 U22491 ( .A1(n19533), .A2(n19845), .B1(n19844), .B2(n19532), .ZN(
        n19531) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19785), .ZN(n19530) );
  OAI211_X1 U22493 ( .C1(n19788), .C2(n19538), .A(n19531), .B(n19530), .ZN(
        P2_U3102) );
  AOI22_X1 U22494 ( .A1(n19533), .A2(n19852), .B1(n19850), .B2(n19532), .ZN(
        n19537) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19535), .B1(
        n19534), .B2(n19791), .ZN(n19536) );
  OAI211_X1 U22496 ( .C1(n19796), .C2(n19538), .A(n19537), .B(n19536), .ZN(
        P2_U3103) );
  NOR2_X1 U22497 ( .A1(n19994), .A2(n19541), .ZN(n19573) );
  NOR3_X1 U22498 ( .A1(n10828), .A2(n19573), .A3(n19798), .ZN(n19545) );
  AOI21_X1 U22499 ( .B1(n19809), .B2(n19549), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19542) );
  AOI22_X1 U22500 ( .A1(n19564), .A2(n19801), .B1(n19800), .B2(n19573), .ZN(
        n19551) );
  NOR2_X1 U22501 ( .A1(n19544), .A2(n19543), .ZN(n19960) );
  INV_X1 U22502 ( .A(n19573), .ZN(n19547) );
  AOI211_X1 U22503 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19547), .A(n19546), 
        .B(n19545), .ZN(n19548) );
  OAI21_X1 U22504 ( .B1(n19549), .B2(n19960), .A(n19548), .ZN(n19566) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19753), .ZN(n19550) );
  OAI211_X1 U22506 ( .C1(n19766), .C2(n19599), .A(n19551), .B(n19550), .ZN(
        P2_U3104) );
  AOI22_X1 U22507 ( .A1(n19564), .A2(n19815), .B1(n19814), .B2(n19573), .ZN(
        n19553) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19767), .ZN(n19552) );
  OAI211_X1 U22509 ( .C1(n19770), .C2(n19599), .A(n19553), .B(n19552), .ZN(
        P2_U3105) );
  AOI22_X1 U22510 ( .A1(n19564), .A2(n19821), .B1(n19820), .B2(n19573), .ZN(
        n19555) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19732), .ZN(n19554) );
  OAI211_X1 U22512 ( .C1(n19735), .C2(n19599), .A(n19555), .B(n19554), .ZN(
        P2_U3106) );
  AOI22_X1 U22513 ( .A1(n19564), .A2(n19827), .B1(n19826), .B2(n19573), .ZN(
        n19557) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19736), .ZN(n19556) );
  OAI211_X1 U22515 ( .C1(n19739), .C2(n19599), .A(n19557), .B(n19556), .ZN(
        P2_U3107) );
  AOI22_X1 U22516 ( .A1(n19564), .A2(n19833), .B1(n9927), .B2(n19573), .ZN(
        n19559) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19777), .ZN(n19558) );
  OAI211_X1 U22518 ( .C1(n19780), .C2(n19599), .A(n19559), .B(n19558), .ZN(
        P2_U3108) );
  AOI22_X1 U22519 ( .A1(n19564), .A2(n19839), .B1(n19838), .B2(n19573), .ZN(
        n19561) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19781), .ZN(n19560) );
  OAI211_X1 U22521 ( .C1(n19784), .C2(n19599), .A(n19561), .B(n19560), .ZN(
        P2_U3109) );
  AOI22_X1 U22522 ( .A1(n19564), .A2(n19845), .B1(n19844), .B2(n19573), .ZN(
        n19563) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19785), .ZN(n19562) );
  OAI211_X1 U22524 ( .C1(n19788), .C2(n19599), .A(n19563), .B(n19562), .ZN(
        P2_U3110) );
  AOI22_X1 U22525 ( .A1(n19564), .A2(n19852), .B1(n19850), .B2(n19573), .ZN(
        n19568) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19791), .ZN(n19567) );
  OAI211_X1 U22527 ( .C1(n19796), .C2(n19599), .A(n19568), .B(n19567), .ZN(
        P2_U3111) );
  NAND2_X1 U22528 ( .A1(n19752), .A2(n19569), .ZN(n19624) );
  NAND2_X1 U22529 ( .A1(n19973), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19661) );
  NOR2_X1 U22530 ( .A1(n19661), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19605) );
  INV_X1 U22531 ( .A(n19605), .ZN(n19608) );
  NOR2_X1 U22532 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19608), .ZN(
        n19594) );
  AOI22_X1 U22533 ( .A1(n19810), .A2(n19625), .B1(n19800), .B2(n19594), .ZN(
        n19581) );
  AOI21_X1 U22534 ( .B1(n19570), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19576) );
  INV_X1 U22535 ( .A(n19599), .ZN(n19571) );
  OAI21_X1 U22536 ( .B1(n19625), .B2(n19571), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19572) );
  NAND2_X1 U22537 ( .A1(n19572), .A2(n19961), .ZN(n19579) );
  INV_X1 U22538 ( .A(n19579), .ZN(n19574) );
  NOR2_X1 U22539 ( .A1(n19594), .A2(n19573), .ZN(n19577) );
  NAND2_X1 U22540 ( .A1(n19574), .A2(n19577), .ZN(n19575) );
  OAI211_X1 U22541 ( .C1(n19594), .C2(n19576), .A(n19575), .B(n19807), .ZN(
        n19596) );
  OAI21_X1 U22542 ( .B1(n10757), .B2(n19594), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19578) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19596), .B1(
        n19801), .B2(n19595), .ZN(n19580) );
  OAI211_X1 U22544 ( .C1(n19813), .C2(n19599), .A(n19581), .B(n19580), .ZN(
        P2_U3112) );
  AOI22_X1 U22545 ( .A1(n19816), .A2(n19625), .B1(n19814), .B2(n19594), .ZN(
        n19583) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19596), .B1(
        n19815), .B2(n19595), .ZN(n19582) );
  OAI211_X1 U22547 ( .C1(n19819), .C2(n19599), .A(n19583), .B(n19582), .ZN(
        P2_U3113) );
  AOI22_X1 U22548 ( .A1(n19822), .A2(n19625), .B1(n19820), .B2(n19594), .ZN(
        n19585) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19596), .B1(
        n19821), .B2(n19595), .ZN(n19584) );
  OAI211_X1 U22550 ( .C1(n19825), .C2(n19599), .A(n19585), .B(n19584), .ZN(
        P2_U3114) );
  AOI22_X1 U22551 ( .A1(n19828), .A2(n19625), .B1(n19826), .B2(n19594), .ZN(
        n19587) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19596), .B1(
        n19827), .B2(n19595), .ZN(n19586) );
  OAI211_X1 U22553 ( .C1(n19831), .C2(n19599), .A(n19587), .B(n19586), .ZN(
        P2_U3115) );
  AOI22_X1 U22554 ( .A1(n19834), .A2(n19625), .B1(n19832), .B2(n19594), .ZN(
        n19589) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19596), .B1(
        n19833), .B2(n19595), .ZN(n19588) );
  OAI211_X1 U22556 ( .C1(n19837), .C2(n19599), .A(n19589), .B(n19588), .ZN(
        P2_U3116) );
  AOI22_X1 U22557 ( .A1(n19840), .A2(n19625), .B1(n19838), .B2(n19594), .ZN(
        n19591) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19596), .B1(
        n19839), .B2(n19595), .ZN(n19590) );
  OAI211_X1 U22559 ( .C1(n19843), .C2(n19599), .A(n19591), .B(n19590), .ZN(
        P2_U3117) );
  AOI22_X1 U22560 ( .A1(n19846), .A2(n19625), .B1(n19844), .B2(n19594), .ZN(
        n19593) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19596), .B1(
        n19845), .B2(n19595), .ZN(n19592) );
  OAI211_X1 U22562 ( .C1(n19849), .C2(n19599), .A(n19593), .B(n19592), .ZN(
        P2_U3118) );
  AOI22_X1 U22563 ( .A1(n19854), .A2(n19625), .B1(n19850), .B2(n19594), .ZN(
        n19598) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19596), .B1(
        n19852), .B2(n19595), .ZN(n19597) );
  OAI211_X1 U22565 ( .C1(n19860), .C2(n19599), .A(n19598), .B(n19597), .ZN(
        P2_U3119) );
  NOR2_X1 U22566 ( .A1(n19600), .A2(n19661), .ZN(n19635) );
  AOI22_X1 U22567 ( .A1(n19753), .A2(n19625), .B1(n19800), .B2(n19635), .ZN(
        n19611) );
  NAND2_X1 U22568 ( .A1(n19963), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19723) );
  OAI21_X1 U22569 ( .B1(n19723), .B2(n19601), .A(n19961), .ZN(n19609) );
  INV_X1 U22570 ( .A(n19635), .ZN(n19602) );
  OAI211_X1 U22571 ( .C1(n19603), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19602), 
        .B(n19756), .ZN(n19604) );
  OAI211_X1 U22572 ( .C1(n19609), .C2(n19605), .A(n19807), .B(n19604), .ZN(
        n19627) );
  OAI21_X1 U22573 ( .B1(n19606), .B2(n19635), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19607) );
  OAI21_X1 U22574 ( .B1(n19609), .B2(n19608), .A(n19607), .ZN(n19626) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19627), .B1(
        n19801), .B2(n19626), .ZN(n19610) );
  OAI211_X1 U22576 ( .C1(n19766), .C2(n19634), .A(n19611), .B(n19610), .ZN(
        P2_U3120) );
  AOI22_X1 U22577 ( .A1(n19767), .A2(n19625), .B1(n19814), .B2(n19635), .ZN(
        n19613) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19627), .B1(
        n19815), .B2(n19626), .ZN(n19612) );
  OAI211_X1 U22579 ( .C1(n19770), .C2(n19634), .A(n19613), .B(n19612), .ZN(
        P2_U3121) );
  AOI22_X1 U22580 ( .A1(n19822), .A2(n19656), .B1(n19820), .B2(n19635), .ZN(
        n19615) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19627), .B1(
        n19821), .B2(n19626), .ZN(n19614) );
  OAI211_X1 U22582 ( .C1(n19825), .C2(n19624), .A(n19615), .B(n19614), .ZN(
        P2_U3122) );
  AOI22_X1 U22583 ( .A1(n19736), .A2(n19625), .B1(n19826), .B2(n19635), .ZN(
        n19617) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19627), .B1(
        n19827), .B2(n19626), .ZN(n19616) );
  OAI211_X1 U22585 ( .C1(n19739), .C2(n19634), .A(n19617), .B(n19616), .ZN(
        P2_U3123) );
  AOI22_X1 U22586 ( .A1(n19834), .A2(n19656), .B1(n19832), .B2(n19635), .ZN(
        n19619) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19627), .B1(
        n19833), .B2(n19626), .ZN(n19618) );
  OAI211_X1 U22588 ( .C1(n19837), .C2(n19624), .A(n19619), .B(n19618), .ZN(
        P2_U3124) );
  AOI22_X1 U22589 ( .A1(n19840), .A2(n19656), .B1(n19838), .B2(n19635), .ZN(
        n19621) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19627), .B1(
        n19839), .B2(n19626), .ZN(n19620) );
  OAI211_X1 U22591 ( .C1(n19843), .C2(n19624), .A(n19621), .B(n19620), .ZN(
        P2_U3125) );
  AOI22_X1 U22592 ( .A1(n19846), .A2(n19656), .B1(n19844), .B2(n19635), .ZN(
        n19623) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19627), .B1(
        n19845), .B2(n19626), .ZN(n19622) );
  OAI211_X1 U22594 ( .C1(n19849), .C2(n19624), .A(n19623), .B(n19622), .ZN(
        P2_U3126) );
  AOI22_X1 U22595 ( .A1(n19791), .A2(n19625), .B1(n19850), .B2(n19635), .ZN(
        n19629) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19627), .B1(
        n19852), .B2(n19626), .ZN(n19628) );
  OAI211_X1 U22597 ( .C1(n19796), .C2(n19634), .A(n19629), .B(n19628), .ZN(
        P2_U3127) );
  INV_X1 U22598 ( .A(n19661), .ZN(n19660) );
  AND2_X1 U22599 ( .A1(n19630), .A2(n19660), .ZN(n19654) );
  OAI21_X1 U22600 ( .B1(n10810), .B2(n19654), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19631) );
  OAI21_X1 U22601 ( .B1(n19661), .B2(n19632), .A(n19631), .ZN(n19655) );
  AOI22_X1 U22602 ( .A1(n19655), .A2(n19801), .B1(n19800), .B2(n19654), .ZN(
        n19641) );
  AOI21_X1 U22603 ( .B1(n19689), .B2(n19634), .A(n19633), .ZN(n19636) );
  NOR2_X1 U22604 ( .A1(n19636), .A2(n19635), .ZN(n19637) );
  AOI211_X1 U22605 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19638), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19637), .ZN(n19639) );
  OAI21_X1 U22606 ( .B1(n19639), .B2(n19654), .A(n19807), .ZN(n19657) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19753), .ZN(n19640) );
  OAI211_X1 U22608 ( .C1(n19766), .C2(n19689), .A(n19641), .B(n19640), .ZN(
        P2_U3128) );
  AOI22_X1 U22609 ( .A1(n19655), .A2(n19815), .B1(n19814), .B2(n19654), .ZN(
        n19643) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19767), .ZN(n19642) );
  OAI211_X1 U22611 ( .C1(n19770), .C2(n19689), .A(n19643), .B(n19642), .ZN(
        P2_U3129) );
  AOI22_X1 U22612 ( .A1(n19655), .A2(n19821), .B1(n19820), .B2(n19654), .ZN(
        n19645) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19732), .ZN(n19644) );
  OAI211_X1 U22614 ( .C1(n19735), .C2(n19689), .A(n19645), .B(n19644), .ZN(
        P2_U3130) );
  AOI22_X1 U22615 ( .A1(n19655), .A2(n19827), .B1(n19826), .B2(n19654), .ZN(
        n19647) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19736), .ZN(n19646) );
  OAI211_X1 U22617 ( .C1(n19739), .C2(n19689), .A(n19647), .B(n19646), .ZN(
        P2_U3131) );
  AOI22_X1 U22618 ( .A1(n19655), .A2(n19833), .B1(n9927), .B2(n19654), .ZN(
        n19649) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19777), .ZN(n19648) );
  OAI211_X1 U22620 ( .C1(n19780), .C2(n19689), .A(n19649), .B(n19648), .ZN(
        P2_U3132) );
  AOI22_X1 U22621 ( .A1(n19655), .A2(n19839), .B1(n19838), .B2(n19654), .ZN(
        n19651) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19781), .ZN(n19650) );
  OAI211_X1 U22623 ( .C1(n19784), .C2(n19689), .A(n19651), .B(n19650), .ZN(
        P2_U3133) );
  AOI22_X1 U22624 ( .A1(n19655), .A2(n19845), .B1(n19844), .B2(n19654), .ZN(
        n19653) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19785), .ZN(n19652) );
  OAI211_X1 U22626 ( .C1(n19788), .C2(n19689), .A(n19653), .B(n19652), .ZN(
        P2_U3134) );
  AOI22_X1 U22627 ( .A1(n19655), .A2(n19852), .B1(n19850), .B2(n19654), .ZN(
        n19659) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19657), .B1(
        n19656), .B2(n19791), .ZN(n19658) );
  OAI211_X1 U22629 ( .C1(n19796), .C2(n19689), .A(n19659), .B(n19658), .ZN(
        P2_U3135) );
  NAND2_X1 U22630 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19660), .ZN(
        n19666) );
  OR2_X1 U22631 ( .A1(n19666), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19664) );
  NOR2_X1 U22632 ( .A1(n19662), .A2(n19661), .ZN(n19684) );
  NOR3_X1 U22633 ( .A1(n19663), .A2(n19684), .A3(n19798), .ZN(n19665) );
  AOI21_X1 U22634 ( .B1(n19798), .B2(n19664), .A(n19665), .ZN(n19685) );
  AOI22_X1 U22635 ( .A1(n19685), .A2(n19801), .B1(n19800), .B2(n19684), .ZN(
        n19671) );
  INV_X1 U22636 ( .A(n19723), .ZN(n19803) );
  NAND2_X1 U22637 ( .A1(n19803), .A2(n19957), .ZN(n19667) );
  AOI21_X1 U22638 ( .B1(n19667), .B2(n19666), .A(n19665), .ZN(n19668) );
  OAI211_X1 U22639 ( .C1(n19684), .C2(n19809), .A(n19668), .B(n19807), .ZN(
        n19686) );
  NOR2_X2 U22640 ( .A1(n19727), .A2(n19669), .ZN(n19716) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19810), .ZN(n19670) );
  OAI211_X1 U22642 ( .C1(n19813), .C2(n19689), .A(n19671), .B(n19670), .ZN(
        P2_U3136) );
  AOI22_X1 U22643 ( .A1(n19685), .A2(n19815), .B1(n19814), .B2(n19684), .ZN(
        n19673) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19816), .ZN(n19672) );
  OAI211_X1 U22645 ( .C1(n19819), .C2(n19689), .A(n19673), .B(n19672), .ZN(
        P2_U3137) );
  AOI22_X1 U22646 ( .A1(n19685), .A2(n19821), .B1(n19820), .B2(n19684), .ZN(
        n19675) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19822), .ZN(n19674) );
  OAI211_X1 U22648 ( .C1(n19825), .C2(n19689), .A(n19675), .B(n19674), .ZN(
        P2_U3138) );
  AOI22_X1 U22649 ( .A1(n19685), .A2(n19827), .B1(n19826), .B2(n19684), .ZN(
        n19677) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19828), .ZN(n19676) );
  OAI211_X1 U22651 ( .C1(n19831), .C2(n19689), .A(n19677), .B(n19676), .ZN(
        P2_U3139) );
  AOI22_X1 U22652 ( .A1(n19685), .A2(n19833), .B1(n9927), .B2(n19684), .ZN(
        n19679) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19834), .ZN(n19678) );
  OAI211_X1 U22654 ( .C1(n19837), .C2(n19689), .A(n19679), .B(n19678), .ZN(
        P2_U3140) );
  AOI22_X1 U22655 ( .A1(n19685), .A2(n19839), .B1(n19838), .B2(n19684), .ZN(
        n19681) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19840), .ZN(n19680) );
  OAI211_X1 U22657 ( .C1(n19843), .C2(n19689), .A(n19681), .B(n19680), .ZN(
        P2_U3141) );
  AOI22_X1 U22658 ( .A1(n19685), .A2(n19845), .B1(n19844), .B2(n19684), .ZN(
        n19683) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19846), .ZN(n19682) );
  OAI211_X1 U22660 ( .C1(n19849), .C2(n19689), .A(n19683), .B(n19682), .ZN(
        P2_U3142) );
  AOI22_X1 U22661 ( .A1(n19685), .A2(n19852), .B1(n19850), .B2(n19684), .ZN(
        n19688) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19686), .B1(
        n19716), .B2(n19854), .ZN(n19687) );
  OAI211_X1 U22663 ( .C1(n19860), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P2_U3143) );
  INV_X1 U22664 ( .A(n19752), .ZN(n19690) );
  INV_X1 U22665 ( .A(n19691), .ZN(n19693) );
  NAND3_X1 U22666 ( .A1(n19984), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19722) );
  NOR2_X1 U22667 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19722), .ZN(
        n19714) );
  OAI21_X1 U22668 ( .B1(n10800), .B2(n19714), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19692) );
  OAI21_X1 U22669 ( .B1(n19693), .B2(n19695), .A(n19692), .ZN(n19715) );
  AOI22_X1 U22670 ( .A1(n19715), .A2(n19801), .B1(n19800), .B2(n19714), .ZN(
        n19701) );
  OAI21_X1 U22671 ( .B1(n19716), .B2(n19744), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19694) );
  OAI21_X1 U22672 ( .B1(n19695), .B2(n19966), .A(n19694), .ZN(n19699) );
  INV_X1 U22673 ( .A(n19714), .ZN(n19696) );
  OAI211_X1 U22674 ( .C1(n19697), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19696), 
        .B(n19756), .ZN(n19698) );
  NAND3_X1 U22675 ( .A1(n19699), .A2(n19807), .A3(n19698), .ZN(n19717) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19753), .ZN(n19700) );
  OAI211_X1 U22677 ( .C1(n19766), .C2(n19751), .A(n19701), .B(n19700), .ZN(
        P2_U3144) );
  AOI22_X1 U22678 ( .A1(n19715), .A2(n19815), .B1(n19814), .B2(n19714), .ZN(
        n19703) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19767), .ZN(n19702) );
  OAI211_X1 U22680 ( .C1(n19770), .C2(n19751), .A(n19703), .B(n19702), .ZN(
        P2_U3145) );
  AOI22_X1 U22681 ( .A1(n19715), .A2(n19821), .B1(n19820), .B2(n19714), .ZN(
        n19705) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19732), .ZN(n19704) );
  OAI211_X1 U22683 ( .C1(n19735), .C2(n19751), .A(n19705), .B(n19704), .ZN(
        P2_U3146) );
  AOI22_X1 U22684 ( .A1(n19715), .A2(n19827), .B1(n19826), .B2(n19714), .ZN(
        n19707) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19736), .ZN(n19706) );
  OAI211_X1 U22686 ( .C1(n19739), .C2(n19751), .A(n19707), .B(n19706), .ZN(
        P2_U3147) );
  AOI22_X1 U22687 ( .A1(n19715), .A2(n19833), .B1(n9927), .B2(n19714), .ZN(
        n19709) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19777), .ZN(n19708) );
  OAI211_X1 U22689 ( .C1(n19780), .C2(n19751), .A(n19709), .B(n19708), .ZN(
        P2_U3148) );
  AOI22_X1 U22690 ( .A1(n19715), .A2(n19839), .B1(n19838), .B2(n19714), .ZN(
        n19711) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19781), .ZN(n19710) );
  OAI211_X1 U22692 ( .C1(n19784), .C2(n19751), .A(n19711), .B(n19710), .ZN(
        P2_U3149) );
  AOI22_X1 U22693 ( .A1(n19715), .A2(n19845), .B1(n19844), .B2(n19714), .ZN(
        n19713) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19785), .ZN(n19712) );
  OAI211_X1 U22695 ( .C1(n19788), .C2(n19751), .A(n19713), .B(n19712), .ZN(
        P2_U3150) );
  AOI22_X1 U22696 ( .A1(n19715), .A2(n19852), .B1(n19850), .B2(n19714), .ZN(
        n19719) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19717), .B1(
        n19716), .B2(n19791), .ZN(n19718) );
  OAI211_X1 U22698 ( .C1(n19796), .C2(n19751), .A(n19719), .B(n19718), .ZN(
        P2_U3151) );
  NOR2_X1 U22699 ( .A1(n19994), .A2(n19722), .ZN(n19755) );
  OAI21_X1 U22700 ( .B1(n10799), .B2(n19755), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19720) );
  OAI21_X1 U22701 ( .B1(n19722), .B2(n19756), .A(n19720), .ZN(n19747) );
  AOI22_X1 U22702 ( .A1(n19747), .A2(n19801), .B1(n19800), .B2(n19755), .ZN(
        n19729) );
  AOI21_X1 U22703 ( .B1(n19721), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19725) );
  OAI21_X1 U22704 ( .B1(n19723), .B2(n19726), .A(n19722), .ZN(n19724) );
  OAI211_X1 U22705 ( .C1(n19755), .C2(n19725), .A(n19724), .B(n19807), .ZN(
        n19748) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19748), .B1(
        n19790), .B2(n19810), .ZN(n19728) );
  OAI211_X1 U22707 ( .C1(n19813), .C2(n19751), .A(n19729), .B(n19728), .ZN(
        P2_U3152) );
  AOI22_X1 U22708 ( .A1(n19747), .A2(n19815), .B1(n19814), .B2(n19755), .ZN(
        n19731) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19748), .B1(
        n19790), .B2(n19816), .ZN(n19730) );
  OAI211_X1 U22710 ( .C1(n19819), .C2(n19751), .A(n19731), .B(n19730), .ZN(
        P2_U3153) );
  AOI22_X1 U22711 ( .A1(n19747), .A2(n19821), .B1(n19820), .B2(n19755), .ZN(
        n19734) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19748), .B1(
        n19744), .B2(n19732), .ZN(n19733) );
  OAI211_X1 U22713 ( .C1(n19735), .C2(n19776), .A(n19734), .B(n19733), .ZN(
        P2_U3154) );
  AOI22_X1 U22714 ( .A1(n19747), .A2(n19827), .B1(n19826), .B2(n19755), .ZN(
        n19738) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19748), .B1(
        n19744), .B2(n19736), .ZN(n19737) );
  OAI211_X1 U22716 ( .C1(n19739), .C2(n19776), .A(n19738), .B(n19737), .ZN(
        P2_U3155) );
  AOI22_X1 U22717 ( .A1(n19747), .A2(n19833), .B1(n9927), .B2(n19755), .ZN(
        n19741) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19748), .B1(
        n19790), .B2(n19834), .ZN(n19740) );
  OAI211_X1 U22719 ( .C1(n19837), .C2(n19751), .A(n19741), .B(n19740), .ZN(
        P2_U3156) );
  AOI22_X1 U22720 ( .A1(n19747), .A2(n19839), .B1(n19838), .B2(n19755), .ZN(
        n19743) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19748), .B1(
        n19790), .B2(n19840), .ZN(n19742) );
  OAI211_X1 U22722 ( .C1(n19843), .C2(n19751), .A(n19743), .B(n19742), .ZN(
        P2_U3157) );
  AOI22_X1 U22723 ( .A1(n19747), .A2(n19845), .B1(n19844), .B2(n19755), .ZN(
        n19746) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19748), .B1(
        n19744), .B2(n19785), .ZN(n19745) );
  OAI211_X1 U22725 ( .C1(n19788), .C2(n19776), .A(n19746), .B(n19745), .ZN(
        P2_U3158) );
  AOI22_X1 U22726 ( .A1(n19747), .A2(n19852), .B1(n19850), .B2(n19755), .ZN(
        n19750) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19748), .B1(
        n19790), .B2(n19854), .ZN(n19749) );
  OAI211_X1 U22728 ( .C1(n19860), .C2(n19751), .A(n19750), .B(n19749), .ZN(
        P2_U3159) );
  AND3_X1 U22729 ( .A1(n19994), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19797), .ZN(n19789) );
  AOI22_X1 U22730 ( .A1(n19753), .A2(n19790), .B1(n19800), .B2(n19789), .ZN(
        n19765) );
  INV_X1 U22731 ( .A(n19859), .ZN(n19773) );
  OAI21_X1 U22732 ( .B1(n19773), .B2(n19790), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19754) );
  NAND2_X1 U22733 ( .A1(n19754), .A2(n19961), .ZN(n19763) );
  NOR2_X1 U22734 ( .A1(n19789), .A2(n19755), .ZN(n19762) );
  INV_X1 U22735 ( .A(n19762), .ZN(n19760) );
  INV_X1 U22736 ( .A(n19789), .ZN(n19757) );
  OAI211_X1 U22737 ( .C1(n19758), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19757), 
        .B(n19756), .ZN(n19759) );
  OAI211_X1 U22738 ( .C1(n19763), .C2(n19760), .A(n19807), .B(n19759), .ZN(
        n19793) );
  OAI21_X1 U22739 ( .B1(n10803), .B2(n19789), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19761) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19793), .B1(
        n19801), .B2(n19792), .ZN(n19764) );
  OAI211_X1 U22741 ( .C1(n19766), .C2(n19859), .A(n19765), .B(n19764), .ZN(
        P2_U3160) );
  AOI22_X1 U22742 ( .A1(n19767), .A2(n19790), .B1(n19814), .B2(n19789), .ZN(
        n19769) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19793), .B1(
        n19815), .B2(n19792), .ZN(n19768) );
  OAI211_X1 U22744 ( .C1(n19770), .C2(n19859), .A(n19769), .B(n19768), .ZN(
        P2_U3161) );
  AOI22_X1 U22745 ( .A1(n19822), .A2(n19773), .B1(n19820), .B2(n19789), .ZN(
        n19772) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19793), .B1(
        n19821), .B2(n19792), .ZN(n19771) );
  OAI211_X1 U22747 ( .C1(n19825), .C2(n19776), .A(n19772), .B(n19771), .ZN(
        P2_U3162) );
  AOI22_X1 U22748 ( .A1(n19828), .A2(n19773), .B1(n19826), .B2(n19789), .ZN(
        n19775) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19793), .B1(
        n19827), .B2(n19792), .ZN(n19774) );
  OAI211_X1 U22750 ( .C1(n19831), .C2(n19776), .A(n19775), .B(n19774), .ZN(
        P2_U3163) );
  AOI22_X1 U22751 ( .A1(n19777), .A2(n19790), .B1(n19832), .B2(n19789), .ZN(
        n19779) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19793), .B1(
        n19833), .B2(n19792), .ZN(n19778) );
  OAI211_X1 U22753 ( .C1(n19780), .C2(n19859), .A(n19779), .B(n19778), .ZN(
        P2_U3164) );
  AOI22_X1 U22754 ( .A1(n19781), .A2(n19790), .B1(n19838), .B2(n19789), .ZN(
        n19783) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19793), .B1(
        n19839), .B2(n19792), .ZN(n19782) );
  OAI211_X1 U22756 ( .C1(n19784), .C2(n19859), .A(n19783), .B(n19782), .ZN(
        P2_U3165) );
  AOI22_X1 U22757 ( .A1(n19785), .A2(n19790), .B1(n19844), .B2(n19789), .ZN(
        n19787) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19793), .B1(
        n19845), .B2(n19792), .ZN(n19786) );
  OAI211_X1 U22759 ( .C1(n19788), .C2(n19859), .A(n19787), .B(n19786), .ZN(
        P2_U3166) );
  AOI22_X1 U22760 ( .A1(n19791), .A2(n19790), .B1(n19850), .B2(n19789), .ZN(
        n19795) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19793), .B1(
        n19852), .B2(n19792), .ZN(n19794) );
  OAI211_X1 U22762 ( .C1(n19796), .C2(n19859), .A(n19795), .B(n19794), .ZN(
        P2_U3167) );
  NAND2_X1 U22763 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19797), .ZN(
        n19805) );
  OR2_X1 U22764 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19805), .ZN(n19799) );
  NOR3_X1 U22765 ( .A1(n10801), .A2(n19851), .A3(n19798), .ZN(n19804) );
  AOI21_X1 U22766 ( .B1(n19798), .B2(n19799), .A(n19804), .ZN(n19853) );
  AOI22_X1 U22767 ( .A1(n19853), .A2(n19801), .B1(n19851), .B2(n19800), .ZN(
        n19812) );
  NAND2_X1 U22768 ( .A1(n19803), .A2(n19802), .ZN(n19806) );
  AOI21_X1 U22769 ( .B1(n19806), .B2(n19805), .A(n19804), .ZN(n19808) );
  OAI211_X1 U22770 ( .C1(n19851), .C2(n19809), .A(n19808), .B(n19807), .ZN(
        n19856) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19810), .ZN(n19811) );
  OAI211_X1 U22772 ( .C1(n19813), .C2(n19859), .A(n19812), .B(n19811), .ZN(
        P2_U3168) );
  AOI22_X1 U22773 ( .A1(n19853), .A2(n19815), .B1(n19851), .B2(n19814), .ZN(
        n19818) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19816), .ZN(n19817) );
  OAI211_X1 U22775 ( .C1(n19819), .C2(n19859), .A(n19818), .B(n19817), .ZN(
        P2_U3169) );
  AOI22_X1 U22776 ( .A1(n19853), .A2(n19821), .B1(n19851), .B2(n19820), .ZN(
        n19824) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19822), .ZN(n19823) );
  OAI211_X1 U22778 ( .C1(n19825), .C2(n19859), .A(n19824), .B(n19823), .ZN(
        P2_U3170) );
  AOI22_X1 U22779 ( .A1(n19853), .A2(n19827), .B1(n19851), .B2(n19826), .ZN(
        n19830) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19828), .ZN(n19829) );
  OAI211_X1 U22781 ( .C1(n19831), .C2(n19859), .A(n19830), .B(n19829), .ZN(
        P2_U3171) );
  AOI22_X1 U22782 ( .A1(n19853), .A2(n19833), .B1(n19851), .B2(n19832), .ZN(
        n19836) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19834), .ZN(n19835) );
  OAI211_X1 U22784 ( .C1(n19837), .C2(n19859), .A(n19836), .B(n19835), .ZN(
        P2_U3172) );
  AOI22_X1 U22785 ( .A1(n19853), .A2(n19839), .B1(n19851), .B2(n19838), .ZN(
        n19842) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19840), .ZN(n19841) );
  OAI211_X1 U22787 ( .C1(n19843), .C2(n19859), .A(n19842), .B(n19841), .ZN(
        P2_U3173) );
  AOI22_X1 U22788 ( .A1(n19853), .A2(n19845), .B1(n19851), .B2(n19844), .ZN(
        n19848) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19846), .ZN(n19847) );
  OAI211_X1 U22790 ( .C1(n19849), .C2(n19859), .A(n19848), .B(n19847), .ZN(
        P2_U3174) );
  AOI22_X1 U22791 ( .A1(n19853), .A2(n19852), .B1(n19851), .B2(n19850), .ZN(
        n19858) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19854), .ZN(n19857) );
  OAI211_X1 U22793 ( .C1(n19860), .C2(n19859), .A(n19858), .B(n19857), .ZN(
        P2_U3175) );
  OAI211_X1 U22794 ( .C1(n19862), .C2(n19861), .A(n19872), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19868) );
  NOR3_X1 U22795 ( .A1(n19872), .A2(n19958), .A3(n19863), .ZN(n19865) );
  OAI21_X1 U22796 ( .B1(n19866), .B2(n19865), .A(n19864), .ZN(n19867) );
  NAND3_X1 U22797 ( .A1(n19869), .A2(n19868), .A3(n19867), .ZN(P2_U3177) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19870), .ZN(
        P2_U3179) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19870), .ZN(
        P2_U3180) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19870), .ZN(
        P2_U3181) );
  AND2_X1 U22801 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19870), .ZN(
        P2_U3182) );
  AND2_X1 U22802 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19870), .ZN(
        P2_U3183) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19870), .ZN(
        P2_U3184) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19870), .ZN(
        P2_U3185) );
  AND2_X1 U22805 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19870), .ZN(
        P2_U3186) );
  AND2_X1 U22806 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19870), .ZN(
        P2_U3187) );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19870), .ZN(
        P2_U3188) );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19870), .ZN(
        P2_U3189) );
  AND2_X1 U22809 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19870), .ZN(
        P2_U3190) );
  AND2_X1 U22810 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19870), .ZN(
        P2_U3191) );
  AND2_X1 U22811 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19870), .ZN(
        P2_U3192) );
  AND2_X1 U22812 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19870), .ZN(
        P2_U3193) );
  AND2_X1 U22813 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19870), .ZN(
        P2_U3194) );
  AND2_X1 U22814 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19870), .ZN(
        P2_U3195) );
  AND2_X1 U22815 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19870), .ZN(
        P2_U3196) );
  AND2_X1 U22816 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19870), .ZN(
        P2_U3197) );
  AND2_X1 U22817 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19870), .ZN(
        P2_U3198) );
  AND2_X1 U22818 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19870), .ZN(
        P2_U3199) );
  AND2_X1 U22819 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19870), .ZN(
        P2_U3200) );
  AND2_X1 U22820 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19870), .ZN(P2_U3201) );
  AND2_X1 U22821 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19870), .ZN(P2_U3202) );
  AND2_X1 U22822 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19870), .ZN(P2_U3203) );
  AND2_X1 U22823 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19870), .ZN(P2_U3204) );
  AND2_X1 U22824 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19870), .ZN(P2_U3205) );
  AND2_X1 U22825 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19870), .ZN(P2_U3206) );
  AND2_X1 U22826 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19870), .ZN(P2_U3207) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19870), .ZN(P2_U3208) );
  OAI21_X1 U22828 ( .B1(n19871), .B2(n19879), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19888) );
  NAND2_X1 U22829 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19872), .ZN(n19886) );
  NAND3_X1 U22830 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19886), .ZN(n19875) );
  AOI211_X1 U22831 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21001), .A(
        n20005), .B(n19873), .ZN(n19874) );
  AOI21_X1 U22832 ( .B1(n19888), .B2(n19875), .A(n19874), .ZN(n19876) );
  INV_X1 U22833 ( .A(n19876), .ZN(P2_U3209) );
  AND2_X1 U22834 ( .A1(n19877), .A2(n19886), .ZN(n19881) );
  NOR2_X1 U22835 ( .A1(HOLD), .A2(n19878), .ZN(n19887) );
  OAI211_X1 U22836 ( .C1(n19887), .C2(n19889), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19879), .ZN(n19880) );
  OAI211_X1 U22837 ( .C1(n19882), .C2(n21001), .A(n19881), .B(n19880), .ZN(
        P2_U3210) );
  OAI22_X1 U22838 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19883), .B1(NA), 
        .B2(n19886), .ZN(n19884) );
  OAI211_X1 U22839 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19884), .ZN(n19885) );
  OAI221_X1 U22840 ( .B1(n19888), .B2(n19887), .C1(n19888), .C2(n19886), .A(
        n19885), .ZN(P2_U3211) );
  OAI222_X1 U22841 ( .A1(n19949), .A2(n19892), .B1(n19891), .B2(n20005), .C1(
        n19890), .C2(n19946), .ZN(P2_U3212) );
  OAI222_X1 U22842 ( .A1(n19949), .A2(n19894), .B1(n19893), .B2(n20005), .C1(
        n19892), .C2(n19946), .ZN(P2_U3213) );
  OAI222_X1 U22843 ( .A1(n19949), .A2(n19896), .B1(n19895), .B2(n20005), .C1(
        n19894), .C2(n19946), .ZN(P2_U3214) );
  OAI222_X1 U22844 ( .A1(n19949), .A2(n19898), .B1(n19897), .B2(n20005), .C1(
        n19896), .C2(n19946), .ZN(P2_U3215) );
  OAI222_X1 U22845 ( .A1(n19949), .A2(n19900), .B1(n19899), .B2(n20005), .C1(
        n19898), .C2(n19946), .ZN(P2_U3216) );
  OAI222_X1 U22846 ( .A1(n19949), .A2(n19902), .B1(n19901), .B2(n20005), .C1(
        n19900), .C2(n19946), .ZN(P2_U3217) );
  INV_X1 U22847 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19904) );
  OAI222_X1 U22848 ( .A1(n19949), .A2(n19904), .B1(n19903), .B2(n20005), .C1(
        n19902), .C2(n19946), .ZN(P2_U3218) );
  OAI222_X1 U22849 ( .A1(n19949), .A2(n19906), .B1(n19905), .B2(n20005), .C1(
        n19904), .C2(n19946), .ZN(P2_U3219) );
  OAI222_X1 U22850 ( .A1(n19949), .A2(n19908), .B1(n19907), .B2(n20005), .C1(
        n19906), .C2(n19946), .ZN(P2_U3220) );
  OAI222_X1 U22851 ( .A1(n19949), .A2(n19910), .B1(n19909), .B2(n20005), .C1(
        n19908), .C2(n19946), .ZN(P2_U3221) );
  OAI222_X1 U22852 ( .A1(n19949), .A2(n19912), .B1(n19911), .B2(n20005), .C1(
        n19910), .C2(n19946), .ZN(P2_U3222) );
  OAI222_X1 U22853 ( .A1(n19949), .A2(n11393), .B1(n19913), .B2(n20005), .C1(
        n19912), .C2(n19946), .ZN(P2_U3223) );
  INV_X1 U22854 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19915) );
  OAI222_X1 U22855 ( .A1(n19949), .A2(n19915), .B1(n19914), .B2(n20005), .C1(
        n11393), .C2(n19946), .ZN(P2_U3224) );
  OAI222_X1 U22856 ( .A1(n19949), .A2(n19917), .B1(n19916), .B2(n20005), .C1(
        n19915), .C2(n19946), .ZN(P2_U3225) );
  OAI222_X1 U22857 ( .A1(n19949), .A2(n19919), .B1(n19918), .B2(n20005), .C1(
        n19917), .C2(n19946), .ZN(P2_U3226) );
  OAI222_X1 U22858 ( .A1(n19949), .A2(n19921), .B1(n19920), .B2(n20005), .C1(
        n19919), .C2(n19946), .ZN(P2_U3227) );
  OAI222_X1 U22859 ( .A1(n19949), .A2(n19923), .B1(n19922), .B2(n20005), .C1(
        n19921), .C2(n19946), .ZN(P2_U3228) );
  OAI222_X1 U22860 ( .A1(n19949), .A2(n19925), .B1(n19924), .B2(n20005), .C1(
        n19923), .C2(n19946), .ZN(P2_U3229) );
  OAI222_X1 U22861 ( .A1(n19949), .A2(n19927), .B1(n19926), .B2(n20005), .C1(
        n19925), .C2(n19946), .ZN(P2_U3230) );
  OAI222_X1 U22862 ( .A1(n19949), .A2(n19929), .B1(n19928), .B2(n20005), .C1(
        n19927), .C2(n19946), .ZN(P2_U3231) );
  OAI222_X1 U22863 ( .A1(n19949), .A2(n15188), .B1(n19930), .B2(n20005), .C1(
        n19929), .C2(n19946), .ZN(P2_U3232) );
  INV_X1 U22864 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19932) );
  OAI222_X1 U22865 ( .A1(n19949), .A2(n19932), .B1(n19931), .B2(n20005), .C1(
        n15188), .C2(n19946), .ZN(P2_U3233) );
  OAI222_X1 U22866 ( .A1(n19949), .A2(n19934), .B1(n19933), .B2(n20005), .C1(
        n19932), .C2(n19946), .ZN(P2_U3234) );
  OAI222_X1 U22867 ( .A1(n19949), .A2(n19936), .B1(n19935), .B2(n20005), .C1(
        n19934), .C2(n19946), .ZN(P2_U3235) );
  OAI222_X1 U22868 ( .A1(n19949), .A2(n19938), .B1(n19937), .B2(n20005), .C1(
        n19936), .C2(n19946), .ZN(P2_U3236) );
  INV_X1 U22869 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19941) );
  OAI222_X1 U22870 ( .A1(n19949), .A2(n19941), .B1(n19939), .B2(n20005), .C1(
        n19938), .C2(n19946), .ZN(P2_U3237) );
  OAI222_X1 U22871 ( .A1(n19946), .A2(n19941), .B1(n19940), .B2(n20005), .C1(
        n19942), .C2(n19949), .ZN(P2_U3238) );
  OAI222_X1 U22872 ( .A1(n19949), .A2(n19944), .B1(n19943), .B2(n20005), .C1(
        n19942), .C2(n19946), .ZN(P2_U3239) );
  INV_X1 U22873 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19947) );
  OAI222_X1 U22874 ( .A1(n19949), .A2(n19947), .B1(n19945), .B2(n20005), .C1(
        n19944), .C2(n19946), .ZN(P2_U3240) );
  INV_X1 U22875 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19948) );
  OAI222_X1 U22876 ( .A1(n19949), .A2(n11194), .B1(n19948), .B2(n20005), .C1(
        n19947), .C2(n19946), .ZN(P2_U3241) );
  OAI22_X1 U22877 ( .A1(n20006), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20005), .ZN(n19950) );
  INV_X1 U22878 ( .A(n19950), .ZN(P2_U3585) );
  MUX2_X1 U22879 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20006), .Z(P2_U3586) );
  OAI22_X1 U22880 ( .A1(n20006), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20005), .ZN(n19951) );
  INV_X1 U22881 ( .A(n19951), .ZN(P2_U3587) );
  OAI22_X1 U22882 ( .A1(n20006), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20005), .ZN(n19952) );
  INV_X1 U22883 ( .A(n19952), .ZN(P2_U3588) );
  OAI21_X1 U22884 ( .B1(n19956), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19954), 
        .ZN(n19953) );
  INV_X1 U22885 ( .A(n19953), .ZN(P2_U3591) );
  OAI21_X1 U22886 ( .B1(n19956), .B2(n19955), .A(n19954), .ZN(P2_U3592) );
  NAND2_X1 U22887 ( .A1(n19957), .A2(n19974), .ZN(n19967) );
  NAND3_X1 U22888 ( .A1(n19981), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19958), 
        .ZN(n19959) );
  NAND2_X1 U22889 ( .A1(n19959), .A2(n19985), .ZN(n19968) );
  NAND2_X1 U22890 ( .A1(n19967), .A2(n19968), .ZN(n19964) );
  AOI222_X1 U22891 ( .A1(n19964), .A2(n19963), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19962), .C1(n19961), .C2(n19960), .ZN(n19965) );
  AOI22_X1 U22892 ( .A1(n19995), .A2(n19966), .B1(n19965), .B2(n19992), .ZN(
        P2_U3602) );
  OAI21_X1 U22893 ( .B1(n19969), .B2(n19968), .A(n19967), .ZN(n19970) );
  AOI21_X1 U22894 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19971), .A(n19970), 
        .ZN(n19972) );
  AOI22_X1 U22895 ( .A1(n19995), .A2(n19973), .B1(n19972), .B2(n19992), .ZN(
        P2_U3603) );
  INV_X1 U22896 ( .A(n19974), .ZN(n19980) );
  INV_X1 U22897 ( .A(n19975), .ZN(n19976) );
  NAND3_X1 U22898 ( .A1(n19981), .A2(n19985), .A3(n19976), .ZN(n19979) );
  NAND2_X1 U22899 ( .A1(n19977), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19978) );
  OAI211_X1 U22900 ( .C1(n19981), .C2(n19980), .A(n19979), .B(n19978), .ZN(
        n19982) );
  INV_X1 U22901 ( .A(n19982), .ZN(n19983) );
  AOI22_X1 U22902 ( .A1(n19995), .A2(n19984), .B1(n19983), .B2(n19992), .ZN(
        P2_U3604) );
  INV_X1 U22903 ( .A(n19985), .ZN(n19987) );
  OAI21_X1 U22904 ( .B1(n19988), .B2(n19987), .A(n19986), .ZN(n19989) );
  AOI21_X1 U22905 ( .B1(n19991), .B2(n19990), .A(n19989), .ZN(n19993) );
  AOI22_X1 U22906 ( .A1(n19995), .A2(n19994), .B1(n19993), .B2(n19992), .ZN(
        P2_U3605) );
  INV_X1 U22907 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19996) );
  AOI22_X1 U22908 ( .A1(n20005), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19996), 
        .B2(n20006), .ZN(P2_U3608) );
  AOI22_X1 U22909 ( .A1(n20000), .A2(n19999), .B1(n19998), .B2(n19997), .ZN(
        n20001) );
  NAND2_X1 U22910 ( .A1(n20002), .A2(n20001), .ZN(n20004) );
  MUX2_X1 U22911 ( .A(P2_MORE_REG_SCAN_IN), .B(n20004), .S(n20003), .Z(
        P2_U3609) );
  OAI22_X1 U22912 ( .A1(n20006), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20005), .ZN(n20007) );
  INV_X1 U22913 ( .A(n20007), .ZN(P2_U3611) );
  AOI21_X1 U22914 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20782), .A(n20776), 
        .ZN(n20778) );
  INV_X1 U22915 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21226) );
  AOI21_X1 U22916 ( .B1(n20778), .B2(n21226), .A(n20887), .ZN(P1_U2802) );
  OAI21_X1 U22917 ( .B1(n20009), .B2(n20008), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20010) );
  OAI21_X1 U22918 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20011), .A(n20010), 
        .ZN(P1_U2803) );
  INV_X1 U22919 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n21053) );
  NOR2_X1 U22920 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20013) );
  NOR2_X1 U22921 ( .A1(n20887), .A2(n20013), .ZN(n20012) );
  AOI22_X1 U22922 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20887), .B1(n21053), 
        .B2(n20012), .ZN(P1_U2804) );
  NOR2_X1 U22923 ( .A1(n20887), .A2(n20778), .ZN(n20829) );
  OAI21_X1 U22924 ( .B1(BS16), .B2(n20013), .A(n20829), .ZN(n20827) );
  OAI21_X1 U22925 ( .B1(n20829), .B2(n21003), .A(n20827), .ZN(P1_U2805) );
  OAI21_X1 U22926 ( .B1(n20015), .B2(n20014), .A(n20155), .ZN(P1_U2806) );
  NOR4_X1 U22927 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20019) );
  NOR4_X1 U22928 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20018) );
  NOR4_X1 U22929 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20017) );
  NOR4_X1 U22930 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20016) );
  NAND4_X1 U22931 ( .A1(n20019), .A2(n20018), .A3(n20017), .A4(n20016), .ZN(
        n20025) );
  NOR4_X1 U22932 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20023) );
  AOI211_X1 U22933 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20022) );
  NOR4_X1 U22934 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20021) );
  NOR4_X1 U22935 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20020) );
  NAND4_X1 U22936 ( .A1(n20023), .A2(n20022), .A3(n20021), .A4(n20020), .ZN(
        n20024) );
  NOR2_X1 U22937 ( .A1(n20025), .A2(n20024), .ZN(n20870) );
  INV_X1 U22938 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20993) );
  NOR3_X1 U22939 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20027) );
  OAI21_X1 U22940 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20027), .A(n20870), .ZN(
        n20026) );
  OAI21_X1 U22941 ( .B1(n20870), .B2(n20993), .A(n20026), .ZN(P1_U2807) );
  INV_X1 U22942 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20828) );
  AOI21_X1 U22943 ( .B1(n20867), .B2(n20828), .A(n20027), .ZN(n20028) );
  INV_X1 U22944 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20978) );
  INV_X1 U22945 ( .A(n20870), .ZN(n20872) );
  AOI22_X1 U22946 ( .A1(n20870), .A2(n20028), .B1(n20978), .B2(n20872), .ZN(
        P1_U2808) );
  OAI21_X1 U22947 ( .B1(n20030), .B2(n20031), .A(n20029), .ZN(n20045) );
  AOI22_X1 U22948 ( .A1(n10462), .A2(n20070), .B1(n20043), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20039) );
  NOR3_X1 U22949 ( .A1(n20032), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n20031), .ZN(
        n20037) );
  INV_X1 U22950 ( .A(n20033), .ZN(n20034) );
  NAND2_X1 U22951 ( .A1(n20073), .A2(n20034), .ZN(n20035) );
  OAI211_X1 U22952 ( .C1(n11881), .C2(n20057), .A(n20035), .B(n20055), .ZN(
        n20036) );
  AOI211_X1 U22953 ( .C1(n20082), .C2(n20047), .A(n20037), .B(n20036), .ZN(
        n20038) );
  OAI211_X1 U22954 ( .C1(n20045), .C2(n21181), .A(n20039), .B(n20038), .ZN(
        P1_U2833) );
  AOI22_X1 U22955 ( .A1(n20070), .A2(n20040), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20069), .ZN(n20052) );
  INV_X1 U22956 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20967) );
  INV_X1 U22957 ( .A(n20041), .ZN(n20042) );
  AOI22_X1 U22958 ( .A1(n20043), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n20042), .B2(
        n20073), .ZN(n20044) );
  OAI21_X1 U22959 ( .B1(n20045), .B2(n20967), .A(n20044), .ZN(n20046) );
  AOI21_X1 U22960 ( .B1(n20048), .B2(n20047), .A(n20046), .ZN(n20051) );
  NAND3_X1 U22961 ( .A1(n20077), .A2(n20049), .A3(n20967), .ZN(n20050) );
  NAND4_X1 U22962 ( .A1(n20052), .A2(n20051), .A3(n20055), .A4(n20050), .ZN(
        P1_U2834) );
  INV_X1 U22963 ( .A(n20053), .ZN(n20054) );
  NAND3_X1 U22964 ( .A1(n20077), .A2(n20951), .A3(n20054), .ZN(n20065) );
  OAI21_X1 U22965 ( .B1(n20057), .B2(n20056), .A(n20055), .ZN(n20061) );
  NOR2_X1 U22966 ( .A1(n20059), .A2(n20058), .ZN(n20060) );
  NOR2_X1 U22967 ( .A1(n20061), .A2(n20060), .ZN(n20064) );
  NAND2_X1 U22968 ( .A1(n20070), .A2(n20084), .ZN(n20063) );
  NAND2_X1 U22969 ( .A1(n20043), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20062) );
  NAND4_X1 U22970 ( .A1(n20065), .A2(n20064), .A3(n20063), .A4(n20062), .ZN(
        n20066) );
  AOI21_X1 U22971 ( .B1(n20085), .B2(n20076), .A(n20066), .ZN(n20067) );
  OAI21_X1 U22972 ( .B1(n20951), .B2(n20068), .A(n20067), .ZN(P1_U2835) );
  AOI222_X1 U22973 ( .A1(n20850), .A2(n20071), .B1(n20070), .B2(n20087), .C1(
        n20069), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20081) );
  INV_X1 U22974 ( .A(n20072), .ZN(n20074) );
  AOI22_X1 U22975 ( .A1(n20043), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20074), .B2(
        n20073), .ZN(n20080) );
  AOI22_X1 U22976 ( .A1(n20090), .A2(n20076), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n20075), .ZN(n20079) );
  INV_X1 U22977 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20786) );
  NAND4_X1 U22978 ( .A1(n20077), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n20786), .ZN(n20078) );
  NAND4_X1 U22979 ( .A1(n20081), .A2(n20080), .A3(n20079), .A4(n20078), .ZN(
        P1_U2837) );
  AOI22_X1 U22980 ( .A1(n20082), .A2(n20089), .B1(n20088), .B2(n10462), .ZN(
        n20083) );
  OAI21_X1 U22981 ( .B1(n20092), .B2(n21021), .A(n20083), .ZN(P1_U2865) );
  AOI22_X1 U22982 ( .A1(n20085), .A2(n20089), .B1(n20088), .B2(n20084), .ZN(
        n20086) );
  OAI21_X1 U22983 ( .B1(n20092), .B2(n21242), .A(n20086), .ZN(P1_U2867) );
  AOI22_X1 U22984 ( .A1(n20090), .A2(n20089), .B1(n20088), .B2(n20087), .ZN(
        n20091) );
  OAI21_X1 U22985 ( .B1(n20092), .B2(n12340), .A(n20091), .ZN(P1_U2869) );
  AOI22_X1 U22986 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20095), .B1(n15907), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20093) );
  OAI21_X1 U22987 ( .B1(n20094), .B2(n20877), .A(n20093), .ZN(P1_U2921) );
  INV_X1 U22988 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20097) );
  AOI22_X1 U22989 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20096) );
  OAI21_X1 U22990 ( .B1(n20097), .B2(n20122), .A(n20096), .ZN(P1_U2922) );
  INV_X1 U22991 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20099) );
  AOI22_X1 U22992 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20098) );
  OAI21_X1 U22993 ( .B1(n20099), .B2(n20122), .A(n20098), .ZN(P1_U2923) );
  INV_X1 U22994 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20101) );
  AOI22_X1 U22995 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20100) );
  OAI21_X1 U22996 ( .B1(n20101), .B2(n20122), .A(n20100), .ZN(P1_U2924) );
  INV_X1 U22997 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20103) );
  AOI22_X1 U22998 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20102) );
  OAI21_X1 U22999 ( .B1(n20103), .B2(n20122), .A(n20102), .ZN(P1_U2925) );
  AOI22_X1 U23000 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20104) );
  OAI21_X1 U23001 ( .B1(n14001), .B2(n20122), .A(n20104), .ZN(P1_U2926) );
  INV_X1 U23002 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20106) );
  AOI22_X1 U23003 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20105) );
  OAI21_X1 U23004 ( .B1(n20106), .B2(n20122), .A(n20105), .ZN(P1_U2927) );
  AOI22_X1 U23005 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20107) );
  OAI21_X1 U23006 ( .B1(n20108), .B2(n20122), .A(n20107), .ZN(P1_U2928) );
  INV_X1 U23007 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U23008 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20109) );
  OAI21_X1 U23009 ( .B1(n20110), .B2(n20122), .A(n20109), .ZN(P1_U2929) );
  AOI22_X1 U23010 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20111) );
  OAI21_X1 U23011 ( .B1(n11870), .B2(n20122), .A(n20111), .ZN(P1_U2930) );
  AOI22_X1 U23012 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20112) );
  OAI21_X1 U23013 ( .B1(n13566), .B2(n20122), .A(n20112), .ZN(P1_U2931) );
  AOI22_X1 U23014 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20113) );
  OAI21_X1 U23015 ( .B1(n20114), .B2(n20122), .A(n20113), .ZN(P1_U2932) );
  AOI22_X1 U23016 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20115) );
  OAI21_X1 U23017 ( .B1(n13462), .B2(n20122), .A(n20115), .ZN(P1_U2933) );
  AOI22_X1 U23018 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20116) );
  OAI21_X1 U23019 ( .B1(n20117), .B2(n20122), .A(n20116), .ZN(P1_U2934) );
  AOI22_X1 U23020 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U23021 ( .B1(n20119), .B2(n20122), .A(n20118), .ZN(P1_U2935) );
  AOI22_X1 U23022 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20120), .B1(n15907), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23023 ( .B1(n20123), .B2(n20122), .A(n20121), .ZN(P1_U2936) );
  AOI22_X1 U23024 ( .A1(n20135), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20134), .ZN(n20125) );
  NAND2_X1 U23025 ( .A1(n20125), .A2(n20124), .ZN(P1_U2961) );
  AOI22_X1 U23026 ( .A1(n20135), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20134), .ZN(n20127) );
  NAND2_X1 U23027 ( .A1(n20127), .A2(n20126), .ZN(P1_U2962) );
  AOI22_X1 U23028 ( .A1(n20135), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20134), .ZN(n20129) );
  NAND2_X1 U23029 ( .A1(n20129), .A2(n20128), .ZN(P1_U2963) );
  AOI22_X1 U23030 ( .A1(n20135), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20134), .ZN(n20131) );
  NAND2_X1 U23031 ( .A1(n20131), .A2(n20130), .ZN(P1_U2964) );
  AOI22_X1 U23032 ( .A1(n20135), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20134), .ZN(n20133) );
  NAND2_X1 U23033 ( .A1(n20133), .A2(n20132), .ZN(P1_U2965) );
  AOI22_X1 U23034 ( .A1(n20135), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20134), .ZN(n20137) );
  NAND2_X1 U23035 ( .A1(n20137), .A2(n20136), .ZN(P1_U2966) );
  OAI21_X1 U23036 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20139), .A(
        n20138), .ZN(n20165) );
  NOR2_X1 U23037 ( .A1(n20140), .A2(n20867), .ZN(n20159) );
  OAI22_X1 U23038 ( .A1(n20143), .A2(n20142), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20141), .ZN(n20144) );
  AOI211_X1 U23039 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20152), .A(
        n20159), .B(n20144), .ZN(n20145) );
  OAI21_X1 U23040 ( .B1(n20155), .B2(n20165), .A(n20145), .ZN(P1_U2998) );
  OAI21_X1 U23041 ( .B1(n20147), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n20146), .ZN(n20175) );
  INV_X1 U23042 ( .A(n20148), .ZN(n20150) );
  AND2_X1 U23043 ( .A1(n20149), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20168) );
  AOI21_X1 U23044 ( .B1(n20150), .B2(n20178), .A(n20168), .ZN(n20154) );
  OAI21_X1 U23045 ( .B1(n20152), .B2(n20151), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20153) );
  OAI211_X1 U23046 ( .C1(n20175), .C2(n20155), .A(n20154), .B(n20153), .ZN(
        P1_U2999) );
  AND3_X1 U23047 ( .A1(n20157), .A2(n20156), .A3(n12328), .ZN(n20158) );
  AOI211_X1 U23048 ( .C1(n20160), .C2(n20169), .A(n20159), .B(n20158), .ZN(
        n20164) );
  AOI21_X1 U23049 ( .B1(n20162), .B2(n20161), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20167) );
  OAI21_X1 U23050 ( .B1(n20171), .B2(n20167), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20163) );
  OAI211_X1 U23051 ( .C1(n20165), .C2(n20176), .A(n20164), .B(n20163), .ZN(
        P1_U3030) );
  INV_X1 U23052 ( .A(n20166), .ZN(n20170) );
  AOI211_X1 U23053 ( .C1(n20170), .C2(n20169), .A(n20168), .B(n20167), .ZN(
        n20174) );
  OAI21_X1 U23054 ( .B1(n20172), .B2(n20171), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20173) );
  OAI211_X1 U23055 ( .C1(n20176), .C2(n20175), .A(n20174), .B(n20173), .ZN(
        P1_U3031) );
  NOR2_X1 U23056 ( .A1(n12265), .A2(n20857), .ZN(P1_U3032) );
  NAND2_X1 U23057 ( .A1(n20178), .A2(n20177), .ZN(n20219) );
  INV_X1 U23058 ( .A(n20219), .ZN(n20224) );
  NAND2_X1 U23059 ( .A1(n20179), .A2(n20178), .ZN(n20218) );
  INV_X1 U23060 ( .A(n20218), .ZN(n20225) );
  AOI22_X1 U23061 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20224), .B1(DATAI_16_), 
        .B2(n20225), .ZN(n20671) );
  AOI22_X2 U23062 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20224), .B1(DATAI_24_), 
        .B2(n20225), .ZN(n20716) );
  NAND2_X1 U23063 ( .A1(n20226), .A2(n11627), .ZN(n20583) );
  NOR3_X1 U23064 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20239) );
  NAND2_X1 U23065 ( .A1(n20866), .A2(n20239), .ZN(n20227) );
  OAI22_X1 U23066 ( .A1(n20735), .A2(n20716), .B1(n20583), .B2(n20227), .ZN(
        n20182) );
  INV_X1 U23067 ( .A(n20182), .ZN(n20194) );
  INV_X1 U23068 ( .A(n20259), .ZN(n20183) );
  OAI21_X1 U23069 ( .B1(n20183), .B2(n20760), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20184) );
  NAND2_X1 U23070 ( .A1(n20184), .A2(n20858), .ZN(n20192) );
  OR2_X1 U23071 ( .A1(n20850), .A2(n20459), .ZN(n20265) );
  NOR2_X1 U23072 ( .A1(n20265), .A2(n20660), .ZN(n20188) );
  NAND2_X1 U23073 ( .A1(n20190), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20661) );
  AND2_X1 U23074 ( .A1(n20342), .A2(n20661), .ZN(n20518) );
  INV_X1 U23075 ( .A(n20461), .ZN(n20185) );
  NAND2_X1 U23076 ( .A1(n20185), .A2(n20520), .ZN(n20337) );
  AOI22_X1 U23077 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20337), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20227), .ZN(n20186) );
  OAI211_X1 U23078 ( .C1(n20192), .C2(n20188), .A(n20518), .B(n20186), .ZN(
        n20232) );
  NOR2_X2 U23079 ( .A1(n20187), .A2(n20236), .ZN(n20705) );
  INV_X1 U23080 ( .A(n20188), .ZN(n20191) );
  OR2_X1 U23081 ( .A1(n20190), .A2(n20189), .ZN(n20522) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20232), .B1(
        n20705), .B2(n20231), .ZN(n20193) );
  OAI211_X1 U23083 ( .C1(n20671), .C2(n20259), .A(n20194), .B(n20193), .ZN(
        P1_U3033) );
  AOI22_X1 U23084 ( .A1(DATAI_17_), .A2(n20225), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20224), .ZN(n20675) );
  AOI22_X2 U23085 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20224), .B1(DATAI_25_), 
        .B2(n20225), .ZN(n20722) );
  NAND2_X1 U23086 ( .A1(n20226), .A2(n11616), .ZN(n20595) );
  OAI22_X1 U23087 ( .A1(n20735), .A2(n20722), .B1(n20595), .B2(n20227), .ZN(
        n20195) );
  INV_X1 U23088 ( .A(n20195), .ZN(n20198) );
  NOR2_X2 U23089 ( .A1(n20196), .A2(n20236), .ZN(n20717) );
  AOI22_X1 U23090 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20232), .B1(
        n20717), .B2(n20231), .ZN(n20197) );
  OAI211_X1 U23091 ( .C1(n20675), .C2(n20259), .A(n20198), .B(n20197), .ZN(
        P1_U3034) );
  INV_X1 U23092 ( .A(DATAI_18_), .ZN(n21198) );
  OAI22_X1 U23093 ( .A1(n20199), .A2(n20219), .B1(n21198), .B2(n20218), .ZN(
        n20639) );
  INV_X1 U23094 ( .A(n20639), .ZN(n20728) );
  NAND2_X1 U23095 ( .A1(n20226), .A2(n11618), .ZN(n20599) );
  OAI22_X1 U23096 ( .A1(n20735), .A2(n20642), .B1(n20599), .B2(n20227), .ZN(
        n20200) );
  INV_X1 U23097 ( .A(n20200), .ZN(n20203) );
  NOR2_X2 U23098 ( .A1(n20201), .A2(n20236), .ZN(n20723) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20232), .B1(
        n20723), .B2(n20231), .ZN(n20202) );
  OAI211_X1 U23100 ( .C1(n20728), .C2(n20259), .A(n20203), .B(n20202), .ZN(
        P1_U3035) );
  INV_X1 U23101 ( .A(DATAI_19_), .ZN(n21005) );
  OAI22_X1 U23102 ( .A1(n15093), .A2(n20219), .B1(n21005), .B2(n20218), .ZN(
        n20643) );
  INV_X1 U23103 ( .A(n20643), .ZN(n20736) );
  AOI22_X1 U23104 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20224), .B1(DATAI_27_), 
        .B2(n20225), .ZN(n20646) );
  NAND2_X1 U23105 ( .A1(n20226), .A2(n20204), .ZN(n20603) );
  OAI22_X1 U23106 ( .A1(n20735), .A2(n20646), .B1(n20603), .B2(n20227), .ZN(
        n20205) );
  INV_X1 U23107 ( .A(n20205), .ZN(n20208) );
  NOR2_X2 U23108 ( .A1(n20206), .A2(n20236), .ZN(n20729) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20232), .B1(
        n20729), .B2(n20231), .ZN(n20207) );
  OAI211_X1 U23110 ( .C1(n20736), .C2(n20259), .A(n20208), .B(n20207), .ZN(
        P1_U3036) );
  INV_X1 U23111 ( .A(DATAI_20_), .ZN(n21024) );
  OAI22_X1 U23112 ( .A1(n21024), .A2(n20218), .B1(n15086), .B2(n20219), .ZN(
        n20739) );
  AOI22_X2 U23113 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20224), .B1(DATAI_28_), 
        .B2(n20225), .ZN(n20742) );
  NAND2_X1 U23114 ( .A1(n20226), .A2(n11609), .ZN(n20607) );
  OAI22_X1 U23115 ( .A1(n20735), .A2(n20742), .B1(n20607), .B2(n20227), .ZN(
        n20209) );
  INV_X1 U23116 ( .A(n20209), .ZN(n20212) );
  NOR2_X2 U23117 ( .A1(n20210), .A2(n20236), .ZN(n20737) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20232), .B1(
        n20737), .B2(n20231), .ZN(n20211) );
  OAI211_X1 U23119 ( .C1(n20683), .C2(n20259), .A(n20212), .B(n20211), .ZN(
        P1_U3037) );
  INV_X1 U23120 ( .A(DATAI_21_), .ZN(n21158) );
  OAI22_X1 U23121 ( .A1(n21158), .A2(n20218), .B1(n15074), .B2(n20219), .ZN(
        n20745) );
  INV_X1 U23122 ( .A(n20745), .ZN(n20687) );
  AOI22_X2 U23123 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20224), .B1(DATAI_29_), 
        .B2(n20225), .ZN(n20748) );
  NAND2_X1 U23124 ( .A1(n20226), .A2(n20213), .ZN(n20539) );
  OAI22_X1 U23125 ( .A1(n20735), .A2(n20748), .B1(n20539), .B2(n20227), .ZN(
        n20214) );
  INV_X1 U23126 ( .A(n20214), .ZN(n20217) );
  NOR2_X2 U23127 ( .A1(n20215), .A2(n20236), .ZN(n20743) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20232), .B1(
        n20743), .B2(n20231), .ZN(n20216) );
  OAI211_X1 U23129 ( .C1(n20687), .C2(n20259), .A(n20217), .B(n20216), .ZN(
        P1_U3038) );
  INV_X1 U23130 ( .A(DATAI_22_), .ZN(n21152) );
  OAI22_X1 U23131 ( .A1(n15067), .A2(n20219), .B1(n21152), .B2(n20218), .ZN(
        n20751) );
  INV_X1 U23132 ( .A(n20751), .ZN(n20691) );
  AOI22_X2 U23133 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20224), .B1(DATAI_30_), 
        .B2(n20225), .ZN(n20754) );
  NAND2_X1 U23134 ( .A1(n20226), .A2(n11540), .ZN(n20615) );
  OAI22_X1 U23135 ( .A1(n20735), .A2(n20754), .B1(n20615), .B2(n20227), .ZN(
        n20220) );
  INV_X1 U23136 ( .A(n20220), .ZN(n20223) );
  NOR2_X2 U23137 ( .A1(n20236), .A2(n20221), .ZN(n20749) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20232), .B1(
        n20749), .B2(n20231), .ZN(n20222) );
  OAI211_X1 U23139 ( .C1(n20691), .C2(n20259), .A(n20223), .B(n20222), .ZN(
        P1_U3039) );
  AOI22_X1 U23140 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20224), .B1(DATAI_23_), 
        .B2(n20225), .ZN(n20699) );
  NAND2_X1 U23141 ( .A1(n20226), .A2(n11554), .ZN(n20620) );
  OAI22_X1 U23142 ( .A1(n20735), .A2(n20765), .B1(n20620), .B2(n20227), .ZN(
        n20228) );
  INV_X1 U23143 ( .A(n20228), .ZN(n20234) );
  INV_X1 U23144 ( .A(n20229), .ZN(n20230) );
  NOR2_X2 U23145 ( .A1(n20236), .A2(n20230), .ZN(n20756) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20232), .B1(
        n20756), .B2(n20231), .ZN(n20233) );
  OAI211_X1 U23147 ( .C1(n20699), .C2(n20259), .A(n20234), .B(n20233), .ZN(
        P1_U3040) );
  INV_X1 U23148 ( .A(n20239), .ZN(n20235) );
  NOR2_X1 U23149 ( .A1(n20866), .A2(n20235), .ZN(n20255) );
  INV_X1 U23150 ( .A(n20265), .ZN(n20300) );
  INV_X1 U23151 ( .A(n20364), .ZN(n20627) );
  AOI21_X1 U23152 ( .B1(n20300), .B2(n20627), .A(n20255), .ZN(n20237) );
  OAI22_X1 U23153 ( .A1(n20237), .A2(n20852), .B1(n20235), .B2(n20703), .ZN(
        n20254) );
  AOI22_X1 U23154 ( .A1(n20706), .A2(n20255), .B1(n20705), .B2(n20254), .ZN(
        n20241) );
  OR2_X1 U23155 ( .A1(n13427), .A2(n21003), .ZN(n20629) );
  OAI211_X1 U23156 ( .C1(n20298), .C2(n20629), .A(n20858), .B(n20237), .ZN(
        n20238) );
  OAI211_X1 U23157 ( .C1(n20858), .C2(n20239), .A(n20710), .B(n20238), .ZN(
        n20256) );
  OR2_X1 U23158 ( .A1(n13427), .A2(n20260), .ZN(n20634) );
  INV_X1 U23159 ( .A(n20671), .ZN(n20713) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20713), .ZN(n20240) );
  OAI211_X1 U23161 ( .C1(n20716), .C2(n20259), .A(n20241), .B(n20240), .ZN(
        P1_U3041) );
  AOI22_X1 U23162 ( .A1(n20718), .A2(n20255), .B1(n20717), .B2(n20254), .ZN(
        n20243) );
  INV_X1 U23163 ( .A(n20675), .ZN(n20719) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20719), .ZN(n20242) );
  OAI211_X1 U23165 ( .C1(n20722), .C2(n20259), .A(n20243), .B(n20242), .ZN(
        P1_U3042) );
  AOI22_X1 U23166 ( .A1(n20724), .A2(n20255), .B1(n20723), .B2(n20254), .ZN(
        n20245) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20639), .ZN(n20244) );
  OAI211_X1 U23168 ( .C1(n20642), .C2(n20259), .A(n20245), .B(n20244), .ZN(
        P1_U3043) );
  AOI22_X1 U23169 ( .A1(n20730), .A2(n20255), .B1(n20729), .B2(n20254), .ZN(
        n20247) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20643), .ZN(n20246) );
  OAI211_X1 U23171 ( .C1(n20646), .C2(n20259), .A(n20247), .B(n20246), .ZN(
        P1_U3044) );
  AOI22_X1 U23172 ( .A1(n20738), .A2(n20255), .B1(n20737), .B2(n20254), .ZN(
        n20249) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20739), .ZN(n20248) );
  OAI211_X1 U23174 ( .C1(n20742), .C2(n20259), .A(n20249), .B(n20248), .ZN(
        P1_U3045) );
  AOI22_X1 U23175 ( .A1(n20744), .A2(n20255), .B1(n20743), .B2(n20254), .ZN(
        n20251) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20745), .ZN(n20250) );
  OAI211_X1 U23177 ( .C1(n20748), .C2(n20259), .A(n20251), .B(n20250), .ZN(
        P1_U3046) );
  AOI22_X1 U23178 ( .A1(n20750), .A2(n20255), .B1(n20749), .B2(n20254), .ZN(
        n20253) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20751), .ZN(n20252) );
  OAI211_X1 U23180 ( .C1(n20754), .C2(n20259), .A(n20253), .B(n20252), .ZN(
        P1_U3047) );
  AOI22_X1 U23181 ( .A1(n20758), .A2(n20255), .B1(n20756), .B2(n20254), .ZN(
        n20258) );
  INV_X1 U23182 ( .A(n20699), .ZN(n20759) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20256), .B1(
        n20262), .B2(n20759), .ZN(n20257) );
  OAI211_X1 U23184 ( .C1(n20765), .C2(n20259), .A(n20258), .B(n20257), .ZN(
        P1_U3048) );
  NAND3_X1 U23185 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20856), .A3(
        n15856), .ZN(n20304) );
  OR2_X1 U23186 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20304), .ZN(
        n20290) );
  OAI22_X1 U23187 ( .A1(n20328), .A2(n20671), .B1(n20583), .B2(n20290), .ZN(
        n20261) );
  INV_X1 U23188 ( .A(n20261), .ZN(n20271) );
  INV_X1 U23189 ( .A(n20328), .ZN(n20263) );
  OAI21_X1 U23190 ( .B1(n20263), .B2(n20262), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20264) );
  NAND2_X1 U23191 ( .A1(n20264), .A2(n20858), .ZN(n20269) );
  NOR2_X1 U23192 ( .A1(n20265), .A2(n20586), .ZN(n20267) );
  OR2_X1 U23193 ( .A1(n20520), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20396) );
  AND2_X1 U23194 ( .A1(n20396), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20393) );
  AOI21_X1 U23195 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20290), .A(n20393), 
        .ZN(n20266) );
  OAI211_X1 U23196 ( .C1(n20269), .C2(n20267), .A(n20518), .B(n20266), .ZN(
        n20294) );
  INV_X1 U23197 ( .A(n20267), .ZN(n20268) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20294), .B1(
        n20705), .B2(n20293), .ZN(n20270) );
  OAI211_X1 U23199 ( .C1(n20716), .C2(n20291), .A(n20271), .B(n20270), .ZN(
        P1_U3049) );
  OAI22_X1 U23200 ( .A1(n20328), .A2(n20675), .B1(n20290), .B2(n20595), .ZN(
        n20272) );
  INV_X1 U23201 ( .A(n20272), .ZN(n20274) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20294), .B1(
        n20717), .B2(n20293), .ZN(n20273) );
  OAI211_X1 U23203 ( .C1(n20722), .C2(n20291), .A(n20274), .B(n20273), .ZN(
        P1_U3050) );
  OAI22_X1 U23204 ( .A1(n20291), .A2(n20642), .B1(n20290), .B2(n20599), .ZN(
        n20275) );
  INV_X1 U23205 ( .A(n20275), .ZN(n20277) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20294), .B1(
        n20723), .B2(n20293), .ZN(n20276) );
  OAI211_X1 U23207 ( .C1(n20728), .C2(n20328), .A(n20277), .B(n20276), .ZN(
        P1_U3051) );
  OAI22_X1 U23208 ( .A1(n20328), .A2(n20736), .B1(n20290), .B2(n20603), .ZN(
        n20278) );
  INV_X1 U23209 ( .A(n20278), .ZN(n20280) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20294), .B1(
        n20729), .B2(n20293), .ZN(n20279) );
  OAI211_X1 U23211 ( .C1(n20646), .C2(n20291), .A(n20280), .B(n20279), .ZN(
        P1_U3052) );
  OAI22_X1 U23212 ( .A1(n20328), .A2(n20683), .B1(n20290), .B2(n20607), .ZN(
        n20281) );
  INV_X1 U23213 ( .A(n20281), .ZN(n20283) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20294), .B1(
        n20737), .B2(n20293), .ZN(n20282) );
  OAI211_X1 U23215 ( .C1(n20742), .C2(n20291), .A(n20283), .B(n20282), .ZN(
        P1_U3053) );
  OAI22_X1 U23216 ( .A1(n20291), .A2(n20748), .B1(n20290), .B2(n20539), .ZN(
        n20284) );
  INV_X1 U23217 ( .A(n20284), .ZN(n20286) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20294), .B1(
        n20743), .B2(n20293), .ZN(n20285) );
  OAI211_X1 U23219 ( .C1(n20687), .C2(n20328), .A(n20286), .B(n20285), .ZN(
        P1_U3054) );
  OAI22_X1 U23220 ( .A1(n20291), .A2(n20754), .B1(n20290), .B2(n20615), .ZN(
        n20287) );
  INV_X1 U23221 ( .A(n20287), .ZN(n20289) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20294), .B1(
        n20749), .B2(n20293), .ZN(n20288) );
  OAI211_X1 U23223 ( .C1(n20691), .C2(n20328), .A(n20289), .B(n20288), .ZN(
        P1_U3055) );
  OAI22_X1 U23224 ( .A1(n20291), .A2(n20765), .B1(n20290), .B2(n20620), .ZN(
        n20292) );
  INV_X1 U23225 ( .A(n20292), .ZN(n20296) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20294), .B1(
        n20756), .B2(n20293), .ZN(n20295) );
  OAI211_X1 U23227 ( .C1(n20699), .C2(n20328), .A(n20296), .B(n20295), .ZN(
        P1_U3056) );
  OR2_X1 U23228 ( .A1(n20553), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20327) );
  OAI22_X1 U23229 ( .A1(n20338), .A2(n20671), .B1(n20583), .B2(n20327), .ZN(
        n20297) );
  INV_X1 U23230 ( .A(n20297), .ZN(n20308) );
  OAI21_X1 U23231 ( .B1(n20298), .B2(n20708), .A(n20858), .ZN(n20306) );
  AND2_X1 U23232 ( .A1(n11685), .A2(n20861), .ZN(n20701) );
  INV_X1 U23233 ( .A(n20327), .ZN(n20299) );
  AOI21_X1 U23234 ( .B1(n20300), .B2(n20701), .A(n20299), .ZN(n20305) );
  INV_X1 U23235 ( .A(n20305), .ZN(n20303) );
  INV_X1 U23236 ( .A(n20710), .ZN(n20301) );
  AOI21_X1 U23237 ( .B1(n20852), .B2(n20304), .A(n20301), .ZN(n20302) );
  OAI21_X1 U23238 ( .B1(n20306), .B2(n20303), .A(n20302), .ZN(n20331) );
  OAI22_X1 U23239 ( .A1(n20306), .A2(n20305), .B1(n20189), .B2(n20304), .ZN(
        n20330) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20331), .B1(
        n20705), .B2(n20330), .ZN(n20307) );
  OAI211_X1 U23241 ( .C1(n20716), .C2(n20328), .A(n20308), .B(n20307), .ZN(
        P1_U3057) );
  OAI22_X1 U23242 ( .A1(n20338), .A2(n20675), .B1(n20595), .B2(n20327), .ZN(
        n20309) );
  INV_X1 U23243 ( .A(n20309), .ZN(n20311) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20331), .B1(
        n20717), .B2(n20330), .ZN(n20310) );
  OAI211_X1 U23245 ( .C1(n20722), .C2(n20328), .A(n20311), .B(n20310), .ZN(
        P1_U3058) );
  OAI22_X1 U23246 ( .A1(n20338), .A2(n20728), .B1(n20327), .B2(n20599), .ZN(
        n20312) );
  INV_X1 U23247 ( .A(n20312), .ZN(n20314) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20331), .B1(
        n20723), .B2(n20330), .ZN(n20313) );
  OAI211_X1 U23249 ( .C1(n20642), .C2(n20328), .A(n20314), .B(n20313), .ZN(
        P1_U3059) );
  OAI22_X1 U23250 ( .A1(n20338), .A2(n20736), .B1(n20603), .B2(n20327), .ZN(
        n20315) );
  INV_X1 U23251 ( .A(n20315), .ZN(n20317) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20331), .B1(
        n20729), .B2(n20330), .ZN(n20316) );
  OAI211_X1 U23253 ( .C1(n20646), .C2(n20328), .A(n20317), .B(n20316), .ZN(
        P1_U3060) );
  OAI22_X1 U23254 ( .A1(n20338), .A2(n20683), .B1(n20607), .B2(n20327), .ZN(
        n20318) );
  INV_X1 U23255 ( .A(n20318), .ZN(n20320) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20331), .B1(
        n20737), .B2(n20330), .ZN(n20319) );
  OAI211_X1 U23257 ( .C1(n20742), .C2(n20328), .A(n20320), .B(n20319), .ZN(
        P1_U3061) );
  OAI22_X1 U23258 ( .A1(n20328), .A2(n20748), .B1(n20539), .B2(n20327), .ZN(
        n20321) );
  INV_X1 U23259 ( .A(n20321), .ZN(n20323) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20331), .B1(
        n20743), .B2(n20330), .ZN(n20322) );
  OAI211_X1 U23261 ( .C1(n20687), .C2(n20338), .A(n20323), .B(n20322), .ZN(
        P1_U3062) );
  OAI22_X1 U23262 ( .A1(n20338), .A2(n20691), .B1(n20327), .B2(n20615), .ZN(
        n20324) );
  INV_X1 U23263 ( .A(n20324), .ZN(n20326) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20331), .B1(
        n20749), .B2(n20330), .ZN(n20325) );
  OAI211_X1 U23265 ( .C1(n20754), .C2(n20328), .A(n20326), .B(n20325), .ZN(
        P1_U3063) );
  OAI22_X1 U23266 ( .A1(n20328), .A2(n20765), .B1(n20327), .B2(n20620), .ZN(
        n20329) );
  INV_X1 U23267 ( .A(n20329), .ZN(n20333) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20331), .B1(
        n20756), .B2(n20330), .ZN(n20332) );
  OAI211_X1 U23269 ( .C1(n20699), .C2(n20338), .A(n20333), .B(n20332), .ZN(
        P1_U3064) );
  INV_X1 U23270 ( .A(n20432), .ZN(n20335) );
  NOR3_X1 U23271 ( .A1(n15856), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20368) );
  INV_X1 U23272 ( .A(n20368), .ZN(n20365) );
  NOR2_X1 U23273 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20365), .ZN(
        n20359) );
  NOR2_X1 U23274 ( .A1(n13398), .A2(n20336), .ZN(n20392) );
  NAND2_X1 U23275 ( .A1(n20392), .A2(n20858), .ZN(n20427) );
  OAI22_X1 U23276 ( .A1(n20427), .A2(n20660), .B1(n20661), .B2(n20337), .ZN(
        n20358) );
  AOI22_X1 U23277 ( .A1(n20706), .A2(n20359), .B1(n20705), .B2(n20358), .ZN(
        n20345) );
  INV_X1 U23278 ( .A(n20392), .ZN(n20341) );
  INV_X1 U23279 ( .A(n20388), .ZN(n20339) );
  OAI21_X1 U23280 ( .B1(n20360), .B2(n20339), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20340) );
  OAI21_X1 U23281 ( .B1(n20660), .B2(n20341), .A(n20340), .ZN(n20343) );
  AND2_X1 U23282 ( .A1(n20342), .A2(n20522), .ZN(n20666) );
  OAI221_X1 U23283 ( .B1(n20359), .B2(n20466), .C1(n20359), .C2(n20343), .A(
        n20666), .ZN(n20361) );
  INV_X1 U23284 ( .A(n20716), .ZN(n20668) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20668), .ZN(n20344) );
  OAI211_X1 U23286 ( .C1(n20671), .C2(n20388), .A(n20345), .B(n20344), .ZN(
        P1_U3065) );
  AOI22_X1 U23287 ( .A1(n20718), .A2(n20359), .B1(n20717), .B2(n20358), .ZN(
        n20347) );
  INV_X1 U23288 ( .A(n20722), .ZN(n20672) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20672), .ZN(n20346) );
  OAI211_X1 U23290 ( .C1(n20675), .C2(n20388), .A(n20347), .B(n20346), .ZN(
        P1_U3066) );
  AOI22_X1 U23291 ( .A1(n20724), .A2(n20359), .B1(n20723), .B2(n20358), .ZN(
        n20349) );
  INV_X1 U23292 ( .A(n20642), .ZN(n20725) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20725), .ZN(n20348) );
  OAI211_X1 U23294 ( .C1(n20728), .C2(n20388), .A(n20349), .B(n20348), .ZN(
        P1_U3067) );
  AOI22_X1 U23295 ( .A1(n20730), .A2(n20359), .B1(n20729), .B2(n20358), .ZN(
        n20351) );
  INV_X1 U23296 ( .A(n20646), .ZN(n20731) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20731), .ZN(n20350) );
  OAI211_X1 U23298 ( .C1(n20736), .C2(n20388), .A(n20351), .B(n20350), .ZN(
        P1_U3068) );
  AOI22_X1 U23299 ( .A1(n20738), .A2(n20359), .B1(n20737), .B2(n20358), .ZN(
        n20353) );
  INV_X1 U23300 ( .A(n20742), .ZN(n20680) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20680), .ZN(n20352) );
  OAI211_X1 U23302 ( .C1(n20683), .C2(n20388), .A(n20353), .B(n20352), .ZN(
        P1_U3069) );
  AOI22_X1 U23303 ( .A1(n20744), .A2(n20359), .B1(n20743), .B2(n20358), .ZN(
        n20355) );
  INV_X1 U23304 ( .A(n20748), .ZN(n20684) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20684), .ZN(n20354) );
  OAI211_X1 U23306 ( .C1(n20687), .C2(n20388), .A(n20355), .B(n20354), .ZN(
        P1_U3070) );
  AOI22_X1 U23307 ( .A1(n20750), .A2(n20359), .B1(n20749), .B2(n20358), .ZN(
        n20357) );
  INV_X1 U23308 ( .A(n20754), .ZN(n20688) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20688), .ZN(n20356) );
  OAI211_X1 U23310 ( .C1(n20691), .C2(n20388), .A(n20357), .B(n20356), .ZN(
        P1_U3071) );
  AOI22_X1 U23311 ( .A1(n20758), .A2(n20359), .B1(n20756), .B2(n20358), .ZN(
        n20363) );
  INV_X1 U23312 ( .A(n20765), .ZN(n20694) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20694), .ZN(n20362) );
  OAI211_X1 U23314 ( .C1(n20699), .C2(n20388), .A(n20363), .B(n20362), .ZN(
        P1_U3072) );
  NOR2_X1 U23315 ( .A1(n20866), .A2(n20365), .ZN(n20384) );
  INV_X1 U23316 ( .A(n20384), .ZN(n20366) );
  OAI222_X1 U23317 ( .A1(n20366), .A2(n20852), .B1(n20703), .B2(n20365), .C1(
        n20364), .C2(n20427), .ZN(n20383) );
  AOI22_X1 U23318 ( .A1(n20706), .A2(n20384), .B1(n20705), .B2(n20383), .ZN(
        n20370) );
  NOR3_X1 U23319 ( .A1(n20432), .A2(n20852), .A3(n20629), .ZN(n20367) );
  OAI21_X1 U23320 ( .B1(n20368), .B2(n20367), .A(n20710), .ZN(n20385) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20713), .ZN(n20369) );
  OAI211_X1 U23322 ( .C1(n20716), .C2(n20388), .A(n20370), .B(n20369), .ZN(
        P1_U3073) );
  AOI22_X1 U23323 ( .A1(n20718), .A2(n20384), .B1(n20717), .B2(n20383), .ZN(
        n20372) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20719), .ZN(n20371) );
  OAI211_X1 U23325 ( .C1(n20722), .C2(n20388), .A(n20372), .B(n20371), .ZN(
        P1_U3074) );
  AOI22_X1 U23326 ( .A1(n20724), .A2(n20384), .B1(n20723), .B2(n20383), .ZN(
        n20374) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20639), .ZN(n20373) );
  OAI211_X1 U23328 ( .C1(n20642), .C2(n20388), .A(n20374), .B(n20373), .ZN(
        P1_U3075) );
  AOI22_X1 U23329 ( .A1(n20730), .A2(n20384), .B1(n20729), .B2(n20383), .ZN(
        n20376) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20643), .ZN(n20375) );
  OAI211_X1 U23331 ( .C1(n20646), .C2(n20388), .A(n20376), .B(n20375), .ZN(
        P1_U3076) );
  AOI22_X1 U23332 ( .A1(n20738), .A2(n20384), .B1(n20737), .B2(n20383), .ZN(
        n20378) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20739), .ZN(n20377) );
  OAI211_X1 U23334 ( .C1(n20742), .C2(n20388), .A(n20378), .B(n20377), .ZN(
        P1_U3077) );
  AOI22_X1 U23335 ( .A1(n20744), .A2(n20384), .B1(n20743), .B2(n20383), .ZN(
        n20380) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20745), .ZN(n20379) );
  OAI211_X1 U23337 ( .C1(n20748), .C2(n20388), .A(n20380), .B(n20379), .ZN(
        P1_U3078) );
  AOI22_X1 U23338 ( .A1(n20750), .A2(n20384), .B1(n20749), .B2(n20383), .ZN(
        n20382) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20751), .ZN(n20381) );
  OAI211_X1 U23340 ( .C1(n20754), .C2(n20388), .A(n20382), .B(n20381), .ZN(
        P1_U3079) );
  AOI22_X1 U23341 ( .A1(n20758), .A2(n20384), .B1(n20756), .B2(n20383), .ZN(
        n20387) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20385), .B1(
        n20390), .B2(n20759), .ZN(n20386) );
  OAI211_X1 U23343 ( .C1(n20765), .C2(n20388), .A(n20387), .B(n20386), .ZN(
        P1_U3080) );
  NOR2_X1 U23344 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20429), .ZN(
        n20413) );
  INV_X1 U23345 ( .A(n20413), .ZN(n20419) );
  OAI22_X1 U23346 ( .A1(n20425), .A2(n20716), .B1(n20583), .B2(n20419), .ZN(
        n20389) );
  INV_X1 U23347 ( .A(n20389), .ZN(n20400) );
  OAI21_X1 U23348 ( .B1(n20451), .B2(n20390), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20391) );
  NAND2_X1 U23349 ( .A1(n20391), .A2(n20858), .ZN(n20398) );
  INV_X1 U23350 ( .A(n20398), .ZN(n20394) );
  NAND2_X1 U23351 ( .A1(n20392), .A2(n20660), .ZN(n20397) );
  AOI21_X1 U23352 ( .B1(n20394), .B2(n20397), .A(n20393), .ZN(n20395) );
  OAI211_X1 U23353 ( .C1(n20413), .C2(n20466), .A(n20666), .B(n20395), .ZN(
        n20422) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20422), .B1(
        n20705), .B2(n20421), .ZN(n20399) );
  OAI211_X1 U23355 ( .C1(n20671), .C2(n20448), .A(n20400), .B(n20399), .ZN(
        P1_U3081) );
  OAI22_X1 U23356 ( .A1(n20448), .A2(n20675), .B1(n20595), .B2(n20419), .ZN(
        n20401) );
  INV_X1 U23357 ( .A(n20401), .ZN(n20403) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20422), .B1(
        n20717), .B2(n20421), .ZN(n20402) );
  OAI211_X1 U23359 ( .C1(n20722), .C2(n20425), .A(n20403), .B(n20402), .ZN(
        P1_U3082) );
  OAI22_X1 U23360 ( .A1(n20425), .A2(n20642), .B1(n20599), .B2(n20419), .ZN(
        n20404) );
  INV_X1 U23361 ( .A(n20404), .ZN(n20406) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20422), .B1(
        n20723), .B2(n20421), .ZN(n20405) );
  OAI211_X1 U23363 ( .C1(n20728), .C2(n20448), .A(n20406), .B(n20405), .ZN(
        P1_U3083) );
  OAI22_X1 U23364 ( .A1(n20448), .A2(n20736), .B1(n20603), .B2(n20419), .ZN(
        n20407) );
  INV_X1 U23365 ( .A(n20407), .ZN(n20409) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20422), .B1(
        n20729), .B2(n20421), .ZN(n20408) );
  OAI211_X1 U23367 ( .C1(n20646), .C2(n20425), .A(n20409), .B(n20408), .ZN(
        P1_U3084) );
  OAI22_X1 U23368 ( .A1(n20425), .A2(n20742), .B1(n20607), .B2(n20419), .ZN(
        n20410) );
  INV_X1 U23369 ( .A(n20410), .ZN(n20412) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20422), .B1(
        n20737), .B2(n20421), .ZN(n20411) );
  OAI211_X1 U23371 ( .C1(n20683), .C2(n20448), .A(n20412), .B(n20411), .ZN(
        P1_U3085) );
  AOI22_X1 U23372 ( .A1(n20451), .A2(n20745), .B1(n20744), .B2(n20413), .ZN(
        n20415) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20422), .B1(
        n20743), .B2(n20421), .ZN(n20414) );
  OAI211_X1 U23374 ( .C1(n20748), .C2(n20425), .A(n20415), .B(n20414), .ZN(
        P1_U3086) );
  OAI22_X1 U23375 ( .A1(n20425), .A2(n20754), .B1(n20615), .B2(n20419), .ZN(
        n20416) );
  INV_X1 U23376 ( .A(n20416), .ZN(n20418) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20422), .B1(
        n20749), .B2(n20421), .ZN(n20417) );
  OAI211_X1 U23378 ( .C1(n20691), .C2(n20448), .A(n20418), .B(n20417), .ZN(
        P1_U3087) );
  OAI22_X1 U23379 ( .A1(n20448), .A2(n20699), .B1(n20620), .B2(n20419), .ZN(
        n20420) );
  INV_X1 U23380 ( .A(n20420), .ZN(n20424) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20422), .B1(
        n20756), .B2(n20421), .ZN(n20423) );
  OAI211_X1 U23382 ( .C1(n20765), .C2(n20425), .A(n20424), .B(n20423), .ZN(
        P1_U3088) );
  INV_X1 U23383 ( .A(n20430), .ZN(n20450) );
  INV_X1 U23384 ( .A(n20701), .ZN(n20428) );
  OAI222_X1 U23385 ( .A1(n20852), .A2(n20430), .B1(n20703), .B2(n20429), .C1(
        n20428), .C2(n20427), .ZN(n20449) );
  AOI22_X1 U23386 ( .A1(n20706), .A2(n20450), .B1(n20705), .B2(n20449), .ZN(
        n20435) );
  OR2_X1 U23387 ( .A1(n20708), .A2(n20852), .ZN(n20431) );
  NOR2_X1 U23388 ( .A1(n20432), .A2(n20431), .ZN(n20849) );
  OAI21_X1 U23389 ( .B1(n20433), .B2(n20849), .A(n20710), .ZN(n20452) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20668), .ZN(n20434) );
  OAI211_X1 U23391 ( .C1(n20671), .C2(n20455), .A(n20435), .B(n20434), .ZN(
        P1_U3089) );
  AOI22_X1 U23392 ( .A1(n20718), .A2(n20450), .B1(n20717), .B2(n20449), .ZN(
        n20437) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20672), .ZN(n20436) );
  OAI211_X1 U23394 ( .C1(n20675), .C2(n20455), .A(n20437), .B(n20436), .ZN(
        P1_U3090) );
  AOI22_X1 U23395 ( .A1(n20724), .A2(n20450), .B1(n20723), .B2(n20449), .ZN(
        n20439) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20725), .ZN(n20438) );
  OAI211_X1 U23397 ( .C1(n20728), .C2(n20455), .A(n20439), .B(n20438), .ZN(
        P1_U3091) );
  AOI22_X1 U23398 ( .A1(n20730), .A2(n20450), .B1(n20729), .B2(n20449), .ZN(
        n20441) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20731), .ZN(n20440) );
  OAI211_X1 U23400 ( .C1(n20736), .C2(n20455), .A(n20441), .B(n20440), .ZN(
        P1_U3092) );
  AOI22_X1 U23401 ( .A1(n20738), .A2(n20450), .B1(n20737), .B2(n20449), .ZN(
        n20443) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20452), .B1(
        n20483), .B2(n20739), .ZN(n20442) );
  OAI211_X1 U23403 ( .C1(n20742), .C2(n20448), .A(n20443), .B(n20442), .ZN(
        P1_U3093) );
  AOI22_X1 U23404 ( .A1(n20744), .A2(n20450), .B1(n20743), .B2(n20449), .ZN(
        n20445) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20452), .B1(
        n20483), .B2(n20745), .ZN(n20444) );
  OAI211_X1 U23406 ( .C1(n20748), .C2(n20448), .A(n20445), .B(n20444), .ZN(
        P1_U3094) );
  AOI22_X1 U23407 ( .A1(n20750), .A2(n20450), .B1(n20749), .B2(n20449), .ZN(
        n20447) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20452), .B1(
        n20483), .B2(n20751), .ZN(n20446) );
  OAI211_X1 U23409 ( .C1(n20754), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        P1_U3095) );
  AOI22_X1 U23410 ( .A1(n20758), .A2(n20450), .B1(n20756), .B2(n20449), .ZN(
        n20454) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20694), .ZN(n20453) );
  OAI211_X1 U23412 ( .C1(n20699), .C2(n20455), .A(n20454), .B(n20453), .ZN(
        P1_U3096) );
  INV_X1 U23413 ( .A(n20456), .ZN(n20457) );
  INV_X1 U23414 ( .A(n20850), .ZN(n20460) );
  NOR3_X1 U23415 ( .A1(n20856), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20490) );
  INV_X1 U23416 ( .A(n20490), .ZN(n20487) );
  NOR2_X1 U23417 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20487), .ZN(
        n20481) );
  AOI21_X1 U23418 ( .B1(n20554), .B2(n20586), .A(n20481), .ZN(n20463) );
  NAND2_X1 U23419 ( .A1(n20461), .A2(n20520), .ZN(n20590) );
  OAI22_X1 U23420 ( .A1(n20463), .A2(n20852), .B1(n20522), .B2(n20590), .ZN(
        n20482) );
  AOI22_X1 U23421 ( .A1(n20705), .A2(n20482), .B1(n20706), .B2(n20481), .ZN(
        n20468) );
  INV_X1 U23422 ( .A(n20512), .ZN(n20462) );
  OAI21_X1 U23423 ( .B1(n20462), .B2(n20483), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20464) );
  NAND2_X1 U23424 ( .A1(n20464), .A2(n20463), .ZN(n20465) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20668), .ZN(n20467) );
  OAI211_X1 U23426 ( .C1(n20671), .C2(n20512), .A(n20468), .B(n20467), .ZN(
        P1_U3097) );
  AOI22_X1 U23427 ( .A1(n20717), .A2(n20482), .B1(n20718), .B2(n20481), .ZN(
        n20470) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20672), .ZN(n20469) );
  OAI211_X1 U23429 ( .C1(n20675), .C2(n20512), .A(n20470), .B(n20469), .ZN(
        P1_U3098) );
  AOI22_X1 U23430 ( .A1(n20723), .A2(n20482), .B1(n20724), .B2(n20481), .ZN(
        n20472) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20725), .ZN(n20471) );
  OAI211_X1 U23432 ( .C1(n20728), .C2(n20512), .A(n20472), .B(n20471), .ZN(
        P1_U3099) );
  AOI22_X1 U23433 ( .A1(n20729), .A2(n20482), .B1(n20730), .B2(n20481), .ZN(
        n20474) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20731), .ZN(n20473) );
  OAI211_X1 U23435 ( .C1(n20736), .C2(n20512), .A(n20474), .B(n20473), .ZN(
        P1_U3100) );
  AOI22_X1 U23436 ( .A1(n20737), .A2(n20482), .B1(n20738), .B2(n20481), .ZN(
        n20476) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20680), .ZN(n20475) );
  OAI211_X1 U23438 ( .C1(n20683), .C2(n20512), .A(n20476), .B(n20475), .ZN(
        P1_U3101) );
  AOI22_X1 U23439 ( .A1(n20743), .A2(n20482), .B1(n20744), .B2(n20481), .ZN(
        n20478) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20684), .ZN(n20477) );
  OAI211_X1 U23441 ( .C1(n20687), .C2(n20512), .A(n20478), .B(n20477), .ZN(
        P1_U3102) );
  AOI22_X1 U23442 ( .A1(n20749), .A2(n20482), .B1(n20750), .B2(n20481), .ZN(
        n20480) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20688), .ZN(n20479) );
  OAI211_X1 U23444 ( .C1(n20691), .C2(n20512), .A(n20480), .B(n20479), .ZN(
        P1_U3103) );
  AOI22_X1 U23445 ( .A1(n20756), .A2(n20482), .B1(n20758), .B2(n20481), .ZN(
        n20486) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20694), .ZN(n20485) );
  OAI211_X1 U23447 ( .C1(n20699), .C2(n20512), .A(n20486), .B(n20485), .ZN(
        P1_U3104) );
  NOR2_X1 U23448 ( .A1(n20866), .A2(n20487), .ZN(n20506) );
  AOI21_X1 U23449 ( .B1(n20554), .B2(n20627), .A(n20506), .ZN(n20488) );
  OAI22_X1 U23450 ( .A1(n20488), .A2(n20852), .B1(n20487), .B2(n20703), .ZN(
        n20507) );
  AOI22_X1 U23451 ( .A1(n20705), .A2(n20507), .B1(n20706), .B2(n20506), .ZN(
        n20493) );
  OAI211_X1 U23452 ( .C1(n20557), .C2(n20629), .A(n20858), .B(n20488), .ZN(
        n20489) );
  OAI211_X1 U23453 ( .C1(n20858), .C2(n20490), .A(n20710), .B(n20489), .ZN(
        n20509) );
  INV_X1 U23454 ( .A(n20634), .ZN(n20491) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20713), .ZN(n20492) );
  OAI211_X1 U23456 ( .C1(n20716), .C2(n20512), .A(n20493), .B(n20492), .ZN(
        P1_U3105) );
  AOI22_X1 U23457 ( .A1(n20717), .A2(n20507), .B1(n20718), .B2(n20506), .ZN(
        n20495) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20719), .ZN(n20494) );
  OAI211_X1 U23459 ( .C1(n20722), .C2(n20512), .A(n20495), .B(n20494), .ZN(
        P1_U3106) );
  AOI22_X1 U23460 ( .A1(n20723), .A2(n20507), .B1(n20724), .B2(n20506), .ZN(
        n20497) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20639), .ZN(n20496) );
  OAI211_X1 U23462 ( .C1(n20642), .C2(n20512), .A(n20497), .B(n20496), .ZN(
        P1_U3107) );
  AOI22_X1 U23463 ( .A1(n20729), .A2(n20507), .B1(n20730), .B2(n20506), .ZN(
        n20499) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20643), .ZN(n20498) );
  OAI211_X1 U23465 ( .C1(n20646), .C2(n20512), .A(n20499), .B(n20498), .ZN(
        P1_U3108) );
  AOI22_X1 U23466 ( .A1(n20737), .A2(n20507), .B1(n20738), .B2(n20506), .ZN(
        n20501) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20739), .ZN(n20500) );
  OAI211_X1 U23468 ( .C1(n20742), .C2(n20512), .A(n20501), .B(n20500), .ZN(
        P1_U3109) );
  AOI22_X1 U23469 ( .A1(n20743), .A2(n20507), .B1(n20744), .B2(n20506), .ZN(
        n20503) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20745), .ZN(n20502) );
  OAI211_X1 U23471 ( .C1(n20748), .C2(n20512), .A(n20503), .B(n20502), .ZN(
        P1_U3110) );
  AOI22_X1 U23472 ( .A1(n20749), .A2(n20507), .B1(n20750), .B2(n20506), .ZN(
        n20505) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20751), .ZN(n20504) );
  OAI211_X1 U23474 ( .C1(n20754), .C2(n20512), .A(n20505), .B(n20504), .ZN(
        P1_U3111) );
  AOI22_X1 U23475 ( .A1(n20756), .A2(n20507), .B1(n20758), .B2(n20506), .ZN(
        n20511) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20759), .ZN(n20510) );
  OAI211_X1 U23477 ( .C1(n20765), .C2(n20512), .A(n20511), .B(n20510), .ZN(
        P1_U3112) );
  NOR3_X1 U23478 ( .A1(n20856), .A2(n20514), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20559) );
  NAND2_X1 U23479 ( .A1(n20866), .A2(n20559), .ZN(n20546) );
  OAI22_X1 U23480 ( .A1(n20581), .A2(n20671), .B1(n20583), .B2(n20546), .ZN(
        n20515) );
  INV_X1 U23481 ( .A(n20515), .ZN(n20526) );
  NAND2_X1 U23482 ( .A1(n20581), .A2(n20547), .ZN(n20516) );
  AOI21_X1 U23483 ( .B1(n20516), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20852), 
        .ZN(n20519) );
  NAND2_X1 U23484 ( .A1(n20554), .A2(n20660), .ZN(n20523) );
  AOI22_X1 U23485 ( .A1(n20519), .A2(n20523), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20546), .ZN(n20517) );
  OAI21_X1 U23486 ( .B1(n20856), .B2(n20520), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20665) );
  NAND3_X1 U23487 ( .A1(n20518), .A2(n20517), .A3(n20665), .ZN(n20550) );
  INV_X1 U23488 ( .A(n20519), .ZN(n20524) );
  INV_X1 U23489 ( .A(n20520), .ZN(n20521) );
  NAND2_X1 U23490 ( .A1(n20521), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20662) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20550), .B1(
        n20705), .B2(n20549), .ZN(n20525) );
  OAI211_X1 U23492 ( .C1(n20716), .C2(n20547), .A(n20526), .B(n20525), .ZN(
        P1_U3113) );
  OAI22_X1 U23493 ( .A1(n20547), .A2(n20722), .B1(n20595), .B2(n20546), .ZN(
        n20527) );
  INV_X1 U23494 ( .A(n20527), .ZN(n20529) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20550), .B1(
        n20717), .B2(n20549), .ZN(n20528) );
  OAI211_X1 U23496 ( .C1(n20675), .C2(n20581), .A(n20529), .B(n20528), .ZN(
        P1_U3114) );
  OAI22_X1 U23497 ( .A1(n20581), .A2(n20728), .B1(n20599), .B2(n20546), .ZN(
        n20530) );
  INV_X1 U23498 ( .A(n20530), .ZN(n20532) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20550), .B1(
        n20723), .B2(n20549), .ZN(n20531) );
  OAI211_X1 U23500 ( .C1(n20642), .C2(n20547), .A(n20532), .B(n20531), .ZN(
        P1_U3115) );
  OAI22_X1 U23501 ( .A1(n20581), .A2(n20736), .B1(n20603), .B2(n20546), .ZN(
        n20533) );
  INV_X1 U23502 ( .A(n20533), .ZN(n20535) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20550), .B1(
        n20729), .B2(n20549), .ZN(n20534) );
  OAI211_X1 U23504 ( .C1(n20646), .C2(n20547), .A(n20535), .B(n20534), .ZN(
        P1_U3116) );
  OAI22_X1 U23505 ( .A1(n20547), .A2(n20742), .B1(n20607), .B2(n20546), .ZN(
        n20536) );
  INV_X1 U23506 ( .A(n20536), .ZN(n20538) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20550), .B1(
        n20737), .B2(n20549), .ZN(n20537) );
  OAI211_X1 U23508 ( .C1(n20683), .C2(n20581), .A(n20538), .B(n20537), .ZN(
        P1_U3117) );
  OAI22_X1 U23509 ( .A1(n20547), .A2(n20748), .B1(n20539), .B2(n20546), .ZN(
        n20540) );
  INV_X1 U23510 ( .A(n20540), .ZN(n20542) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20550), .B1(
        n20743), .B2(n20549), .ZN(n20541) );
  OAI211_X1 U23512 ( .C1(n20687), .C2(n20581), .A(n20542), .B(n20541), .ZN(
        P1_U3118) );
  OAI22_X1 U23513 ( .A1(n20547), .A2(n20754), .B1(n20615), .B2(n20546), .ZN(
        n20543) );
  INV_X1 U23514 ( .A(n20543), .ZN(n20545) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20550), .B1(
        n20749), .B2(n20549), .ZN(n20544) );
  OAI211_X1 U23516 ( .C1(n20691), .C2(n20581), .A(n20545), .B(n20544), .ZN(
        P1_U3119) );
  OAI22_X1 U23517 ( .A1(n20547), .A2(n20765), .B1(n20620), .B2(n20546), .ZN(
        n20548) );
  INV_X1 U23518 ( .A(n20548), .ZN(n20552) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20550), .B1(
        n20756), .B2(n20549), .ZN(n20551) );
  OAI211_X1 U23520 ( .C1(n20699), .C2(n20581), .A(n20552), .B(n20551), .ZN(
        P1_U3120) );
  AOI21_X1 U23521 ( .B1(n20554), .B2(n20701), .A(n10455), .ZN(n20556) );
  INV_X1 U23522 ( .A(n20559), .ZN(n20555) );
  OAI22_X1 U23523 ( .A1(n20556), .A2(n20852), .B1(n20555), .B2(n20703), .ZN(
        n20576) );
  AOI22_X1 U23524 ( .A1(n20705), .A2(n20576), .B1(n20706), .B2(n10455), .ZN(
        n20562) );
  OAI211_X1 U23525 ( .C1(n20557), .C2(n20708), .A(n20858), .B(n20556), .ZN(
        n20558) );
  OAI211_X1 U23526 ( .C1(n20858), .C2(n20559), .A(n20710), .B(n20558), .ZN(
        n20578) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20713), .ZN(n20561) );
  OAI211_X1 U23528 ( .C1(n20716), .C2(n20581), .A(n20562), .B(n20561), .ZN(
        P1_U3121) );
  AOI22_X1 U23529 ( .A1(n20717), .A2(n20576), .B1(n20718), .B2(n10455), .ZN(
        n20564) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20719), .ZN(n20563) );
  OAI211_X1 U23531 ( .C1(n20722), .C2(n20581), .A(n20564), .B(n20563), .ZN(
        P1_U3122) );
  AOI22_X1 U23532 ( .A1(n20723), .A2(n20576), .B1(n20724), .B2(n10455), .ZN(
        n20566) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20639), .ZN(n20565) );
  OAI211_X1 U23534 ( .C1(n20642), .C2(n20581), .A(n20566), .B(n20565), .ZN(
        P1_U3123) );
  AOI22_X1 U23535 ( .A1(n20729), .A2(n20576), .B1(n20730), .B2(n10455), .ZN(
        n20569) );
  INV_X1 U23536 ( .A(n20581), .ZN(n20567) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20578), .B1(
        n20567), .B2(n20731), .ZN(n20568) );
  OAI211_X1 U23538 ( .C1(n20736), .C2(n20626), .A(n20569), .B(n20568), .ZN(
        P1_U3124) );
  AOI22_X1 U23539 ( .A1(n20737), .A2(n20576), .B1(n20738), .B2(n10455), .ZN(
        n20571) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20739), .ZN(n20570) );
  OAI211_X1 U23541 ( .C1(n20742), .C2(n20581), .A(n20571), .B(n20570), .ZN(
        P1_U3125) );
  AOI22_X1 U23542 ( .A1(n20743), .A2(n20576), .B1(n20744), .B2(n10455), .ZN(
        n20573) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20745), .ZN(n20572) );
  OAI211_X1 U23544 ( .C1(n20748), .C2(n20581), .A(n20573), .B(n20572), .ZN(
        P1_U3126) );
  AOI22_X1 U23545 ( .A1(n20749), .A2(n20576), .B1(n20750), .B2(n10455), .ZN(
        n20575) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20751), .ZN(n20574) );
  OAI211_X1 U23547 ( .C1(n20754), .C2(n20581), .A(n20575), .B(n20574), .ZN(
        P1_U3127) );
  AOI22_X1 U23548 ( .A1(n20756), .A2(n20576), .B1(n20758), .B2(n10455), .ZN(
        n20580) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20759), .ZN(n20579) );
  OAI211_X1 U23550 ( .C1(n20765), .C2(n20581), .A(n20580), .B(n20579), .ZN(
        P1_U3128) );
  NOR3_X1 U23551 ( .A1(n15856), .A2(n20856), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20633) );
  NAND2_X1 U23552 ( .A1(n20866), .A2(n20633), .ZN(n20619) );
  OAI22_X1 U23553 ( .A1(n20658), .A2(n20671), .B1(n20583), .B2(n20619), .ZN(
        n20584) );
  INV_X1 U23554 ( .A(n20584), .ZN(n20594) );
  INV_X1 U23555 ( .A(n20590), .ZN(n20588) );
  NAND2_X1 U23556 ( .A1(n20626), .A2(n20658), .ZN(n20585) );
  AOI21_X1 U23557 ( .B1(n20585), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20852), 
        .ZN(n20589) );
  NOR2_X1 U23558 ( .A1(n13398), .A2(n10037), .ZN(n20702) );
  NAND2_X1 U23559 ( .A1(n20702), .A2(n20586), .ZN(n20591) );
  AOI22_X1 U23560 ( .A1(n20589), .A2(n20591), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20619), .ZN(n20587) );
  OAI211_X1 U23561 ( .C1(n20588), .C2(n20189), .A(n20666), .B(n20587), .ZN(
        n20623) );
  INV_X1 U23562 ( .A(n20589), .ZN(n20592) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20623), .B1(
        n20705), .B2(n20622), .ZN(n20593) );
  OAI211_X1 U23564 ( .C1(n20716), .C2(n20626), .A(n20594), .B(n20593), .ZN(
        P1_U3129) );
  OAI22_X1 U23565 ( .A1(n20658), .A2(n20675), .B1(n20595), .B2(n20619), .ZN(
        n20596) );
  INV_X1 U23566 ( .A(n20596), .ZN(n20598) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20623), .B1(
        n20717), .B2(n20622), .ZN(n20597) );
  OAI211_X1 U23568 ( .C1(n20722), .C2(n20626), .A(n20598), .B(n20597), .ZN(
        P1_U3130) );
  OAI22_X1 U23569 ( .A1(n20658), .A2(n20728), .B1(n20599), .B2(n20619), .ZN(
        n20600) );
  INV_X1 U23570 ( .A(n20600), .ZN(n20602) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20623), .B1(
        n20723), .B2(n20622), .ZN(n20601) );
  OAI211_X1 U23572 ( .C1(n20642), .C2(n20626), .A(n20602), .B(n20601), .ZN(
        P1_U3131) );
  OAI22_X1 U23573 ( .A1(n20658), .A2(n20736), .B1(n20603), .B2(n20619), .ZN(
        n20604) );
  INV_X1 U23574 ( .A(n20604), .ZN(n20606) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20623), .B1(
        n20729), .B2(n20622), .ZN(n20605) );
  OAI211_X1 U23576 ( .C1(n20646), .C2(n20626), .A(n20606), .B(n20605), .ZN(
        P1_U3132) );
  OAI22_X1 U23577 ( .A1(n20658), .A2(n20683), .B1(n20607), .B2(n20619), .ZN(
        n20608) );
  INV_X1 U23578 ( .A(n20608), .ZN(n20610) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20623), .B1(
        n20737), .B2(n20622), .ZN(n20609) );
  OAI211_X1 U23580 ( .C1(n20742), .C2(n20626), .A(n20610), .B(n20609), .ZN(
        P1_U3133) );
  INV_X1 U23581 ( .A(n20658), .ZN(n20612) );
  INV_X1 U23582 ( .A(n20619), .ZN(n20611) );
  AOI22_X1 U23583 ( .A1(n20612), .A2(n20745), .B1(n20744), .B2(n20611), .ZN(
        n20614) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20623), .B1(
        n20743), .B2(n20622), .ZN(n20613) );
  OAI211_X1 U23585 ( .C1(n20748), .C2(n20626), .A(n20614), .B(n20613), .ZN(
        P1_U3134) );
  OAI22_X1 U23586 ( .A1(n20658), .A2(n20691), .B1(n20615), .B2(n20619), .ZN(
        n20616) );
  INV_X1 U23587 ( .A(n20616), .ZN(n20618) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20623), .B1(
        n20749), .B2(n20622), .ZN(n20617) );
  OAI211_X1 U23589 ( .C1(n20754), .C2(n20626), .A(n20618), .B(n20617), .ZN(
        P1_U3135) );
  OAI22_X1 U23590 ( .A1(n20658), .A2(n20699), .B1(n20620), .B2(n20619), .ZN(
        n20621) );
  INV_X1 U23591 ( .A(n20621), .ZN(n20625) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20623), .B1(
        n20756), .B2(n20622), .ZN(n20624) );
  OAI211_X1 U23593 ( .C1(n20765), .C2(n20626), .A(n20625), .B(n20624), .ZN(
        P1_U3136) );
  INV_X1 U23594 ( .A(n20633), .ZN(n20628) );
  NOR2_X1 U23595 ( .A1(n20866), .A2(n20628), .ZN(n20654) );
  AOI21_X1 U23596 ( .B1(n20702), .B2(n20627), .A(n20654), .ZN(n20630) );
  OAI22_X1 U23597 ( .A1(n20630), .A2(n20852), .B1(n20628), .B2(n20703), .ZN(
        n20653) );
  AOI22_X1 U23598 ( .A1(n20706), .A2(n20654), .B1(n20705), .B2(n20653), .ZN(
        n20636) );
  NOR2_X1 U23599 ( .A1(n20709), .A2(n20629), .ZN(n20848) );
  INV_X1 U23600 ( .A(n20848), .ZN(n20631) );
  NAND2_X1 U23601 ( .A1(n20631), .A2(n20630), .ZN(n20632) );
  OAI221_X1 U23602 ( .B1(n20858), .B2(n20633), .C1(n20852), .C2(n20632), .A(
        n20710), .ZN(n20655) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20713), .ZN(n20635) );
  OAI211_X1 U23604 ( .C1(n20716), .C2(n20658), .A(n20636), .B(n20635), .ZN(
        P1_U3137) );
  AOI22_X1 U23605 ( .A1(n20718), .A2(n20654), .B1(n20717), .B2(n20653), .ZN(
        n20638) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20719), .ZN(n20637) );
  OAI211_X1 U23607 ( .C1(n20722), .C2(n20658), .A(n20638), .B(n20637), .ZN(
        P1_U3138) );
  AOI22_X1 U23608 ( .A1(n20724), .A2(n20654), .B1(n20723), .B2(n20653), .ZN(
        n20641) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20639), .ZN(n20640) );
  OAI211_X1 U23610 ( .C1(n20642), .C2(n20658), .A(n20641), .B(n20640), .ZN(
        P1_U3139) );
  AOI22_X1 U23611 ( .A1(n20730), .A2(n20654), .B1(n20729), .B2(n20653), .ZN(
        n20645) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20643), .ZN(n20644) );
  OAI211_X1 U23613 ( .C1(n20646), .C2(n20658), .A(n20645), .B(n20644), .ZN(
        P1_U3140) );
  AOI22_X1 U23614 ( .A1(n20738), .A2(n20654), .B1(n20737), .B2(n20653), .ZN(
        n20648) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20739), .ZN(n20647) );
  OAI211_X1 U23616 ( .C1(n20742), .C2(n20658), .A(n20648), .B(n20647), .ZN(
        P1_U3141) );
  AOI22_X1 U23617 ( .A1(n20744), .A2(n20654), .B1(n20743), .B2(n20653), .ZN(
        n20650) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20745), .ZN(n20649) );
  OAI211_X1 U23619 ( .C1(n20748), .C2(n20658), .A(n20650), .B(n20649), .ZN(
        P1_U3142) );
  AOI22_X1 U23620 ( .A1(n20750), .A2(n20654), .B1(n20749), .B2(n20653), .ZN(
        n20652) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20751), .ZN(n20651) );
  OAI211_X1 U23622 ( .C1(n20754), .C2(n20658), .A(n20652), .B(n20651), .ZN(
        P1_U3143) );
  AOI22_X1 U23623 ( .A1(n20758), .A2(n20654), .B1(n20756), .B2(n20653), .ZN(
        n20657) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20655), .B1(
        n20695), .B2(n20759), .ZN(n20656) );
  OAI211_X1 U23625 ( .C1(n20765), .C2(n20658), .A(n20657), .B(n20656), .ZN(
        P1_U3144) );
  INV_X1 U23626 ( .A(n20712), .ZN(n20704) );
  NOR2_X1 U23627 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20704), .ZN(
        n20693) );
  NAND2_X1 U23628 ( .A1(n20702), .A2(n20660), .ZN(n20663) );
  OAI22_X1 U23629 ( .A1(n20663), .A2(n20852), .B1(n20662), .B2(n20661), .ZN(
        n20692) );
  AOI22_X1 U23630 ( .A1(n20706), .A2(n20693), .B1(n20705), .B2(n20692), .ZN(
        n20670) );
  INV_X1 U23631 ( .A(n20764), .ZN(n20732) );
  OAI21_X1 U23632 ( .B1(n20732), .B2(n20695), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20664) );
  AOI21_X1 U23633 ( .B1(n20664), .B2(n20663), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20667) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20668), .ZN(n20669) );
  OAI211_X1 U23635 ( .C1(n20671), .C2(n20764), .A(n20670), .B(n20669), .ZN(
        P1_U3145) );
  AOI22_X1 U23636 ( .A1(n20718), .A2(n20693), .B1(n20717), .B2(n20692), .ZN(
        n20674) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20672), .ZN(n20673) );
  OAI211_X1 U23638 ( .C1(n20675), .C2(n20764), .A(n20674), .B(n20673), .ZN(
        P1_U3146) );
  AOI22_X1 U23639 ( .A1(n20724), .A2(n20693), .B1(n20723), .B2(n20692), .ZN(
        n20677) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20725), .ZN(n20676) );
  OAI211_X1 U23641 ( .C1(n20728), .C2(n20764), .A(n20677), .B(n20676), .ZN(
        P1_U3147) );
  AOI22_X1 U23642 ( .A1(n20730), .A2(n20693), .B1(n20729), .B2(n20692), .ZN(
        n20679) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20731), .ZN(n20678) );
  OAI211_X1 U23644 ( .C1(n20736), .C2(n20764), .A(n20679), .B(n20678), .ZN(
        P1_U3148) );
  AOI22_X1 U23645 ( .A1(n20738), .A2(n20693), .B1(n20737), .B2(n20692), .ZN(
        n20682) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20680), .ZN(n20681) );
  OAI211_X1 U23647 ( .C1(n20683), .C2(n20764), .A(n20682), .B(n20681), .ZN(
        P1_U3149) );
  AOI22_X1 U23648 ( .A1(n20744), .A2(n20693), .B1(n20743), .B2(n20692), .ZN(
        n20686) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20684), .ZN(n20685) );
  OAI211_X1 U23650 ( .C1(n20687), .C2(n20764), .A(n20686), .B(n20685), .ZN(
        P1_U3150) );
  AOI22_X1 U23651 ( .A1(n20750), .A2(n20693), .B1(n20749), .B2(n20692), .ZN(
        n20690) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20688), .ZN(n20689) );
  OAI211_X1 U23653 ( .C1(n20691), .C2(n20764), .A(n20690), .B(n20689), .ZN(
        P1_U3151) );
  AOI22_X1 U23654 ( .A1(n20758), .A2(n20693), .B1(n20756), .B2(n20692), .ZN(
        n20698) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20696), .B1(
        n20695), .B2(n20694), .ZN(n20697) );
  OAI211_X1 U23656 ( .C1(n20699), .C2(n20764), .A(n20698), .B(n20697), .ZN(
        P1_U3152) );
  INV_X1 U23657 ( .A(n20700), .ZN(n20757) );
  AOI21_X1 U23658 ( .B1(n20702), .B2(n20701), .A(n20757), .ZN(n20707) );
  OAI22_X1 U23659 ( .A1(n20707), .A2(n20852), .B1(n20704), .B2(n20703), .ZN(
        n20755) );
  AOI22_X1 U23660 ( .A1(n20706), .A2(n20757), .B1(n20705), .B2(n20755), .ZN(
        n20715) );
  OAI21_X1 U23661 ( .B1(n20709), .B2(n20708), .A(n20707), .ZN(n20711) );
  OAI221_X1 U23662 ( .B1(n20858), .B2(n20712), .C1(n20852), .C2(n20711), .A(
        n20710), .ZN(n20761) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20713), .ZN(n20714) );
  OAI211_X1 U23664 ( .C1(n20716), .C2(n20764), .A(n20715), .B(n20714), .ZN(
        P1_U3153) );
  AOI22_X1 U23665 ( .A1(n20718), .A2(n20757), .B1(n20717), .B2(n20755), .ZN(
        n20721) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20719), .ZN(n20720) );
  OAI211_X1 U23667 ( .C1(n20722), .C2(n20764), .A(n20721), .B(n20720), .ZN(
        P1_U3154) );
  AOI22_X1 U23668 ( .A1(n20724), .A2(n20757), .B1(n20723), .B2(n20755), .ZN(
        n20727) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20761), .B1(
        n20732), .B2(n20725), .ZN(n20726) );
  OAI211_X1 U23670 ( .C1(n20728), .C2(n20735), .A(n20727), .B(n20726), .ZN(
        P1_U3155) );
  AOI22_X1 U23671 ( .A1(n20730), .A2(n20757), .B1(n20729), .B2(n20755), .ZN(
        n20734) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20761), .B1(
        n20732), .B2(n20731), .ZN(n20733) );
  OAI211_X1 U23673 ( .C1(n20736), .C2(n20735), .A(n20734), .B(n20733), .ZN(
        P1_U3156) );
  AOI22_X1 U23674 ( .A1(n20738), .A2(n20757), .B1(n20737), .B2(n20755), .ZN(
        n20741) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20739), .ZN(n20740) );
  OAI211_X1 U23676 ( .C1(n20742), .C2(n20764), .A(n20741), .B(n20740), .ZN(
        P1_U3157) );
  AOI22_X1 U23677 ( .A1(n20744), .A2(n20757), .B1(n20743), .B2(n20755), .ZN(
        n20747) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20745), .ZN(n20746) );
  OAI211_X1 U23679 ( .C1(n20748), .C2(n20764), .A(n20747), .B(n20746), .ZN(
        P1_U3158) );
  AOI22_X1 U23680 ( .A1(n20750), .A2(n20757), .B1(n20749), .B2(n20755), .ZN(
        n20753) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20751), .ZN(n20752) );
  OAI211_X1 U23682 ( .C1(n20754), .C2(n20764), .A(n20753), .B(n20752), .ZN(
        P1_U3159) );
  AOI22_X1 U23683 ( .A1(n20758), .A2(n20757), .B1(n20756), .B2(n20755), .ZN(
        n20763) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20759), .ZN(n20762) );
  OAI211_X1 U23685 ( .C1(n20765), .C2(n20764), .A(n20763), .B(n20762), .ZN(
        P1_U3160) );
  OAI221_X1 U23686 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20768), .C1(n20703), 
        .C2(n20767), .A(n20766), .ZN(P1_U3163) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20769), .ZN(
        P1_U3164) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20769), .ZN(
        P1_U3165) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20769), .ZN(
        P1_U3166) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20769), .ZN(
        P1_U3167) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20769), .ZN(
        P1_U3168) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20769), .ZN(
        P1_U3169) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20769), .ZN(
        P1_U3170) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20769), .ZN(
        P1_U3171) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20769), .ZN(
        P1_U3172) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20769), .ZN(
        P1_U3173) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20769), .ZN(
        P1_U3174) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20769), .ZN(
        P1_U3175) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20769), .ZN(
        P1_U3176) );
  AND2_X1 U23700 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20769), .ZN(
        P1_U3177) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20769), .ZN(
        P1_U3178) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20769), .ZN(
        P1_U3179) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20769), .ZN(
        P1_U3180) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20769), .ZN(
        P1_U3181) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20769), .ZN(
        P1_U3182) );
  AND2_X1 U23706 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20769), .ZN(
        P1_U3183) );
  AND2_X1 U23707 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20769), .ZN(
        P1_U3184) );
  AND2_X1 U23708 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20769), .ZN(
        P1_U3185) );
  AND2_X1 U23709 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20769), .ZN(P1_U3186) );
  AND2_X1 U23710 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20769), .ZN(P1_U3187) );
  AND2_X1 U23711 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20769), .ZN(P1_U3188) );
  AND2_X1 U23712 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20769), .ZN(P1_U3189) );
  AND2_X1 U23713 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20769), .ZN(P1_U3190) );
  AND2_X1 U23714 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20769), .ZN(P1_U3191) );
  AND2_X1 U23715 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20769), .ZN(P1_U3192) );
  AND2_X1 U23716 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20769), .ZN(P1_U3193) );
  AOI21_X1 U23717 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20876), .A(n20776), 
        .ZN(n20781) );
  NOR2_X1 U23718 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20770) );
  NOR2_X1 U23719 ( .A1(n20770), .A2(n21001), .ZN(n20771) );
  AOI211_X1 U23720 ( .C1(NA), .C2(n20776), .A(n20771), .B(n20971), .ZN(n20772)
         );
  OAI22_X1 U23721 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20781), .B1(n20887), 
        .B2(n20772), .ZN(P1_U3194) );
  NOR2_X1 U23722 ( .A1(NA), .A2(n20971), .ZN(n20775) );
  AOI21_X1 U23723 ( .B1(NA), .B2(n20773), .A(n20782), .ZN(n20774) );
  AOI21_X1 U23724 ( .B1(n20775), .B2(P1_STATE_REG_0__SCAN_IN), .A(n20774), 
        .ZN(n20780) );
  NOR3_X1 U23725 ( .A1(NA), .A2(n20776), .A3(n20880), .ZN(n20777) );
  OAI22_X1 U23726 ( .A1(n20778), .A2(n20777), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20971), .ZN(n20779) );
  OAI22_X1 U23727 ( .A1(n20781), .A2(n20780), .B1(n21001), .B2(n20779), .ZN(
        P1_U3196) );
  INV_X1 U23728 ( .A(n20887), .ZN(n20888) );
  NOR2_X1 U23729 ( .A1(n20782), .A2(n20888), .ZN(n20820) );
  INV_X1 U23730 ( .A(n20820), .ZN(n20799) );
  INV_X1 U23731 ( .A(n20799), .ZN(n20815) );
  AOI222_X1 U23732 ( .A1(n20812), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20815), .ZN(n20783) );
  INV_X1 U23733 ( .A(n20783), .ZN(P1_U3197) );
  INV_X1 U23734 ( .A(n20812), .ZN(n20802) );
  INV_X1 U23735 ( .A(n20802), .ZN(n20819) );
  AOI222_X1 U23736 ( .A1(n20815), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20819), .ZN(n20784) );
  INV_X1 U23737 ( .A(n20784), .ZN(P1_U3198) );
  OAI222_X1 U23738 ( .A1(n20799), .A2(n20786), .B1(n20785), .B2(n20887), .C1(
        n21170), .C2(n20802), .ZN(P1_U3199) );
  AOI222_X1 U23739 ( .A1(n20815), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20819), .ZN(n20787) );
  INV_X1 U23740 ( .A(n20787), .ZN(P1_U3200) );
  AOI222_X1 U23741 ( .A1(n20815), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20819), .ZN(n20788) );
  INV_X1 U23742 ( .A(n20788), .ZN(P1_U3201) );
  AOI222_X1 U23743 ( .A1(n20815), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20819), .ZN(n20789) );
  INV_X1 U23744 ( .A(n20789), .ZN(P1_U3202) );
  AOI222_X1 U23745 ( .A1(n20820), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20819), .ZN(n20790) );
  INV_X1 U23746 ( .A(n20790), .ZN(P1_U3203) );
  AOI222_X1 U23747 ( .A1(n20812), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20815), .ZN(n20791) );
  INV_X1 U23748 ( .A(n20791), .ZN(P1_U3204) );
  AOI222_X1 U23749 ( .A1(n20815), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20819), .ZN(n20792) );
  INV_X1 U23750 ( .A(n20792), .ZN(P1_U3205) );
  AOI222_X1 U23751 ( .A1(n20820), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20819), .ZN(n20793) );
  INV_X1 U23752 ( .A(n20793), .ZN(P1_U3206) );
  AOI222_X1 U23753 ( .A1(n20820), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20819), .ZN(n20794) );
  INV_X1 U23754 ( .A(n20794), .ZN(P1_U3207) );
  AOI222_X1 U23755 ( .A1(n20815), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20819), .ZN(n20795) );
  INV_X1 U23756 ( .A(n20795), .ZN(P1_U3208) );
  AOI222_X1 U23757 ( .A1(n20812), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20815), .ZN(n20796) );
  INV_X1 U23758 ( .A(n20796), .ZN(P1_U3209) );
  AOI222_X1 U23759 ( .A1(n20812), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20815), .ZN(n20797) );
  INV_X1 U23760 ( .A(n20797), .ZN(P1_U3210) );
  AOI22_X1 U23761 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20888), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20812), .ZN(n20798) );
  OAI21_X1 U23762 ( .B1(n20800), .B2(n20799), .A(n20798), .ZN(P1_U3211) );
  AOI22_X1 U23763 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20888), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20820), .ZN(n20801) );
  OAI21_X1 U23764 ( .B1(n21244), .B2(n20802), .A(n20801), .ZN(P1_U3212) );
  AOI222_X1 U23765 ( .A1(n20819), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20815), .ZN(n20803) );
  INV_X1 U23766 ( .A(n20803), .ZN(P1_U3213) );
  AOI222_X1 U23767 ( .A1(n20815), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20819), .ZN(n20804) );
  INV_X1 U23768 ( .A(n20804), .ZN(P1_U3214) );
  AOI222_X1 U23769 ( .A1(n20812), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20815), .ZN(n20805) );
  INV_X1 U23770 ( .A(n20805), .ZN(P1_U3215) );
  AOI222_X1 U23771 ( .A1(n20819), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20815), .ZN(n20806) );
  INV_X1 U23772 ( .A(n20806), .ZN(P1_U3216) );
  AOI222_X1 U23773 ( .A1(n20812), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20820), .ZN(n20807) );
  INV_X1 U23774 ( .A(n20807), .ZN(P1_U3217) );
  AOI222_X1 U23775 ( .A1(n20820), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20819), .ZN(n20808) );
  INV_X1 U23776 ( .A(n20808), .ZN(P1_U3218) );
  AOI222_X1 U23777 ( .A1(n20819), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20815), .ZN(n20809) );
  INV_X1 U23778 ( .A(n20809), .ZN(P1_U3219) );
  AOI222_X1 U23779 ( .A1(n20819), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20815), .ZN(n20810) );
  INV_X1 U23780 ( .A(n20810), .ZN(P1_U3220) );
  AOI222_X1 U23781 ( .A1(n20815), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20819), .ZN(n20811) );
  INV_X1 U23782 ( .A(n20811), .ZN(P1_U3221) );
  AOI222_X1 U23783 ( .A1(n20812), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20815), .ZN(n20813) );
  INV_X1 U23784 ( .A(n20813), .ZN(P1_U3222) );
  AOI222_X1 U23785 ( .A1(n20815), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20814), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20819), .ZN(n20816) );
  INV_X1 U23786 ( .A(n20816), .ZN(P1_U3223) );
  AOI222_X1 U23787 ( .A1(n20820), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20819), .ZN(n20817) );
  INV_X1 U23788 ( .A(n20817), .ZN(P1_U3224) );
  AOI222_X1 U23789 ( .A1(n20820), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20819), .ZN(n20818) );
  INV_X1 U23790 ( .A(n20818), .ZN(P1_U3225) );
  AOI222_X1 U23791 ( .A1(n20820), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20888), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20819), .ZN(n20821) );
  INV_X1 U23792 ( .A(n20821), .ZN(P1_U3226) );
  OAI22_X1 U23793 ( .A1(n20888), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20887), .ZN(n20822) );
  INV_X1 U23794 ( .A(n20822), .ZN(P1_U3458) );
  OAI22_X1 U23795 ( .A1(n20888), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20887), .ZN(n20823) );
  INV_X1 U23796 ( .A(n20823), .ZN(P1_U3459) );
  OAI22_X1 U23797 ( .A1(n20888), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20887), .ZN(n20824) );
  INV_X1 U23798 ( .A(n20824), .ZN(P1_U3460) );
  OAI22_X1 U23799 ( .A1(n20888), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20887), .ZN(n20825) );
  INV_X1 U23800 ( .A(n20825), .ZN(P1_U3461) );
  OAI21_X1 U23801 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20829), .A(n20827), 
        .ZN(n20826) );
  INV_X1 U23802 ( .A(n20826), .ZN(P1_U3464) );
  OAI21_X1 U23803 ( .B1(n20829), .B2(n20828), .A(n20827), .ZN(P1_U3465) );
  INV_X1 U23804 ( .A(n20830), .ZN(n20832) );
  OAI22_X1 U23805 ( .A1(n20832), .A2(n20837), .B1(n20831), .B2(n20841), .ZN(
        n20833) );
  MUX2_X1 U23806 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20833), .S(
        n20844), .Z(P1_U3469) );
  INV_X1 U23807 ( .A(n20834), .ZN(n20839) );
  INV_X1 U23808 ( .A(n20835), .ZN(n20836) );
  OAI222_X1 U23809 ( .A1(n20841), .A2(n20840), .B1(n20839), .B2(n20838), .C1(
        n20837), .C2(n20836), .ZN(n20843) );
  OAI22_X1 U23810 ( .A1(n20844), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20843), .B2(n20842), .ZN(n20845) );
  INV_X1 U23811 ( .A(n20845), .ZN(P1_U3472) );
  AOI211_X1 U23812 ( .C1(n20846), .C2(n21003), .A(n20848), .B(n20847), .ZN(
        n20853) );
  AOI21_X1 U23813 ( .B1(n20860), .B2(n20850), .A(n20849), .ZN(n20851) );
  OAI21_X1 U23814 ( .B1(n20853), .B2(n20852), .A(n20851), .ZN(n20854) );
  NAND2_X1 U23815 ( .A1(n20854), .A2(n20857), .ZN(n20855) );
  OAI21_X1 U23816 ( .B1(n20857), .B2(n20856), .A(n20855), .ZN(P1_U3475) );
  INV_X1 U23817 ( .A(n20857), .ZN(n20865) );
  AOI22_X1 U23818 ( .A1(n20861), .A2(n20860), .B1(n20859), .B2(n20858), .ZN(
        n20864) );
  NOR2_X1 U23819 ( .A1(n20865), .A2(n20862), .ZN(n20863) );
  AOI22_X1 U23820 ( .A1(n20866), .A2(n20865), .B1(n20864), .B2(n20863), .ZN(
        P1_U3478) );
  AOI21_X1 U23821 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20868) );
  AOI22_X1 U23822 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20868), .B2(n20867), .ZN(n20869) );
  INV_X1 U23823 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21219) );
  AOI22_X1 U23824 ( .A1(n20870), .A2(n20869), .B1(n21219), .B2(n20872), .ZN(
        P1_U3481) );
  INV_X1 U23825 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21058) );
  INV_X1 U23826 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21247) );
  NOR2_X1 U23827 ( .A1(n20872), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U23828 ( .A1(n21058), .A2(n20872), .B1(n21247), .B2(n20871), .ZN(
        P1_U3482) );
  AOI22_X1 U23829 ( .A1(n20887), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21056), 
        .B2(n20888), .ZN(P1_U3483) );
  INV_X1 U23830 ( .A(n20873), .ZN(n20874) );
  OAI211_X1 U23831 ( .C1(n20877), .C2(n20876), .A(n20875), .B(n20874), .ZN(
        n20886) );
  INV_X1 U23832 ( .A(n20878), .ZN(n20882) );
  AOI21_X1 U23833 ( .B1(n10434), .B2(n21003), .A(n20879), .ZN(n20881) );
  OAI211_X1 U23834 ( .C1(n20882), .C2(n20881), .A(n20880), .B(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20883) );
  NAND3_X1 U23835 ( .A1(n20886), .A2(n20884), .A3(n20883), .ZN(n20885) );
  OAI21_X1 U23836 ( .B1(n20886), .B2(n20971), .A(n20885), .ZN(P1_U3485) );
  OAI22_X1 U23837 ( .A1(n20888), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20887), .ZN(n20889) );
  INV_X1 U23838 ( .A(n20889), .ZN(P1_U3486) );
  INV_X1 U23839 ( .A(DATAI_4_), .ZN(n21270) );
  XNOR2_X1 U23840 ( .A(n21152), .B(keyinput_g10), .ZN(n20896) );
  AOI22_X1 U23841 ( .A1(DATAI_29_), .A2(keyinput_g3), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_g102), .ZN(n20890) );
  OAI221_X1 U23842 ( .B1(DATAI_29_), .B2(keyinput_g3), .C1(
        P1_EBX_REG_13__SCAN_IN), .C2(keyinput_g102), .A(n20890), .ZN(n20895)
         );
  AOI22_X1 U23843 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(keyinput_g82), .ZN(n20891) );
  OAI221_X1 U23844 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_g82), .A(n20891), .ZN(n20894) );
  AOI22_X1 U23845 ( .A1(DATAI_10_), .A2(keyinput_g22), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(keyinput_g86), .ZN(n20892) );
  OAI221_X1 U23846 ( .B1(DATAI_10_), .B2(keyinput_g22), .C1(
        P1_EBX_REG_29__SCAN_IN), .C2(keyinput_g86), .A(n20892), .ZN(n20893) );
  NOR4_X1 U23847 ( .A1(n20896), .A2(n20895), .A3(n20894), .A4(n20893), .ZN(
        n20924) );
  AOI22_X1 U23848 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n20897) );
  OAI221_X1 U23849 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_g85), .A(n20897), .ZN(n20904) );
  AOI22_X1 U23850 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput_g80), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_g126), .ZN(n20898) );
  OAI221_X1 U23851 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput_g80), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_g126), .A(n20898), .ZN(n20903)
         );
  AOI22_X1 U23852 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(keyinput_g90), .ZN(n20899) );
  OAI221_X1 U23853 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(
        P1_EBX_REG_25__SCAN_IN), .C2(keyinput_g90), .A(n20899), .ZN(n20902) );
  AOI22_X1 U23854 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_g59), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .ZN(n20900) );
  OAI221_X1 U23855 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .C1(
        P1_EBX_REG_11__SCAN_IN), .C2(keyinput_g104), .A(n20900), .ZN(n20901)
         );
  NOR4_X1 U23856 ( .A1(n20904), .A2(n20903), .A3(n20902), .A4(n20901), .ZN(
        n20923) );
  AOI22_X1 U23857 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_g72), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput_g84), .ZN(n20905) );
  OAI221_X1 U23858 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_g72), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_g84), .A(n20905), .ZN(n20912) );
  AOI22_X1 U23859 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        DATAI_30_), .B2(keyinput_g2), .ZN(n20906) );
  OAI221_X1 U23860 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_30_), .C2(keyinput_g2), .A(n20906), .ZN(n20911) );
  AOI22_X1 U23861 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(keyinput_g93), .ZN(n20907) );
  OAI221_X1 U23862 ( .B1(DATAI_11_), .B2(keyinput_g21), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput_g93), .A(n20907), .ZN(n20910) );
  AOI22_X1 U23863 ( .A1(BS16), .A2(keyinput_g35), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(keyinput_g74), .ZN(n20908) );
  OAI221_X1 U23864 ( .B1(BS16), .B2(keyinput_g35), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(keyinput_g74), .A(n20908), .ZN(n20909) );
  NOR4_X1 U23865 ( .A1(n20912), .A2(n20911), .A3(n20910), .A4(n20909), .ZN(
        n20922) );
  AOI22_X1 U23866 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput_g68), .B1(
        P1_EBX_REG_28__SCAN_IN), .B2(keyinput_g87), .ZN(n20913) );
  OAI221_X1 U23867 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput_g68), .C1(
        P1_EBX_REG_28__SCAN_IN), .C2(keyinput_g87), .A(n20913), .ZN(n20920) );
  AOI22_X1 U23868 ( .A1(NA), .A2(keyinput_g34), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(keyinput_g81), .ZN(n20914) );
  OAI221_X1 U23869 ( .B1(NA), .B2(keyinput_g34), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(keyinput_g81), .A(n20914), .ZN(n20919) );
  AOI22_X1 U23870 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(keyinput_g119), .ZN(n20915) );
  OAI221_X1 U23871 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(
        P1_EAX_REG_28__SCAN_IN), .C2(keyinput_g119), .A(n20915), .ZN(n20918)
         );
  AOI22_X1 U23872 ( .A1(DATAI_16_), .A2(keyinput_g16), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n20916) );
  OAI221_X1 U23873 ( .B1(DATAI_16_), .B2(keyinput_g16), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n20916), .ZN(n20917)
         );
  NOR4_X1 U23874 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  NAND4_X1 U23875 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n21070) );
  AOI22_X1 U23876 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .ZN(n20925) );
  OAI221_X1 U23877 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_REIP_REG_8__SCAN_IN), .C2(keyinput_g75), .A(n20925), .ZN(n20932) );
  AOI22_X1 U23878 ( .A1(DATAI_25_), .A2(keyinput_g7), .B1(
        P1_EBX_REG_27__SCAN_IN), .B2(keyinput_g88), .ZN(n20926) );
  OAI221_X1 U23879 ( .B1(DATAI_25_), .B2(keyinput_g7), .C1(
        P1_EBX_REG_27__SCAN_IN), .C2(keyinput_g88), .A(n20926), .ZN(n20931) );
  AOI22_X1 U23880 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_g61), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(keyinput_g117), .ZN(n20927) );
  OAI221_X1 U23881 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_g117), .A(n20927), .ZN(n20930)
         );
  AOI22_X1 U23882 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_g63), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(keyinput_g98), .ZN(n20928) );
  OAI221_X1 U23883 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput_g98), .A(n20928), .ZN(n20929) );
  NOR4_X1 U23884 ( .A1(n20932), .A2(n20931), .A3(n20930), .A4(n20929), .ZN(
        n20964) );
  AOI22_X1 U23885 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(keyinput_g69), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(keyinput_g107), .ZN(n20933) );
  OAI221_X1 U23886 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(keyinput_g69), .C1(
        P1_EBX_REG_8__SCAN_IN), .C2(keyinput_g107), .A(n20933), .ZN(n20940) );
  AOI22_X1 U23887 ( .A1(DATAI_23_), .A2(keyinput_g9), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .ZN(n20934) );
  OAI221_X1 U23888 ( .B1(DATAI_23_), .B2(keyinput_g9), .C1(
        P1_REIP_REG_4__SCAN_IN), .C2(keyinput_g79), .A(n20934), .ZN(n20939) );
  AOI22_X1 U23889 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(keyinput_g99), .ZN(n20935) );
  OAI221_X1 U23890 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        P1_EBX_REG_16__SCAN_IN), .C2(keyinput_g99), .A(n20935), .ZN(n20938) );
  AOI22_X1 U23891 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_g71), .ZN(n20936) );
  OAI221_X1 U23892 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput_g71), .A(n20936), .ZN(n20937)
         );
  NOR4_X1 U23893 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20963) );
  AOI22_X1 U23894 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_g67), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_g125), .ZN(n20941) );
  OAI221_X1 U23895 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_g67), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_g125), .A(n20941), .ZN(n20948)
         );
  AOI22_X1 U23896 ( .A1(DATAI_12_), .A2(keyinput_g20), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(keyinput_g95), .ZN(n20942) );
  OAI221_X1 U23897 ( .B1(DATAI_12_), .B2(keyinput_g20), .C1(
        P1_EBX_REG_20__SCAN_IN), .C2(keyinput_g95), .A(n20942), .ZN(n20947) );
  AOI22_X1 U23898 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(keyinput_g70), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_g66), .ZN(n20943) );
  OAI221_X1 U23899 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(keyinput_g70), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(keyinput_g66), .A(n20943), .ZN(n20946)
         );
  AOI22_X1 U23900 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(keyinput_g96), .ZN(n20944) );
  OAI221_X1 U23901 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        P1_EBX_REG_19__SCAN_IN), .C2(keyinput_g96), .A(n20944), .ZN(n20945) );
  NOR4_X1 U23902 ( .A1(n20948), .A2(n20947), .A3(n20946), .A4(n20945), .ZN(
        n20962) );
  INV_X1 U23903 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n20950) );
  AOI22_X1 U23904 ( .A1(n20951), .A2(keyinput_g78), .B1(n20950), .B2(
        keyinput_g116), .ZN(n20949) );
  OAI221_X1 U23905 ( .B1(n20951), .B2(keyinput_g78), .C1(n20950), .C2(
        keyinput_g116), .A(n20949), .ZN(n20960) );
  AOI22_X1 U23906 ( .A1(n12136), .A2(keyinput_g124), .B1(keyinput_g0), .B2(
        n21205), .ZN(n20952) );
  OAI221_X1 U23907 ( .B1(n12136), .B2(keyinput_g124), .C1(n21205), .C2(
        keyinput_g0), .A(n20952), .ZN(n20959) );
  AOI22_X1 U23908 ( .A1(n21153), .A2(keyinput_g55), .B1(keyinput_g26), .B2(
        n13655), .ZN(n20953) );
  OAI221_X1 U23909 ( .B1(n21153), .B2(keyinput_g55), .C1(n13655), .C2(
        keyinput_g26), .A(n20953), .ZN(n20958) );
  INV_X1 U23910 ( .A(DATAI_31_), .ZN(n20956) );
  AOI22_X1 U23911 ( .A1(n20956), .A2(keyinput_g1), .B1(keyinput_g91), .B2(
        n20955), .ZN(n20954) );
  OAI221_X1 U23912 ( .B1(n20956), .B2(keyinput_g1), .C1(n20955), .C2(
        keyinput_g91), .A(n20954), .ZN(n20957) );
  NOR4_X1 U23913 ( .A1(n20960), .A2(n20959), .A3(n20958), .A4(n20957), .ZN(
        n20961) );
  NAND4_X1 U23914 ( .A1(n20964), .A2(n20963), .A3(n20962), .A4(n20961), .ZN(
        n21069) );
  AOI22_X1 U23915 ( .A1(n20967), .A2(keyinput_g77), .B1(keyinput_g64), .B2(
        n20966), .ZN(n20965) );
  OAI221_X1 U23916 ( .B1(n20967), .B2(keyinput_g77), .C1(n20966), .C2(
        keyinput_g64), .A(n20965), .ZN(n20975) );
  INV_X1 U23917 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n21164) );
  AOI22_X1 U23918 ( .A1(n21164), .A2(keyinput_g94), .B1(keyinput_g113), .B2(
        n10158), .ZN(n20968) );
  OAI221_X1 U23919 ( .B1(n21164), .B2(keyinput_g94), .C1(n10158), .C2(
        keyinput_g113), .A(n20968), .ZN(n20974) );
  AOI22_X1 U23920 ( .A1(n21219), .A2(keyinput_g50), .B1(n13617), .B2(
        keyinput_g25), .ZN(n20969) );
  OAI221_X1 U23921 ( .B1(n21219), .B2(keyinput_g50), .C1(n13617), .C2(
        keyinput_g25), .A(n20969), .ZN(n20973) );
  INV_X1 U23922 ( .A(READY2), .ZN(n21179) );
  AOI22_X1 U23923 ( .A1(n21179), .A2(keyinput_g37), .B1(keyinput_g43), .B2(
        n20971), .ZN(n20970) );
  OAI221_X1 U23924 ( .B1(n21179), .B2(keyinput_g37), .C1(n20971), .C2(
        keyinput_g43), .A(n20970), .ZN(n20972) );
  NOR4_X1 U23925 ( .A1(n20975), .A2(n20974), .A3(n20973), .A4(n20972), .ZN(
        n21015) );
  AOI22_X1 U23926 ( .A1(n12340), .A2(keyinput_g112), .B1(n21184), .B2(
        keyinput_g52), .ZN(n20976) );
  OAI221_X1 U23927 ( .B1(n12340), .B2(keyinput_g112), .C1(n21184), .C2(
        keyinput_g52), .A(n20976), .ZN(n20988) );
  AOI22_X1 U23928 ( .A1(n20979), .A2(keyinput_g105), .B1(keyinput_g51), .B2(
        n20978), .ZN(n20977) );
  OAI221_X1 U23929 ( .B1(n20979), .B2(keyinput_g105), .C1(n20978), .C2(
        keyinput_g51), .A(n20977), .ZN(n20987) );
  INV_X1 U23930 ( .A(DATAI_0_), .ZN(n20981) );
  AOI22_X1 U23931 ( .A1(n20982), .A2(keyinput_g111), .B1(keyinput_g32), .B2(
        n20981), .ZN(n20980) );
  OAI221_X1 U23932 ( .B1(n20982), .B2(keyinput_g111), .C1(n20981), .C2(
        keyinput_g32), .A(n20980), .ZN(n20986) );
  INV_X1 U23933 ( .A(DATAI_26_), .ZN(n20984) );
  AOI22_X1 U23934 ( .A1(n20984), .A2(keyinput_g6), .B1(keyinput_g83), .B2(
        n21247), .ZN(n20983) );
  OAI221_X1 U23935 ( .B1(n20984), .B2(keyinput_g6), .C1(n21247), .C2(
        keyinput_g83), .A(n20983), .ZN(n20985) );
  NOR4_X1 U23936 ( .A1(n20988), .A2(n20987), .A3(n20986), .A4(n20985), .ZN(
        n21014) );
  AOI22_X1 U23937 ( .A1(n20990), .A2(keyinput_g121), .B1(keyinput_g18), .B2(
        n21245), .ZN(n20989) );
  OAI221_X1 U23938 ( .B1(n20990), .B2(keyinput_g121), .C1(n21245), .C2(
        keyinput_g18), .A(n20989), .ZN(n20999) );
  INV_X1 U23939 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21217) );
  AOI22_X1 U23940 ( .A1(n21217), .A2(keyinput_g40), .B1(n12176), .B2(
        keyinput_g122), .ZN(n20991) );
  OAI221_X1 U23941 ( .B1(n21217), .B2(keyinput_g40), .C1(n12176), .C2(
        keyinput_g122), .A(n20991), .ZN(n20998) );
  AOI22_X1 U23942 ( .A1(n20993), .A2(keyinput_g49), .B1(n14676), .B2(
        keyinput_g60), .ZN(n20992) );
  OAI221_X1 U23943 ( .B1(n20993), .B2(keyinput_g49), .C1(n14676), .C2(
        keyinput_g60), .A(n20992), .ZN(n20997) );
  AOI22_X1 U23944 ( .A1(n20995), .A2(keyinput_g115), .B1(keyinput_g24), .B2(
        n21188), .ZN(n20994) );
  OAI221_X1 U23945 ( .B1(n20995), .B2(keyinput_g115), .C1(n21188), .C2(
        keyinput_g24), .A(n20994), .ZN(n20996) );
  NOR4_X1 U23946 ( .A1(n20999), .A2(n20998), .A3(n20997), .A4(n20996), .ZN(
        n21013) );
  AOI22_X1 U23947 ( .A1(n10161), .A2(keyinput_g109), .B1(keyinput_g33), .B2(
        n21001), .ZN(n21000) );
  OAI221_X1 U23948 ( .B1(n10161), .B2(keyinput_g109), .C1(n21001), .C2(
        keyinput_g33), .A(n21000), .ZN(n21011) );
  AOI22_X1 U23949 ( .A1(n21003), .A2(keyinput_g44), .B1(keyinput_g120), .B2(
        n12211), .ZN(n21002) );
  OAI221_X1 U23950 ( .B1(n21003), .B2(keyinput_g44), .C1(n12211), .C2(
        keyinput_g120), .A(n21002), .ZN(n21010) );
  AOI22_X1 U23951 ( .A1(n12248), .A2(keyinput_g118), .B1(keyinput_g13), .B2(
        n21005), .ZN(n21004) );
  OAI221_X1 U23952 ( .B1(n12248), .B2(keyinput_g118), .C1(n21005), .C2(
        keyinput_g13), .A(n21004), .ZN(n21009) );
  AOI22_X1 U23953 ( .A1(n21007), .A2(keyinput_g73), .B1(n21187), .B2(
        keyinput_g54), .ZN(n21006) );
  OAI221_X1 U23954 ( .B1(n21007), .B2(keyinput_g73), .C1(n21187), .C2(
        keyinput_g54), .A(n21006), .ZN(n21008) );
  NOR4_X1 U23955 ( .A1(n21011), .A2(n21010), .A3(n21009), .A4(n21008), .ZN(
        n21012) );
  NAND4_X1 U23956 ( .A1(n21015), .A2(n21014), .A3(n21013), .A4(n21012), .ZN(
        n21068) );
  INV_X1 U23957 ( .A(DATAI_3_), .ZN(n21017) );
  AOI22_X1 U23958 ( .A1(n21017), .A2(keyinput_g29), .B1(n21212), .B2(
        keyinput_g89), .ZN(n21016) );
  OAI221_X1 U23959 ( .B1(n21017), .B2(keyinput_g29), .C1(n21212), .C2(
        keyinput_g89), .A(n21016), .ZN(n21028) );
  AOI22_X1 U23960 ( .A1(n21019), .A2(keyinput_g123), .B1(keyinput_g110), .B2(
        n21242), .ZN(n21018) );
  OAI221_X1 U23961 ( .B1(n21019), .B2(keyinput_g123), .C1(n21242), .C2(
        keyinput_g110), .A(n21018), .ZN(n21027) );
  AOI22_X1 U23962 ( .A1(n21022), .A2(keyinput_g23), .B1(n21021), .B2(
        keyinput_g108), .ZN(n21020) );
  OAI221_X1 U23963 ( .B1(n21022), .B2(keyinput_g23), .C1(n21021), .C2(
        keyinput_g108), .A(n21020), .ZN(n21026) );
  AOI22_X1 U23964 ( .A1(n21235), .A2(keyinput_g114), .B1(keyinput_g12), .B2(
        n21024), .ZN(n21023) );
  OAI221_X1 U23965 ( .B1(n21235), .B2(keyinput_g114), .C1(n21024), .C2(
        keyinput_g12), .A(n21023), .ZN(n21025) );
  NOR4_X1 U23966 ( .A1(n21028), .A2(n21027), .A3(n21026), .A4(n21025), .ZN(
        n21066) );
  AOI22_X1 U23967 ( .A1(n21227), .A2(keyinput_g106), .B1(n10167), .B2(
        keyinput_g103), .ZN(n21029) );
  OAI221_X1 U23968 ( .B1(n21227), .B2(keyinput_g106), .C1(n10167), .C2(
        keyinput_g103), .A(n21029), .ZN(n21038) );
  AOI22_X1 U23969 ( .A1(n21229), .A2(keyinput_g65), .B1(n21214), .B2(
        keyinput_g92), .ZN(n21030) );
  OAI221_X1 U23970 ( .B1(n21229), .B2(keyinput_g65), .C1(n21214), .C2(
        keyinput_g92), .A(n21030), .ZN(n21037) );
  INV_X1 U23971 ( .A(DATAI_27_), .ZN(n21032) );
  INV_X1 U23972 ( .A(DATAI_28_), .ZN(n21185) );
  AOI22_X1 U23973 ( .A1(n21032), .A2(keyinput_g5), .B1(n21185), .B2(
        keyinput_g4), .ZN(n21031) );
  OAI221_X1 U23974 ( .B1(n21032), .B2(keyinput_g5), .C1(n21185), .C2(
        keyinput_g4), .A(n21031), .ZN(n21036) );
  INV_X1 U23975 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21034) );
  AOI22_X1 U23976 ( .A1(n12374), .A2(keyinput_g100), .B1(keyinput_g58), .B2(
        n21034), .ZN(n21033) );
  OAI221_X1 U23977 ( .B1(n12374), .B2(keyinput_g100), .C1(n21034), .C2(
        keyinput_g58), .A(n21033), .ZN(n21035) );
  NOR4_X1 U23978 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21065) );
  AOI22_X1 U23979 ( .A1(n12872), .A2(keyinput_g53), .B1(keyinput_g14), .B2(
        n21198), .ZN(n21039) );
  OAI221_X1 U23980 ( .B1(n12872), .B2(keyinput_g53), .C1(n21198), .C2(
        keyinput_g14), .A(n21039), .ZN(n21051) );
  INV_X1 U23981 ( .A(READY1), .ZN(n21216) );
  AOI22_X1 U23982 ( .A1(n21041), .A2(keyinput_g45), .B1(n21216), .B2(
        keyinput_g36), .ZN(n21040) );
  OAI221_X1 U23983 ( .B1(n21041), .B2(keyinput_g45), .C1(n21216), .C2(
        keyinput_g36), .A(n21040), .ZN(n21050) );
  INV_X1 U23984 ( .A(DATAI_2_), .ZN(n21044) );
  AOI22_X1 U23985 ( .A1(n21044), .A2(keyinput_g30), .B1(n21043), .B2(
        keyinput_g97), .ZN(n21042) );
  OAI221_X1 U23986 ( .B1(n21044), .B2(keyinput_g30), .C1(n21043), .C2(
        keyinput_g97), .A(n21042), .ZN(n21049) );
  INV_X1 U23987 ( .A(DATAI_1_), .ZN(n21046) );
  AOI22_X1 U23988 ( .A1(n21047), .A2(keyinput_g19), .B1(keyinput_g31), .B2(
        n21046), .ZN(n21045) );
  OAI221_X1 U23989 ( .B1(n21047), .B2(keyinput_g19), .C1(n21046), .C2(
        keyinput_g31), .A(n21045), .ZN(n21048) );
  NOR4_X1 U23990 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21064) );
  INV_X1 U23991 ( .A(DATAI_5_), .ZN(n21204) );
  AOI22_X1 U23992 ( .A1(n21053), .A2(keyinput_g42), .B1(n21204), .B2(
        keyinput_g27), .ZN(n21052) );
  OAI221_X1 U23993 ( .B1(n21053), .B2(keyinput_g42), .C1(n21204), .C2(
        keyinput_g27), .A(n21052), .ZN(n21062) );
  AOI22_X1 U23994 ( .A1(n21220), .A2(keyinput_g56), .B1(n21181), .B2(
        keyinput_g76), .ZN(n21054) );
  OAI221_X1 U23995 ( .B1(n21220), .B2(keyinput_g56), .C1(n21181), .C2(
        keyinput_g76), .A(n21054), .ZN(n21061) );
  INV_X1 U23996 ( .A(DATAI_24_), .ZN(n21155) );
  AOI22_X1 U23997 ( .A1(n21056), .A2(keyinput_g47), .B1(n21155), .B2(
        keyinput_g8), .ZN(n21055) );
  OAI221_X1 U23998 ( .B1(n21056), .B2(keyinput_g47), .C1(n21155), .C2(
        keyinput_g8), .A(n21055), .ZN(n21060) );
  AOI22_X1 U23999 ( .A1(n21058), .A2(keyinput_g48), .B1(n13586), .B2(
        keyinput_g17), .ZN(n21057) );
  OAI221_X1 U24000 ( .B1(n21058), .B2(keyinput_g48), .C1(n13586), .C2(
        keyinput_g17), .A(n21057), .ZN(n21059) );
  NOR4_X1 U24001 ( .A1(n21062), .A2(n21061), .A3(n21060), .A4(n21059), .ZN(
        n21063) );
  NAND4_X1 U24002 ( .A1(n21066), .A2(n21065), .A3(n21064), .A4(n21063), .ZN(
        n21067) );
  NOR4_X1 U24003 ( .A1(n21070), .A2(n21069), .A3(n21068), .A4(n21067), .ZN(
        n21269) );
  OAI22_X1 U24004 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_f88), .B1(
        keyinput_f33), .B2(HOLD), .ZN(n21071) );
  AOI221_X1 U24005 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_f88), .C1(HOLD), 
        .C2(keyinput_f33), .A(n21071), .ZN(n21078) );
  OAI22_X1 U24006 ( .A1(DATAI_3_), .A2(keyinput_f29), .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_f47), .ZN(n21072) );
  AOI221_X1 U24007 ( .B1(DATAI_3_), .B2(keyinput_f29), .C1(keyinput_f47), .C2(
        P1_W_R_N_REG_SCAN_IN), .A(n21072), .ZN(n21077) );
  OAI22_X1 U24008 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_f58), .B1(
        DATAI_29_), .B2(keyinput_f3), .ZN(n21073) );
  AOI221_X1 U24009 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .C1(
        keyinput_f3), .C2(DATAI_29_), .A(n21073), .ZN(n21076) );
  OAI22_X1 U24010 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_f112), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(keyinput_f80), .ZN(n21074) );
  AOI221_X1 U24011 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_f112), .C1(
        keyinput_f80), .C2(P1_REIP_REG_3__SCAN_IN), .A(n21074), .ZN(n21075) );
  NAND4_X1 U24012 ( .A1(n21078), .A2(n21077), .A3(n21076), .A4(n21075), .ZN(
        n21106) );
  OAI22_X1 U24013 ( .A1(DATAI_20_), .A2(keyinput_f12), .B1(keyinput_f49), .B2(
        P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21079) );
  AOI221_X1 U24014 ( .B1(DATAI_20_), .B2(keyinput_f12), .C1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_f49), .A(n21079), .ZN(
        n21086) );
  OAI22_X1 U24015 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f26), .B2(DATAI_6_), .ZN(n21080) );
  AOI221_X1 U24016 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .C1(
        DATAI_6_), .C2(keyinput_f26), .A(n21080), .ZN(n21085) );
  OAI22_X1 U24017 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_f120), .B1(
        keyinput_f105), .B2(P1_EBX_REG_10__SCAN_IN), .ZN(n21081) );
  AOI221_X1 U24018 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .C1(
        P1_EBX_REG_10__SCAN_IN), .C2(keyinput_f105), .A(n21081), .ZN(n21084)
         );
  OAI22_X1 U24019 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_f87), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(keyinput_f82), .ZN(n21082) );
  AOI221_X1 U24020 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_f87), .C1(
        keyinput_f82), .C2(P1_REIP_REG_1__SCAN_IN), .A(n21082), .ZN(n21083) );
  NAND4_X1 U24021 ( .A1(n21086), .A2(n21085), .A3(n21084), .A4(n21083), .ZN(
        n21105) );
  OAI22_X1 U24022 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_f116), .B1(
        keyinput_f97), .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n21087) );
  AOI221_X1 U24023 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_f116), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_f97), .A(n21087), .ZN(n21094) );
  OAI22_X1 U24024 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_f75), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_f48), .ZN(n21088) );
  AOI221_X1 U24025 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_f75), .C1(
        keyinput_f48), .C2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21088), .ZN(
        n21093) );
  OAI22_X1 U24026 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(NA), 
        .B2(keyinput_f34), .ZN(n21089) );
  AOI221_X1 U24027 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f34), .C2(NA), .A(n21089), .ZN(n21092) );
  OAI22_X1 U24028 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_f123), .B1(
        keyinput_f115), .B2(P1_EBX_REG_0__SCAN_IN), .ZN(n21090) );
  AOI221_X1 U24029 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .C1(
        P1_EBX_REG_0__SCAN_IN), .C2(keyinput_f115), .A(n21090), .ZN(n21091) );
  NAND4_X1 U24030 ( .A1(n21094), .A2(n21093), .A3(n21092), .A4(n21091), .ZN(
        n21104) );
  OAI22_X1 U24031 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput_f77), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(keyinput_f78), .ZN(n21095) );
  AOI221_X1 U24032 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput_f77), .C1(
        keyinput_f78), .C2(P1_REIP_REG_5__SCAN_IN), .A(n21095), .ZN(n21102) );
  OAI22_X1 U24033 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_f103), .B1(
        keyinput_f72), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n21096) );
  AOI221_X1 U24034 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .C1(
        P1_REIP_REG_11__SCAN_IN), .C2(keyinput_f72), .A(n21096), .ZN(n21101)
         );
  OAI22_X1 U24035 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_f67), .B1(
        keyinput_f16), .B2(DATAI_16_), .ZN(n21097) );
  AOI221_X1 U24036 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .C1(
        DATAI_16_), .C2(keyinput_f16), .A(n21097), .ZN(n21100) );
  OAI22_X1 U24037 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput_f127), .B1(
        keyinput_f31), .B2(DATAI_1_), .ZN(n21098) );
  AOI221_X1 U24038 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput_f127), .C1(
        DATAI_1_), .C2(keyinput_f31), .A(n21098), .ZN(n21099) );
  NAND4_X1 U24039 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21103) );
  NOR4_X1 U24040 ( .A1(n21106), .A2(n21105), .A3(n21104), .A4(n21103), .ZN(
        n21265) );
  OAI22_X1 U24041 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        keyinput_f109), .B2(P1_EBX_REG_6__SCAN_IN), .ZN(n21107) );
  AOI221_X1 U24042 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        P1_EBX_REG_6__SCAN_IN), .C2(keyinput_f109), .A(n21107), .ZN(n21114) );
  OAI22_X1 U24043 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_f122), .B1(BS16), 
        .B2(keyinput_f35), .ZN(n21108) );
  AOI221_X1 U24044 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_f122), .C1(
        keyinput_f35), .C2(BS16), .A(n21108), .ZN(n21113) );
  OAI22_X1 U24045 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        keyinput_f38), .B2(P1_READREQUEST_REG_SCAN_IN), .ZN(n21109) );
  AOI221_X1 U24046 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_f38), .A(n21109), .ZN(n21112) );
  OAI22_X1 U24047 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(keyinput_f70), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(keyinput_f73), .ZN(n21110) );
  AOI221_X1 U24048 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(keyinput_f70), .C1(
        keyinput_f73), .C2(P1_REIP_REG_10__SCAN_IN), .A(n21110), .ZN(n21111)
         );
  NAND4_X1 U24049 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21263) );
  OAI22_X1 U24050 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(keyinput_f121), .B1(
        keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .ZN(n21115) );
  AOI221_X1 U24051 ( .B1(P1_EAX_REG_26__SCAN_IN), .B2(keyinput_f121), .C1(
        P1_M_IO_N_REG_SCAN_IN), .C2(keyinput_f41), .A(n21115), .ZN(n21141) );
  INV_X1 U24052 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21121) );
  OAI22_X1 U24053 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(keyinput_f108), .B1(
        keyinput_f59), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n21116) );
  AOI221_X1 U24054 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(keyinput_f108), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_f59), .A(n21116), .ZN(n21119)
         );
  OAI22_X1 U24055 ( .A1(DATAI_13_), .A2(keyinput_f19), .B1(keyinput_f43), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21117) );
  AOI221_X1 U24056 ( .B1(DATAI_13_), .B2(keyinput_f19), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f43), .A(n21117), .ZN(
        n21118) );
  OAI211_X1 U24057 ( .C1(n21121), .C2(keyinput_f81), .A(n21119), .B(n21118), 
        .ZN(n21120) );
  AOI21_X1 U24058 ( .B1(n21121), .B2(keyinput_f81), .A(n21120), .ZN(n21140) );
  AOI22_X1 U24059 ( .A1(DATAI_2_), .A2(keyinput_f30), .B1(DATAI_25_), .B2(
        keyinput_f7), .ZN(n21122) );
  OAI221_X1 U24060 ( .B1(DATAI_2_), .B2(keyinput_f30), .C1(DATAI_25_), .C2(
        keyinput_f7), .A(n21122), .ZN(n21129) );
  AOI22_X1 U24061 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(keyinput_f102), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(keyinput_f96), .ZN(n21123) );
  OAI221_X1 U24062 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(keyinput_f102), .C1(
        P1_EBX_REG_19__SCAN_IN), .C2(keyinput_f96), .A(n21123), .ZN(n21128) );
  AOI22_X1 U24063 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .ZN(n21124) );
  OAI221_X1 U24064 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(P1_REIP_REG_21__SCAN_IN), .C2(keyinput_f62), .A(n21124), .ZN(
        n21127) );
  AOI22_X1 U24065 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(DATAI_31_), .B2(
        keyinput_f1), .ZN(n21125) );
  OAI221_X1 U24066 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(DATAI_31_), .C2(
        keyinput_f1), .A(n21125), .ZN(n21126) );
  NOR4_X1 U24067 ( .A1(n21129), .A2(n21128), .A3(n21127), .A4(n21126), .ZN(
        n21139) );
  AOI22_X1 U24068 ( .A1(DATAI_0_), .A2(keyinput_f32), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n21130) );
  OAI221_X1 U24069 ( .B1(DATAI_0_), .B2(keyinput_f32), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n21130), .ZN(n21137)
         );
  AOI22_X1 U24070 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_f71), .ZN(n21131) );
  OAI221_X1 U24071 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput_f71), .A(n21131), .ZN(n21136)
         );
  AOI22_X1 U24072 ( .A1(DATAI_27_), .A2(keyinput_f5), .B1(
        P1_EBX_REG_24__SCAN_IN), .B2(keyinput_f91), .ZN(n21132) );
  OAI221_X1 U24073 ( .B1(DATAI_27_), .B2(keyinput_f5), .C1(
        P1_EBX_REG_24__SCAN_IN), .C2(keyinput_f91), .A(n21132), .ZN(n21135) );
  AOI22_X1 U24074 ( .A1(DATAI_12_), .A2(keyinput_f20), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(keyinput_f98), .ZN(n21133) );
  OAI221_X1 U24075 ( .B1(DATAI_12_), .B2(keyinput_f20), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput_f98), .A(n21133), .ZN(n21134) );
  NOR4_X1 U24076 ( .A1(n21137), .A2(n21136), .A3(n21135), .A4(n21134), .ZN(
        n21138) );
  NAND4_X1 U24077 ( .A1(n21141), .A2(n21140), .A3(n21139), .A4(n21138), .ZN(
        n21262) );
  AOI22_X1 U24078 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(keyinput_f68), .ZN(n21142) );
  OAI221_X1 U24079 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        P1_REIP_REG_15__SCAN_IN), .C2(keyinput_f68), .A(n21142), .ZN(n21149)
         );
  AOI22_X1 U24080 ( .A1(DATAI_17_), .A2(keyinput_f15), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(keyinput_f64), .ZN(n21143) );
  OAI221_X1 U24081 ( .B1(DATAI_17_), .B2(keyinput_f15), .C1(
        P1_REIP_REG_19__SCAN_IN), .C2(keyinput_f64), .A(n21143), .ZN(n21148)
         );
  AOI22_X1 U24082 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .ZN(n21144) );
  OAI221_X1 U24083 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_f61), .A(n21144), .ZN(n21147)
         );
  AOI22_X1 U24084 ( .A1(DATAI_23_), .A2(keyinput_f9), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(keyinput_f95), .ZN(n21145) );
  OAI221_X1 U24085 ( .B1(DATAI_23_), .B2(keyinput_f9), .C1(
        P1_EBX_REG_20__SCAN_IN), .C2(keyinput_f95), .A(n21145), .ZN(n21146) );
  NOR4_X1 U24086 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21196) );
  AOI22_X1 U24087 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n21150) );
  OAI221_X1 U24088 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        P1_FLUSH_REG_SCAN_IN), .C2(keyinput_f46), .A(n21150), .ZN(n21162) );
  AOI22_X1 U24089 ( .A1(n21153), .A2(keyinput_f55), .B1(keyinput_f10), .B2(
        n21152), .ZN(n21151) );
  OAI221_X1 U24090 ( .B1(n21153), .B2(keyinput_f55), .C1(n21152), .C2(
        keyinput_f10), .A(n21151), .ZN(n21161) );
  AOI22_X1 U24091 ( .A1(n12248), .A2(keyinput_f118), .B1(keyinput_f8), .B2(
        n21155), .ZN(n21154) );
  OAI221_X1 U24092 ( .B1(n12248), .B2(keyinput_f118), .C1(n21155), .C2(
        keyinput_f8), .A(n21154), .ZN(n21160) );
  AOI22_X1 U24093 ( .A1(n21158), .A2(keyinput_f11), .B1(n21157), .B2(
        keyinput_f126), .ZN(n21156) );
  OAI221_X1 U24094 ( .B1(n21158), .B2(keyinput_f11), .C1(n21157), .C2(
        keyinput_f126), .A(n21156), .ZN(n21159) );
  NOR4_X1 U24095 ( .A1(n21162), .A2(n21161), .A3(n21160), .A4(n21159), .ZN(
        n21195) );
  AOI22_X1 U24096 ( .A1(n21165), .A2(keyinput_f86), .B1(keyinput_f94), .B2(
        n21164), .ZN(n21163) );
  OAI221_X1 U24097 ( .B1(n21165), .B2(keyinput_f86), .C1(n21164), .C2(
        keyinput_f94), .A(n21163), .ZN(n21176) );
  AOI22_X1 U24098 ( .A1(n21168), .A2(keyinput_f93), .B1(keyinput_f84), .B2(
        n21167), .ZN(n21166) );
  OAI221_X1 U24099 ( .B1(n21168), .B2(keyinput_f93), .C1(n21167), .C2(
        keyinput_f84), .A(n21166), .ZN(n21175) );
  AOI22_X1 U24100 ( .A1(n10158), .A2(keyinput_f113), .B1(keyinput_f79), .B2(
        n21170), .ZN(n21169) );
  OAI221_X1 U24101 ( .B1(n10158), .B2(keyinput_f113), .C1(n21170), .C2(
        keyinput_f79), .A(n21169), .ZN(n21174) );
  AOI22_X1 U24102 ( .A1(n21172), .A2(keyinput_f63), .B1(n12872), .B2(
        keyinput_f53), .ZN(n21171) );
  OAI221_X1 U24103 ( .B1(n21172), .B2(keyinput_f63), .C1(n12872), .C2(
        keyinput_f53), .A(n21171), .ZN(n21173) );
  NOR4_X1 U24104 ( .A1(n21176), .A2(n21175), .A3(n21174), .A4(n21173), .ZN(
        n21194) );
  AOI22_X1 U24105 ( .A1(n21179), .A2(keyinput_f37), .B1(n21178), .B2(
        keyinput_f125), .ZN(n21177) );
  OAI221_X1 U24106 ( .B1(n21179), .B2(keyinput_f37), .C1(n21178), .C2(
        keyinput_f125), .A(n21177), .ZN(n21192) );
  AOI22_X1 U24107 ( .A1(n21182), .A2(keyinput_f21), .B1(n21181), .B2(
        keyinput_f76), .ZN(n21180) );
  OAI221_X1 U24108 ( .B1(n21182), .B2(keyinput_f21), .C1(n21181), .C2(
        keyinput_f76), .A(n21180), .ZN(n21191) );
  AOI22_X1 U24109 ( .A1(n21185), .A2(keyinput_f4), .B1(n21184), .B2(
        keyinput_f52), .ZN(n21183) );
  OAI221_X1 U24110 ( .B1(n21185), .B2(keyinput_f4), .C1(n21184), .C2(
        keyinput_f52), .A(n21183), .ZN(n21190) );
  AOI22_X1 U24111 ( .A1(n21188), .A2(keyinput_f24), .B1(n21187), .B2(
        keyinput_f54), .ZN(n21186) );
  OAI221_X1 U24112 ( .B1(n21188), .B2(keyinput_f24), .C1(n21187), .C2(
        keyinput_f54), .A(n21186), .ZN(n21189) );
  NOR4_X1 U24113 ( .A1(n21192), .A2(n21191), .A3(n21190), .A4(n21189), .ZN(
        n21193) );
  NAND4_X1 U24114 ( .A1(n21196), .A2(n21195), .A3(n21194), .A4(n21193), .ZN(
        n21261) );
  AOI22_X1 U24115 ( .A1(n21199), .A2(keyinput_f57), .B1(keyinput_f14), .B2(
        n21198), .ZN(n21197) );
  OAI221_X1 U24116 ( .B1(n21199), .B2(keyinput_f57), .C1(n21198), .C2(
        keyinput_f14), .A(n21197), .ZN(n21209) );
  AOI22_X1 U24117 ( .A1(n12374), .A2(keyinput_f100), .B1(n21201), .B2(
        keyinput_f119), .ZN(n21200) );
  OAI221_X1 U24118 ( .B1(n12374), .B2(keyinput_f100), .C1(n21201), .C2(
        keyinput_f119), .A(n21200), .ZN(n21208) );
  AOI22_X1 U24119 ( .A1(n13586), .A2(keyinput_f17), .B1(n12136), .B2(
        keyinput_f124), .ZN(n21202) );
  OAI221_X1 U24120 ( .B1(n13586), .B2(keyinput_f17), .C1(n12136), .C2(
        keyinput_f124), .A(n21202), .ZN(n21207) );
  AOI22_X1 U24121 ( .A1(n21205), .A2(keyinput_f0), .B1(n21204), .B2(
        keyinput_f27), .ZN(n21203) );
  OAI221_X1 U24122 ( .B1(n21205), .B2(keyinput_f0), .C1(n21204), .C2(
        keyinput_f27), .A(n21203), .ZN(n21206) );
  NOR4_X1 U24123 ( .A1(n21209), .A2(n21208), .A3(n21207), .A4(n21206), .ZN(
        n21259) );
  AOI22_X1 U24124 ( .A1(n21212), .A2(keyinput_f89), .B1(keyinput_f90), .B2(
        n21211), .ZN(n21210) );
  OAI221_X1 U24125 ( .B1(n21212), .B2(keyinput_f89), .C1(n21211), .C2(
        keyinput_f90), .A(n21210), .ZN(n21224) );
  AOI22_X1 U24126 ( .A1(n10164), .A2(keyinput_f107), .B1(n21214), .B2(
        keyinput_f92), .ZN(n21213) );
  OAI221_X1 U24127 ( .B1(n10164), .B2(keyinput_f107), .C1(n21214), .C2(
        keyinput_f92), .A(n21213), .ZN(n21223) );
  AOI22_X1 U24128 ( .A1(n21217), .A2(keyinput_f40), .B1(n21216), .B2(
        keyinput_f36), .ZN(n21215) );
  OAI221_X1 U24129 ( .B1(n21217), .B2(keyinput_f40), .C1(n21216), .C2(
        keyinput_f36), .A(n21215), .ZN(n21222) );
  AOI22_X1 U24130 ( .A1(n21220), .A2(keyinput_f56), .B1(keyinput_f50), .B2(
        n21219), .ZN(n21218) );
  OAI221_X1 U24131 ( .B1(n21220), .B2(keyinput_f56), .C1(n21219), .C2(
        keyinput_f50), .A(n21218), .ZN(n21221) );
  NOR4_X1 U24132 ( .A1(n21224), .A2(n21223), .A3(n21222), .A4(n21221), .ZN(
        n21258) );
  AOI22_X1 U24133 ( .A1(n21227), .A2(keyinput_f106), .B1(keyinput_f39), .B2(
        n21226), .ZN(n21225) );
  OAI221_X1 U24134 ( .B1(n21227), .B2(keyinput_f106), .C1(n21226), .C2(
        keyinput_f39), .A(n21225), .ZN(n21239) );
  AOI22_X1 U24135 ( .A1(n21230), .A2(keyinput_f104), .B1(keyinput_f65), .B2(
        n21229), .ZN(n21228) );
  OAI221_X1 U24136 ( .B1(n21230), .B2(keyinput_f104), .C1(n21229), .C2(
        keyinput_f65), .A(n21228), .ZN(n21238) );
  AOI22_X1 U24137 ( .A1(n13617), .A2(keyinput_f25), .B1(n21232), .B2(
        keyinput_f69), .ZN(n21231) );
  OAI221_X1 U24138 ( .B1(n13617), .B2(keyinput_f25), .C1(n21232), .C2(
        keyinput_f69), .A(n21231), .ZN(n21237) );
  AOI22_X1 U24139 ( .A1(n21235), .A2(keyinput_f114), .B1(keyinput_f22), .B2(
        n21234), .ZN(n21233) );
  OAI221_X1 U24140 ( .B1(n21235), .B2(keyinput_f114), .C1(n21234), .C2(
        keyinput_f22), .A(n21233), .ZN(n21236) );
  NOR4_X1 U24141 ( .A1(n21239), .A2(n21238), .A3(n21237), .A4(n21236), .ZN(
        n21257) );
  INV_X1 U24142 ( .A(DATAI_30_), .ZN(n21241) );
  AOI22_X1 U24143 ( .A1(n21242), .A2(keyinput_f110), .B1(keyinput_f2), .B2(
        n21241), .ZN(n21240) );
  OAI221_X1 U24144 ( .B1(n21242), .B2(keyinput_f110), .C1(n21241), .C2(
        keyinput_f2), .A(n21240), .ZN(n21255) );
  AOI22_X1 U24145 ( .A1(n21245), .A2(keyinput_f18), .B1(n21244), .B2(
        keyinput_f66), .ZN(n21243) );
  OAI221_X1 U24146 ( .B1(n21245), .B2(keyinput_f18), .C1(n21244), .C2(
        keyinput_f66), .A(n21243), .ZN(n21254) );
  AOI22_X1 U24147 ( .A1(n21248), .A2(keyinput_f99), .B1(keyinput_f83), .B2(
        n21247), .ZN(n21246) );
  OAI221_X1 U24148 ( .B1(n21248), .B2(keyinput_f99), .C1(n21247), .C2(
        keyinput_f83), .A(n21246), .ZN(n21253) );
  AOI22_X1 U24149 ( .A1(n21251), .A2(keyinput_f74), .B1(n21250), .B2(
        keyinput_f117), .ZN(n21249) );
  OAI221_X1 U24150 ( .B1(n21251), .B2(keyinput_f74), .C1(n21250), .C2(
        keyinput_f117), .A(n21249), .ZN(n21252) );
  NOR4_X1 U24151 ( .A1(n21255), .A2(n21254), .A3(n21253), .A4(n21252), .ZN(
        n21256) );
  NAND4_X1 U24152 ( .A1(n21259), .A2(n21258), .A3(n21257), .A4(n21256), .ZN(
        n21260) );
  NOR4_X1 U24153 ( .A1(n21263), .A2(n21262), .A3(n21261), .A4(n21260), .ZN(
        n21264) );
  AOI22_X1 U24154 ( .A1(n21265), .A2(n21264), .B1(keyinput_f28), .B2(DATAI_4_), 
        .ZN(n21266) );
  OAI21_X1 U24155 ( .B1(keyinput_f28), .B2(DATAI_4_), .A(n21266), .ZN(n21267)
         );
  OAI21_X1 U24156 ( .B1(n21270), .B2(keyinput_g28), .A(n21267), .ZN(n21268) );
  AOI211_X1 U24157 ( .C1(n21270), .C2(keyinput_g28), .A(n21269), .B(n21268), 
        .ZN(n21272) );
  AOI22_X1 U24158 ( .A1(n16641), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16643), .ZN(n21271) );
  XNOR2_X1 U24159 ( .A(n21272), .B(n21271), .ZN(U355) );
  CLKBUF_X3 U14663 ( .A(n11668), .Z(n12063) );
  BUF_X1 U11464 ( .A(n12105), .Z(n12084) );
  BUF_X2 U11247 ( .A(n12327), .Z(n12404) );
  CLKBUF_X1 U11264 ( .A(n11668), .Z(n12541) );
  AND2_X1 U11273 ( .A1(n13377), .A2(n11488), .ZN(n11600) );
  CLKBUF_X1 U11274 ( .A(n11096), .Z(n11138) );
  OR2_X1 U11286 ( .A1(n15176), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9950) );
  CLKBUF_X1 U11295 ( .A(n11622), .Z(n14846) );
  CLKBUF_X1 U11297 ( .A(n12617), .Z(n20456) );
  CLKBUF_X1 U12707 ( .A(n14364), .Z(n14378) );
  INV_X1 U12932 ( .A(n10501), .ZN(n9801) );
endmodule

