

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916;

  NAND2_X1 U2304 ( .A1(n3593), .A2(n3594), .ZN(n3595) );
  AOI21_X1 U2305 ( .B1(n3189), .B2(n3188), .A(n3187), .ZN(n3203) );
  CLKBUF_X2 U2306 ( .A(n2881), .Z(n3075) );
  AND2_X2 U2308 ( .A1(n3162), .A2(n3163), .ZN(n3302) );
  NAND2_X1 U2309 ( .A1(n2517), .A2(n2516), .ZN(n2271) );
  NOR2_X1 U2310 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2504)
         );
  NOR4_X1 U2312 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4386), .ZN(n4158)
         );
  OAI22_X1 U2313 ( .A1(n4736), .A2(n4733), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3619), .ZN(n3600) );
  OR2_X1 U2314 ( .A1(n4221), .A2(n4220), .ZN(n4243) );
  INV_X1 U2315 ( .A(n2273), .ZN(n3837) );
  OAI211_X1 U2316 ( .C1(n3166), .C2(n2278), .A(n3165), .B(n2495), .ZN(n3189)
         );
  NAND2_X1 U2317 ( .A1(n2517), .A2(n2516), .ZN(n2525) );
  OR2_X1 U2318 ( .A1(n4257), .A2(n4256), .ZN(n2443) );
  INV_X1 U2319 ( .A(IR_REG_31__SCAN_IN), .ZN(n3113) );
  XNOR2_X1 U2320 ( .A(n2623), .B(IR_REG_30__SCAN_IN), .ZN(n4648) );
  AND2_X1 U2321 ( .A1(n2323), .A2(n2288), .ZN(n2269) );
  NOR2_X2 U2322 ( .A1(n3208), .A2(n2294), .ZN(n3210) );
  NAND4_X2 U2323 ( .A1(n3039), .A2(n3038), .A3(n3037), .A4(n3036), .ZN(n4299)
         );
  NAND2_X1 U2324 ( .A1(n2517), .A2(n2516), .ZN(n2270) );
  NOR2_X2 U2325 ( .A1(n3026), .A2(n2420), .ZN(n2416) );
  NOR2_X2 U2326 ( .A1(n3212), .A2(n3213), .ZN(n3238) );
  AND2_X4 U2327 ( .A1(n4648), .A2(n2842), .ZN(n2879) );
  OAI22_X2 U2328 ( .A1(n3423), .A2(n3422), .B1(n3421), .B2(n3420), .ZN(n3465)
         );
  AND2_X2 U2329 ( .A1(n2332), .A2(n2331), .ZN(n3423) );
  CLKBUF_X1 U2330 ( .A(n3302), .Z(n2272) );
  NOR2_X2 U2331 ( .A1(n4669), .A2(n3291), .ZN(n4680) );
  XNOR2_X2 U2332 ( .A(n2406), .B(IR_REG_2__SCAN_IN), .ZN(n3143) );
  INV_X1 U2333 ( .A(n2273), .ZN(n2279) );
  AND2_X1 U2334 ( .A1(n3184), .A2(n3163), .ZN(n2287) );
  AND2_X1 U2335 ( .A1(n2443), .A2(n2442), .ZN(n4758) );
  NOR2_X1 U2336 ( .A1(n3600), .A2(n4224), .ZN(n4216) );
  AOI221_X1 U2337 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_122), .C1(n2831), 
        .C2(n2729), .A(n2728), .ZN(n2730) );
  NAND2_X1 U2338 ( .A1(n4284), .A2(n4280), .ZN(n3092) );
  AOI221_X1 U2339 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_58), .C1(n2831), .C2(
        n2830), .A(n2829), .ZN(n2832) );
  NOR2_X1 U2340 ( .A1(n4306), .A2(n3853), .ZN(n4284) );
  NAND2_X1 U2341 ( .A1(n2453), .A2(n2452), .ZN(n2457) );
  OR2_X1 U2342 ( .A1(n4337), .A2(n3024), .ZN(n4314) );
  NOR2_X2 U2343 ( .A1(n3242), .A2(n3241), .ZN(n3948) );
  AND2_X1 U2344 ( .A1(n3004), .A2(REG3_REG_24__SCAN_IN), .ZN(n3016) );
  OAI22_X1 U2345 ( .A1(n3337), .A2(n2898), .B1(n3390), .B2(n3338), .ZN(n3388)
         );
  INV_X1 U2346 ( .A(n2275), .ZN(n2276) );
  INV_X1 U2347 ( .A(n2275), .ZN(n2277) );
  INV_X1 U2348 ( .A(n2287), .ZN(n2275) );
  INV_X1 U2349 ( .A(n3184), .ZN(n3162) );
  NAND2_X1 U2350 ( .A1(n4070), .A2(n4067), .ZN(n4128) );
  NAND2_X1 U2351 ( .A1(n2286), .A2(n2877), .ZN(n4190) );
  NAND2_X1 U2352 ( .A1(n2290), .A2(n2885), .ZN(n4188) );
  NAND2_X1 U2353 ( .A1(n2608), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  NAND4_X1 U2354 ( .A1(n2867), .A2(n2866), .A3(n2865), .A4(n2864), .ZN(n4187)
         );
  AND2_X1 U2355 ( .A1(n3221), .A2(REG2_REG_4__SCAN_IN), .ZN(n3285) );
  CLKBUF_X1 U2356 ( .A(n3284), .Z(n3286) );
  INV_X1 U2357 ( .A(n3256), .ZN(n3737) );
  NAND3_X1 U2358 ( .A1(n4650), .A2(n4649), .A3(n3106), .ZN(n3163) );
  NAND2_X1 U2359 ( .A1(n2390), .A2(IR_REG_31__SCAN_IN), .ZN(n2623) );
  XNOR2_X1 U2360 ( .A(n2614), .B(IR_REG_21__SCAN_IN), .ZN(n4157) );
  OR2_X1 U2361 ( .A1(n2630), .A2(n2309), .ZN(n2517) );
  NOR2_X1 U2362 ( .A1(n2491), .A2(IR_REG_21__SCAN_IN), .ZN(n2490) );
  OR2_X1 U2363 ( .A1(n2492), .A2(IR_REG_25__SCAN_IN), .ZN(n2491) );
  AND2_X1 U2364 ( .A1(n2568), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  AND2_X1 U2365 ( .A1(n2496), .A2(n2503), .ZN(n2450) );
  AND2_X1 U2366 ( .A1(n2502), .A2(n2831), .ZN(n2496) );
  AND4_X1 U2367 ( .A1(n2506), .A2(n2504), .A3(n2505), .A4(n2507), .ZN(n2449)
         );
  NOR2_X1 U2368 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2506)
         );
  NOR2_X1 U2369 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2503)
         );
  NOR2_X1 U2370 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2505)
         );
  NOR2_X1 U2371 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2567)
         );
  NOR2_X2 U2372 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2519)
         );
  NAND2_X4 U2373 ( .A1(n2287), .A2(n3164), .ZN(n3827) );
  INV_X2 U2374 ( .A(IR_REG_3__SCAN_IN), .ZN(n2831) );
  NAND2_X1 U2375 ( .A1(n4246), .A2(n4247), .ZN(n4253) );
  NOR2_X2 U2376 ( .A1(n2570), .A2(n2569), .ZN(n2574) );
  XNOR2_X2 U2377 ( .A(n2610), .B(n2609), .ZN(n3046) );
  BUF_X2 U2378 ( .A(n3046), .Z(n2619) );
  INV_X1 U2379 ( .A(n2272), .ZN(n2278) );
  AND2_X1 U2380 ( .A1(n3162), .A2(n3163), .ZN(n2280) );
  AND2_X1 U2381 ( .A1(n3162), .A2(n3163), .ZN(n2281) );
  OAI21_X2 U2382 ( .B1(n3747), .B2(n2462), .A(n2459), .ZN(n2333) );
  AOI21_X2 U2383 ( .B1(n2269), .B2(n3585), .A(n3584), .ZN(n3747) );
  INV_X2 U2384 ( .A(n3855), .ZN(n3835) );
  AOI21_X1 U2385 ( .B1(n2424), .B2(n4376), .A(n2422), .ZN(n2421) );
  INV_X1 U2386 ( .A(n4379), .ZN(n2422) );
  INV_X1 U2387 ( .A(IR_REG_26__SCAN_IN), .ZN(n2335) );
  NOR2_X1 U2388 ( .A1(n2489), .A2(n3937), .ZN(n2487) );
  OAI21_X1 U2389 ( .B1(n2480), .B2(n3570), .A(n2479), .ZN(n2478) );
  INV_X1 U2390 ( .A(n3567), .ZN(n2479) );
  NAND2_X1 U2391 ( .A1(n3744), .A2(n3745), .ZN(n2469) );
  NOR2_X1 U2392 ( .A1(n2412), .A2(n3033), .ZN(n2411) );
  INV_X1 U2393 ( .A(n2413), .ZN(n2412) );
  NAND2_X1 U2394 ( .A1(n2361), .A2(n2360), .ZN(n4342) );
  INV_X1 U2395 ( .A(n4361), .ZN(n2361) );
  NAND2_X1 U2396 ( .A1(n4187), .A2(n3304), .ZN(n2434) );
  OR2_X1 U2397 ( .A1(n3194), .A2(n3359), .ZN(n4070) );
  NOR2_X1 U2398 ( .A1(n2440), .A2(n2439), .ZN(n4823) );
  AND2_X1 U2399 ( .A1(n4835), .A2(n3396), .ZN(n2439) );
  NOR2_X1 U2400 ( .A1(n3388), .A2(n2441), .ZN(n2440) );
  AND2_X1 U2401 ( .A1(n4185), .A2(n3347), .ZN(n2441) );
  AOI21_X1 U2402 ( .B1(n2464), .B2(n2466), .A(n2308), .ZN(n2463) );
  INV_X1 U2403 ( .A(n2470), .ZN(n2464) );
  NAND2_X1 U2404 ( .A1(n3365), .A2(n2287), .ZN(n3190) );
  AND2_X1 U2405 ( .A1(n3365), .A2(n2281), .ZN(n3193) );
  OR2_X1 U2406 ( .A1(n4694), .A2(n4695), .ZN(n2405) );
  NAND2_X1 U2407 ( .A1(n4253), .A2(n2316), .ZN(n4257) );
  NAND2_X1 U2408 ( .A1(n4361), .A2(n2356), .ZN(n2351) );
  OAI21_X1 U2409 ( .B1(n4361), .B2(n2355), .A(n2352), .ZN(n4296) );
  AOI21_X1 U2410 ( .B1(n2354), .B2(n2353), .A(n4303), .ZN(n2352) );
  INV_X1 U2411 ( .A(n2356), .ZN(n2353) );
  NAND2_X1 U2412 ( .A1(n2417), .A2(n2419), .ZN(n4358) );
  NOR2_X1 U2413 ( .A1(n4263), .A2(n4264), .ZN(n4760) );
  OAI21_X1 U2414 ( .B1(n3837), .B2(n3483), .A(n2318), .ZN(n3424) );
  NAND2_X1 U2415 ( .A1(n2276), .A2(n3500), .ZN(n2318) );
  NAND2_X1 U2416 ( .A1(n2486), .A2(n2282), .ZN(n2485) );
  INV_X1 U2417 ( .A(n2487), .ZN(n2486) );
  NAND2_X1 U2418 ( .A1(n3746), .A2(n2471), .ZN(n2470) );
  INV_X1 U2419 ( .A(n3744), .ZN(n2471) );
  NOR2_X1 U2421 ( .A1(n2416), .A2(n3033), .ZN(n2409) );
  NOR2_X1 U2422 ( .A1(n2358), .A2(n4110), .ZN(n2356) );
  NAND2_X1 U2423 ( .A1(n4130), .A2(n4108), .ZN(n2357) );
  AND2_X1 U2424 ( .A1(n2381), .A2(n4099), .ZN(n2380) );
  INV_X1 U2425 ( .A(n4140), .ZN(n2371) );
  INV_X1 U2426 ( .A(n2304), .ZN(n2364) );
  NAND2_X1 U2427 ( .A1(n2433), .A2(n2432), .ZN(n2431) );
  NOR2_X1 U2428 ( .A1(n4150), .A2(n2428), .ZN(n2427) );
  INV_X1 U2429 ( .A(n2430), .ZN(n2428) );
  NAND2_X1 U2430 ( .A1(n3239), .A2(n3325), .ZN(n2430) );
  NAND2_X1 U2431 ( .A1(n3321), .A2(n2431), .ZN(n2429) );
  OR2_X1 U2432 ( .A1(n4188), .A2(n3256), .ZN(n4071) );
  NOR2_X1 U2433 ( .A1(n3832), .A2(n3839), .ZN(n2342) );
  NAND2_X1 U2434 ( .A1(n4456), .A2(n4415), .ZN(n2338) );
  AND2_X1 U2435 ( .A1(n4121), .A2(n2306), .ZN(n2437) );
  NAND2_X1 U2436 ( .A1(n2330), .A2(IR_REG_31__SCAN_IN), .ZN(n2607) );
  OR2_X1 U2437 ( .A1(n2611), .A2(IR_REG_22__SCAN_IN), .ZN(n2330) );
  AND4_X1 U2438 ( .A1(n2567), .A2(n2510), .A3(n2509), .A4(n2508), .ZN(n2511)
         );
  NOR2_X1 U2439 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2510)
         );
  NOR2_X1 U2440 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2509)
         );
  INV_X1 U2441 ( .A(IR_REG_13__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U2442 ( .A1(n2329), .A2(n2328), .ZN(n2327) );
  OAI22_X1 U2443 ( .A1(n3540), .A2(n3837), .B1(n2275), .B2(n3962), .ZN(n3466)
         );
  INV_X1 U2444 ( .A(n2469), .ZN(n2467) );
  NOR2_X1 U2445 ( .A1(n2488), .A2(n2489), .ZN(n3830) );
  OR2_X1 U2446 ( .A1(n3886), .A2(n3888), .ZN(n3895) );
  NAND2_X1 U2447 ( .A1(n3513), .A2(n2289), .ZN(n2477) );
  NOR2_X1 U2448 ( .A1(n3569), .A2(n2322), .ZN(n2321) );
  INV_X1 U2449 ( .A(n2480), .ZN(n2322) );
  NOR2_X1 U2450 ( .A1(n2478), .A2(n2476), .ZN(n2475) );
  INV_X1 U2451 ( .A(n3474), .ZN(n2476) );
  NAND2_X1 U2452 ( .A1(n2302), .A2(n2474), .ZN(n2473) );
  INV_X1 U2453 ( .A(n2478), .ZN(n2474) );
  XNOR2_X1 U2454 ( .A(n3207), .B(n3835), .ZN(n3211) );
  NAND2_X1 U2455 ( .A1(n2280), .A2(n4188), .ZN(n3206) );
  NAND2_X1 U2456 ( .A1(n2466), .A2(n3927), .ZN(n2462) );
  INV_X1 U2457 ( .A(n2460), .ZN(n2459) );
  OAI21_X1 U2458 ( .B1(n2463), .B2(n2461), .A(n2310), .ZN(n2460) );
  NAND2_X1 U2459 ( .A1(n3344), .A2(n2456), .ZN(n2455) );
  INV_X1 U2460 ( .A(n3307), .ZN(n2456) );
  AND2_X1 U2461 ( .A1(n2874), .A2(REG3_REG_0__SCAN_IN), .ZN(n2875) );
  NOR2_X1 U2462 ( .A1(n4648), .A2(n2626), .ZN(n2880) );
  XNOR2_X1 U2463 ( .A(n3143), .B(n3137), .ZN(n4207) );
  NOR2_X1 U2464 ( .A1(n3219), .A2(n2445), .ZN(n3284) );
  AND2_X1 U2465 ( .A1(n3220), .A2(n3144), .ZN(n2445) );
  NAND2_X1 U2466 ( .A1(n4664), .A2(n3274), .ZN(n3276) );
  OR2_X1 U2467 ( .A1(n2548), .A2(IR_REG_9__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U2468 ( .A1(n2447), .A2(n2446), .ZN(n3293) );
  OR2_X1 U2469 ( .A1(n3292), .A2(REG2_REG_7__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U2470 ( .A1(n4680), .A2(n2448), .ZN(n2447) );
  NAND2_X1 U2471 ( .A1(n3292), .A2(REG2_REG_7__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U2472 ( .A1(n2405), .A2(n2293), .ZN(n2404) );
  XNOR2_X1 U2473 ( .A(n3595), .B(n4865), .ZN(n4706) );
  NAND2_X1 U2474 ( .A1(n2402), .A2(n2401), .ZN(n3612) );
  NAND2_X1 U2475 ( .A1(n2404), .A2(REG1_REG_9__SCAN_IN), .ZN(n2401) );
  OAI21_X1 U2476 ( .B1(n2404), .B2(REG1_REG_9__SCAN_IN), .A(n2403), .ZN(n2402)
         );
  OAI21_X1 U2477 ( .B1(n4714), .B2(n2305), .A(n3615), .ZN(n3617) );
  OR2_X1 U2478 ( .A1(n4712), .A2(REG1_REG_11__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U2479 ( .A1(n4718), .A2(n3597), .ZN(n3598) );
  NAND2_X1 U2480 ( .A1(n2393), .A2(n2392), .ZN(n4235) );
  NAND2_X1 U2481 ( .A1(n4223), .A2(REG1_REG_15__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U2482 ( .A1(n4231), .A2(n2394), .ZN(n2393) );
  INV_X1 U2483 ( .A(n4233), .ZN(n2394) );
  AOI21_X1 U2484 ( .B1(n2416), .B2(n2414), .A(n2300), .ZN(n2413) );
  INV_X1 U2485 ( .A(n2418), .ZN(n2414) );
  AND2_X1 U2486 ( .A1(n3016), .A2(n3015), .ZN(n3027) );
  INV_X1 U2487 ( .A(n4405), .ZN(n4362) );
  OAI21_X1 U2488 ( .B1(n3629), .B2(n2375), .A(n2298), .ZN(n3070) );
  INV_X1 U2489 ( .A(n2376), .ZN(n2375) );
  NOR2_X1 U2490 ( .A1(n4547), .A2(n4444), .ZN(n2982) );
  NAND2_X1 U2491 ( .A1(n4032), .A2(n3059), .ZN(n2372) );
  AND4_X1 U2492 ( .A1(n2920), .A2(n2919), .A3(n2918), .A4(n2917), .ZN(n3652)
         );
  NAND2_X1 U2493 ( .A1(n3054), .A2(n4052), .ZN(n3451) );
  NAND2_X1 U2494 ( .A1(n4849), .A2(n2905), .ZN(n3491) );
  NAND2_X1 U2495 ( .A1(n2391), .A2(n4081), .ZN(n4831) );
  NAND2_X1 U2496 ( .A1(n3389), .A2(n4079), .ZN(n2391) );
  AND2_X1 U2497 ( .A1(n4916), .A2(n3121), .ZN(n4838) );
  AOI21_X1 U2498 ( .B1(n4128), .B2(n3354), .A(n2878), .ZN(n3253) );
  NAND2_X1 U2499 ( .A1(n2525), .A2(n2522), .ZN(n2523) );
  OR2_X1 U2500 ( .A1(n2584), .A2(n4270), .ZN(n4509) );
  INV_X1 U2501 ( .A(n3092), .ZN(n2583) );
  AND2_X1 U2502 ( .A1(n2589), .A2(n4649), .ZN(n3116) );
  INV_X1 U2503 ( .A(IR_REG_28__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U2504 ( .A1(n2513), .A2(n2490), .ZN(n2632) );
  NAND2_X1 U2505 ( .A1(n2514), .A2(n2493), .ZN(n2492) );
  NAND2_X1 U2506 ( .A1(n2457), .A2(n3408), .ZN(n2332) );
  NAND2_X1 U2507 ( .A1(n3410), .A2(n3409), .ZN(n2331) );
  INV_X1 U2508 ( .A(n3483), .ZN(n4837) );
  AND2_X1 U2509 ( .A1(n3132), .A2(n3131), .ZN(n3146) );
  XNOR2_X1 U2510 ( .A(n3284), .B(n4655), .ZN(n3221) );
  XNOR2_X1 U2511 ( .A(n3276), .B(n3275), .ZN(n4675) );
  NAND2_X1 U2512 ( .A1(n4675), .A2(REG1_REG_6__SCAN_IN), .ZN(n4674) );
  XNOR2_X1 U2513 ( .A(n3293), .B(n4856), .ZN(n4699) );
  NAND2_X1 U2514 ( .A1(n3297), .A2(n3296), .ZN(n3593) );
  XNOR2_X1 U2515 ( .A(n3598), .B(n4892), .ZN(n4730) );
  NAND2_X1 U2516 ( .A1(n4730), .A2(REG2_REG_12__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U2517 ( .A1(n3620), .A2(REG1_REG_14__SCAN_IN), .ZN(n4226) );
  AOI21_X1 U2518 ( .B1(n4257), .B2(n4256), .A(n4771), .ZN(n4262) );
  INV_X1 U2519 ( .A(n4729), .ZN(n4771) );
  NAND2_X1 U2520 ( .A1(n4759), .A2(REG2_REG_18__SCAN_IN), .ZN(n2442) );
  XNOR2_X1 U2521 ( .A(n2398), .B(n4762), .ZN(n2397) );
  NAND2_X1 U2522 ( .A1(n2400), .A2(n2399), .ZN(n2398) );
  NAND2_X1 U2523 ( .A1(n4759), .A2(REG1_REG_18__SCAN_IN), .ZN(n2399) );
  AND2_X1 U2524 ( .A1(n3146), .A2(n4168), .ZN(n4769) );
  NAND2_X1 U2525 ( .A1(n4279), .A2(n2348), .ZN(n2347) );
  OR2_X1 U2526 ( .A1(n4433), .A2(n4280), .ZN(n2348) );
  INV_X1 U2527 ( .A(n4462), .ZN(n4826) );
  OAI21_X1 U2528 ( .B1(n4284), .B2(n4280), .A(n3092), .ZN(n4276) );
  INV_X1 U2529 ( .A(n2529), .ZN(n2350) );
  INV_X1 U2530 ( .A(n3527), .ZN(n2481) );
  OAI22_X1 U2531 ( .A1(n4362), .A2(n3837), .B1(n4395), .B2(n2275), .ZN(n3814)
         );
  AND2_X1 U2532 ( .A1(n3475), .A2(n3476), .ZN(n3474) );
  INV_X1 U2533 ( .A(n3927), .ZN(n2461) );
  INV_X1 U2534 ( .A(n3174), .ZN(n3176) );
  AND3_X1 U2535 ( .A1(n3158), .A2(n3157), .A3(n3156), .ZN(n3174) );
  OR2_X1 U2536 ( .A1(n4299), .A2(n4288), .ZN(n4019) );
  AND2_X1 U2537 ( .A1(n2424), .A2(n2423), .ZN(n2418) );
  NAND2_X1 U2538 ( .A1(n2376), .A2(n2374), .ZN(n2373) );
  INV_X1 U2539 ( .A(n2379), .ZN(n2374) );
  NOR2_X1 U2540 ( .A1(n4103), .A2(n2377), .ZN(n2376) );
  INV_X1 U2541 ( .A(n4100), .ZN(n2377) );
  AND2_X1 U2542 ( .A1(n2380), .A2(n4123), .ZN(n2379) );
  NOR2_X1 U2543 ( .A1(n3751), .A2(n3586), .ZN(n2345) );
  INV_X1 U2544 ( .A(n4566), .ZN(n3769) );
  NAND2_X1 U2545 ( .A1(n3691), .A2(n2343), .ZN(n3625) );
  NOR2_X1 U2546 ( .A1(n2344), .A2(n3757), .ZN(n2343) );
  INV_X1 U2547 ( .A(n2345), .ZN(n2344) );
  AND2_X1 U2548 ( .A1(n4832), .A2(n3396), .ZN(n2341) );
  INV_X1 U2549 ( .A(n3364), .ZN(n3166) );
  OR2_X1 U2550 ( .A1(n2551), .A2(IR_REG_10__SCAN_IN), .ZN(n2552) );
  INV_X1 U2551 ( .A(IR_REG_6__SCAN_IN), .ZN(n2543) );
  AOI21_X1 U2552 ( .B1(n2455), .B2(n2315), .A(n3409), .ZN(n2452) );
  NAND2_X1 U2553 ( .A1(n3945), .A2(n2315), .ZN(n2453) );
  OR2_X1 U2554 ( .A1(n2990), .A2(n3983), .ZN(n2996) );
  OAI21_X1 U2555 ( .B1(n2279), .B2(n3652), .A(n2319), .ZN(n3467) );
  NAND2_X1 U2556 ( .A1(n2276), .A2(n2320), .ZN(n2319) );
  OAI21_X1 U2557 ( .B1(n3837), .B2(n3239), .A(n2317), .ZN(n3240) );
  NAND2_X1 U2558 ( .A1(n2277), .A2(n2432), .ZN(n2317) );
  OAI22_X1 U2559 ( .A1(n3494), .A2(n3837), .B1(n4832), .B2(n2275), .ZN(n3412)
         );
  OR2_X1 U2560 ( .A1(n2984), .A2(n2805), .ZN(n2990) );
  NAND2_X1 U2561 ( .A1(n2481), .A2(n2313), .ZN(n2480) );
  OAI22_X1 U2562 ( .A1(n3666), .A2(n3837), .B1(n3635), .B2(n2275), .ZN(n3529)
         );
  AOI21_X1 U2563 ( .B1(n2299), .B2(n2485), .A(n2283), .ZN(n2482) );
  NOR2_X1 U2564 ( .A1(n2485), .A2(n3830), .ZN(n2484) );
  NOR2_X1 U2565 ( .A1(n2945), .A2(n3921), .ZN(n2954) );
  OR2_X1 U2566 ( .A1(n2928), .A2(n3531), .ZN(n2930) );
  OR2_X1 U2567 ( .A1(n2930), .A2(n3579), .ZN(n2937) );
  NAND2_X1 U2568 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  INV_X1 U2569 ( .A(n3509), .ZN(n3511) );
  OAI22_X1 U2570 ( .A1(n4835), .A2(n3837), .B1(n3396), .B2(n2275), .ZN(n3346)
         );
  NAND2_X1 U2571 ( .A1(n2326), .A2(n2324), .ZN(n2329) );
  AND2_X1 U2572 ( .A1(n2482), .A2(n2325), .ZN(n2324) );
  INV_X1 U2573 ( .A(n3906), .ZN(n2325) );
  NOR2_X1 U2574 ( .A1(n2937), .A2(n2936), .ZN(n2943) );
  NAND2_X1 U2575 ( .A1(n2943), .A2(REG3_REG_15__SCAN_IN), .ZN(n2945) );
  AND2_X1 U2576 ( .A1(n3753), .A2(n3752), .ZN(n4904) );
  NAND2_X1 U2577 ( .A1(n3747), .A2(n2470), .ZN(n2468) );
  AND4_X1 U2578 ( .A1(n2857), .A2(n2856), .A3(n2855), .A4(n2854), .ZN(n3540)
         );
  NAND2_X1 U2579 ( .A1(n3141), .A2(n4191), .ZN(n4204) );
  NAND2_X1 U2580 ( .A1(n4205), .A2(n4204), .ZN(n4203) );
  AOI22_X1 U2581 ( .A1(n3140), .A2(n4206), .B1(REG1_REG_2__SCAN_IN), .B2(n2527), .ZN(n3223) );
  AOI21_X1 U2582 ( .B1(REG2_REG_5__SCAN_IN), .B2(n3288), .A(n4659), .ZN(n3290)
         );
  INV_X1 U2583 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U2584 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  NAND2_X1 U2585 ( .A1(n4760), .A2(n4761), .ZN(n2400) );
  XNOR2_X1 U2586 ( .A(n4290), .B(n2386), .ZN(n2385) );
  INV_X1 U2587 ( .A(n4289), .ZN(n2386) );
  NAND2_X1 U2588 ( .A1(n2410), .A2(n2407), .ZN(n4282) );
  AOI21_X1 U2589 ( .B1(n2409), .B2(n2413), .A(n2408), .ZN(n2407) );
  NOR2_X1 U2590 ( .A1(n4011), .A2(n4517), .ZN(n2408) );
  NAND2_X1 U2591 ( .A1(n4342), .A2(n4108), .ZN(n4320) );
  NAND2_X1 U2592 ( .A1(n2378), .A2(n4100), .ZN(n4423) );
  NAND2_X1 U2593 ( .A1(n3629), .A2(n2379), .ZN(n2378) );
  NAND2_X1 U2594 ( .A1(n3629), .A2(n2380), .ZN(n4440) );
  AOI21_X1 U2595 ( .B1(n3699), .B2(n2961), .A(n2960), .ZN(n4500) );
  NAND2_X1 U2596 ( .A1(n3629), .A2(n4099), .ZN(n4468) );
  OAI21_X1 U2597 ( .B1(n4032), .B2(n2370), .A(n2367), .ZN(n3631) );
  AOI21_X1 U2598 ( .B1(n2369), .B2(n4139), .A(n2368), .ZN(n2367) );
  INV_X1 U2599 ( .A(n4029), .ZN(n2368) );
  NAND2_X1 U2600 ( .A1(n3631), .A2(n3630), .ZN(n3629) );
  INV_X1 U2601 ( .A(n4571), .ZN(n3757) );
  NAND2_X1 U2602 ( .A1(n3691), .A2(n2345), .ZN(n3723) );
  AOI21_X1 U2603 ( .B1(n2437), .B2(n2285), .A(n2307), .ZN(n2436) );
  NAND2_X1 U2604 ( .A1(n2921), .A2(REG3_REG_11__SCAN_IN), .ZN(n2928) );
  NAND2_X1 U2605 ( .A1(n3055), .A2(n4057), .ZN(n3649) );
  NAND2_X1 U2606 ( .A1(n3538), .A2(n4060), .ZN(n3055) );
  OAI21_X1 U2607 ( .B1(n3451), .B2(n4084), .A(n4086), .ZN(n3538) );
  NOR2_X1 U2608 ( .A1(n2908), .A2(n2852), .ZN(n2915) );
  OAI21_X1 U2609 ( .B1(n4831), .B2(n3053), .A(n4053), .ZN(n3492) );
  INV_X1 U2610 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3431) );
  NOR2_X1 U2611 ( .A1(n2364), .A2(n2363), .ZN(n2362) );
  INV_X1 U2612 ( .A(n4078), .ZN(n2363) );
  NAND2_X1 U2613 ( .A1(n2893), .A2(REG3_REG_5__SCAN_IN), .ZN(n2892) );
  INV_X1 U2614 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3349) );
  NOR2_X1 U2615 ( .A1(n2892), .A2(n3349), .ZN(n2899) );
  OAI21_X1 U2616 ( .B1(n2427), .B2(n2426), .A(n2425), .ZN(n3337) );
  INV_X1 U2617 ( .A(n2434), .ZN(n2426) );
  NAND2_X1 U2618 ( .A1(n3321), .A2(n2295), .ZN(n2425) );
  NAND2_X1 U2619 ( .A1(n2429), .A2(n2430), .ZN(n3378) );
  NAND2_X1 U2620 ( .A1(n4071), .A2(n4074), .ZN(n4120) );
  INV_X1 U2621 ( .A(n4128), .ZN(n3356) );
  NOR2_X1 U2622 ( .A1(n3092), .A2(n4047), .ZN(n4270) );
  NAND2_X1 U2623 ( .A1(n4367), .A2(n2314), .ZN(n4306) );
  NAND2_X1 U2624 ( .A1(n4367), .A2(n2342), .ZN(n4328) );
  NAND2_X1 U2625 ( .A1(n4548), .A2(n4395), .ZN(n2337) );
  NOR2_X1 U2626 ( .A1(n4394), .A2(n3823), .ZN(n4367) );
  NOR2_X1 U2627 ( .A1(n4479), .A2(n4444), .ZN(n4454) );
  OR2_X1 U2628 ( .A1(n4478), .A2(n3783), .ZN(n4479) );
  NOR2_X1 U2629 ( .A1(n3625), .A2(n3769), .ZN(n4489) );
  NAND2_X1 U2630 ( .A1(n3691), .A2(n4583), .ZN(n3725) );
  INV_X1 U2631 ( .A(n3574), .ZN(n3677) );
  AND2_X1 U2632 ( .A1(n3678), .A2(n3677), .ZN(n3691) );
  NOR2_X1 U2633 ( .A1(n3645), .A2(n3556), .ZN(n3678) );
  INV_X1 U2634 ( .A(n3556), .ZN(n3635) );
  NAND2_X1 U2635 ( .A1(n2438), .A2(n2437), .ZN(n3647) );
  AND2_X1 U2636 ( .A1(n2438), .A2(n2306), .ZN(n3648) );
  OR2_X1 U2637 ( .A1(n3537), .A2(n2285), .ZN(n2438) );
  OR2_X1 U2638 ( .A1(n3644), .A2(n3514), .ZN(n3645) );
  NAND2_X1 U2639 ( .A1(n3536), .A2(n3539), .ZN(n3644) );
  AND2_X1 U2640 ( .A1(n3502), .A2(n3962), .ZN(n3536) );
  AND2_X1 U2641 ( .A1(n3397), .A2(n2340), .ZN(n3502) );
  AND2_X1 U2642 ( .A1(n2341), .A2(n3493), .ZN(n2340) );
  NAND2_X1 U2643 ( .A1(n3397), .A2(n2341), .ZN(n4821) );
  NAND2_X1 U2644 ( .A1(n4823), .A2(n4830), .ZN(n4849) );
  INV_X1 U2645 ( .A(n3347), .ZN(n3396) );
  NAND2_X1 U2646 ( .A1(n3397), .A2(n3396), .ZN(n4820) );
  OR2_X1 U2647 ( .A1(n3332), .A2(n3304), .ZN(n3373) );
  NOR2_X1 U2648 ( .A1(n3373), .A2(n3438), .ZN(n3397) );
  NOR2_X1 U2649 ( .A1(n3366), .A2(n3737), .ZN(n3331) );
  INV_X1 U2650 ( .A(n4406), .ZN(n4834) );
  NAND2_X1 U2651 ( .A1(n2301), .A2(n2528), .ZN(n3256) );
  NAND2_X1 U2652 ( .A1(n2525), .A2(n2786), .ZN(n2528) );
  AND3_X1 U2653 ( .A1(n3088), .A2(n3087), .A3(n3086), .ZN(n3096) );
  INV_X1 U2654 ( .A(IR_REG_7__SCAN_IN), .ZN(n2544) );
  NOR2_X1 U2655 ( .A1(n2519), .A2(n3113), .ZN(n2406) );
  NAND2_X1 U2656 ( .A1(n2521), .A2(n2520), .ZN(n4194) );
  AOI21_X1 U2657 ( .B1(n3867), .B2(n3868), .A(n4016), .ZN(n3870) );
  NOR2_X1 U2658 ( .A1(n3992), .A2(n3780), .ZN(n3782) );
  NOR2_X1 U2659 ( .A1(n3855), .A2(n3186), .ZN(n3187) );
  INV_X1 U2660 ( .A(n3185), .ZN(n3186) );
  NAND2_X1 U2661 ( .A1(n2477), .A2(n2480), .ZN(n3568) );
  NOR2_X1 U2662 ( .A1(n3945), .A2(n3307), .ZN(n3345) );
  OAI21_X1 U2663 ( .B1(n3747), .B2(n2465), .A(n2463), .ZN(n3929) );
  AOI21_X1 U2664 ( .B1(n3879), .B2(n3828), .A(n3829), .ZN(n3936) );
  INV_X1 U2665 ( .A(n4370), .ZN(n3942) );
  NAND2_X1 U2666 ( .A1(n2477), .A2(n2321), .ZN(n2323) );
  NAND2_X1 U2667 ( .A1(n3513), .A2(n3512), .ZN(n3528) );
  OAI21_X1 U2668 ( .B1(n3945), .B2(n2455), .A(n2315), .ZN(n2454) );
  INV_X1 U2669 ( .A(n4897), .ZN(n3994) );
  INV_X1 U2670 ( .A(n4896), .ZN(n3995) );
  INV_X1 U2671 ( .A(n4912), .ZN(n4014) );
  OR2_X1 U2672 ( .A1(n3195), .A2(n4916), .ZN(n4896) );
  NAND4_X1 U2673 ( .A1(n3032), .A2(n3031), .A3(n3030), .A4(n3029), .ZN(n4324)
         );
  NAND4_X1 U2674 ( .A1(n3021), .A2(n3020), .A3(n3019), .A4(n3018), .ZN(n4347)
         );
  NAND4_X1 U2675 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .ZN(n4405)
         );
  NAND4_X1 U2676 ( .A1(n2995), .A2(n2994), .A3(n2993), .A4(n2992), .ZN(n4425)
         );
  NAND4_X1 U2677 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n4547)
         );
  INV_X1 U2678 ( .A(n3666), .ZN(n4180) );
  INV_X1 U2679 ( .A(n3540), .ZN(n4183) );
  NAND4_X1 U2680 ( .A1(n2904), .A2(n2903), .A3(n2902), .A4(n2901), .ZN(n4184)
         );
  NAND2_X1 U2681 ( .A1(n2881), .A2(REG1_REG_1__SCAN_IN), .ZN(n2868) );
  NOR2_X1 U2682 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  XNOR2_X1 U2683 ( .A(n4194), .B(REG2_REG_1__SCAN_IN), .ZN(n4193) );
  NAND2_X1 U2684 ( .A1(n4193), .A2(n4192), .ZN(n4191) );
  NOR2_X1 U2685 ( .A1(n3285), .A2(n2444), .ZN(n4661) );
  NOR2_X1 U2686 ( .A1(n3286), .A2(n3270), .ZN(n2444) );
  NAND2_X1 U2687 ( .A1(n4674), .A2(n3277), .ZN(n4689) );
  NAND2_X1 U2688 ( .A1(n2395), .A2(n4690), .ZN(n4688) );
  OR2_X1 U2689 ( .A1(n4689), .A2(n2396), .ZN(n2395) );
  AND2_X1 U2690 ( .A1(n3292), .A2(REG1_REG_7__SCAN_IN), .ZN(n2396) );
  INV_X1 U2691 ( .A(n4680), .ZN(n4679) );
  INV_X1 U2692 ( .A(n2405), .ZN(n4693) );
  NAND2_X1 U2693 ( .A1(n4698), .A2(n3294), .ZN(n3297) );
  INV_X1 U2694 ( .A(n2404), .ZN(n3610) );
  NAND2_X1 U2695 ( .A1(n4703), .A2(n3614), .ZN(n4714) );
  XNOR2_X1 U2696 ( .A(n3617), .B(n4892), .ZN(n4724) );
  AND2_X1 U2697 ( .A1(n3146), .A2(n3145), .ZN(n4729) );
  NAND2_X1 U2698 ( .A1(n4728), .A2(n3599), .ZN(n4736) );
  NAND2_X1 U2699 ( .A1(n4226), .A2(n4227), .ZN(n4231) );
  AND2_X1 U2700 ( .A1(n2384), .A2(n2382), .ZN(n4515) );
  NOR2_X1 U2701 ( .A1(n4291), .A2(n2383), .ZN(n2382) );
  NAND2_X1 U2702 ( .A1(n2385), .A2(n4449), .ZN(n2384) );
  AND2_X1 U2703 ( .A1(n4292), .A2(n4838), .ZN(n2383) );
  OAI21_X1 U2704 ( .B1(n4420), .B2(n2415), .A(n2413), .ZN(n4304) );
  NAND2_X1 U2705 ( .A1(n2351), .A2(n2354), .ZN(n4298) );
  AND2_X1 U2706 ( .A1(n3034), .A2(n3028), .ZN(n4302) );
  XNOR2_X1 U2707 ( .A(n4318), .B(n4317), .ZN(n4528) );
  NAND2_X1 U2708 ( .A1(n4316), .A2(n4315), .ZN(n4318) );
  NAND2_X1 U2709 ( .A1(n2372), .A2(n2369), .ZN(n3729) );
  NAND2_X1 U2710 ( .A1(n2372), .A2(n4027), .ZN(n3728) );
  AND4_X1 U2711 ( .A1(n2912), .A2(n2911), .A3(n2910), .A4(n2909), .ZN(n3483)
         );
  INV_X1 U2712 ( .A(n4122), .ZN(n2365) );
  NAND2_X1 U2713 ( .A1(n3051), .A2(n4078), .ZN(n2366) );
  INV_X1 U2714 ( .A(n4883), .ZN(n4870) );
  AOI211_X1 U2715 ( .C1(n4406), .C2(n4299), .A(n3081), .B(n4278), .ZN(n3082)
         );
  OAI211_X1 U2716 ( .C1(n4516), .C2(n4845), .A(n4515), .B(n4514), .ZN(n4602)
         );
  NAND2_X1 U2717 ( .A1(n3117), .A2(n3159), .ZN(n4658) );
  AND2_X1 U2718 ( .A1(n2621), .A2(n2389), .ZN(n2388) );
  XNOR2_X1 U2719 ( .A(n2588), .B(IR_REG_26__SCAN_IN), .ZN(n4649) );
  XNOR2_X1 U2720 ( .A(n2586), .B(IR_REG_25__SCAN_IN), .ZN(n3106) );
  XNOR2_X1 U2721 ( .A(n2585), .B(IR_REG_24__SCAN_IN), .ZN(n4650) );
  INV_X1 U2722 ( .A(n2618), .ZN(n4651) );
  INV_X1 U2723 ( .A(n3292), .ZN(n4817) );
  AOI21_X1 U2724 ( .B1(n2443), .B2(n4262), .A(n4261), .ZN(n4267) );
  AOI21_X1 U2725 ( .B1(n2397), .B2(n4769), .A(n4768), .ZN(n4770) );
  OR2_X1 U2726 ( .A1(n2643), .A2(n2642), .ZN(n2841) );
  NAND2_X1 U2727 ( .A1(n2349), .A2(n2346), .ZN(U3354) );
  OAI21_X1 U2728 ( .B1(n4277), .B2(n4278), .A(n4826), .ZN(n2349) );
  AOI21_X1 U2729 ( .B1(n4281), .B2(n4305), .A(n2347), .ZN(n2346) );
  OR2_X1 U2730 ( .A1(n3937), .A2(n2488), .ZN(n2282) );
  NAND2_X1 U2731 ( .A1(n3979), .A2(n3819), .ZN(n3879) );
  NAND2_X1 U2732 ( .A1(n2558), .A2(n2296), .ZN(n2611) );
  AND2_X1 U2733 ( .A1(n2483), .A2(n3830), .ZN(n2283) );
  AND2_X1 U2734 ( .A1(n3500), .A2(n4837), .ZN(n2284) );
  AND2_X1 U2735 ( .A1(n3539), .A2(n3652), .ZN(n2285) );
  NAND2_X1 U2736 ( .A1(n4489), .A2(n4490), .ZN(n4478) );
  INV_X1 U2737 ( .A(n2336), .ZN(n4393) );
  INV_X1 U2738 ( .A(n3611), .ZN(n2403) );
  NOR3_X1 U2739 ( .A1(n4479), .A2(n3800), .A3(n4444), .ZN(n4414) );
  INV_X1 U2740 ( .A(n4395), .ZN(n4388) );
  NAND2_X1 U2741 ( .A1(n2468), .A2(n2469), .ZN(n3915) );
  CLKBUF_X3 U2742 ( .A(n2880), .Z(n2887) );
  AND2_X1 U2743 ( .A1(n2873), .A2(n2872), .ZN(n2286) );
  INV_X1 U2744 ( .A(n3819), .ZN(n2483) );
  OAI22_X1 U2745 ( .A1(n2333), .A2(n3782), .B1(n3781), .B2(n3991), .ZN(n3886)
         );
  AND2_X1 U2746 ( .A1(n4347), .A2(n4524), .ZN(n4110) );
  INV_X1 U2747 ( .A(n4110), .ZN(n2359) );
  OAI21_X1 U2748 ( .B1(n2271), .B2(n2524), .A(n2523), .ZN(n3359) );
  AND2_X1 U2749 ( .A1(n2472), .A2(n2473), .ZN(n2288) );
  XNOR2_X1 U2750 ( .A(n2625), .B(n2389), .ZN(n2842) );
  AND2_X1 U2751 ( .A1(n2481), .A2(n3512), .ZN(n2289) );
  AND3_X1 U2752 ( .A1(n2884), .A2(n2883), .A3(n2882), .ZN(n2290) );
  NOR2_X1 U2753 ( .A1(n4648), .A2(n2842), .ZN(n2881) );
  AND2_X1 U2754 ( .A1(n4648), .A2(n2626), .ZN(n2874) );
  INV_X1 U2755 ( .A(n4108), .ZN(n2358) );
  INV_X1 U2756 ( .A(IR_REG_2__SCAN_IN), .ZN(n2526) );
  INV_X1 U2757 ( .A(n3828), .ZN(n2488) );
  AND2_X1 U2758 ( .A1(n3879), .A2(n3830), .ZN(n2291) );
  INV_X1 U2759 ( .A(n2513), .ZN(n2613) );
  OR2_X1 U2760 ( .A1(n2611), .A2(n2492), .ZN(n2292) );
  OR2_X1 U2761 ( .A1(n4702), .A2(n4688), .ZN(n2293) );
  INV_X1 U2762 ( .A(n2416), .ZN(n2415) );
  AND2_X1 U2763 ( .A1(n3209), .A2(n4188), .ZN(n2294) );
  AND2_X1 U2764 ( .A1(n2431), .A2(n2434), .ZN(n2295) );
  AND2_X1 U2765 ( .A1(n2511), .A2(n2512), .ZN(n2296) );
  INV_X1 U2766 ( .A(n3003), .ZN(n2423) );
  INV_X1 U2767 ( .A(n4130), .ZN(n2360) );
  AND2_X1 U2768 ( .A1(n2357), .A2(n4112), .ZN(n2297) );
  INV_X1 U2769 ( .A(n2420), .ZN(n2419) );
  NOR2_X1 U2770 ( .A1(n2421), .A2(n3003), .ZN(n2420) );
  AND4_X1 U2771 ( .A1(n2891), .A2(n2890), .A3(n2889), .A4(n2888), .ZN(n3239)
         );
  INV_X1 U2772 ( .A(n3239), .ZN(n2433) );
  INV_X1 U2773 ( .A(n2355), .ZN(n2354) );
  NOR2_X1 U2774 ( .A1(n2297), .A2(n4110), .ZN(n2355) );
  AND2_X1 U2775 ( .A1(n4037), .A2(n2373), .ZN(n2298) );
  OR2_X1 U2776 ( .A1(n2487), .A2(n2483), .ZN(n2299) );
  OR2_X1 U2777 ( .A1(n2499), .A2(n2498), .ZN(n2300) );
  INV_X1 U2778 ( .A(IR_REG_21__SCAN_IN), .ZN(n2512) );
  INV_X1 U2779 ( .A(n4303), .ZN(n4297) );
  OR2_X1 U2780 ( .A1(n2525), .A2(n2527), .ZN(n2301) );
  NAND2_X1 U2781 ( .A1(n2289), .A2(n3569), .ZN(n2302) );
  OR2_X1 U2782 ( .A1(n3163), .A2(n3167), .ZN(n2303) );
  AOI22_X1 U2784 ( .A1(n4185), .A2(n3854), .B1(n2273), .B2(n3347), .ZN(n3406)
         );
  INV_X1 U2785 ( .A(IR_REG_29__SCAN_IN), .ZN(n2389) );
  INV_X1 U2786 ( .A(n3539), .ZN(n2320) );
  NAND2_X1 U2787 ( .A1(n4186), .A2(n3338), .ZN(n2304) );
  AND2_X1 U2788 ( .A1(n4712), .A2(REG1_REG_11__SCAN_IN), .ZN(n2305) );
  OR2_X1 U2789 ( .A1(n2558), .A2(n3113), .ZN(n2562) );
  INV_X1 U2790 ( .A(IR_REG_22__SCAN_IN), .ZN(n2493) );
  MUX2_X1 U2791 ( .A(n4224), .B(n2560), .S(n2271), .Z(n4583) );
  NAND2_X1 U2792 ( .A1(n2320), .A2(n4182), .ZN(n2306) );
  AND2_X1 U2793 ( .A1(n3651), .A2(n2927), .ZN(n2307) );
  NOR3_X1 U2794 ( .A1(n4479), .A2(n2338), .A3(n2337), .ZN(n2339) );
  NOR3_X1 U2795 ( .A1(n4479), .A2(n2338), .A3(n3800), .ZN(n2336) );
  INV_X1 U2796 ( .A(n2370), .ZN(n2369) );
  NAND2_X1 U2797 ( .A1(n2371), .A2(n4027), .ZN(n2370) );
  INV_X1 U2798 ( .A(n2466), .ZN(n2465) );
  NOR2_X1 U2799 ( .A1(n3765), .A2(n2467), .ZN(n2466) );
  NAND2_X1 U2800 ( .A1(n3764), .A2(n3913), .ZN(n2308) );
  NAND2_X1 U2801 ( .A1(n4367), .A2(n4350), .ZN(n4327) );
  INV_X1 U2802 ( .A(n3493), .ZN(n3500) );
  AND2_X1 U2803 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2309)
         );
  NAND2_X1 U2804 ( .A1(n2617), .A2(n4879), .ZN(n4889) );
  OR2_X1 U2805 ( .A1(n3773), .A2(n3772), .ZN(n2310) );
  NOR2_X1 U2806 ( .A1(n2458), .A2(n3948), .ZN(n3945) );
  INV_X1 U2807 ( .A(n4456), .ZN(n4444) );
  NAND2_X1 U2808 ( .A1(n2525), .A2(DATAI_21_), .ZN(n4548) );
  AND2_X1 U2809 ( .A1(n2429), .A2(n2427), .ZN(n2311) );
  NOR2_X1 U2810 ( .A1(n2451), .A2(n2534), .ZN(n2312) );
  NAND4_X1 U2811 ( .A1(n2871), .A2(n2870), .A3(n2869), .A4(n2868), .ZN(n3194)
         );
  INV_X1 U2812 ( .A(n4840), .ZN(n4449) );
  MUX2_X1 U2813 ( .A(n3222), .B(n2530), .S(n2271), .Z(n3325) );
  INV_X1 U2814 ( .A(n3325), .ZN(n2432) );
  XNOR2_X1 U2815 ( .A(n3201), .B(n3202), .ZN(n3204) );
  NAND2_X1 U2816 ( .A1(n2334), .A2(IR_REG_31__SCAN_IN), .ZN(n2630) );
  OAI22_X1 U2817 ( .A1(n3204), .A2(n3203), .B1(n3202), .B2(n3201), .ZN(n3212)
         );
  AND2_X1 U2818 ( .A1(n3520), .A2(n3519), .ZN(n2313) );
  AND2_X1 U2819 ( .A1(n2342), .A2(n4517), .ZN(n2314) );
  NAND2_X1 U2820 ( .A1(n3312), .A2(n3311), .ZN(n2315) );
  OR2_X1 U2821 ( .A1(n4653), .A2(REG2_REG_17__SCAN_IN), .ZN(n2316) );
  INV_X1 U2822 ( .A(IR_REG_4__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2823 ( .A1(n2326), .A2(n2482), .ZN(n3904) );
  OR2_X2 U2824 ( .A1(n3979), .A2(n2484), .ZN(n2326) );
  INV_X1 U2825 ( .A(n2329), .ZN(n4003) );
  OAI21_X1 U2826 ( .B1(n4004), .B2(n2327), .A(n4005), .ZN(n3867) );
  INV_X1 U2827 ( .A(n4007), .ZN(n2328) );
  AND2_X2 U2828 ( .A1(n2558), .A2(n2511), .ZN(n2513) );
  INV_X1 U2829 ( .A(n2333), .ZN(n3990) );
  NAND3_X1 U2830 ( .A1(n2513), .A2(n2335), .A3(n2490), .ZN(n2334) );
  INV_X1 U2831 ( .A(n2339), .ZN(n4394) );
  NAND2_X1 U2832 ( .A1(n2350), .A2(n2496), .ZN(n2534) );
  AND3_X2 U2833 ( .A1(n2449), .A2(n2450), .A3(n2350), .ZN(n2558) );
  NAND2_X1 U2834 ( .A1(n3051), .A2(n2362), .ZN(n3052) );
  XNOR2_X1 U2835 ( .A(n2366), .B(n2365), .ZN(n3339) );
  INV_X1 U2836 ( .A(n4035), .ZN(n2381) );
  NAND2_X1 U2837 ( .A1(n2281), .A2(n3194), .ZN(n3191) );
  AND2_X1 U2838 ( .A1(n2490), .A2(n2388), .ZN(n2387) );
  NAND2_X1 U2839 ( .A1(n2387), .A2(n2513), .ZN(n2390) );
  NAND3_X1 U2840 ( .A1(n2513), .A2(n2490), .A3(n2621), .ZN(n2624) );
  NAND2_X1 U2841 ( .A1(n4296), .A2(n4018), .ZN(n4290) );
  NAND2_X1 U2842 ( .A1(n4420), .A2(n2411), .ZN(n2410) );
  NAND2_X1 U2843 ( .A1(n4420), .A2(n2418), .ZN(n2417) );
  AND2_X1 U2844 ( .A1(n4403), .A2(n4377), .ZN(n2424) );
  NAND2_X1 U2845 ( .A1(n3537), .A2(n2437), .ZN(n2435) );
  NAND2_X1 U2846 ( .A1(n2435), .A2(n2436), .ZN(n3551) );
  NAND4_X1 U2847 ( .A1(n2503), .A2(n2506), .A3(n2504), .A4(n2505), .ZN(n2451)
         );
  INV_X1 U2848 ( .A(n2454), .ZN(n3410) );
  OR2_X1 U2849 ( .A1(n3946), .A2(n3947), .ZN(n2458) );
  NAND2_X1 U2850 ( .A1(n3958), .A2(n3474), .ZN(n3513) );
  NAND2_X1 U2851 ( .A1(n3958), .A2(n2475), .ZN(n2472) );
  INV_X1 U2852 ( .A(n3829), .ZN(n2489) );
  AOI21_X2 U2853 ( .B1(n3194), .B2(n3209), .A(n3193), .ZN(n3202) );
  NAND2_X1 U2854 ( .A1(n3359), .A2(n3194), .ZN(n4067) );
  OAI21_X1 U2855 ( .B1(n3100), .B2(n3091), .A(n3090), .ZN(n3094) );
  NAND2_X1 U2856 ( .A1(n2880), .A2(REG0_REG_1__SCAN_IN), .ZN(n2869) );
  NAND2_X1 U2857 ( .A1(n2624), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U2858 ( .A1(n3191), .A2(n3190), .ZN(n3192) );
  NAND2_X1 U2859 ( .A1(n3211), .A2(n3210), .ZN(n3236) );
  AOI21_X2 U2860 ( .B1(n3685), .B2(n2953), .A(n2952), .ZN(n3624) );
  OR2_X1 U2861 ( .A1(n2840), .A2(n2839), .ZN(n2494) );
  INV_X1 U2862 ( .A(n3289), .ZN(n3275) );
  INV_X1 U2863 ( .A(n4234), .ZN(n4914) );
  INV_X1 U2864 ( .A(n4855), .ZN(n3099) );
  INV_X1 U2865 ( .A(n4852), .ZN(n3091) );
  OR2_X1 U2866 ( .A1(n3163), .A2(n4774), .ZN(n2495) );
  NAND4_X1 U2867 ( .A1(n2926), .A2(n2925), .A3(n2924), .A4(n2923), .ZN(n4181)
         );
  INV_X1 U2868 ( .A(n4184), .ZN(n3494) );
  AND2_X1 U2869 ( .A1(n3185), .A2(n2303), .ZN(n2497) );
  AND2_X1 U2870 ( .A1(n4518), .A2(n4524), .ZN(n2498) );
  NOR2_X1 U2871 ( .A1(n3025), .A2(n4315), .ZN(n2499) );
  INV_X1 U2872 ( .A(n3143), .ZN(n2527) );
  INV_X1 U2873 ( .A(n3651), .ZN(n3514) );
  OR2_X1 U2874 ( .A1(n4276), .A2(n4646), .ZN(n2500) );
  OR2_X1 U2875 ( .A1(n4276), .A2(n4591), .ZN(n2501) );
  INV_X1 U2876 ( .A(n3827), .ZN(n3209) );
  INV_X1 U2877 ( .A(IR_REG_19__SCAN_IN), .ZN(n2508) );
  AND2_X1 U2878 ( .A1(n4341), .A2(n4131), .ZN(n4108) );
  OR2_X1 U2879 ( .A1(n3822), .A2(n3821), .ZN(n3828) );
  AND2_X1 U2880 ( .A1(n3069), .A2(n3068), .ZN(n4037) );
  NOR2_X1 U2881 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2514)
         );
  INV_X1 U2882 ( .A(n3407), .ZN(n3408) );
  INV_X1 U2883 ( .A(n4181), .ZN(n2927) );
  INV_X1 U2884 ( .A(n4047), .ZN(n2582) );
  AND2_X1 U2885 ( .A1(n2636), .A2(n2633), .ZN(n2621) );
  INV_X1 U2886 ( .A(n4194), .ZN(n2524) );
  INV_X1 U2887 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2852) );
  INV_X1 U2888 ( .A(n3222), .ZN(n3144) );
  OR2_X1 U2889 ( .A1(n4324), .A2(n4517), .ZN(n4018) );
  OR2_X1 U2890 ( .A1(n3024), .A2(n3023), .ZN(n4315) );
  NAND2_X1 U2891 ( .A1(n2962), .A2(REG3_REG_18__SCAN_IN), .ZN(n2968) );
  OR2_X1 U2892 ( .A1(n4178), .A2(n4583), .ZN(n4027) );
  NAND2_X1 U2893 ( .A1(n4184), .A2(n4819), .ZN(n2905) );
  NOR2_X1 U2894 ( .A1(n2583), .A2(n2582), .ZN(n2584) );
  AND2_X1 U2895 ( .A1(n4652), .A2(n3175), .ZN(n4443) );
  NOR2_X1 U2896 ( .A1(n2996), .A2(n3881), .ZN(n3004) );
  NOR2_X1 U2897 ( .A1(n2968), .A2(n3889), .ZN(n2975) );
  INV_X1 U2898 ( .A(n4190), .ZN(n3196) );
  INV_X1 U2899 ( .A(n4347), .ZN(n4518) );
  AND2_X1 U2900 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2954), .ZN(n2962) );
  NAND2_X1 U2901 ( .A1(n3980), .A2(n3981), .ZN(n3979) );
  AND2_X1 U2902 ( .A1(n2879), .A2(REG2_REG_0__SCAN_IN), .ZN(n2876) );
  XNOR2_X1 U2903 ( .A(n3220), .B(n3144), .ZN(n3147) );
  OR2_X1 U2904 ( .A1(n3034), .A2(n3861), .ZN(n4275) );
  OR2_X1 U2905 ( .A1(n4425), .A2(n4415), .ZN(n4385) );
  INV_X1 U2906 ( .A(n4175), .ZN(n4491) );
  INV_X1 U2907 ( .A(n4901), .ZN(n3751) );
  NOR2_X1 U2908 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  AND2_X1 U2909 ( .A1(n2915), .A2(REG3_REG_10__SCAN_IN), .ZN(n2921) );
  OR2_X1 U2910 ( .A1(n2906), .A2(n3431), .ZN(n2908) );
  AND2_X1 U2911 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2893) );
  INV_X1 U2912 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3089) );
  INV_X1 U2913 ( .A(n4480), .ZN(n3783) );
  AND2_X1 U2914 ( .A1(n4051), .A2(n3074), .ZN(n4840) );
  AND2_X1 U2915 ( .A1(n2618), .A2(n4155), .ZN(n3175) );
  AND4_X1 U2916 ( .A1(n2934), .A2(n2933), .A3(n2932), .A4(n2931), .ZN(n3666)
         );
  NOR2_X1 U2917 ( .A1(n4236), .A2(n4754), .ZN(n4240) );
  AND2_X1 U2918 ( .A1(n4275), .A2(n3035), .ZN(n4283) );
  AOI22_X1 U2919 ( .A1(n3551), .A2(n2935), .B1(n3635), .B2(n3666), .ZN(n3665)
         );
  NAND2_X1 U2920 ( .A1(n2899), .A2(REG3_REG_7__SCAN_IN), .ZN(n2906) );
  INV_X1 U2921 ( .A(n4879), .ZN(n4866) );
  NAND2_X1 U2922 ( .A1(n3091), .A2(n3089), .ZN(n3090) );
  AND2_X1 U2923 ( .A1(n2592), .A2(n2591), .ZN(n3157) );
  NAND2_X1 U2924 ( .A1(n4452), .A2(n4786), .ZN(n4587) );
  INV_X1 U2925 ( .A(n3157), .ZN(n3095) );
  AND2_X1 U2926 ( .A1(n3163), .A2(n3102), .ZN(n3159) );
  AND2_X1 U2927 ( .A1(n3131), .A2(n3130), .ZN(n4764) );
  OR2_X1 U2928 ( .A1(n3195), .A2(n3228), .ZN(n4897) );
  OR2_X1 U2929 ( .A1(n3173), .A2(n3172), .ZN(n4016) );
  NAND4_X1 U2930 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n4364)
         );
  NAND4_X1 U2931 ( .A1(n2851), .A2(n2850), .A3(n2849), .A4(n2848), .ZN(n4179)
         );
  INV_X1 U2932 ( .A(n3652), .ZN(n4182) );
  INV_X1 U2933 ( .A(n4856), .ZN(n4702) );
  NAND2_X1 U2934 ( .A1(n4826), .A2(n2620), .ZN(n4883) );
  OR2_X1 U2935 ( .A1(n2616), .A2(n4786), .ZN(n4879) );
  INV_X1 U2936 ( .A(n4305), .ZN(n4502) );
  NAND2_X1 U2937 ( .A1(n4855), .A2(n3093), .ZN(n4646) );
  INV_X1 U2938 ( .A(n4766), .ZN(n4829) );
  INV_X1 U2939 ( .A(n4712), .ZN(n4877) );
  XNOR2_X1 U2940 ( .A(n2841), .B(n2494), .ZN(U3261) );
  INV_X2 U2941 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2942 ( .A1(n2519), .A2(n2526), .ZN(n2529) );
  INV_X1 U2943 ( .A(IR_REG_27__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U2944 ( .A1(n2636), .A2(n2631), .ZN(n2515) );
  NAND2_X1 U2945 ( .A1(n2630), .A2(n2515), .ZN(n2516) );
  MUX2_X1 U2946 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2270), .Z(n3364) );
  NAND2_X1 U2947 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2518)
         );
  MUX2_X1 U2948 ( .A(IR_REG_31__SCAN_IN), .B(n2518), .S(IR_REG_1__SCAN_IN), 
        .Z(n2521) );
  INV_X1 U2949 ( .A(n2519), .ZN(n2520) );
  INV_X1 U2950 ( .A(DATAI_1_), .ZN(n2522) );
  NAND2_X1 U2951 ( .A1(n3166), .A2(n3359), .ZN(n3366) );
  INV_X1 U2952 ( .A(DATAI_2_), .ZN(n2786) );
  NAND2_X1 U2953 ( .A1(n2529), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  XNOR2_X1 U2954 ( .A(n2531), .B(n2831), .ZN(n3222) );
  INV_X1 U2955 ( .A(DATAI_3_), .ZN(n2530) );
  NAND2_X1 U2956 ( .A1(n3331), .A2(n3325), .ZN(n3332) );
  NAND2_X1 U2957 ( .A1(n2531), .A2(n2831), .ZN(n2532) );
  NAND2_X1 U2958 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  XNOR2_X1 U2959 ( .A(n2533), .B(IR_REG_4__SCAN_IN), .ZN(n4655) );
  MUX2_X1 U2960 ( .A(n4655), .B(DATAI_4_), .S(n2525), .Z(n3304) );
  NAND2_X1 U2961 ( .A1(n2534), .A2(IR_REG_31__SCAN_IN), .ZN(n2535) );
  XNOR2_X1 U2962 ( .A(n2535), .B(IR_REG_5__SCAN_IN), .ZN(n3288) );
  MUX2_X1 U2963 ( .A(n3288), .B(DATAI_5_), .S(n2525), .Z(n3438) );
  NOR2_X1 U2964 ( .A1(n2534), .A2(IR_REG_5__SCAN_IN), .ZN(n2546) );
  OR2_X1 U2965 ( .A1(n2546), .A2(n3113), .ZN(n2536) );
  XNOR2_X1 U2966 ( .A(n2536), .B(IR_REG_6__SCAN_IN), .ZN(n3289) );
  MUX2_X1 U2967 ( .A(n3289), .B(DATAI_6_), .S(n2271), .Z(n3347) );
  NAND2_X1 U2968 ( .A1(n2546), .A2(n2543), .ZN(n2537) );
  NAND2_X1 U2969 ( .A1(n2537), .A2(IR_REG_31__SCAN_IN), .ZN(n2538) );
  XNOR2_X1 U2970 ( .A(n2538), .B(IR_REG_7__SCAN_IN), .ZN(n3292) );
  MUX2_X1 U2971 ( .A(n4817), .B(n4816), .S(n2271), .Z(n4832) );
  INV_X1 U2972 ( .A(n4832), .ZN(n4819) );
  NAND2_X1 U2973 ( .A1(n2538), .A2(n2544), .ZN(n2539) );
  NAND2_X1 U2974 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  XNOR2_X1 U2975 ( .A(n2540), .B(IR_REG_8__SCAN_IN), .ZN(n4856) );
  INV_X1 U2976 ( .A(DATAI_8_), .ZN(n2541) );
  MUX2_X1 U2977 ( .A(n4702), .B(n2541), .S(n2525), .Z(n3493) );
  INV_X1 U2978 ( .A(IR_REG_8__SCAN_IN), .ZN(n2542) );
  AND3_X1 U2979 ( .A1(n2544), .A2(n2543), .A3(n2542), .ZN(n2545) );
  NAND2_X1 U2980 ( .A1(n2546), .A2(n2545), .ZN(n2548) );
  NAND2_X1 U2981 ( .A1(n2548), .A2(IR_REG_31__SCAN_IN), .ZN(n2547) );
  MUX2_X1 U2982 ( .A(IR_REG_31__SCAN_IN), .B(n2547), .S(IR_REG_9__SCAN_IN), 
        .Z(n2549) );
  NAND2_X1 U2983 ( .A1(n2549), .A2(n2551), .ZN(n3611) );
  MUX2_X1 U2984 ( .A(n3611), .B(n2779), .S(n2270), .Z(n3962) );
  NAND2_X1 U2985 ( .A1(n2551), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  XNOR2_X1 U2986 ( .A(n2550), .B(IR_REG_10__SCAN_IN), .ZN(n3613) );
  INV_X1 U2987 ( .A(n3613), .ZN(n4865) );
  INV_X1 U2988 ( .A(DATAI_10_), .ZN(n4864) );
  MUX2_X1 U2989 ( .A(n4865), .B(n4864), .S(n2271), .Z(n3539) );
  NAND2_X1 U2990 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  XNOR2_X1 U2991 ( .A(n2554), .B(IR_REG_11__SCAN_IN), .ZN(n4712) );
  MUX2_X1 U2992 ( .A(n4877), .B(n4876), .S(n2525), .Z(n3651) );
  INV_X1 U2993 ( .A(IR_REG_11__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U2994 ( .A1(n2554), .A2(n2553), .ZN(n2555) );
  NAND2_X1 U2995 ( .A1(n2555), .A2(IR_REG_31__SCAN_IN), .ZN(n2556) );
  XNOR2_X1 U2996 ( .A(n2556), .B(IR_REG_12__SCAN_IN), .ZN(n3616) );
  MUX2_X1 U2997 ( .A(n3616), .B(DATAI_12_), .S(n2270), .Z(n3556) );
  OR2_X1 U2998 ( .A1(n2312), .A2(n3113), .ZN(n2557) );
  XNOR2_X1 U2999 ( .A(n2557), .B(IR_REG_13__SCAN_IN), .ZN(n3619) );
  MUX2_X1 U3000 ( .A(n3619), .B(DATAI_13_), .S(n2270), .Z(n3574) );
  INV_X1 U3001 ( .A(IR_REG_14__SCAN_IN), .ZN(n2559) );
  XNOR2_X1 U3002 ( .A(n2562), .B(n2559), .ZN(n4224) );
  INV_X1 U3003 ( .A(DATAI_14_), .ZN(n2560) );
  NAND2_X1 U3004 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U3005 ( .A1(n2562), .A2(n2561), .ZN(n2570) );
  OR2_X1 U3006 ( .A1(n2570), .A2(IR_REG_15__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U3007 ( .A1(n2570), .A2(IR_REG_15__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U3008 ( .A1(n2565), .A2(n2563), .ZN(n4232) );
  INV_X1 U3009 ( .A(DATAI_15_), .ZN(n2564) );
  MUX2_X1 U3010 ( .A(n4232), .B(n2564), .S(n2525), .Z(n4901) );
  NAND2_X1 U3011 ( .A1(n2565), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  XNOR2_X1 U3012 ( .A(n2566), .B(IR_REG_16__SCAN_IN), .ZN(n4234) );
  INV_X1 U3013 ( .A(DATAI_16_), .ZN(n4913) );
  MUX2_X1 U3014 ( .A(n4914), .B(n4913), .S(n2525), .Z(n4571) );
  INV_X1 U3015 ( .A(n2567), .ZN(n2568) );
  INV_X1 U3016 ( .A(IR_REG_17__SCAN_IN), .ZN(n2571) );
  XNOR2_X1 U3017 ( .A(n2574), .B(n2571), .ZN(n4241) );
  INV_X1 U3018 ( .A(DATAI_17_), .ZN(n2572) );
  MUX2_X1 U3019 ( .A(n4241), .B(n2572), .S(n2271), .Z(n4566) );
  NAND2_X1 U3020 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U3021 ( .A1(n2574), .A2(n2573), .ZN(n2575) );
  XNOR2_X1 U3022 ( .A(n2575), .B(IR_REG_18__SCAN_IN), .ZN(n4268) );
  INV_X1 U3023 ( .A(DATAI_18_), .ZN(n2764) );
  MUX2_X1 U3024 ( .A(n4268), .B(n2764), .S(n2270), .Z(n4490) );
  INV_X1 U3025 ( .A(n2575), .ZN(n2577) );
  NAND2_X1 U3026 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U3027 ( .A1(n2577), .A2(n2576), .ZN(n2579) );
  INV_X1 U3028 ( .A(n2579), .ZN(n2578) );
  NAND2_X1 U3029 ( .A1(n2578), .A2(n2508), .ZN(n2608) );
  NAND2_X1 U3030 ( .A1(n2579), .A2(IR_REG_19__SCAN_IN), .ZN(n2580) );
  NAND2_X2 U3031 ( .A1(n2608), .A2(n2580), .ZN(n4766) );
  INV_X1 U3032 ( .A(DATAI_19_), .ZN(n2581) );
  MUX2_X1 U3033 ( .A(n4766), .B(n2581), .S(n2525), .Z(n4480) );
  NAND2_X1 U3034 ( .A1(n2271), .A2(DATAI_20_), .ZN(n4456) );
  NAND2_X1 U3035 ( .A1(n2271), .A2(DATAI_22_), .ZN(n4415) );
  NAND2_X1 U3036 ( .A1(n2270), .A2(DATAI_23_), .ZN(n4395) );
  NAND2_X1 U3037 ( .A1(n2525), .A2(DATAI_24_), .ZN(n4369) );
  INV_X1 U3038 ( .A(n4369), .ZN(n3823) );
  NAND2_X1 U3039 ( .A1(n2271), .A2(DATAI_25_), .ZN(n4350) );
  NAND2_X1 U3040 ( .A1(n2271), .A2(DATAI_26_), .ZN(n4524) );
  INV_X1 U3041 ( .A(n4524), .ZN(n3832) );
  NAND2_X1 U3042 ( .A1(n2525), .A2(DATAI_27_), .ZN(n4517) );
  INV_X1 U3043 ( .A(n4517), .ZN(n3845) );
  NAND2_X1 U3044 ( .A1(n2525), .A2(DATAI_28_), .ZN(n4288) );
  INV_X1 U3045 ( .A(n4288), .ZN(n3853) );
  NAND2_X1 U3046 ( .A1(n2270), .A2(DATAI_29_), .ZN(n4280) );
  AND2_X1 U3047 ( .A1(n2271), .A2(DATAI_30_), .ZN(n4047) );
  INV_X1 U3048 ( .A(IR_REG_23__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U3049 ( .A1(n2607), .A2(n2606), .ZN(n2605) );
  NAND2_X1 U3050 ( .A1(n2605), .A2(IR_REG_31__SCAN_IN), .ZN(n2585) );
  INV_X1 U3051 ( .A(n4650), .ZN(n2590) );
  NAND2_X1 U3052 ( .A1(n2292), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  INV_X1 U3053 ( .A(n3106), .ZN(n2603) );
  NAND2_X1 U3054 ( .A1(n2590), .A2(n2603), .ZN(n2587) );
  MUX2_X1 U3055 ( .A(n2590), .B(n2587), .S(B_REG_SCAN_IN), .Z(n2589) );
  NAND2_X1 U3056 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  INV_X1 U3057 ( .A(D_REG_0__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U3058 ( .A1(n3116), .A2(n3119), .ZN(n2592) );
  INV_X1 U3059 ( .A(n4649), .ZN(n2604) );
  NAND2_X1 U3060 ( .A1(n2604), .A2(n2590), .ZN(n2591) );
  NOR4_X1 U3061 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2596) );
  NOR4_X1 U3062 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2595) );
  NOR4_X1 U3063 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2594) );
  NOR4_X1 U3064 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2593) );
  NAND4_X1 U3065 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n2602)
         );
  NOR2_X1 U3066 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_30__SCAN_IN), .ZN(n2600)
         );
  NOR4_X1 U3067 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2599) );
  NOR4_X1 U3068 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2598) );
  NOR4_X1 U3069 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2597) );
  NAND4_X1 U3070 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n2601)
         );
  OAI21_X1 U3071 ( .B1(n2602), .B2(n2601), .A(n3116), .ZN(n3087) );
  NAND2_X1 U3072 ( .A1(n2604), .A2(n2603), .ZN(n3123) );
  AND2_X1 U3073 ( .A1(n3087), .A2(n3123), .ZN(n3158) );
  OAI21_X1 U3074 ( .B1(n2607), .B2(n2606), .A(n2605), .ZN(n3244) );
  AND2_X1 U3075 ( .A1(n3244), .A2(STATE_REG_SCAN_IN), .ZN(n3102) );
  INV_X1 U3076 ( .A(IR_REG_20__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U3077 ( .A1(n2619), .A2(n4766), .ZN(n3169) );
  NAND2_X1 U3078 ( .A1(n2611), .A2(IR_REG_31__SCAN_IN), .ZN(n2612) );
  XNOR2_X1 U3079 ( .A(n2612), .B(n2493), .ZN(n2618) );
  NAND2_X1 U3080 ( .A1(n2613), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  AND2_X1 U3081 ( .A1(n4651), .A2(n4157), .ZN(n3121) );
  NAND2_X1 U3082 ( .A1(n3169), .A2(n3121), .ZN(n3243) );
  NAND2_X1 U3083 ( .A1(n3159), .A2(n3243), .ZN(n3084) );
  INV_X1 U3084 ( .A(n3084), .ZN(n3178) );
  INV_X1 U3085 ( .A(D_REG_1__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U3086 ( .A1(n3116), .A2(n2615), .ZN(n3156) );
  NAND4_X1 U3087 ( .A1(n3095), .A2(n3158), .A3(n3178), .A4(n3156), .ZN(n2617)
         );
  INV_X1 U3088 ( .A(n4157), .ZN(n4155) );
  NAND2_X1 U3089 ( .A1(n3159), .A2(n4155), .ZN(n2616) );
  AND2_X1 U3090 ( .A1(n2619), .A2(n4829), .ZN(n4777) );
  NAND2_X1 U3091 ( .A1(n4777), .A2(n2618), .ZN(n4786) );
  AND2_X2 U3092 ( .A1(n2619), .A2(n3175), .ZN(n3093) );
  NAND2_X1 U3093 ( .A1(n3093), .A2(n4766), .ZN(n3164) );
  INV_X1 U3094 ( .A(n3164), .ZN(n2620) );
  NOR2_X1 U3095 ( .A1(n4509), .A2(n4883), .ZN(n2643) );
  INV_X1 U3096 ( .A(n2619), .ZN(n4652) );
  INV_X2 U3097 ( .A(n4443), .ZN(n4833) );
  NOR2_X1 U3098 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2633)
         );
  NAND2_X1 U3099 ( .A1(n3075), .A2(REG1_REG_31__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3100 ( .A1(n2879), .A2(REG2_REG_31__SCAN_IN), .ZN(n2628) );
  INV_X1 U3101 ( .A(n2842), .ZN(n2626) );
  NAND2_X1 U3102 ( .A1(n2887), .A2(REG0_REG_31__SCAN_IN), .ZN(n2627) );
  NAND3_X1 U3103 ( .A1(n2629), .A2(n2628), .A3(n2627), .ZN(n4173) );
  INV_X1 U3104 ( .A(n4173), .ZN(n4048) );
  XNOR2_X1 U3105 ( .A(n2630), .B(n2631), .ZN(n4168) );
  INV_X1 U3106 ( .A(B_REG_SCAN_IN), .ZN(n2638) );
  INV_X1 U3107 ( .A(n2632), .ZN(n2634) );
  AND2_X1 U3108 ( .A1(n2634), .A2(n2633), .ZN(n2635) );
  OR2_X1 U3109 ( .A1(n2635), .A2(n3113), .ZN(n2637) );
  XNOR2_X1 U3110 ( .A(n2637), .B(n2636), .ZN(n4916) );
  OAI21_X1 U3111 ( .B1(n4168), .B2(n2638), .A(n4838), .ZN(n3079) );
  NOR2_X1 U3112 ( .A1(n4048), .A2(n3079), .ZN(n4271) );
  INV_X1 U3113 ( .A(n4271), .ZN(n2639) );
  OAI21_X1 U3114 ( .B1(n2582), .B2(n4833), .A(n2639), .ZN(n4598) );
  NAND2_X1 U3115 ( .A1(n4598), .A2(n4889), .ZN(n2641) );
  NAND2_X1 U3116 ( .A1(n4462), .A2(REG2_REG_30__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3117 ( .A1(n2641), .A2(n2640), .ZN(n2642) );
  AOI22_X1 U3118 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_125), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_124), .ZN(n2644) );
  OAI221_X1 U3119 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_124), .A(n2644), .ZN(n2734) );
  INV_X1 U3120 ( .A(keyinput_123), .ZN(n2731) );
  INV_X1 U3121 ( .A(keyinput_122), .ZN(n2729) );
  INV_X1 U3122 ( .A(keyinput_113), .ZN(n2716) );
  INV_X1 U3123 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3939) );
  INV_X1 U3124 ( .A(keyinput_112), .ZN(n2714) );
  INV_X1 U3125 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3930) );
  INV_X1 U3126 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3908) );
  OAI22_X1 U3127 ( .A1(n3531), .A2(keyinput_108), .B1(n3908), .B2(keyinput_109), .ZN(n2645) );
  AOI221_X1 U3128 ( .B1(n3531), .B2(keyinput_108), .C1(keyinput_109), .C2(
        n3908), .A(n2645), .ZN(n2712) );
  INV_X1 U3129 ( .A(keyinput_107), .ZN(n2708) );
  INV_X1 U3130 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2805) );
  OAI22_X1 U3131 ( .A1(n3431), .A2(keyinput_105), .B1(keyinput_104), .B2(
        REG3_REG_28__SCAN_IN), .ZN(n2646) );
  AOI221_X1 U3132 ( .B1(n3431), .B2(keyinput_105), .C1(REG3_REG_28__SCAN_IN), 
        .C2(keyinput_104), .A(n2646), .ZN(n2705) );
  INV_X1 U3133 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3889) );
  INV_X1 U3134 ( .A(keyinput_103), .ZN(n2703) );
  XOR2_X1 U3135 ( .A(DATAI_0_), .B(keyinput_95), .Z(n2701) );
  INV_X1 U3136 ( .A(DATAI_7_), .ZN(n4816) );
  INV_X1 U3137 ( .A(DATAI_6_), .ZN(n4808) );
  OAI22_X1 U3138 ( .A1(n4816), .A2(keyinput_88), .B1(n4808), .B2(keyinput_89), 
        .ZN(n2647) );
  AOI221_X1 U3139 ( .B1(n4816), .B2(keyinput_88), .C1(keyinput_89), .C2(n4808), 
        .A(n2647), .ZN(n2683) );
  INV_X1 U3140 ( .A(keyinput_86), .ZN(n2681) );
  INV_X1 U3141 ( .A(DATAI_9_), .ZN(n2779) );
  INV_X1 U3142 ( .A(keyinput_85), .ZN(n2679) );
  INV_X1 U3143 ( .A(keyinput_84), .ZN(n2677) );
  INV_X1 U3144 ( .A(DATAI_11_), .ZN(n4876) );
  INV_X1 U3145 ( .A(keyinput_83), .ZN(n2675) );
  INV_X1 U3146 ( .A(DATAI_12_), .ZN(n4891) );
  INV_X1 U3147 ( .A(keyinput_82), .ZN(n2673) );
  INV_X1 U31480 ( .A(DATAI_13_), .ZN(n4893) );
  OAI22_X1 U31490 ( .A1(n4913), .A2(keyinput_79), .B1(keyinput_80), .B2(
        DATAI_15_), .ZN(n2648) );
  AOI221_X1 U3150 ( .B1(n4913), .B2(keyinput_79), .C1(DATAI_15_), .C2(
        keyinput_80), .A(n2648), .ZN(n2671) );
  OAI22_X1 U3151 ( .A1(DATAI_17_), .A2(keyinput_78), .B1(keyinput_81), .B2(
        DATAI_14_), .ZN(n2649) );
  AOI221_X1 U3152 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(DATAI_14_), .C2(
        keyinput_81), .A(n2649), .ZN(n2670) );
  INV_X1 U3153 ( .A(keyinput_77), .ZN(n2668) );
  INV_X1 U3154 ( .A(DATAI_21_), .ZN(n3104) );
  INV_X1 U3155 ( .A(keyinput_73), .ZN(n2662) );
  INV_X1 U3156 ( .A(DATAI_22_), .ZN(n2757) );
  AOI22_X1 U3157 ( .A1(DATAI_24_), .A2(keyinput_71), .B1(DATAI_25_), .B2(
        keyinput_70), .ZN(n2650) );
  OAI221_X1 U3158 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(DATAI_25_), .C2(
        keyinput_70), .A(n2650), .ZN(n2659) );
  INV_X1 U3159 ( .A(DATAI_26_), .ZN(n2751) );
  INV_X1 U3160 ( .A(keyinput_69), .ZN(n2657) );
  INV_X1 U3161 ( .A(DATAI_29_), .ZN(n3110) );
  INV_X1 U3162 ( .A(DATAI_28_), .ZN(n4915) );
  AOI22_X1 U3163 ( .A1(n3110), .A2(keyinput_66), .B1(keyinput_67), .B2(n4915), 
        .ZN(n2651) );
  OAI221_X1 U3164 ( .B1(n3110), .B2(keyinput_66), .C1(n4915), .C2(keyinput_67), 
        .A(n2651), .ZN(n2654) );
  OAI22_X1 U3165 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        DATAI_31_), .ZN(n2652) );
  AOI221_X1 U3166 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n2652), .ZN(n2653) );
  OAI22_X1 U3167 ( .A1(n2654), .A2(n2653), .B1(keyinput_68), .B2(DATAI_27_), 
        .ZN(n2655) );
  AOI21_X1 U3168 ( .B1(keyinput_68), .B2(DATAI_27_), .A(n2655), .ZN(n2656) );
  AOI221_X1 U3169 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(n2751), .C2(n2657), 
        .A(n2656), .ZN(n2658) );
  OAI22_X1 U3170 ( .A1(n2659), .A2(n2658), .B1(keyinput_72), .B2(DATAI_23_), 
        .ZN(n2660) );
  AOI21_X1 U3171 ( .B1(keyinput_72), .B2(DATAI_23_), .A(n2660), .ZN(n2661) );
  AOI221_X1 U3172 ( .B1(DATAI_22_), .B2(n2662), .C1(n2757), .C2(keyinput_73), 
        .A(n2661), .ZN(n2665) );
  INV_X1 U3173 ( .A(DATAI_20_), .ZN(n2759) );
  AOI22_X1 U3174 ( .A1(n2759), .A2(keyinput_75), .B1(keyinput_76), .B2(n2581), 
        .ZN(n2663) );
  OAI221_X1 U3175 ( .B1(n2759), .B2(keyinput_75), .C1(n2581), .C2(keyinput_76), 
        .A(n2663), .ZN(n2664) );
  AOI211_X1 U3176 ( .C1(n3104), .C2(keyinput_74), .A(n2665), .B(n2664), .ZN(
        n2666) );
  OAI21_X1 U3177 ( .B1(n3104), .B2(keyinput_74), .A(n2666), .ZN(n2667) );
  OAI221_X1 U3178 ( .B1(DATAI_18_), .B2(keyinput_77), .C1(n2764), .C2(n2668), 
        .A(n2667), .ZN(n2669) );
  NAND3_X1 U3179 ( .A1(n2671), .A2(n2670), .A3(n2669), .ZN(n2672) );
  OAI221_X1 U3180 ( .B1(DATAI_13_), .B2(n2673), .C1(n4893), .C2(keyinput_82), 
        .A(n2672), .ZN(n2674) );
  OAI221_X1 U3181 ( .B1(DATAI_12_), .B2(n2675), .C1(n4891), .C2(keyinput_83), 
        .A(n2674), .ZN(n2676) );
  OAI221_X1 U3182 ( .B1(DATAI_11_), .B2(n2677), .C1(n4876), .C2(keyinput_84), 
        .A(n2676), .ZN(n2678) );
  OAI221_X1 U3183 ( .B1(DATAI_10_), .B2(n2679), .C1(n4864), .C2(keyinput_85), 
        .A(n2678), .ZN(n2680) );
  OAI221_X1 U3184 ( .B1(DATAI_9_), .B2(n2681), .C1(n2779), .C2(keyinput_86), 
        .A(n2680), .ZN(n2682) );
  OAI211_X1 U3185 ( .C1(DATAI_8_), .C2(keyinput_87), .A(n2683), .B(n2682), 
        .ZN(n2684) );
  AOI21_X1 U3186 ( .B1(DATAI_8_), .B2(keyinput_87), .A(n2684), .ZN(n2687) );
  INV_X1 U3187 ( .A(DATAI_5_), .ZN(n4806) );
  AOI22_X1 U3188 ( .A1(DATAI_4_), .A2(keyinput_91), .B1(n4806), .B2(
        keyinput_90), .ZN(n2685) );
  OAI221_X1 U3189 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(n4806), .C2(
        keyinput_90), .A(n2685), .ZN(n2686) );
  OAI22_X1 U3190 ( .A1(n2687), .A2(n2686), .B1(DATAI_3_), .B2(keyinput_92), 
        .ZN(n2688) );
  AOI21_X1 U3191 ( .B1(DATAI_3_), .B2(keyinput_92), .A(n2688), .ZN(n2691) );
  XNOR2_X1 U3192 ( .A(n2786), .B(keyinput_93), .ZN(n2690) );
  XNOR2_X1 U3193 ( .A(keyinput_94), .B(n2522), .ZN(n2689) );
  OR3_X1 U3194 ( .A1(n2691), .A2(n2690), .A3(n2689), .ZN(n2700) );
  INV_X1 U3195 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2936) );
  OAI22_X1 U3196 ( .A1(n2936), .A2(keyinput_99), .B1(keyinput_101), .B2(
        REG3_REG_10__SCAN_IN), .ZN(n2692) );
  AOI221_X1 U3197 ( .B1(n2936), .B2(keyinput_99), .C1(REG3_REG_10__SCAN_IN), 
        .C2(keyinput_101), .A(n2692), .ZN(n2699) );
  INV_X1 U3198 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3871) );
  INV_X1 U3199 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U3200 ( .A1(n3871), .A2(keyinput_98), .B1(n4793), .B2(keyinput_102), 
        .ZN(n2693) );
  OAI221_X1 U3201 ( .B1(n3871), .B2(keyinput_98), .C1(n4793), .C2(keyinput_102), .A(n2693), .ZN(n2697) );
  INV_X1 U3202 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3413) );
  OAI22_X1 U3203 ( .A1(n3413), .A2(keyinput_97), .B1(keyinput_100), .B2(
        REG3_REG_23__SCAN_IN), .ZN(n2694) );
  AOI221_X1 U3204 ( .B1(n3413), .B2(keyinput_97), .C1(REG3_REG_23__SCAN_IN), 
        .C2(keyinput_100), .A(n2694), .ZN(n2695) );
  OAI21_X1 U3205 ( .B1(keyinput_96), .B2(STATE_REG_SCAN_IN), .A(n2695), .ZN(
        n2696) );
  AOI211_X1 U3206 ( .C1(keyinput_96), .C2(STATE_REG_SCAN_IN), .A(n2697), .B(
        n2696), .ZN(n2698) );
  OAI211_X1 U3207 ( .C1(n2701), .C2(n2700), .A(n2699), .B(n2698), .ZN(n2702)
         );
  OAI221_X1 U3208 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_103), .C1(n3889), 
        .C2(n2703), .A(n2702), .ZN(n2704) );
  AOI22_X1 U3209 ( .A1(n2705), .A2(n2704), .B1(keyinput_106), .B2(
        REG3_REG_1__SCAN_IN), .ZN(n2706) );
  OAI21_X1 U32100 ( .B1(keyinput_106), .B2(REG3_REG_1__SCAN_IN), .A(n2706), 
        .ZN(n2707) );
  OAI221_X1 U32110 ( .B1(REG3_REG_21__SCAN_IN), .B2(n2708), .C1(n2805), .C2(
        keyinput_107), .A(n2707), .ZN(n2711) );
  INV_X1 U32120 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3921) );
  INV_X1 U32130 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U32140 ( .A1(n3921), .A2(keyinput_110), .B1(n3314), .B2(
        keyinput_111), .ZN(n2709) );
  OAI221_X1 U32150 ( .B1(n3921), .B2(keyinput_110), .C1(n3314), .C2(
        keyinput_111), .A(n2709), .ZN(n2710) );
  AOI21_X1 U32160 ( .B1(n2712), .B2(n2711), .A(n2710), .ZN(n2713) );
  AOI221_X1 U32170 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2714), .C1(n3930), .C2(
        keyinput_112), .A(n2713), .ZN(n2715) );
  AOI221_X1 U32180 ( .B1(REG3_REG_24__SCAN_IN), .B2(n2716), .C1(n3939), .C2(
        keyinput_113), .A(n2715), .ZN(n2722) );
  INV_X1 U32190 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2718) );
  INV_X1 U32200 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U32210 ( .A1(n2718), .A2(keyinput_116), .B1(n3974), .B2(
        keyinput_117), .ZN(n2717) );
  OAI221_X1 U32220 ( .B1(n2718), .B2(keyinput_116), .C1(n3974), .C2(
        keyinput_117), .A(n2717), .ZN(n2721) );
  INV_X1 U32230 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U32240 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_115), .B1(n3218), 
        .B2(keyinput_114), .ZN(n2719) );
  OAI221_X1 U32250 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_115), .C1(n3218), 
        .C2(keyinput_114), .A(n2719), .ZN(n2720) );
  NOR3_X1 U32260 ( .A1(n2722), .A2(n2721), .A3(n2720), .ZN(n2727) );
  INV_X1 U32270 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3579) );
  INV_X1 U32280 ( .A(IR_REG_1__SCAN_IN), .ZN(n2822) );
  AOI22_X1 U32290 ( .A1(n3579), .A2(keyinput_118), .B1(n2822), .B2(
        keyinput_120), .ZN(n2723) );
  OAI221_X1 U32300 ( .B1(n3579), .B2(keyinput_118), .C1(n2822), .C2(
        keyinput_120), .A(n2723), .ZN(n2726) );
  AOI22_X1 U32310 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_121), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_119), .ZN(n2724) );
  OAI221_X1 U32320 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_121), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_119), .A(n2724), .ZN(n2725) );
  NOR3_X1 U32330 ( .A1(n2727), .A2(n2726), .A3(n2725), .ZN(n2728) );
  AOI221_X1 U32340 ( .B1(IR_REG_4__SCAN_IN), .B2(n2731), .C1(n2502), .C2(
        keyinput_123), .A(n2730), .ZN(n2733) );
  NAND2_X1 U32350 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_126), .ZN(n2732) );
  OAI221_X1 U32360 ( .B1(n2734), .B2(n2733), .C1(IR_REG_7__SCAN_IN), .C2(
        keyinput_126), .A(n2732), .ZN(n2736) );
  AOI21_X1 U32370 ( .B1(keyinput_127), .B2(n2736), .A(keyinput_63), .ZN(n2738)
         );
  INV_X1 U32380 ( .A(keyinput_127), .ZN(n2735) );
  AOI21_X1 U32390 ( .B1(n2736), .B2(n2735), .A(IR_REG_8__SCAN_IN), .ZN(n2737)
         );
  AOI22_X1 U32400 ( .A1(IR_REG_8__SCAN_IN), .A2(n2738), .B1(keyinput_63), .B2(
        n2737), .ZN(n2840) );
  INV_X1 U32410 ( .A(keyinput_59), .ZN(n2833) );
  INV_X1 U32420 ( .A(keyinput_58), .ZN(n2830) );
  XOR2_X1 U32430 ( .A(keyinput_49), .B(REG3_REG_24__SCAN_IN), .Z(n2819) );
  INV_X1 U32440 ( .A(keyinput_48), .ZN(n2815) );
  XNOR2_X1 U32450 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n2808) );
  INV_X1 U32460 ( .A(DATAI_0_), .ZN(n4773) );
  AOI22_X1 U32470 ( .A1(DATAI_4_), .A2(keyinput_27), .B1(n4806), .B2(
        keyinput_26), .ZN(n2739) );
  OAI221_X1 U32480 ( .B1(DATAI_4_), .B2(keyinput_27), .C1(n4806), .C2(
        keyinput_26), .A(n2739), .ZN(n2784) );
  OAI22_X1 U32490 ( .A1(DATAI_7_), .A2(keyinput_24), .B1(DATAI_6_), .B2(
        keyinput_25), .ZN(n2740) );
  AOI221_X1 U32500 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(keyinput_25), .C2(
        DATAI_6_), .A(n2740), .ZN(n2781) );
  INV_X1 U32510 ( .A(keyinput_22), .ZN(n2778) );
  INV_X1 U32520 ( .A(keyinput_21), .ZN(n2776) );
  INV_X1 U32530 ( .A(keyinput_20), .ZN(n2774) );
  INV_X1 U32540 ( .A(keyinput_19), .ZN(n2772) );
  INV_X1 U32550 ( .A(keyinput_18), .ZN(n2770) );
  OAI22_X1 U32560 ( .A1(n2564), .A2(keyinput_16), .B1(keyinput_14), .B2(
        DATAI_17_), .ZN(n2741) );
  AOI221_X1 U32570 ( .B1(n2564), .B2(keyinput_16), .C1(DATAI_17_), .C2(
        keyinput_14), .A(n2741), .ZN(n2768) );
  OAI22_X1 U32580 ( .A1(DATAI_16_), .A2(keyinput_15), .B1(keyinput_17), .B2(
        DATAI_14_), .ZN(n2742) );
  AOI221_X1 U32590 ( .B1(DATAI_16_), .B2(keyinput_15), .C1(DATAI_14_), .C2(
        keyinput_17), .A(n2742), .ZN(n2767) );
  INV_X1 U32600 ( .A(keyinput_13), .ZN(n2765) );
  INV_X1 U32610 ( .A(keyinput_9), .ZN(n2756) );
  INV_X1 U32620 ( .A(DATAI_25_), .ZN(n3108) );
  AOI22_X1 U32630 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(n3108), .B2(
        keyinput_6), .ZN(n2743) );
  OAI221_X1 U32640 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(n3108), .C2(
        keyinput_6), .A(n2743), .ZN(n2753) );
  INV_X1 U32650 ( .A(keyinput_5), .ZN(n2750) );
  INV_X1 U32660 ( .A(DATAI_27_), .ZN(n3112) );
  AOI22_X1 U32670 ( .A1(DATAI_29_), .A2(keyinput_2), .B1(n4915), .B2(
        keyinput_3), .ZN(n2744) );
  OAI221_X1 U32680 ( .B1(DATAI_29_), .B2(keyinput_2), .C1(n4915), .C2(
        keyinput_3), .A(n2744), .ZN(n2747) );
  OAI22_X1 U32690 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        DATAI_31_), .ZN(n2745) );
  AOI221_X1 U32700 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n2745), .ZN(n2746) );
  OAI22_X1 U32710 ( .A1(keyinput_4), .A2(n3112), .B1(n2747), .B2(n2746), .ZN(
        n2748) );
  AOI21_X1 U32720 ( .B1(keyinput_4), .B2(n3112), .A(n2748), .ZN(n2749) );
  AOI221_X1 U32730 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n2751), .C2(n2750), 
        .A(n2749), .ZN(n2752) );
  OAI22_X1 U32740 ( .A1(n2753), .A2(n2752), .B1(keyinput_8), .B2(DATAI_23_), 
        .ZN(n2754) );
  AOI21_X1 U32750 ( .B1(keyinput_8), .B2(DATAI_23_), .A(n2754), .ZN(n2755) );
  AOI221_X1 U32760 ( .B1(DATAI_22_), .B2(keyinput_9), .C1(n2757), .C2(n2756), 
        .A(n2755), .ZN(n2761) );
  AOI22_X1 U32770 ( .A1(DATAI_21_), .A2(keyinput_10), .B1(n2759), .B2(
        keyinput_11), .ZN(n2758) );
  OAI221_X1 U32780 ( .B1(DATAI_21_), .B2(keyinput_10), .C1(n2759), .C2(
        keyinput_11), .A(n2758), .ZN(n2760) );
  AOI211_X1 U32790 ( .C1(DATAI_19_), .C2(keyinput_12), .A(n2761), .B(n2760), 
        .ZN(n2762) );
  OAI21_X1 U32800 ( .B1(DATAI_19_), .B2(keyinput_12), .A(n2762), .ZN(n2763) );
  OAI221_X1 U32810 ( .B1(DATAI_18_), .B2(n2765), .C1(n2764), .C2(keyinput_13), 
        .A(n2763), .ZN(n2766) );
  NAND3_X1 U32820 ( .A1(n2768), .A2(n2767), .A3(n2766), .ZN(n2769) );
  OAI221_X1 U32830 ( .B1(DATAI_13_), .B2(n2770), .C1(n4893), .C2(keyinput_18), 
        .A(n2769), .ZN(n2771) );
  OAI221_X1 U32840 ( .B1(DATAI_12_), .B2(n2772), .C1(n4891), .C2(keyinput_19), 
        .A(n2771), .ZN(n2773) );
  OAI221_X1 U32850 ( .B1(DATAI_11_), .B2(keyinput_20), .C1(n4876), .C2(n2774), 
        .A(n2773), .ZN(n2775) );
  OAI221_X1 U32860 ( .B1(DATAI_10_), .B2(keyinput_21), .C1(n4864), .C2(n2776), 
        .A(n2775), .ZN(n2777) );
  OAI221_X1 U32870 ( .B1(DATAI_9_), .B2(keyinput_22), .C1(n2779), .C2(n2778), 
        .A(n2777), .ZN(n2780) );
  OAI211_X1 U32880 ( .C1(DATAI_8_), .C2(keyinput_23), .A(n2781), .B(n2780), 
        .ZN(n2782) );
  AOI21_X1 U32890 ( .B1(DATAI_8_), .B2(keyinput_23), .A(n2782), .ZN(n2783) );
  OAI22_X1 U32900 ( .A1(keyinput_28), .A2(n2530), .B1(n2784), .B2(n2783), .ZN(
        n2785) );
  AOI21_X1 U32910 ( .B1(keyinput_28), .B2(n2530), .A(n2785), .ZN(n2790) );
  XNOR2_X1 U32920 ( .A(n2786), .B(keyinput_29), .ZN(n2789) );
  AND2_X1 U32930 ( .A1(keyinput_31), .A2(n4773), .ZN(n2788) );
  XNOR2_X1 U32940 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n2787) );
  NOR4_X1 U32950 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(n2791)
         );
  OAI21_X1 U32960 ( .B1(n4773), .B2(keyinput_31), .A(n2791), .ZN(n2801) );
  XOR2_X1 U32970 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_38), .Z(n2798) );
  INV_X1 U32980 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U32990 ( .A1(n3477), .A2(keyinput_37), .B1(U3149), .B2(keyinput_32), 
        .ZN(n2792) );
  OAI221_X1 U33000 ( .B1(n3477), .B2(keyinput_37), .C1(U3149), .C2(keyinput_32), .A(n2792), .ZN(n2797) );
  AOI22_X1 U33010 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_35), .B1(n3871), 
        .B2(keyinput_34), .ZN(n2793) );
  OAI221_X1 U33020 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_35), .C1(n3871), 
        .C2(keyinput_34), .A(n2793), .ZN(n2796) );
  AOI22_X1 U33030 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_36), .B1(n3413), 
        .B2(keyinput_33), .ZN(n2794) );
  OAI221_X1 U33040 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_36), .C1(n3413), 
        .C2(keyinput_33), .A(n2794), .ZN(n2795) );
  NOR4_X1 U33050 ( .A1(n2798), .A2(n2797), .A3(n2796), .A4(n2795), .ZN(n2800)
         );
  NOR2_X1 U33060 ( .A1(n3889), .A2(keyinput_39), .ZN(n2799) );
  AOI221_X1 U33070 ( .B1(n2801), .B2(n2800), .C1(keyinput_39), .C2(n3889), .A(
        n2799), .ZN(n2804) );
  AOI22_X1 U33080 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_40), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput_41), .ZN(n2802) );
  OAI221_X1 U33090 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_40), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput_41), .A(n2802), .ZN(n2803) );
  OR2_X1 U33100 ( .A1(n2804), .A2(n2803), .ZN(n2807) );
  INV_X1 U33110 ( .A(keyinput_43), .ZN(n2806) );
  AOI222_X1 U33120 ( .A1(n2808), .A2(n2807), .B1(n2806), .B2(n2805), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_43), .ZN(n2813) );
  AOI22_X1 U33130 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_44), .B1(n3908), 
        .B2(keyinput_45), .ZN(n2809) );
  OAI221_X1 U33140 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_44), .C1(n3908), 
        .C2(keyinput_45), .A(n2809), .ZN(n2812) );
  OAI22_X1 U33150 ( .A1(n3314), .A2(keyinput_47), .B1(keyinput_46), .B2(
        REG3_REG_16__SCAN_IN), .ZN(n2810) );
  AOI221_X1 U33160 ( .B1(n3314), .B2(keyinput_47), .C1(REG3_REG_16__SCAN_IN), 
        .C2(keyinput_46), .A(n2810), .ZN(n2811) );
  OAI21_X1 U33170 ( .B1(n2813), .B2(n2812), .A(n2811), .ZN(n2814) );
  OAI221_X1 U33180 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2815), .C1(n3930), .C2(
        keyinput_48), .A(n2814), .ZN(n2818) );
  AOI22_X1 U33190 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_52), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput_53), .ZN(n2816) );
  OAI221_X1 U33200 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_52), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_53), .A(n2816), .ZN(n2817) );
  AOI21_X1 U33210 ( .B1(n2819), .B2(n2818), .A(n2817), .ZN(n2828) );
  OAI22_X1 U33220 ( .A1(n2852), .A2(keyinput_51), .B1(keyinput_50), .B2(
        REG3_REG_4__SCAN_IN), .ZN(n2820) );
  AOI221_X1 U33230 ( .B1(n2852), .B2(keyinput_51), .C1(REG3_REG_4__SCAN_IN), 
        .C2(keyinput_50), .A(n2820), .ZN(n2827) );
  INV_X1 U33240 ( .A(IR_REG_0__SCAN_IN), .ZN(n4774) );
  AOI22_X1 U33250 ( .A1(n4774), .A2(keyinput_55), .B1(keyinput_54), .B2(n3579), 
        .ZN(n2821) );
  OAI221_X1 U33260 ( .B1(n4774), .B2(keyinput_55), .C1(n3579), .C2(keyinput_54), .A(n2821), .ZN(n2826) );
  XOR2_X1 U33270 ( .A(n2822), .B(keyinput_56), .Z(n2824) );
  XNOR2_X1 U33280 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n2823) );
  NAND2_X1 U33290 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  AOI211_X1 U33300 ( .C1(n2828), .C2(n2827), .A(n2826), .B(n2825), .ZN(n2829)
         );
  AOI221_X1 U33310 ( .B1(IR_REG_4__SCAN_IN), .B2(n2833), .C1(n2502), .C2(
        keyinput_59), .A(n2832), .ZN(n2837) );
  XOR2_X1 U33320 ( .A(keyinput_61), .B(n2543), .Z(n2835) );
  XNOR2_X1 U33330 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n2834) );
  NAND2_X1 U33340 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  OAI22_X1 U33350 ( .A1(n2837), .A2(n2836), .B1(IR_REG_7__SCAN_IN), .B2(
        keyinput_62), .ZN(n2838) );
  AOI21_X1 U33360 ( .B1(keyinput_62), .B2(IR_REG_7__SCAN_IN), .A(n2838), .ZN(
        n2839) );
  NAND2_X1 U33370 ( .A1(n2887), .A2(REG0_REG_16__SCAN_IN), .ZN(n2846) );
  NAND2_X1 U33380 ( .A1(n2879), .A2(REG2_REG_16__SCAN_IN), .ZN(n2845) );
  AOI21_X1 U33390 ( .B1(n2945), .B2(n3921), .A(n2954), .ZN(n3923) );
  NAND2_X1 U33400 ( .A1(n2998), .A2(n3923), .ZN(n2844) );
  NAND2_X1 U33410 ( .A1(n3075), .A2(REG1_REG_16__SCAN_IN), .ZN(n2843) );
  NAND4_X1 U33420 ( .A1(n2846), .A2(n2845), .A3(n2844), .A4(n2843), .ZN(n4176)
         );
  INV_X1 U33430 ( .A(n4176), .ZN(n4898) );
  NAND2_X1 U33440 ( .A1(n2887), .A2(REG0_REG_13__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U33450 ( .A1(n2879), .A2(REG2_REG_13__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U33460 ( .A1(n2930), .A2(n3579), .ZN(n2847) );
  AND2_X1 U33470 ( .A1(n2937), .A2(n2847), .ZN(n3679) );
  NAND2_X1 U33480 ( .A1(n2998), .A2(n3679), .ZN(n2849) );
  NAND2_X1 U33490 ( .A1(n3075), .A2(REG1_REG_13__SCAN_IN), .ZN(n2848) );
  INV_X1 U33500 ( .A(n3962), .ZN(n3456) );
  NAND2_X1 U33510 ( .A1(n2887), .A2(REG0_REG_9__SCAN_IN), .ZN(n2857) );
  NAND2_X1 U33520 ( .A1(n2879), .A2(REG2_REG_9__SCAN_IN), .ZN(n2856) );
  AND2_X1 U3353 ( .A1(n2908), .A2(n2852), .ZN(n2853) );
  NOR2_X1 U33540 ( .A1(n2915), .A2(n2853), .ZN(n3965) );
  NAND2_X1 U3355 ( .A1(n2874), .A2(n3965), .ZN(n2855) );
  NAND2_X1 U3356 ( .A1(n3075), .A2(REG1_REG_9__SCAN_IN), .ZN(n2854) );
  NAND2_X1 U3357 ( .A1(n2887), .A2(REG0_REG_6__SCAN_IN), .ZN(n2862) );
  NAND2_X1 U3358 ( .A1(n2879), .A2(REG2_REG_6__SCAN_IN), .ZN(n2861) );
  AND2_X1 U3359 ( .A1(n2892), .A2(n3349), .ZN(n2858) );
  NOR2_X1 U3360 ( .A1(n2899), .A2(n2858), .ZN(n4809) );
  NAND2_X1 U3361 ( .A1(n2874), .A2(n4809), .ZN(n2860) );
  NAND2_X1 U3362 ( .A1(n3075), .A2(REG1_REG_6__SCAN_IN), .ZN(n2859) );
  NAND4_X1 U3363 ( .A1(n2862), .A2(n2861), .A3(n2860), .A4(n2859), .ZN(n4185)
         );
  INV_X1 U3364 ( .A(n4185), .ZN(n4835) );
  NAND2_X1 U3365 ( .A1(n2887), .A2(REG0_REG_4__SCAN_IN), .ZN(n2867) );
  NAND2_X1 U3366 ( .A1(n2879), .A2(REG2_REG_4__SCAN_IN), .ZN(n2866) );
  NOR2_X1 U3367 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2863) );
  NOR2_X1 U3368 ( .A1(n2893), .A2(n2863), .ZN(n3954) );
  NAND2_X1 U3369 ( .A1(n2874), .A2(n3954), .ZN(n2865) );
  NAND2_X1 U3370 ( .A1(n2881), .A2(REG1_REG_4__SCAN_IN), .ZN(n2864) );
  NAND2_X1 U3371 ( .A1(n2879), .A2(REG2_REG_1__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3372 ( .A1(n2874), .A2(REG3_REG_1__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U3373 ( .A1(n2880), .A2(REG0_REG_0__SCAN_IN), .ZN(n2873) );
  NAND2_X1 U3374 ( .A1(n2881), .A2(REG1_REG_0__SCAN_IN), .ZN(n2872) );
  AND2_X1 U3375 ( .A1(n4190), .A2(n3364), .ZN(n3354) );
  INV_X1 U3376 ( .A(n3359), .ZN(n3365) );
  AND2_X1 U3377 ( .A1(n3365), .A2(n3194), .ZN(n2878) );
  NAND2_X1 U3378 ( .A1(n2879), .A2(REG2_REG_2__SCAN_IN), .ZN(n2884) );
  NAND2_X1 U3379 ( .A1(n2880), .A2(REG0_REG_2__SCAN_IN), .ZN(n2883) );
  NAND2_X1 U3380 ( .A1(n2881), .A2(REG1_REG_2__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3381 ( .A1(n2874), .A2(REG3_REG_2__SCAN_IN), .ZN(n2885) );
  NAND2_X1 U3382 ( .A1(n4188), .A2(n3256), .ZN(n4074) );
  NAND2_X1 U3383 ( .A1(n3253), .A2(n4120), .ZN(n3255) );
  OR2_X1 U3384 ( .A1(n4188), .A2(n3737), .ZN(n2886) );
  NAND2_X1 U3385 ( .A1(n3255), .A2(n2886), .ZN(n3321) );
  NAND2_X1 U3386 ( .A1(n2887), .A2(REG0_REG_3__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3387 ( .A1(n2879), .A2(REG2_REG_3__SCAN_IN), .ZN(n2890) );
  NAND2_X1 U3388 ( .A1(n2874), .A2(n4793), .ZN(n2889) );
  NAND2_X1 U3389 ( .A1(n3075), .A2(REG1_REG_3__SCAN_IN), .ZN(n2888) );
  XNOR2_X1 U3390 ( .A(n4187), .B(n3304), .ZN(n4150) );
  NAND2_X1 U3391 ( .A1(n2887), .A2(REG0_REG_5__SCAN_IN), .ZN(n2897) );
  NAND2_X1 U3392 ( .A1(n2879), .A2(REG2_REG_5__SCAN_IN), .ZN(n2896) );
  OAI21_X1 U3393 ( .B1(n2893), .B2(REG3_REG_5__SCAN_IN), .A(n2892), .ZN(n3440)
         );
  INV_X1 U3394 ( .A(n3440), .ZN(n3317) );
  NAND2_X1 U3395 ( .A1(n2874), .A2(n3317), .ZN(n2895) );
  NAND2_X1 U3396 ( .A1(n3075), .A2(REG1_REG_5__SCAN_IN), .ZN(n2894) );
  NAND4_X1 U3397 ( .A1(n2897), .A2(n2896), .A3(n2895), .A4(n2894), .ZN(n4186)
         );
  NOR2_X1 U3398 ( .A1(n4186), .A2(n3438), .ZN(n2898) );
  INV_X1 U3399 ( .A(n4186), .ZN(n3390) );
  INV_X1 U3400 ( .A(n3438), .ZN(n3338) );
  NAND2_X1 U3401 ( .A1(n2887), .A2(REG0_REG_7__SCAN_IN), .ZN(n2904) );
  NAND2_X1 U3402 ( .A1(n2879), .A2(REG2_REG_7__SCAN_IN), .ZN(n2903) );
  OR2_X1 U3403 ( .A1(n2899), .A2(REG3_REG_7__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U3404 ( .A1(n2906), .A2(n2900), .ZN(n4844) );
  INV_X1 U3405 ( .A(n4844), .ZN(n3415) );
  NAND2_X1 U3406 ( .A1(n2874), .A2(n3415), .ZN(n2902) );
  NAND2_X1 U3407 ( .A1(n3075), .A2(REG1_REG_7__SCAN_IN), .ZN(n2901) );
  OR2_X1 U3408 ( .A1(n4184), .A2(n4832), .ZN(n4082) );
  NAND2_X1 U3409 ( .A1(n4184), .A2(n4832), .ZN(n4053) );
  NAND2_X1 U3410 ( .A1(n4082), .A2(n4053), .ZN(n4830) );
  NAND2_X1 U3411 ( .A1(n2887), .A2(REG0_REG_8__SCAN_IN), .ZN(n2912) );
  NAND2_X1 U3412 ( .A1(n2879), .A2(REG2_REG_8__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3413 ( .A1(n2906), .A2(n3431), .ZN(n2907) );
  AND2_X1 U3414 ( .A1(n2908), .A2(n2907), .ZN(n4858) );
  NAND2_X1 U3415 ( .A1(n2874), .A2(n4858), .ZN(n2910) );
  NAND2_X1 U3416 ( .A1(n3075), .A2(REG1_REG_8__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U3417 ( .A1(n3483), .A2(n3493), .ZN(n2913) );
  AOI21_X1 U3418 ( .B1(n3491), .B2(n2913), .A(n2284), .ZN(n3449) );
  OAI21_X1 U3419 ( .B1(n3540), .B2(n3962), .A(n3449), .ZN(n2914) );
  OAI21_X1 U3420 ( .B1(n3456), .B2(n4183), .A(n2914), .ZN(n3537) );
  NAND2_X1 U3421 ( .A1(n2887), .A2(REG0_REG_10__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3422 ( .A1(n2879), .A2(REG2_REG_10__SCAN_IN), .ZN(n2919) );
  NOR2_X1 U3423 ( .A1(n2915), .A2(REG3_REG_10__SCAN_IN), .ZN(n2916) );
  NOR2_X1 U3424 ( .A1(n2921), .A2(n2916), .ZN(n4867) );
  NAND2_X1 U3425 ( .A1(n2874), .A2(n4867), .ZN(n2918) );
  NAND2_X1 U3426 ( .A1(n3075), .A2(REG1_REG_10__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U3427 ( .A1(n2887), .A2(REG0_REG_11__SCAN_IN), .ZN(n2926) );
  NAND2_X1 U3428 ( .A1(n2879), .A2(REG2_REG_11__SCAN_IN), .ZN(n2925) );
  OR2_X1 U3429 ( .A1(n2921), .A2(REG3_REG_11__SCAN_IN), .ZN(n2922) );
  NAND2_X1 U3430 ( .A1(n2928), .A2(n2922), .ZN(n4880) );
  INV_X1 U3431 ( .A(n4880), .ZN(n3523) );
  NAND2_X1 U3432 ( .A1(n2874), .A2(n3523), .ZN(n2924) );
  NAND2_X1 U3433 ( .A1(n3075), .A2(REG1_REG_11__SCAN_IN), .ZN(n2923) );
  OR2_X1 U3434 ( .A1(n4181), .A2(n3651), .ZN(n3552) );
  NAND2_X1 U3435 ( .A1(n4181), .A2(n3651), .ZN(n3554) );
  NAND2_X1 U3436 ( .A1(n3552), .A2(n3554), .ZN(n4121) );
  NAND2_X1 U3437 ( .A1(n2887), .A2(REG0_REG_12__SCAN_IN), .ZN(n2934) );
  NAND2_X1 U3438 ( .A1(n2879), .A2(REG2_REG_12__SCAN_IN), .ZN(n2933) );
  NAND2_X1 U3439 ( .A1(n2928), .A2(n3531), .ZN(n2929) );
  AND2_X1 U3440 ( .A1(n2930), .A2(n2929), .ZN(n3558) );
  NAND2_X1 U3441 ( .A1(n2998), .A2(n3558), .ZN(n2932) );
  NAND2_X1 U3442 ( .A1(n3075), .A2(REG1_REG_12__SCAN_IN), .ZN(n2931) );
  NAND2_X1 U3443 ( .A1(n4180), .A2(n3556), .ZN(n2935) );
  OAI21_X1 U3444 ( .B1(n3574), .B2(n4179), .A(n3665), .ZN(n3685) );
  NAND2_X1 U3445 ( .A1(n2887), .A2(REG0_REG_14__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3446 ( .A1(n2879), .A2(REG2_REG_14__SCAN_IN), .ZN(n2941) );
  AND2_X1 U3447 ( .A1(n2937), .A2(n2936), .ZN(n2938) );
  NOR2_X1 U3448 ( .A1(n2943), .A2(n2938), .ZN(n3692) );
  NAND2_X1 U3449 ( .A1(n2998), .A2(n3692), .ZN(n2940) );
  NAND2_X1 U3450 ( .A1(n3075), .A2(REG1_REG_14__SCAN_IN), .ZN(n2939) );
  NAND4_X1 U3451 ( .A1(n2942), .A2(n2941), .A3(n2940), .A4(n2939), .ZN(n4178)
         );
  NAND2_X1 U3452 ( .A1(n4178), .A2(n4583), .ZN(n4028) );
  NAND2_X1 U3453 ( .A1(n4027), .A2(n4028), .ZN(n4139) );
  INV_X1 U3454 ( .A(n4139), .ZN(n3059) );
  NAND2_X1 U3455 ( .A1(n2887), .A2(REG0_REG_15__SCAN_IN), .ZN(n2950) );
  NAND2_X1 U3456 ( .A1(n2879), .A2(REG2_REG_15__SCAN_IN), .ZN(n2949) );
  OR2_X1 U3457 ( .A1(n2943), .A2(REG3_REG_15__SCAN_IN), .ZN(n2944) );
  NAND2_X1 U34580 ( .A1(n2945), .A2(n2944), .ZN(n4911) );
  INV_X1 U34590 ( .A(n4911), .ZN(n2946) );
  NAND2_X1 U3460 ( .A1(n2998), .A2(n2946), .ZN(n2948) );
  NAND2_X1 U3461 ( .A1(n3075), .A2(REG1_REG_15__SCAN_IN), .ZN(n2947) );
  NAND4_X1 U3462 ( .A1(n2950), .A2(n2949), .A3(n2948), .A4(n2947), .ZN(n4177)
         );
  INV_X1 U3463 ( .A(n4177), .ZN(n4572) );
  NOR2_X1 U3464 ( .A1(n4572), .A2(n4901), .ZN(n2951) );
  INV_X1 U3465 ( .A(n4179), .ZN(n4584) );
  NOR2_X1 U3466 ( .A1(n4584), .A2(n3677), .ZN(n3686) );
  NOR3_X1 U34670 ( .A1(n3059), .A2(n2951), .A3(n3686), .ZN(n2953) );
  INV_X1 U3468 ( .A(n4583), .ZN(n3586) );
  OR2_X1 U34690 ( .A1(n4178), .A2(n3586), .ZN(n3720) );
  OAI22_X1 U3470 ( .A1(n2951), .A2(n3720), .B1(n3751), .B2(n4177), .ZN(n2952)
         );
  OR2_X1 U34710 ( .A1(n4176), .A2(n4571), .ZN(n4096) );
  NAND2_X1 U3472 ( .A1(n4176), .A2(n4571), .ZN(n4099) );
  NAND2_X1 U34730 ( .A1(n4096), .A2(n4099), .ZN(n4141) );
  NAND2_X1 U3474 ( .A1(n3624), .A2(n4141), .ZN(n3623) );
  OAI21_X1 U34750 ( .B1(n4898), .B2(n4571), .A(n3623), .ZN(n3699) );
  NAND2_X1 U3476 ( .A1(n2887), .A2(REG0_REG_17__SCAN_IN), .ZN(n2959) );
  NAND2_X1 U34770 ( .A1(n2879), .A2(REG2_REG_17__SCAN_IN), .ZN(n2958) );
  NOR2_X1 U3478 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2954), .ZN(n2955) );
  NOR2_X1 U34790 ( .A1(n2962), .A2(n2955), .ZN(n3932) );
  NAND2_X1 U3480 ( .A1(n2998), .A2(n3932), .ZN(n2957) );
  NAND2_X1 U34810 ( .A1(n3075), .A2(REG1_REG_17__SCAN_IN), .ZN(n2956) );
  NAND4_X1 U3482 ( .A1(n2959), .A2(n2958), .A3(n2957), .A4(n2956), .ZN(n4175)
         );
  NAND2_X1 U34830 ( .A1(n4491), .A2(n4566), .ZN(n2961) );
  NOR2_X1 U3484 ( .A1(n4491), .A2(n4566), .ZN(n2960) );
  NAND2_X1 U34850 ( .A1(n2887), .A2(REG0_REG_18__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3486 ( .A1(n2879), .A2(REG2_REG_18__SCAN_IN), .ZN(n2965) );
  OAI21_X1 U34870 ( .B1(n2962), .B2(REG3_REG_18__SCAN_IN), .A(n2968), .ZN(
        n4497) );
  INV_X1 U3488 ( .A(n4497), .ZN(n3999) );
  NAND2_X1 U34890 ( .A1(n2998), .A2(n3999), .ZN(n2964) );
  NAND2_X1 U3490 ( .A1(n3075), .A2(REG1_REG_18__SCAN_IN), .ZN(n2963) );
  NAND4_X1 U34910 ( .A1(n2966), .A2(n2965), .A3(n2964), .A4(n2963), .ZN(n4174)
         );
  OR2_X1 U3492 ( .A1(n4174), .A2(n4490), .ZN(n4469) );
  NAND2_X1 U34930 ( .A1(n4174), .A2(n4490), .ZN(n4470) );
  NAND2_X1 U3494 ( .A1(n4469), .A2(n4470), .ZN(n4499) );
  NAND2_X1 U34950 ( .A1(n4500), .A2(n4499), .ZN(n4498) );
  INV_X1 U3496 ( .A(n4174), .ZN(n4474) );
  NAND2_X1 U34970 ( .A1(n4474), .A2(n4490), .ZN(n2967) );
  NAND2_X1 U3498 ( .A1(n4498), .A2(n2967), .ZN(n4464) );
  NAND2_X1 U34990 ( .A1(n2887), .A2(REG0_REG_19__SCAN_IN), .ZN(n2973) );
  NAND2_X1 U3500 ( .A1(n2879), .A2(REG2_REG_19__SCAN_IN), .ZN(n2972) );
  AND2_X1 U35010 ( .A1(n2968), .A2(n3889), .ZN(n2969) );
  NOR2_X1 U3502 ( .A1(n2975), .A2(n2969), .ZN(n4482) );
  NAND2_X1 U35030 ( .A1(n2998), .A2(n4482), .ZN(n2971) );
  NAND2_X1 U3504 ( .A1(n3075), .A2(REG1_REG_19__SCAN_IN), .ZN(n2970) );
  NAND4_X1 U35050 ( .A1(n2973), .A2(n2972), .A3(n2971), .A4(n2970), .ZN(n4496)
         );
  NAND2_X1 U35060 ( .A1(n4496), .A2(n3783), .ZN(n2974) );
  INV_X1 U35070 ( .A(n4496), .ZN(n4447) );
  AOI22_X1 U35080 ( .A1(n4464), .A2(n2974), .B1(n4447), .B2(n4480), .ZN(n4438)
         );
  INV_X1 U35090 ( .A(n4438), .ZN(n2983) );
  NAND2_X1 U35100 ( .A1(n2887), .A2(REG0_REG_20__SCAN_IN), .ZN(n2980) );
  NAND2_X1 U35110 ( .A1(n2879), .A2(REG2_REG_20__SCAN_IN), .ZN(n2979) );
  NAND2_X1 U35120 ( .A1(n2975), .A2(REG3_REG_20__SCAN_IN), .ZN(n2984) );
  OR2_X1 U35130 ( .A1(n2975), .A2(REG3_REG_20__SCAN_IN), .ZN(n2976) );
  AND2_X1 U35140 ( .A1(n2984), .A2(n2976), .ZN(n4458) );
  NAND2_X1 U35150 ( .A1(n2998), .A2(n4458), .ZN(n2978) );
  NAND2_X1 U35160 ( .A1(n3075), .A2(REG1_REG_20__SCAN_IN), .ZN(n2977) );
  NAND2_X1 U35170 ( .A1(n4547), .A2(n4444), .ZN(n2981) );
  OAI21_X2 U35180 ( .B1(n2983), .B2(n2982), .A(n2981), .ZN(n4420) );
  NAND2_X1 U35190 ( .A1(n2887), .A2(REG0_REG_21__SCAN_IN), .ZN(n2989) );
  NAND2_X1 U35200 ( .A1(n2879), .A2(REG2_REG_21__SCAN_IN), .ZN(n2988) );
  NAND2_X1 U35210 ( .A1(n2984), .A2(n2805), .ZN(n2985) );
  AND2_X1 U35220 ( .A1(n2990), .A2(n2985), .ZN(n4429) );
  NAND2_X1 U35230 ( .A1(n2998), .A2(n4429), .ZN(n2987) );
  NAND2_X1 U35240 ( .A1(n3075), .A2(REG1_REG_21__SCAN_IN), .ZN(n2986) );
  NAND4_X1 U35250 ( .A1(n2989), .A2(n2988), .A3(n2987), .A4(n2986), .ZN(n4445)
         );
  INV_X1 U35260 ( .A(n4548), .ZN(n3800) );
  AND2_X1 U35270 ( .A1(n4445), .A2(n3800), .ZN(n4376) );
  NAND2_X1 U35280 ( .A1(n2879), .A2(REG2_REG_22__SCAN_IN), .ZN(n2995) );
  NAND2_X1 U35290 ( .A1(n3075), .A2(REG1_REG_22__SCAN_IN), .ZN(n2994) );
  INV_X1 U35300 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U35310 ( .A1(n2990), .A2(n3983), .ZN(n2991) );
  NAND2_X1 U35320 ( .A1(n2996), .A2(n2991), .ZN(n4411) );
  INV_X1 U35330 ( .A(n4411), .ZN(n3987) );
  NAND2_X1 U35340 ( .A1(n2998), .A2(n3987), .ZN(n2993) );
  NAND2_X1 U35350 ( .A1(n2887), .A2(REG0_REG_22__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U35360 ( .A1(n4425), .A2(n4415), .ZN(n3066) );
  NAND2_X1 U35370 ( .A1(n4385), .A2(n3066), .ZN(n4403) );
  INV_X1 U35380 ( .A(n4445), .ZN(n3984) );
  NAND2_X1 U35390 ( .A1(n3984), .A2(n4548), .ZN(n4377) );
  INV_X1 U35400 ( .A(n4415), .ZN(n3811) );
  NAND2_X1 U35410 ( .A1(n4425), .A2(n3811), .ZN(n4379) );
  NAND2_X1 U35420 ( .A1(n2887), .A2(REG0_REG_23__SCAN_IN), .ZN(n3002) );
  NAND2_X1 U35430 ( .A1(n2879), .A2(REG2_REG_23__SCAN_IN), .ZN(n3001) );
  INV_X1 U35440 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3881) );
  AND2_X1 U35450 ( .A1(n2996), .A2(n3881), .ZN(n2997) );
  NOR2_X1 U35460 ( .A1(n3004), .A2(n2997), .ZN(n4396) );
  NAND2_X1 U35470 ( .A1(n2998), .A2(n4396), .ZN(n3000) );
  NAND2_X1 U35480 ( .A1(n3075), .A2(REG1_REG_23__SCAN_IN), .ZN(n2999) );
  NOR2_X1 U35490 ( .A1(n4405), .A2(n4388), .ZN(n3003) );
  NOR2_X1 U35500 ( .A1(n4362), .A2(n4395), .ZN(n4357) );
  NAND2_X1 U35510 ( .A1(n2887), .A2(REG0_REG_24__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U35520 ( .A1(n2879), .A2(REG2_REG_24__SCAN_IN), .ZN(n3008) );
  NOR2_X1 U35530 ( .A1(n3004), .A2(REG3_REG_24__SCAN_IN), .ZN(n3005) );
  OR2_X1 U35540 ( .A1(n3016), .A2(n3005), .ZN(n4370) );
  NAND2_X1 U35550 ( .A1(n2998), .A2(n3942), .ZN(n3007) );
  NAND2_X1 U35560 ( .A1(n3075), .A2(REG1_REG_24__SCAN_IN), .ZN(n3006) );
  NAND4_X1 U35570 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n4389)
         );
  INV_X1 U35580 ( .A(n4389), .ZN(n4345) );
  NOR2_X1 U35590 ( .A1(n4345), .A2(n4369), .ZN(n3010) );
  OR2_X1 U35600 ( .A1(n4357), .A2(n3010), .ZN(n4337) );
  NAND2_X1 U35610 ( .A1(n2879), .A2(REG2_REG_25__SCAN_IN), .ZN(n3014) );
  NAND2_X1 U35620 ( .A1(n3075), .A2(REG1_REG_25__SCAN_IN), .ZN(n3013) );
  XNOR2_X1 U35630 ( .A(n3016), .B(n3908), .ZN(n4352) );
  NAND2_X1 U35640 ( .A1(n2998), .A2(n4352), .ZN(n3012) );
  NAND2_X1 U35650 ( .A1(n2887), .A2(REG0_REG_25__SCAN_IN), .ZN(n3011) );
  INV_X1 U35660 ( .A(n4350), .ZN(n3839) );
  AND2_X1 U35670 ( .A1(n4364), .A2(n3839), .ZN(n3024) );
  NAND2_X1 U35680 ( .A1(n2887), .A2(REG0_REG_26__SCAN_IN), .ZN(n3021) );
  NAND2_X1 U35690 ( .A1(n2879), .A2(REG2_REG_26__SCAN_IN), .ZN(n3020) );
  AND2_X1 U35700 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n3015) );
  AOI21_X1 U35710 ( .B1(n3016), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n3017) );
  NOR2_X1 U35720 ( .A1(n3027), .A2(n3017), .ZN(n4330) );
  NAND2_X1 U35730 ( .A1(n2998), .A2(n4330), .ZN(n3019) );
  NAND2_X1 U35740 ( .A1(n3075), .A2(REG1_REG_26__SCAN_IN), .ZN(n3018) );
  NOR2_X1 U35750 ( .A1(n4518), .A2(n4524), .ZN(n3025) );
  OR2_X1 U35760 ( .A1(n4314), .A2(n3025), .ZN(n3026) );
  OR2_X1 U35770 ( .A1(n4364), .A2(n3839), .ZN(n3022) );
  NAND2_X1 U35780 ( .A1(n4345), .A2(n4369), .ZN(n4338) );
  AND2_X1 U35790 ( .A1(n3022), .A2(n4338), .ZN(n3023) );
  NAND2_X1 U35800 ( .A1(n2879), .A2(REG2_REG_27__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U35810 ( .A1(n3075), .A2(REG1_REG_27__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U3582 ( .A1(n3027), .A2(REG3_REG_27__SCAN_IN), .ZN(n3034) );
  OR2_X1 U3583 ( .A1(n3027), .A2(REG3_REG_27__SCAN_IN), .ZN(n3028) );
  NAND2_X1 U3584 ( .A1(n2998), .A2(n4302), .ZN(n3030) );
  NAND2_X1 U3585 ( .A1(n2887), .A2(REG0_REG_27__SCAN_IN), .ZN(n3029) );
  NOR2_X1 U3586 ( .A1(n4324), .A2(n3845), .ZN(n3033) );
  INV_X1 U3587 ( .A(n4324), .ZN(n4011) );
  NAND2_X1 U3588 ( .A1(n2879), .A2(REG2_REG_28__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U3589 ( .A1(n2887), .A2(REG0_REG_28__SCAN_IN), .ZN(n3038) );
  INV_X1 U3590 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U3591 ( .A1(n3034), .A2(n3861), .ZN(n3035) );
  NAND2_X1 U3592 ( .A1(n2998), .A2(n4283), .ZN(n3037) );
  NAND2_X1 U3593 ( .A1(n3075), .A2(REG1_REG_28__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3594 ( .A1(n4299), .A2(n4288), .ZN(n4020) );
  NAND2_X1 U3595 ( .A1(n4019), .A2(n4020), .ZN(n4289) );
  AOI22_X1 U3596 ( .A1(n4282), .A2(n4289), .B1(n3853), .B2(n4299), .ZN(n3045)
         );
  NAND2_X1 U3597 ( .A1(n2887), .A2(REG0_REG_29__SCAN_IN), .ZN(n3044) );
  NAND2_X1 U3598 ( .A1(n2879), .A2(REG2_REG_29__SCAN_IN), .ZN(n3043) );
  INV_X1 U3599 ( .A(n4275), .ZN(n3040) );
  NAND2_X1 U3600 ( .A1(n2998), .A2(n3040), .ZN(n3042) );
  NAND2_X1 U3601 ( .A1(n3075), .A2(REG1_REG_29__SCAN_IN), .ZN(n3041) );
  NAND4_X1 U3602 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n4292)
         );
  XNOR2_X1 U3603 ( .A(n4292), .B(n4280), .ZN(n4152) );
  XNOR2_X1 U3604 ( .A(n3045), .B(n4152), .ZN(n4281) );
  NAND2_X2 U3605 ( .A1(n3046), .A2(n4157), .ZN(n3184) );
  XNOR2_X1 U3606 ( .A(n3184), .B(n4651), .ZN(n3047) );
  NAND2_X1 U3607 ( .A1(n3047), .A2(n4766), .ZN(n4452) );
  NAND2_X1 U3608 ( .A1(n4281), .A2(n4587), .ZN(n3083) );
  INV_X1 U3609 ( .A(n3121), .ZN(n3170) );
  NOR2_X1 U3610 ( .A1(n4916), .A2(n3170), .ZN(n4406) );
  NOR2_X1 U3611 ( .A1(n4280), .A2(n4833), .ZN(n3081) );
  OR2_X1 U3612 ( .A1(n4190), .A2(n3166), .ZN(n3153) );
  INV_X1 U3613 ( .A(n3153), .ZN(n4069) );
  NAND2_X1 U3614 ( .A1(n3356), .A2(n4069), .ZN(n3355) );
  NAND2_X1 U3615 ( .A1(n3355), .A2(n4070), .ZN(n3049) );
  INV_X1 U3616 ( .A(n4120), .ZN(n3048) );
  NAND2_X1 U3617 ( .A1(n3049), .A2(n3048), .ZN(n3259) );
  NAND2_X1 U3618 ( .A1(n3259), .A2(n4071), .ZN(n3322) );
  OR2_X1 U3619 ( .A1(n2433), .A2(n3325), .ZN(n3375) );
  NAND2_X1 U3620 ( .A1(n2433), .A2(n3325), .ZN(n4073) );
  NAND2_X1 U3621 ( .A1(n3375), .A2(n4073), .ZN(n4125) );
  INV_X1 U3622 ( .A(n4125), .ZN(n3323) );
  NAND2_X1 U3623 ( .A1(n3322), .A2(n3323), .ZN(n3376) );
  INV_X1 U3624 ( .A(n3304), .ZN(n3951) );
  OR2_X1 U3625 ( .A1(n4187), .A2(n3951), .ZN(n3050) );
  AND2_X1 U3626 ( .A1(n3375), .A2(n3050), .ZN(n4076) );
  NAND2_X1 U3627 ( .A1(n3376), .A2(n4076), .ZN(n3051) );
  NAND2_X1 U3628 ( .A1(n4187), .A2(n3951), .ZN(n4078) );
  OR2_X1 U3629 ( .A1(n4186), .A2(n3338), .ZN(n4055) );
  NAND2_X1 U3630 ( .A1(n3052), .A2(n4055), .ZN(n3389) );
  NAND2_X1 U3631 ( .A1(n4185), .A2(n3396), .ZN(n4079) );
  OR2_X1 U3632 ( .A1(n4185), .A2(n3396), .ZN(n4081) );
  INV_X1 U3633 ( .A(n4082), .ZN(n3053) );
  OR2_X1 U3634 ( .A1(n4837), .A2(n3493), .ZN(n4085) );
  NAND2_X1 U3635 ( .A1(n3492), .A2(n4085), .ZN(n3054) );
  NAND2_X1 U3636 ( .A1(n4837), .A2(n3493), .ZN(n4052) );
  AND2_X1 U3637 ( .A1(n4183), .A2(n3962), .ZN(n4084) );
  OR2_X1 U3638 ( .A1(n4183), .A2(n3962), .ZN(n4086) );
  NAND2_X1 U3639 ( .A1(n4182), .A2(n3539), .ZN(n4060) );
  OR2_X1 U3640 ( .A1(n4182), .A2(n3539), .ZN(n4057) );
  NAND2_X1 U3641 ( .A1(n4180), .A2(n3635), .ZN(n3667) );
  NAND2_X1 U3642 ( .A1(n4179), .A2(n3677), .ZN(n3662) );
  AND2_X1 U3643 ( .A1(n3667), .A2(n3662), .ZN(n3057) );
  AND2_X1 U3644 ( .A1(n3057), .A2(n3554), .ZN(n4061) );
  NAND2_X1 U3645 ( .A1(n3649), .A2(n4061), .ZN(n3058) );
  OR2_X1 U3646 ( .A1(n4180), .A2(n3635), .ZN(n3669) );
  NAND2_X1 U3647 ( .A1(n3552), .A2(n3669), .ZN(n3056) );
  NOR2_X1 U3648 ( .A1(n4179), .A2(n3677), .ZN(n3664) );
  AOI21_X1 U3649 ( .B1(n3057), .B2(n3056), .A(n3664), .ZN(n4063) );
  NAND2_X1 U3650 ( .A1(n3058), .A2(n4063), .ZN(n4032) );
  OR2_X1 U3651 ( .A1(n4177), .A2(n4901), .ZN(n4030) );
  NAND2_X1 U3652 ( .A1(n4177), .A2(n4901), .ZN(n4029) );
  NAND2_X1 U3653 ( .A1(n4030), .A2(n4029), .ZN(n4140) );
  INV_X1 U3654 ( .A(n4141), .ZN(n3630) );
  NAND2_X1 U3655 ( .A1(n4496), .A2(n4480), .ZN(n3060) );
  AND2_X1 U3656 ( .A1(n4470), .A2(n3060), .ZN(n3063) );
  NAND2_X1 U3657 ( .A1(n4175), .A2(n4566), .ZN(n4465) );
  NAND2_X1 U3658 ( .A1(n3063), .A2(n4465), .ZN(n4035) );
  NAND2_X1 U3659 ( .A1(n4547), .A2(n4456), .ZN(n4123) );
  INV_X1 U3660 ( .A(n4123), .ZN(n4034) );
  OR2_X1 U3661 ( .A1(n4175), .A2(n4566), .ZN(n4466) );
  NAND2_X1 U3662 ( .A1(n4469), .A2(n4466), .ZN(n3062) );
  NOR2_X1 U3663 ( .A1(n4496), .A2(n4480), .ZN(n3061) );
  AOI21_X1 U3664 ( .B1(n3063), .B2(n3062), .A(n3061), .ZN(n4439) );
  OR2_X1 U3665 ( .A1(n4547), .A2(n4456), .ZN(n4124) );
  NAND2_X1 U3666 ( .A1(n4439), .A2(n4124), .ZN(n3064) );
  NAND2_X1 U3667 ( .A1(n3064), .A2(n4123), .ZN(n4100) );
  OR2_X1 U3668 ( .A1(n4445), .A2(n4548), .ZN(n4382) );
  NAND2_X1 U3669 ( .A1(n4385), .A2(n4382), .ZN(n4103) );
  NAND2_X1 U3670 ( .A1(n4405), .A2(n4395), .ZN(n3065) );
  NAND2_X1 U3671 ( .A1(n3066), .A2(n3065), .ZN(n4107) );
  INV_X1 U3672 ( .A(n4107), .ZN(n3069) );
  NAND2_X1 U3673 ( .A1(n4445), .A2(n4548), .ZN(n4384) );
  INV_X1 U3674 ( .A(n4384), .ZN(n3067) );
  NAND2_X1 U3675 ( .A1(n3067), .A2(n4385), .ZN(n3068) );
  OR2_X1 U3676 ( .A1(n4405), .A2(n4395), .ZN(n4025) );
  NAND2_X1 U3677 ( .A1(n3070), .A2(n4025), .ZN(n4361) );
  NOR2_X1 U3678 ( .A1(n4389), .A2(n4369), .ZN(n4130) );
  NAND2_X1 U3679 ( .A1(n4389), .A2(n4369), .ZN(n4341) );
  NAND2_X1 U3680 ( .A1(n4364), .A2(n4350), .ZN(n4131) );
  OR2_X1 U3681 ( .A1(n4364), .A2(n4350), .ZN(n4319) );
  OR2_X1 U3682 ( .A1(n4347), .A2(n4524), .ZN(n4149) );
  NAND2_X1 U3683 ( .A1(n4319), .A2(n4149), .ZN(n4041) );
  INV_X1 U3684 ( .A(n4041), .ZN(n4112) );
  NAND2_X1 U3685 ( .A1(n4324), .A2(n4517), .ZN(n4113) );
  NAND2_X1 U3686 ( .A1(n4018), .A2(n4113), .ZN(n4303) );
  INV_X1 U3687 ( .A(n4019), .ZN(n3071) );
  AOI21_X1 U3688 ( .B1(n4290), .B2(n4020), .A(n3071), .ZN(n3073) );
  INV_X1 U3689 ( .A(n4152), .ZN(n3072) );
  XNOR2_X1 U3690 ( .A(n3073), .B(n3072), .ZN(n3080) );
  NAND2_X1 U3691 ( .A1(n4652), .A2(n4157), .ZN(n4051) );
  NAND2_X1 U3692 ( .A1(n4829), .A2(n4651), .ZN(n3074) );
  NAND2_X1 U3693 ( .A1(n3075), .A2(REG1_REG_30__SCAN_IN), .ZN(n3078) );
  NAND2_X1 U3694 ( .A1(n2879), .A2(REG2_REG_30__SCAN_IN), .ZN(n3077) );
  NAND2_X1 U3695 ( .A1(n2887), .A2(REG0_REG_30__SCAN_IN), .ZN(n3076) );
  AND3_X1 U3696 ( .A1(n3078), .A2(n3077), .A3(n3076), .ZN(n4022) );
  OAI22_X1 U3697 ( .A1(n3080), .A2(n4840), .B1(n4022), .B2(n3079), .ZN(n4278)
         );
  NAND2_X1 U3698 ( .A1(n3083), .A2(n3082), .ZN(n3100) );
  NOR2_X1 U3699 ( .A1(n4786), .A2(n4157), .ZN(n3085) );
  NOR2_X1 U3700 ( .A1(n3085), .A2(n3084), .ZN(n3088) );
  NAND2_X1 U3701 ( .A1(n3156), .A2(n3123), .ZN(n3086) );
  AND2_X2 U3702 ( .A1(n3096), .A2(n3157), .ZN(n4852) );
  NAND2_X1 U3703 ( .A1(n4852), .A2(n3093), .ZN(n4591) );
  NAND2_X1 U3704 ( .A1(n3094), .A2(n2501), .ZN(U3547) );
  AND2_X2 U3705 ( .A1(n3096), .A2(n3095), .ZN(n4855) );
  INV_X1 U3706 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3707 ( .A1(n3099), .A2(n3097), .ZN(n3098) );
  OAI21_X1 U3708 ( .B1(n3100), .B2(n3099), .A(n3098), .ZN(n3101) );
  NAND2_X1 U3709 ( .A1(n3101), .A2(n2500), .ZN(U3515) );
  INV_X1 U3710 ( .A(n3102), .ZN(n4166) );
  OR2_X2 U3711 ( .A1(n3163), .A2(n4166), .ZN(n4189) );
  INV_X1 U3712 ( .A(n4189), .ZN(U4043) );
  NAND2_X1 U3713 ( .A1(n4157), .A2(STATE_REG_SCAN_IN), .ZN(n3103) );
  OAI21_X1 U3714 ( .B1(STATE_REG_SCAN_IN), .B2(n3104), .A(n3103), .ZN(U3331)
         );
  INV_X1 U3715 ( .A(n4232), .ZN(n4223) );
  NAND2_X1 U3716 ( .A1(n4223), .A2(STATE_REG_SCAN_IN), .ZN(n3105) );
  OAI21_X1 U3717 ( .B1(STATE_REG_SCAN_IN), .B2(n2564), .A(n3105), .ZN(U3337)
         );
  NAND2_X1 U3718 ( .A1(n3106), .A2(STATE_REG_SCAN_IN), .ZN(n3107) );
  OAI21_X1 U3719 ( .B1(STATE_REG_SCAN_IN), .B2(n3108), .A(n3107), .ZN(U3327)
         );
  NAND2_X1 U3720 ( .A1(n2626), .A2(STATE_REG_SCAN_IN), .ZN(n3109) );
  OAI21_X1 U3721 ( .B1(STATE_REG_SCAN_IN), .B2(n3110), .A(n3109), .ZN(U3323)
         );
  INV_X1 U3722 ( .A(n4168), .ZN(n3128) );
  NAND2_X1 U3723 ( .A1(n3128), .A2(STATE_REG_SCAN_IN), .ZN(n3111) );
  OAI21_X1 U3724 ( .B1(STATE_REG_SCAN_IN), .B2(n3112), .A(n3111), .ZN(U3325)
         );
  INV_X1 U3725 ( .A(DATAI_31_), .ZN(n3115) );
  OR4_X1 U3726 ( .A1(n2390), .A2(IR_REG_30__SCAN_IN), .A3(n3113), .A4(U3149), 
        .ZN(n3114) );
  OAI21_X1 U3727 ( .B1(STATE_REG_SCAN_IN), .B2(n3115), .A(n3114), .ZN(U3321)
         );
  INV_X1 U3728 ( .A(n3116), .ZN(n3117) );
  NOR3_X1 U3729 ( .A1(n4166), .A2(n4649), .A3(n4650), .ZN(n3118) );
  AOI21_X1 U3730 ( .B1(n4658), .B2(n3119), .A(n3118), .ZN(U3458) );
  OR2_X1 U3731 ( .A1(n3244), .A2(U3149), .ZN(n4656) );
  INV_X1 U3732 ( .A(n4656), .ZN(n3120) );
  OR2_X1 U3733 ( .A1(n3159), .A2(n3120), .ZN(n3131) );
  NAND2_X1 U3734 ( .A1(n3244), .A2(n3121), .ZN(n3122) );
  NAND2_X1 U3735 ( .A1(n2271), .A2(n3122), .ZN(n3130) );
  NOR2_X1 U3736 ( .A1(n4764), .A2(U4043), .ZN(U3148) );
  INV_X1 U3737 ( .A(n4658), .ZN(n3125) );
  NAND2_X1 U3738 ( .A1(n3125), .A2(n3123), .ZN(n3124) );
  OAI21_X1 U3739 ( .B1(n3125), .B2(n2615), .A(n3124), .ZN(U3459) );
  NAND2_X1 U3740 ( .A1(n4189), .A2(DATAO_REG_30__SCAN_IN), .ZN(n3126) );
  OAI21_X1 U3741 ( .B1(n4022), .B2(n4189), .A(n3126), .ZN(U3580) );
  NOR2_X1 U3742 ( .A1(n4168), .A2(REG2_REG_0__SCAN_IN), .ZN(n3127) );
  NOR2_X1 U3743 ( .A1(n4916), .A2(n3127), .ZN(n3231) );
  OAI21_X1 U3744 ( .B1(REG1_REG_0__SCAN_IN), .B2(n3128), .A(n3231), .ZN(n3129)
         );
  MUX2_X1 U3745 ( .A(n3231), .B(n3129), .S(n4774), .Z(n3136) );
  INV_X1 U3746 ( .A(n3130), .ZN(n3132) );
  INV_X1 U3747 ( .A(n3146), .ZN(n3135) );
  AOI22_X1 U3748 ( .A1(n4764), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3134) );
  INV_X1 U3749 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3167) );
  NAND3_X1 U3750 ( .A1(n4769), .A2(IR_REG_0__SCAN_IN), .A3(n3167), .ZN(n3133)
         );
  OAI211_X1 U3751 ( .C1(n3136), .C2(n3135), .A(n3134), .B(n3133), .ZN(U3240)
         );
  AND2_X1 U3752 ( .A1(n3146), .A2(n4916), .ZN(n4682) );
  INV_X1 U3753 ( .A(n4682), .ZN(n4767) );
  INV_X1 U3754 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3137) );
  INV_X1 U3755 ( .A(n4207), .ZN(n3140) );
  NAND2_X1 U3756 ( .A1(n2524), .A2(REG1_REG_1__SCAN_IN), .ZN(n3139) );
  INV_X1 U3757 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U3758 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n4195) );
  AOI21_X1 U3759 ( .B1(n4194), .B2(n4790), .A(n4195), .ZN(n3138) );
  NAND2_X1 U3760 ( .A1(n3139), .A2(n3138), .ZN(n4198) );
  NAND2_X1 U3761 ( .A1(n4198), .A2(n3139), .ZN(n4206) );
  XNOR2_X1 U3762 ( .A(n3223), .B(n3222), .ZN(n3225) );
  XNOR2_X1 U3763 ( .A(n3225), .B(REG1_REG_3__SCAN_IN), .ZN(n3150) );
  INV_X1 U3764 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3148) );
  INV_X1 U3765 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3142) );
  MUX2_X1 U3766 ( .A(n3142), .B(REG2_REG_2__SCAN_IN), .S(n3143), .Z(n4205) );
  AND2_X1 U3767 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4192)
         );
  NAND2_X1 U3768 ( .A1(n2524), .A2(REG2_REG_1__SCAN_IN), .ZN(n3141) );
  OAI21_X1 U3769 ( .B1(n3143), .B2(n3142), .A(n4203), .ZN(n3220) );
  NOR2_X1 U3770 ( .A1(n3147), .A2(n3148), .ZN(n3219) );
  NOR2_X1 U3771 ( .A1(n4916), .A2(n4168), .ZN(n3145) );
  AOI211_X1 U3772 ( .C1(n3148), .C2(n3147), .A(n3219), .B(n4771), .ZN(n3149)
         );
  AOI21_X1 U3773 ( .B1(n4769), .B2(n3150), .A(n3149), .ZN(n3152) );
  NOR2_X1 U3774 ( .A1(STATE_REG_SCAN_IN), .A2(n4793), .ZN(n3249) );
  AOI21_X1 U3775 ( .B1(n4764), .B2(ADDR_REG_3__SCAN_IN), .A(n3249), .ZN(n3151)
         );
  OAI211_X1 U3776 ( .C1(n3222), .C2(n4767), .A(n3152), .B(n3151), .ZN(U3243)
         );
  INV_X1 U3777 ( .A(n4786), .ZN(n4802) );
  NAND2_X1 U3778 ( .A1(n4190), .A2(n3166), .ZN(n4068) );
  NAND2_X1 U3779 ( .A1(n3153), .A2(n4068), .ZN(n4781) );
  AND2_X1 U3780 ( .A1(n3364), .A2(n3175), .ZN(n4780) );
  INV_X1 U3781 ( .A(n3194), .ZN(n3257) );
  INV_X1 U3782 ( .A(n4838), .ZN(n3689) );
  INV_X1 U3783 ( .A(n4452), .ZN(n3650) );
  OAI21_X1 U3784 ( .B1(n3650), .B2(n4449), .A(n4781), .ZN(n3154) );
  OAI21_X1 U3785 ( .B1(n3257), .B2(n3689), .A(n3154), .ZN(n4778) );
  AOI211_X1 U3786 ( .C1(n4802), .C2(n4781), .A(n4780), .B(n4778), .ZN(n4776)
         );
  NAND2_X1 U3787 ( .A1(n3091), .A2(REG1_REG_0__SCAN_IN), .ZN(n3155) );
  OAI21_X1 U3788 ( .B1(n4776), .B2(n3091), .A(n3155), .ZN(U3518) );
  INV_X1 U3789 ( .A(n3159), .ZN(n3160) );
  NOR2_X1 U3790 ( .A1(n3176), .A2(n3160), .ZN(n3180) );
  NAND2_X1 U3791 ( .A1(n4766), .A2(n4651), .ZN(n4167) );
  NOR2_X1 U3792 ( .A1(n3184), .A2(n4167), .ZN(n3161) );
  NAND2_X1 U3793 ( .A1(n3180), .A2(n3161), .ZN(n3195) );
  INV_X1 U3794 ( .A(n4916), .ZN(n3228) );
  NAND2_X1 U3795 ( .A1(n3209), .A2(n4190), .ZN(n3165) );
  NAND2_X1 U3796 ( .A1(n4190), .A2(n2274), .ZN(n3168) );
  NAND2_X1 U3797 ( .A1(n3364), .A2(n2287), .ZN(n3185) );
  NAND2_X1 U3798 ( .A1(n3168), .A2(n2497), .ZN(n3188) );
  XOR2_X1 U3799 ( .A(n3189), .B(n3188), .Z(n3227) );
  INV_X1 U3800 ( .A(n3180), .ZN(n3173) );
  NAND2_X1 U3801 ( .A1(n3169), .A2(n3175), .ZN(n3171) );
  NAND2_X1 U3802 ( .A1(n3171), .A2(n3170), .ZN(n3172) );
  INV_X1 U3803 ( .A(n4016), .ZN(n4907) );
  NAND2_X1 U3804 ( .A1(n3227), .A2(n4907), .ZN(n3183) );
  NOR3_X1 U3805 ( .A1(n3174), .A2(U3149), .A3(n4833), .ZN(n3246) );
  INV_X1 U3806 ( .A(n3246), .ZN(n3179) );
  INV_X1 U3807 ( .A(n3175), .ZN(n3177) );
  OAI21_X1 U3808 ( .B1(n3177), .B2(n4766), .A(n3176), .ZN(n3245) );
  NAND3_X1 U3809 ( .A1(n3179), .A2(n3178), .A3(n3245), .ZN(n3214) );
  NAND2_X1 U3810 ( .A1(n3180), .A2(n4443), .ZN(n3181) );
  NAND2_X1 U3811 ( .A1(n3181), .A2(n4879), .ZN(n3315) );
  AOI22_X1 U3812 ( .A1(n3214), .A2(REG3_REG_0__SCAN_IN), .B1(n3315), .B2(n3364), .ZN(n3182) );
  OAI211_X1 U3813 ( .C1(n3257), .C2(n4897), .A(n3183), .B(n3182), .ZN(U3229)
         );
  NAND2_X4 U3814 ( .A1(n3184), .A2(n4167), .ZN(n3855) );
  XNOR2_X1 U3815 ( .A(n3192), .B(n3835), .ZN(n3201) );
  XNOR2_X1 U3816 ( .A(n3203), .B(n3204), .ZN(n3200) );
  INV_X2 U3817 ( .A(n3315), .ZN(n3996) );
  NOR2_X1 U3818 ( .A1(n3996), .A2(n3359), .ZN(n3198) );
  INV_X1 U3819 ( .A(n4188), .ZN(n3328) );
  OAI22_X1 U3820 ( .A1(n3196), .A2(n4896), .B1(n4897), .B2(n3328), .ZN(n3197)
         );
  AOI211_X1 U3821 ( .C1(REG3_REG_1__SCAN_IN), .C2(n3214), .A(n3198), .B(n3197), 
        .ZN(n3199) );
  OAI21_X1 U3822 ( .B1(n3200), .B2(n4016), .A(n3199), .ZN(U3219) );
  NAND2_X1 U3823 ( .A1(n3737), .A2(n2287), .ZN(n3205) );
  NAND2_X1 U3824 ( .A1(n3206), .A2(n3205), .ZN(n3207) );
  NOR2_X1 U3825 ( .A1(n3256), .A2(n2279), .ZN(n3208) );
  OAI21_X1 U3826 ( .B1(n3211), .B2(n3210), .A(n3236), .ZN(n3213) );
  AOI21_X1 U3827 ( .B1(n3212), .B2(n3213), .A(n3238), .ZN(n3217) );
  AOI22_X1 U3828 ( .A1(n3214), .A2(REG3_REG_2__SCAN_IN), .B1(n3315), .B2(n3737), .ZN(n3216) );
  AOI22_X1 U3829 ( .A1(n3994), .A2(n2433), .B1(n3995), .B2(n3194), .ZN(n3215)
         );
  OAI211_X1 U3830 ( .C1(n3217), .C2(n4016), .A(n3216), .B(n3215), .ZN(U3234)
         );
  INV_X1 U3831 ( .A(n4655), .ZN(n3270) );
  NOR2_X1 U3832 ( .A1(STATE_REG_SCAN_IN), .A2(n3218), .ZN(n3952) );
  OAI21_X1 U3833 ( .B1(REG2_REG_4__SCAN_IN), .B2(n3221), .A(n4729), .ZN(n3233)
         );
  INV_X1 U3834 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3224) );
  OAI22_X1 U3835 ( .A1(n3225), .A2(n3224), .B1(n3223), .B2(n3222), .ZN(n3269)
         );
  XNOR2_X1 U3836 ( .A(n3269), .B(n4655), .ZN(n3273) );
  XNOR2_X1 U3837 ( .A(n3273), .B(REG1_REG_4__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U3838 ( .A1(n4769), .A2(n3226), .ZN(n3232) );
  NAND2_X1 U3839 ( .A1(n3227), .A2(n4168), .ZN(n3229) );
  OAI211_X1 U3840 ( .C1(n4192), .C2(n4168), .A(n3229), .B(n3228), .ZN(n3230)
         );
  OAI211_X1 U3841 ( .C1(IR_REG_0__SCAN_IN), .C2(n3231), .A(n3230), .B(U4043), 
        .ZN(n4214) );
  OAI211_X1 U3842 ( .C1(n3285), .C2(n3233), .A(n3232), .B(n4214), .ZN(n3234)
         );
  AOI211_X1 U3843 ( .C1(n4764), .C2(ADDR_REG_4__SCAN_IN), .A(n3952), .B(n3234), 
        .ZN(n3235) );
  OAI21_X1 U3844 ( .B1(n4767), .B2(n3270), .A(n3235), .ZN(U3244) );
  INV_X1 U3845 ( .A(n3236), .ZN(n3237) );
  NOR2_X2 U3846 ( .A1(n3238), .A2(n3237), .ZN(n3242) );
  XNOR2_X1 U3847 ( .A(n3240), .B(n3855), .ZN(n3301) );
  OAI22_X1 U3848 ( .A1(n3239), .A2(n3827), .B1(n3837), .B2(n3325), .ZN(n3300)
         );
  XNOR2_X1 U3849 ( .A(n3301), .B(n3300), .ZN(n3241) );
  AOI21_X1 U3850 ( .B1(n3242), .B2(n3241), .A(n3948), .ZN(n3252) );
  AOI22_X1 U3851 ( .A1(n3995), .A2(n4188), .B1(n3994), .B2(n4187), .ZN(n3251)
         );
  NAND4_X1 U3852 ( .A1(n3245), .A2(n3163), .A3(n3244), .A4(n3243), .ZN(n3247)
         );
  AOI21_X1 U3853 ( .B1(STATE_REG_SCAN_IN), .B2(n3247), .A(n3246), .ZN(n4912)
         );
  NOR2_X1 U3854 ( .A1(n3996), .A2(n3325), .ZN(n3248) );
  AOI211_X1 U3855 ( .C1(n4014), .C2(n4793), .A(n3249), .B(n3248), .ZN(n3250)
         );
  OAI211_X1 U3856 ( .C1(n3252), .C2(n4016), .A(n3251), .B(n3250), .ZN(U3215)
         );
  OR2_X1 U3857 ( .A1(n3253), .A2(n4120), .ZN(n3254) );
  NAND2_X1 U3858 ( .A1(n3255), .A2(n3254), .ZN(n3735) );
  OAI22_X1 U3859 ( .A1(n3257), .A2(n4834), .B1(n3256), .B2(n4833), .ZN(n3263)
         );
  NAND3_X1 U3860 ( .A1(n3355), .A2(n4120), .A3(n4070), .ZN(n3258) );
  NAND2_X1 U3861 ( .A1(n3259), .A2(n3258), .ZN(n3260) );
  NAND2_X1 U3862 ( .A1(n3260), .A2(n4449), .ZN(n3262) );
  NAND2_X1 U3863 ( .A1(n3735), .A2(n3650), .ZN(n3261) );
  OAI211_X1 U3864 ( .C1(n3239), .C2(n3689), .A(n3262), .B(n3261), .ZN(n3734)
         );
  AOI211_X1 U3865 ( .C1(n4802), .C2(n3735), .A(n3263), .B(n3734), .ZN(n3267)
         );
  INV_X1 U3866 ( .A(n4591), .ZN(n4510) );
  AND2_X1 U3867 ( .A1(n3366), .A2(n3737), .ZN(n3264) );
  NOR2_X1 U3868 ( .A1(n3331), .A2(n3264), .ZN(n3736) );
  AOI22_X1 U3869 ( .A1(n4510), .A2(n3736), .B1(REG1_REG_2__SCAN_IN), .B2(n3091), .ZN(n3265) );
  OAI21_X1 U3870 ( .B1(n3267), .B2(n3091), .A(n3265), .ZN(U3520) );
  INV_X1 U3871 ( .A(n4646), .ZN(n4596) );
  AOI22_X1 U3872 ( .A1(n4596), .A2(n3736), .B1(REG0_REG_2__SCAN_IN), .B2(n3099), .ZN(n3266) );
  OAI21_X1 U3873 ( .B1(n3267), .B2(n3099), .A(n3266), .ZN(U3471) );
  INV_X1 U3874 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3268) );
  INV_X1 U3875 ( .A(n3288), .ZN(n4807) );
  AOI22_X1 U3876 ( .A1(n3288), .A2(REG1_REG_5__SCAN_IN), .B1(n3268), .B2(n4807), .ZN(n4666) );
  INV_X1 U3877 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3272) );
  INV_X1 U3878 ( .A(n3269), .ZN(n3271) );
  OAI22_X1 U3879 ( .A1(n3273), .A2(n3272), .B1(n3271), .B2(n3270), .ZN(n4665)
         );
  NAND2_X1 U3880 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U3881 ( .A1(n3288), .A2(REG1_REG_5__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U3882 ( .A1(n3289), .A2(n3276), .ZN(n3277) );
  INV_X1 U3883 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U3884 ( .A1(n4817), .A2(n4851), .ZN(n4690) );
  INV_X1 U3885 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4695) );
  XNOR2_X1 U3886 ( .A(n4702), .B(n4688), .ZN(n4694) );
  INV_X1 U3887 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3278) );
  MUX2_X1 U3888 ( .A(REG1_REG_9__SCAN_IN), .B(n3278), .S(n3611), .Z(n3280) );
  OAI21_X1 U3889 ( .B1(n3610), .B2(n3280), .A(n4769), .ZN(n3279) );
  AOI21_X1 U3890 ( .B1(n3610), .B2(n3280), .A(n3279), .ZN(n3283) );
  NOR2_X1 U3891 ( .A1(STATE_REG_SCAN_IN), .A2(n2852), .ZN(n3963) );
  AOI21_X1 U3892 ( .B1(n4764), .B2(ADDR_REG_9__SCAN_IN), .A(n3963), .ZN(n3281)
         );
  OAI21_X1 U3893 ( .B1(n4767), .B2(n3611), .A(n3281), .ZN(n3282) );
  NOR2_X1 U3894 ( .A1(n3283), .A2(n3282), .ZN(n3299) );
  NAND2_X1 U3895 ( .A1(n3288), .A2(REG2_REG_5__SCAN_IN), .ZN(n3287) );
  OAI21_X1 U3896 ( .B1(n3288), .B2(REG2_REG_5__SCAN_IN), .A(n3287), .ZN(n4660)
         );
  NOR2_X1 U3897 ( .A1(n4661), .A2(n4660), .ZN(n4659) );
  NOR2_X1 U3898 ( .A1(n3290), .A2(n3275), .ZN(n3291) );
  INV_X1 U3899 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4671) );
  XNOR2_X1 U3900 ( .A(n3290), .B(n3275), .ZN(n4670) );
  NOR2_X1 U3901 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  OR2_X1 U3902 ( .A1(n4702), .A2(n3293), .ZN(n3294) );
  NAND2_X1 U3903 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4699), .ZN(n4698) );
  INV_X1 U3904 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3295) );
  MUX2_X1 U3905 ( .A(n3295), .B(REG2_REG_9__SCAN_IN), .S(n3611), .Z(n3296) );
  OAI211_X1 U3906 ( .C1(n3297), .C2(n3296), .A(n3593), .B(n4729), .ZN(n3298)
         );
  NAND2_X1 U3907 ( .A1(n3299), .A2(n3298), .ZN(U3249) );
  NOR2_X1 U3908 ( .A1(n3301), .A2(n3300), .ZN(n3947) );
  AOI22_X1 U3909 ( .A1(n4187), .A2(n2274), .B1(n2277), .B2(n3304), .ZN(n3303)
         );
  XNOR2_X1 U3910 ( .A(n3303), .B(n3855), .ZN(n3306) );
  INV_X2 U3911 ( .A(n3827), .ZN(n3854) );
  AOI22_X1 U3912 ( .A1(n4187), .A2(n3854), .B1(n2274), .B2(n3304), .ZN(n3305)
         );
  XNOR2_X1 U3913 ( .A(n3306), .B(n3305), .ZN(n3946) );
  NOR2_X1 U3914 ( .A1(n3306), .A2(n3305), .ZN(n3307) );
  NAND2_X1 U3915 ( .A1(n4186), .A2(n2273), .ZN(n3309) );
  NAND2_X1 U3916 ( .A1(n3438), .A2(n2277), .ZN(n3308) );
  NAND2_X1 U3917 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  XNOR2_X1 U3918 ( .A(n3310), .B(n3835), .ZN(n3312) );
  AOI22_X1 U3919 ( .A1(n4186), .A2(n3854), .B1(n2274), .B2(n3438), .ZN(n3311)
         );
  OR2_X1 U3920 ( .A1(n3312), .A2(n3311), .ZN(n3344) );
  NAND2_X1 U3921 ( .A1(n2315), .A2(n3344), .ZN(n3313) );
  XNOR2_X1 U3922 ( .A(n3345), .B(n3313), .ZN(n3320) );
  AOI22_X1 U3923 ( .A1(n3994), .A2(n4185), .B1(n3995), .B2(n4187), .ZN(n3319)
         );
  NOR2_X1 U3924 ( .A1(STATE_REG_SCAN_IN), .A2(n3314), .ZN(n4662) );
  NOR2_X1 U3925 ( .A1(n3996), .A2(n3338), .ZN(n3316) );
  AOI211_X1 U3926 ( .C1(n4014), .C2(n3317), .A(n4662), .B(n3316), .ZN(n3318)
         );
  OAI211_X1 U3927 ( .C1(n3320), .C2(n4016), .A(n3319), .B(n3318), .ZN(U3224)
         );
  XNOR2_X1 U3928 ( .A(n3321), .B(n4125), .ZN(n4795) );
  OAI21_X1 U3929 ( .B1(n3323), .B2(n3322), .A(n3376), .ZN(n3324) );
  NAND2_X1 U3930 ( .A1(n3324), .A2(n4449), .ZN(n3327) );
  AOI22_X1 U3931 ( .A1(n4187), .A2(n4838), .B1(n4443), .B2(n2432), .ZN(n3326)
         );
  OAI211_X1 U3932 ( .C1(n3328), .C2(n4834), .A(n3327), .B(n3326), .ZN(n3329)
         );
  AOI21_X1 U3933 ( .B1(n3650), .B2(n4795), .A(n3329), .ZN(n4798) );
  INV_X1 U3934 ( .A(n4798), .ZN(n3330) );
  AOI21_X1 U3935 ( .B1(n4802), .B2(n4795), .A(n3330), .ZN(n3336) );
  INV_X1 U3936 ( .A(n3331), .ZN(n3333) );
  INV_X1 U3937 ( .A(n3332), .ZN(n3374) );
  AOI21_X1 U3938 ( .B1(n2432), .B2(n3333), .A(n3374), .ZN(n4794) );
  AOI22_X1 U3939 ( .A1(n4794), .A2(n4596), .B1(REG0_REG_3__SCAN_IN), .B2(n3099), .ZN(n3334) );
  OAI21_X1 U3940 ( .B1(n3336), .B2(n3099), .A(n3334), .ZN(U3473) );
  AOI22_X1 U3941 ( .A1(n4794), .A2(n4510), .B1(REG1_REG_3__SCAN_IN), .B2(n3091), .ZN(n3335) );
  OAI21_X1 U3942 ( .B1(n3336), .B2(n3091), .A(n3335), .ZN(U3521) );
  NAND2_X1 U3943 ( .A1(n2304), .A2(n4055), .ZN(n4122) );
  XNOR2_X1 U3944 ( .A(n3337), .B(n4122), .ZN(n3436) );
  INV_X1 U3945 ( .A(n4187), .ZN(n3444) );
  OAI22_X1 U3946 ( .A1(n3444), .A2(n4834), .B1(n3338), .B2(n4833), .ZN(n3340)
         );
  OAI22_X1 U3947 ( .A1(n3339), .A2(n4840), .B1(n4835), .B2(n3689), .ZN(n3446)
         );
  AOI211_X1 U3948 ( .C1(n3436), .C2(n4587), .A(n3340), .B(n3446), .ZN(n3343)
         );
  AOI21_X1 U3949 ( .B1(n3438), .B2(n3373), .A(n3397), .ZN(n3439) );
  AOI22_X1 U3950 ( .A1(n3439), .A2(n4596), .B1(REG0_REG_5__SCAN_IN), .B2(n3099), .ZN(n3341) );
  OAI21_X1 U3951 ( .B1(n3343), .B2(n3099), .A(n3341), .ZN(U3477) );
  AOI22_X1 U3952 ( .A1(n3439), .A2(n4510), .B1(REG1_REG_5__SCAN_IN), .B2(n3091), .ZN(n3342) );
  OAI21_X1 U3953 ( .B1(n3343), .B2(n3091), .A(n3342), .ZN(U3523) );
  XOR2_X1 U3954 ( .A(n3855), .B(n3346), .Z(n3407) );
  XNOR2_X1 U3955 ( .A(n3407), .B(n3409), .ZN(n3348) );
  XNOR2_X1 U3956 ( .A(n3410), .B(n3348), .ZN(n3353) );
  AOI22_X1 U3957 ( .A1(n3994), .A2(n4184), .B1(n3995), .B2(n4186), .ZN(n3352)
         );
  NOR2_X1 U3958 ( .A1(STATE_REG_SCAN_IN), .A2(n3349), .ZN(n4672) );
  NOR2_X1 U3959 ( .A1(n3996), .A2(n3396), .ZN(n3350) );
  AOI211_X1 U3960 ( .C1(n4014), .C2(n4809), .A(n4672), .B(n3350), .ZN(n3351)
         );
  OAI211_X1 U3961 ( .C1(n3353), .C2(n4016), .A(n3352), .B(n3351), .ZN(U3236)
         );
  XNOR2_X1 U3962 ( .A(n4128), .B(n3354), .ZN(n4787) );
  OAI21_X1 U3963 ( .B1(n3356), .B2(n4069), .A(n3355), .ZN(n3361) );
  NAND2_X1 U3964 ( .A1(n4190), .A2(n4406), .ZN(n3358) );
  NAND2_X1 U3965 ( .A1(n4188), .A2(n4838), .ZN(n3357) );
  OAI211_X1 U3966 ( .C1(n4833), .C2(n3359), .A(n3358), .B(n3357), .ZN(n3360)
         );
  AOI21_X1 U3967 ( .B1(n3361), .B2(n4449), .A(n3360), .ZN(n3362) );
  OAI21_X1 U3968 ( .B1(n4787), .B2(n4452), .A(n3362), .ZN(n4789) );
  INV_X1 U3969 ( .A(n4789), .ZN(n3372) );
  INV_X2 U3970 ( .A(n4889), .ZN(n4462) );
  INV_X1 U3971 ( .A(n4787), .ZN(n3370) );
  OR2_X1 U3972 ( .A1(n3184), .A2(n4766), .ZN(n3437) );
  INV_X1 U3973 ( .A(n3437), .ZN(n3363) );
  AND2_X1 U3974 ( .A1(n4889), .A2(n3363), .ZN(n4871) );
  NAND2_X1 U3975 ( .A1(n3365), .A2(n3364), .ZN(n3367) );
  NAND2_X1 U3976 ( .A1(n3367), .A2(n3366), .ZN(n4785) );
  AOI22_X1 U3977 ( .A1(n4462), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4866), .ZN(n3368) );
  OAI21_X1 U3978 ( .B1(n4883), .B2(n4785), .A(n3368), .ZN(n3369) );
  AOI21_X1 U3979 ( .B1(n3370), .B2(n4871), .A(n3369), .ZN(n3371) );
  OAI21_X1 U3980 ( .B1(n3372), .B2(n4462), .A(n3371), .ZN(U3289) );
  OAI211_X1 U3981 ( .C1(n3374), .C2(n3951), .A(n3093), .B(n3373), .ZN(n4799)
         );
  NOR2_X1 U3982 ( .A1(n4799), .A2(n4829), .ZN(n3384) );
  NAND2_X1 U3983 ( .A1(n3376), .A2(n3375), .ZN(n3377) );
  XOR2_X1 U3984 ( .A(n4150), .B(n3377), .Z(n3383) );
  OAI22_X1 U3985 ( .A1(n3239), .A2(n4834), .B1(n3951), .B2(n4833), .ZN(n3381)
         );
  AND2_X1 U3986 ( .A1(n3378), .A2(n4150), .ZN(n3379) );
  OR2_X1 U3987 ( .A1(n2311), .A2(n3379), .ZN(n3385) );
  NOR2_X1 U3988 ( .A1(n3385), .A2(n4452), .ZN(n3380) );
  AOI211_X1 U3989 ( .C1(n4838), .C2(n4186), .A(n3381), .B(n3380), .ZN(n3382)
         );
  OAI21_X1 U3990 ( .B1(n4840), .B2(n3383), .A(n3382), .ZN(n4800) );
  AOI211_X1 U3991 ( .C1(n4866), .C2(n3954), .A(n3384), .B(n4800), .ZN(n3387)
         );
  INV_X1 U3992 ( .A(n3385), .ZN(n4803) );
  AOI22_X1 U3993 ( .A1(n4803), .A2(n4871), .B1(REG2_REG_4__SCAN_IN), .B2(n4462), .ZN(n3386) );
  OAI21_X1 U3994 ( .B1(n3387), .B2(n4462), .A(n3386), .ZN(U3286) );
  NAND2_X1 U3995 ( .A1(n4081), .A2(n4079), .ZN(n4126) );
  XOR2_X1 U3996 ( .A(n4126), .B(n3388), .Z(n4812) );
  INV_X1 U3997 ( .A(n4812), .ZN(n3395) );
  XNOR2_X1 U3998 ( .A(n3389), .B(n4126), .ZN(n3393) );
  OAI22_X1 U3999 ( .A1(n3390), .A2(n4834), .B1(n4833), .B2(n3396), .ZN(n3391)
         );
  AOI21_X1 U4000 ( .B1(n4838), .B2(n4184), .A(n3391), .ZN(n3392) );
  OAI21_X1 U4001 ( .B1(n3393), .B2(n4840), .A(n3392), .ZN(n3394) );
  AOI21_X1 U4002 ( .B1(n4812), .B2(n3650), .A(n3394), .ZN(n4815) );
  OAI21_X1 U4003 ( .B1(n4786), .B2(n3395), .A(n4815), .ZN(n3404) );
  OR2_X1 U4004 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  NAND2_X1 U4005 ( .A1(n4820), .A2(n3398), .ZN(n4810) );
  INV_X1 U4006 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3399) );
  OAI22_X1 U4007 ( .A1(n4810), .A2(n4591), .B1(n4852), .B2(n3399), .ZN(n3400)
         );
  AOI21_X1 U4008 ( .B1(n3404), .B2(n4852), .A(n3400), .ZN(n3401) );
  INV_X1 U4009 ( .A(n3401), .ZN(U3524) );
  INV_X1 U4010 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3402) );
  OAI22_X1 U4011 ( .A1(n4810), .A2(n4646), .B1(n4855), .B2(n3402), .ZN(n3403)
         );
  AOI21_X1 U4012 ( .B1(n3404), .B2(n4855), .A(n3403), .ZN(n3405) );
  INV_X1 U4013 ( .A(n3405), .ZN(U3479) );
  INV_X1 U4014 ( .A(n3406), .ZN(n3409) );
  NOR2_X1 U4015 ( .A1(n4832), .A2(n3837), .ZN(n3411) );
  AOI21_X1 U4016 ( .B1(n4184), .B2(n3854), .A(n3411), .ZN(n3421) );
  XNOR2_X1 U4017 ( .A(n3412), .B(n3855), .ZN(n3419) );
  XOR2_X1 U4018 ( .A(n3421), .B(n3419), .Z(n3422) );
  XNOR2_X1 U4019 ( .A(n3423), .B(n3422), .ZN(n3418) );
  AOI22_X1 U4020 ( .A1(n3995), .A2(n4185), .B1(n3994), .B2(n4837), .ZN(n3417)
         );
  NOR2_X1 U4021 ( .A1(STATE_REG_SCAN_IN), .A2(n3413), .ZN(n4687) );
  NOR2_X1 U4022 ( .A1(n3996), .A2(n4832), .ZN(n3414) );
  AOI211_X1 U4023 ( .C1(n4014), .C2(n3415), .A(n4687), .B(n3414), .ZN(n3416)
         );
  OAI211_X1 U4024 ( .C1(n3418), .C2(n4016), .A(n3417), .B(n3416), .ZN(U3210)
         );
  INV_X1 U4025 ( .A(n3419), .ZN(n3420) );
  XNOR2_X1 U4026 ( .A(n3424), .B(n3835), .ZN(n3428) );
  OR2_X1 U4027 ( .A1(n3483), .A2(n3827), .ZN(n3426) );
  NAND2_X1 U4028 ( .A1(n3500), .A2(n2273), .ZN(n3425) );
  AND2_X1 U4029 ( .A1(n3426), .A2(n3425), .ZN(n3427) );
  NOR2_X1 U4030 ( .A1(n3428), .A2(n3427), .ZN(n3464) );
  NAND2_X1 U4031 ( .A1(n3428), .A2(n3427), .ZN(n3463) );
  INV_X1 U4032 ( .A(n3463), .ZN(n3429) );
  NOR2_X1 U4033 ( .A1(n3464), .A2(n3429), .ZN(n3430) );
  XNOR2_X1 U4034 ( .A(n3465), .B(n3430), .ZN(n3435) );
  AOI22_X1 U4035 ( .A1(n3994), .A2(n4183), .B1(n3995), .B2(n4184), .ZN(n3434)
         );
  NOR2_X1 U4036 ( .A1(STATE_REG_SCAN_IN), .A2(n3431), .ZN(n4696) );
  NOR2_X1 U4037 ( .A1(n3996), .A2(n3493), .ZN(n3432) );
  AOI211_X1 U4038 ( .C1(n4014), .C2(n4858), .A(n4696), .B(n3432), .ZN(n3433)
         );
  OAI211_X1 U4039 ( .C1(n3435), .C2(n4016), .A(n3434), .B(n3433), .ZN(U3218)
         );
  INV_X1 U4040 ( .A(n3436), .ZN(n3448) );
  NAND2_X1 U4041 ( .A1(n4452), .A2(n3437), .ZN(n4824) );
  AND2_X1 U4042 ( .A1(n4889), .A2(n4824), .ZN(n4305) );
  AND2_X1 U40430 ( .A1(n4889), .A2(n4406), .ZN(n4430) );
  INV_X1 U4044 ( .A(n4430), .ZN(n3459) );
  NAND2_X1 U4045 ( .A1(n4826), .A2(n4443), .ZN(n4433) );
  INV_X1 U4046 ( .A(n4433), .ZN(n3738) );
  AOI22_X1 U4047 ( .A1(n3439), .A2(n4870), .B1(n3438), .B2(n3738), .ZN(n3443)
         );
  NOR2_X1 U4048 ( .A1(n3440), .A2(n4879), .ZN(n3441) );
  AOI21_X1 U4049 ( .B1(n4462), .B2(REG2_REG_5__SCAN_IN), .A(n3441), .ZN(n3442)
         );
  OAI211_X1 U4050 ( .C1(n3444), .C2(n3459), .A(n3443), .B(n3442), .ZN(n3445)
         );
  AOI21_X1 U4051 ( .B1(n3446), .B2(n4889), .A(n3445), .ZN(n3447) );
  OAI21_X1 U4052 ( .B1(n3448), .B2(n4502), .A(n3447), .ZN(U3285) );
  INV_X1 U4053 ( .A(n4084), .ZN(n3450) );
  NAND2_X1 U4054 ( .A1(n3450), .A2(n4086), .ZN(n4127) );
  XNOR2_X1 U4055 ( .A(n3449), .B(n4127), .ZN(n3486) );
  INV_X1 U4056 ( .A(n3486), .ZN(n3462) );
  XOR2_X1 U4057 ( .A(n4127), .B(n3451), .Z(n3452) );
  OAI22_X1 U4058 ( .A1(n3452), .A2(n4840), .B1(n3652), .B2(n3689), .ZN(n3485)
         );
  INV_X1 U4059 ( .A(n3502), .ZN(n3453) );
  AOI21_X1 U4060 ( .B1(n3456), .B2(n3453), .A(n3536), .ZN(n3488) );
  NAND2_X1 U4061 ( .A1(n3488), .A2(n4870), .ZN(n3458) );
  INV_X1 U4062 ( .A(n3965), .ZN(n3454) );
  OAI22_X1 U4063 ( .A1(n4826), .A2(n3295), .B1(n3454), .B2(n4879), .ZN(n3455)
         );
  AOI21_X1 U4064 ( .B1(n3456), .B2(n3738), .A(n3455), .ZN(n3457) );
  OAI211_X1 U4065 ( .C1(n3483), .C2(n3459), .A(n3458), .B(n3457), .ZN(n3460)
         );
  AOI21_X1 U4066 ( .B1(n3485), .B2(n4889), .A(n3460), .ZN(n3461) );
  OAI21_X1 U4067 ( .B1(n3462), .B2(n4502), .A(n3461), .ZN(U3281) );
  OAI21_X1 U4068 ( .B1(n3465), .B2(n3464), .A(n3463), .ZN(n3959) );
  OAI22_X1 U4069 ( .A1(n3540), .A2(n3827), .B1(n3837), .B2(n3962), .ZN(n3471)
         );
  XNOR2_X1 U4070 ( .A(n3466), .B(n3855), .ZN(n3470) );
  XOR2_X1 U4071 ( .A(n3471), .B(n3470), .Z(n3960) );
  NAND2_X1 U4072 ( .A1(n3959), .A2(n3960), .ZN(n3958) );
  XNOR2_X1 U4073 ( .A(n3467), .B(n3835), .ZN(n3509) );
  OR2_X1 U4074 ( .A1(n3652), .A2(n3827), .ZN(n3469) );
  NAND2_X1 U4075 ( .A1(n2320), .A2(n2274), .ZN(n3468) );
  NAND2_X1 U4076 ( .A1(n3469), .A2(n3468), .ZN(n3510) );
  XNOR2_X1 U4077 ( .A(n3509), .B(n3510), .ZN(n3475) );
  INV_X1 U4078 ( .A(n3470), .ZN(n3473) );
  INV_X1 U4079 ( .A(n3471), .ZN(n3472) );
  NAND2_X1 U4080 ( .A1(n3473), .A2(n3472), .ZN(n3476) );
  NAND2_X1 U4081 ( .A1(n3513), .A2(n4907), .ZN(n3482) );
  AOI21_X1 U4082 ( .B1(n3958), .B2(n3476), .A(n3475), .ZN(n3481) );
  AOI22_X1 U4083 ( .A1(n3995), .A2(n4183), .B1(n3994), .B2(n4181), .ZN(n3480)
         );
  NOR2_X1 U4084 ( .A1(STATE_REG_SCAN_IN), .A2(n3477), .ZN(n4710) );
  NOR2_X1 U4085 ( .A1(n3996), .A2(n3539), .ZN(n3478) );
  AOI211_X1 U4086 ( .C1(n4014), .C2(n4867), .A(n4710), .B(n3478), .ZN(n3479)
         );
  OAI211_X1 U4087 ( .C1(n3482), .C2(n3481), .A(n3480), .B(n3479), .ZN(U3214)
         );
  OAI22_X1 U4088 ( .A1(n3483), .A2(n4834), .B1(n4833), .B2(n3962), .ZN(n3484)
         );
  AOI211_X1 U4089 ( .C1(n3486), .C2(n4587), .A(n3485), .B(n3484), .ZN(n3490)
         );
  AOI22_X1 U4090 ( .A1(n3488), .A2(n4510), .B1(REG1_REG_9__SCAN_IN), .B2(n3091), .ZN(n3487) );
  OAI21_X1 U4091 ( .B1(n3490), .B2(n3091), .A(n3487), .ZN(U3527) );
  AOI22_X1 U4092 ( .A1(n3488), .A2(n4596), .B1(REG0_REG_9__SCAN_IN), .B2(n3099), .ZN(n3489) );
  OAI21_X1 U4093 ( .B1(n3490), .B2(n3099), .A(n3489), .ZN(U3485) );
  NAND2_X1 U4094 ( .A1(n4085), .A2(n4052), .ZN(n4132) );
  XOR2_X1 U4095 ( .A(n4132), .B(n3491), .Z(n4860) );
  INV_X1 U4096 ( .A(n4860), .ZN(n3499) );
  XOR2_X1 U4097 ( .A(n4132), .B(n3492), .Z(n3497) );
  OAI22_X1 U4098 ( .A1(n3494), .A2(n4834), .B1(n3493), .B2(n4833), .ZN(n3495)
         );
  AOI21_X1 U4099 ( .B1(n4838), .B2(n4183), .A(n3495), .ZN(n3496) );
  OAI21_X1 U4100 ( .B1(n3497), .B2(n4840), .A(n3496), .ZN(n3498) );
  AOI21_X1 U4101 ( .B1(n4860), .B2(n3650), .A(n3498), .ZN(n4863) );
  OAI21_X1 U4102 ( .B1(n4786), .B2(n3499), .A(n4863), .ZN(n3505) );
  NAND2_X1 U4103 ( .A1(n3505), .A2(n4852), .ZN(n3504) );
  AND2_X1 U4104 ( .A1(n4821), .A2(n3500), .ZN(n3501) );
  NOR2_X1 U4105 ( .A1(n3502), .A2(n3501), .ZN(n4859) );
  NAND2_X1 U4106 ( .A1(n4859), .A2(n4510), .ZN(n3503) );
  OAI211_X1 U4107 ( .C1(n4852), .C2(n4695), .A(n3504), .B(n3503), .ZN(U3526)
         );
  INV_X1 U4108 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U4109 ( .A1(n3505), .A2(n4855), .ZN(n3507) );
  NAND2_X1 U4110 ( .A1(n4859), .A2(n4596), .ZN(n3506) );
  OAI211_X1 U4111 ( .C1(n4855), .C2(n3508), .A(n3507), .B(n3506), .ZN(U3483)
         );
  NAND2_X1 U4112 ( .A1(n4181), .A2(n2273), .ZN(n3516) );
  NAND2_X1 U4113 ( .A1(n3514), .A2(n2276), .ZN(n3515) );
  NAND2_X1 U4114 ( .A1(n3516), .A2(n3515), .ZN(n3517) );
  XNOR2_X1 U4115 ( .A(n3517), .B(n3835), .ZN(n3520) );
  NOR2_X1 U4116 ( .A1(n3651), .A2(n3837), .ZN(n3518) );
  AOI21_X1 U4117 ( .B1(n4181), .B2(n3854), .A(n3518), .ZN(n3519) );
  NOR2_X1 U4118 ( .A1(n3520), .A2(n3519), .ZN(n3527) );
  NOR2_X1 U4119 ( .A1(n3527), .A2(n2313), .ZN(n3521) );
  XNOR2_X1 U4120 ( .A(n3528), .B(n3521), .ZN(n3526) );
  AOI22_X1 U4121 ( .A1(n3995), .A2(n4182), .B1(n3994), .B2(n4180), .ZN(n3525)
         );
  AND2_X1 U4122 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4716) );
  NOR2_X1 U4123 ( .A1(n3996), .A2(n3651), .ZN(n3522) );
  AOI211_X1 U4124 ( .C1(n4014), .C2(n3523), .A(n4716), .B(n3522), .ZN(n3524)
         );
  OAI211_X1 U4125 ( .C1(n3526), .C2(n4016), .A(n3525), .B(n3524), .ZN(U3233)
         );
  XOR2_X1 U4126 ( .A(n3855), .B(n3529), .Z(n3567) );
  AOI22_X1 U4127 ( .A1(n4180), .A2(n3854), .B1(n2273), .B2(n3556), .ZN(n3569)
         );
  XNOR2_X1 U4128 ( .A(n3567), .B(n3569), .ZN(n3530) );
  XNOR2_X1 U4129 ( .A(n3568), .B(n3530), .ZN(n3535) );
  AOI22_X1 U4130 ( .A1(n3995), .A2(n4181), .B1(n3994), .B2(n4179), .ZN(n3534)
         );
  NOR2_X1 U4131 ( .A1(STATE_REG_SCAN_IN), .A2(n3531), .ZN(n4726) );
  NOR2_X1 U4132 ( .A1(n3996), .A2(n3635), .ZN(n3532) );
  AOI211_X1 U4133 ( .C1(n4014), .C2(n3558), .A(n4726), .B(n3532), .ZN(n3533)
         );
  OAI211_X1 U4134 ( .C1(n3535), .C2(n4016), .A(n3534), .B(n3533), .ZN(U3221)
         );
  OAI21_X1 U4135 ( .B1(n3536), .B2(n3539), .A(n3644), .ZN(n4868) );
  INV_X1 U4136 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4137 ( .A1(n4057), .A2(n4060), .ZN(n4133) );
  XNOR2_X1 U4138 ( .A(n3537), .B(n4133), .ZN(n4872) );
  XNOR2_X1 U4139 ( .A(n3538), .B(n4133), .ZN(n3543) );
  OAI22_X1 U4140 ( .A1(n3540), .A2(n4834), .B1(n3539), .B2(n4833), .ZN(n3541)
         );
  AOI21_X1 U4141 ( .B1(n4838), .B2(n4181), .A(n3541), .ZN(n3542) );
  OAI21_X1 U4142 ( .B1(n3543), .B2(n4840), .A(n3542), .ZN(n3544) );
  AOI21_X1 U4143 ( .B1(n4872), .B2(n3650), .A(n3544), .ZN(n4875) );
  INV_X1 U4144 ( .A(n4875), .ZN(n3545) );
  AOI21_X1 U4145 ( .B1(n4802), .B2(n4872), .A(n3545), .ZN(n3548) );
  MUX2_X1 U4146 ( .A(n3546), .B(n3548), .S(n4855), .Z(n3547) );
  OAI21_X1 U4147 ( .B1(n4868), .B2(n4646), .A(n3547), .ZN(U3487) );
  INV_X1 U4148 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3549) );
  MUX2_X1 U4149 ( .A(n3549), .B(n3548), .S(n4852), .Z(n3550) );
  OAI21_X1 U4150 ( .B1(n4868), .B2(n4591), .A(n3550), .ZN(U3528) );
  NAND2_X1 U4151 ( .A1(n3669), .A2(n3667), .ZN(n4138) );
  XNOR2_X1 U4152 ( .A(n3551), .B(n4138), .ZN(n3638) );
  INV_X1 U4153 ( .A(n3638), .ZN(n3566) );
  INV_X1 U4154 ( .A(n3552), .ZN(n3553) );
  AOI21_X1 U4155 ( .B1(n3649), .B2(n3554), .A(n3553), .ZN(n3670) );
  XOR2_X1 U4156 ( .A(n4138), .B(n3670), .Z(n3555) );
  OAI22_X1 U4157 ( .A1(n3555), .A2(n4840), .B1(n4584), .B2(n3689), .ZN(n3637)
         );
  AND2_X1 U4158 ( .A1(n3645), .A2(n3556), .ZN(n3557) );
  OR2_X1 U4159 ( .A1(n3557), .A2(n3678), .ZN(n3643) );
  INV_X1 U4160 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3560) );
  INV_X1 U4161 ( .A(n3558), .ZN(n3559) );
  OAI22_X1 U4162 ( .A1(n4826), .A2(n3560), .B1(n3559), .B2(n4879), .ZN(n3562)
         );
  NOR2_X1 U4163 ( .A1(n4433), .A2(n3635), .ZN(n3561) );
  AOI211_X1 U4164 ( .C1(n4430), .C2(n4181), .A(n3562), .B(n3561), .ZN(n3563)
         );
  OAI21_X1 U4165 ( .B1(n3643), .B2(n4883), .A(n3563), .ZN(n3564) );
  AOI21_X1 U4166 ( .B1(n3637), .B2(n4889), .A(n3564), .ZN(n3565) );
  OAI21_X1 U4167 ( .B1(n3566), .B2(n4502), .A(n3565), .ZN(U3278) );
  INV_X1 U4168 ( .A(n3569), .ZN(n3570) );
  NAND2_X1 U4169 ( .A1(n4179), .A2(n2274), .ZN(n3572) );
  NAND2_X1 U4170 ( .A1(n3574), .A2(n2277), .ZN(n3571) );
  NAND2_X1 U4171 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  XNOR2_X1 U4172 ( .A(n3573), .B(n3835), .ZN(n3576) );
  AOI22_X1 U4173 ( .A1(n4179), .A2(n3854), .B1(n2274), .B2(n3574), .ZN(n3575)
         );
  AND2_X1 U4174 ( .A1(n3576), .A2(n3575), .ZN(n3584) );
  INV_X1 U4175 ( .A(n3584), .ZN(n3577) );
  OR2_X1 U4176 ( .A1(n3576), .A2(n3575), .ZN(n3585) );
  NAND2_X1 U4177 ( .A1(n3577), .A2(n3585), .ZN(n3578) );
  XNOR2_X1 U4178 ( .A(n2269), .B(n3578), .ZN(n3583) );
  AOI22_X1 U4179 ( .A1(n3994), .A2(n4178), .B1(n3995), .B2(n4180), .ZN(n3582)
         );
  NOR2_X1 U4180 ( .A1(STATE_REG_SCAN_IN), .A2(n3579), .ZN(n4745) );
  NOR2_X1 U4181 ( .A1(n3996), .A2(n3677), .ZN(n3580) );
  AOI211_X1 U4182 ( .C1(n4014), .C2(n3679), .A(n4745), .B(n3580), .ZN(n3581)
         );
  OAI211_X1 U4183 ( .C1(n3583), .C2(n4016), .A(n3582), .B(n3581), .ZN(U3231)
         );
  AOI22_X1 U4184 ( .A1(n4178), .A2(n2274), .B1(n2276), .B2(n3586), .ZN(n3587)
         );
  XOR2_X1 U4185 ( .A(n3855), .B(n3587), .Z(n3744) );
  INV_X1 U4186 ( .A(n4178), .ZN(n4895) );
  OAI22_X1 U4187 ( .A1(n4895), .A2(n3827), .B1(n3837), .B2(n4583), .ZN(n3745)
         );
  INV_X1 U4188 ( .A(n3745), .ZN(n3746) );
  XNOR2_X1 U4189 ( .A(n3744), .B(n3746), .ZN(n3588) );
  XNOR2_X1 U4190 ( .A(n3747), .B(n3588), .ZN(n3592) );
  NAND2_X1 U4191 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3605) );
  OAI21_X1 U4192 ( .B1(n3996), .B2(n4583), .A(n3605), .ZN(n3590) );
  OAI22_X1 U4193 ( .A1(n4572), .A2(n4897), .B1(n4896), .B2(n4584), .ZN(n3589)
         );
  AOI211_X1 U4194 ( .C1(n4014), .C2(n3692), .A(n3590), .B(n3589), .ZN(n3591)
         );
  OAI21_X1 U4195 ( .B1(n3592), .B2(n4016), .A(n3591), .ZN(U3212) );
  INV_X1 U4196 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4197 ( .A1(n4712), .A2(REG2_REG_11__SCAN_IN), .ZN(n3597) );
  INV_X1 U4198 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4878) );
  AOI22_X1 U4199 ( .A1(n4712), .A2(REG2_REG_11__SCAN_IN), .B1(n4878), .B2(
        n4877), .ZN(n4720) );
  NAND2_X1 U4200 ( .A1(n2403), .A2(REG2_REG_9__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4201 ( .A1(n3613), .A2(n3595), .ZN(n3596) );
  NAND2_X1 U4202 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U4203 ( .A1(n3596), .A2(n4705), .ZN(n4719) );
  NAND2_X1 U4204 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U4205 ( .A1(n3616), .A2(n3598), .ZN(n3599) );
  INV_X1 U4206 ( .A(n3619), .ZN(n4894) );
  INV_X1 U4207 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4734) );
  NOR2_X1 U4208 ( .A1(n4894), .A2(n4734), .ZN(n4733) );
  INV_X1 U4209 ( .A(n4216), .ZN(n3602) );
  NAND2_X1 U4210 ( .A1(n3600), .A2(n4224), .ZN(n3601) );
  NOR2_X1 U4211 ( .A1(n3603), .A2(n3604), .ZN(n4215) );
  AOI211_X1 U4212 ( .C1(n3604), .C2(n3603), .A(n4215), .B(n4771), .ZN(n3609)
         );
  INV_X1 U4213 ( .A(n3605), .ZN(n3606) );
  AOI21_X1 U4214 ( .B1(n4764), .B2(ADDR_REG_14__SCAN_IN), .A(n3606), .ZN(n3607) );
  OAI21_X1 U4215 ( .B1(n4767), .B2(n4224), .A(n3607), .ZN(n3608) );
  NOR2_X1 U4216 ( .A1(n3609), .A2(n3608), .ZN(n3622) );
  NAND2_X1 U4217 ( .A1(n3613), .A2(n3612), .ZN(n3614) );
  XOR2_X1 U4218 ( .A(n3613), .B(n3612), .Z(n4704) );
  NAND2_X1 U4219 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4704), .ZN(n4703) );
  INV_X1 U4220 ( .A(n3616), .ZN(n4892) );
  NOR2_X1 U4221 ( .A1(n3617), .A2(n4892), .ZN(n3618) );
  INV_X1 U4222 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4725) );
  NOR2_X1 U4223 ( .A1(n4725), .A2(n4724), .ZN(n4723) );
  NOR2_X1 U4224 ( .A1(n3618), .A2(n4723), .ZN(n4741) );
  NAND2_X1 U4225 ( .A1(n3619), .A2(REG1_REG_13__SCAN_IN), .ZN(n4739) );
  NOR2_X1 U4226 ( .A1(n3619), .A2(REG1_REG_13__SCAN_IN), .ZN(n4737) );
  AOI21_X1 U4227 ( .B1(n4741), .B2(n4739), .A(n4737), .ZN(n4225) );
  XNOR2_X1 U4228 ( .A(n4225), .B(n4224), .ZN(n3620) );
  OAI211_X1 U4229 ( .C1(n3620), .C2(REG1_REG_14__SCAN_IN), .A(n4769), .B(n4226), .ZN(n3621) );
  NAND2_X1 U4230 ( .A1(n3622), .A2(n3621), .ZN(U3254) );
  OAI21_X1 U4231 ( .B1(n3624), .B2(n4141), .A(n3623), .ZN(n4577) );
  INV_X1 U4232 ( .A(n3625), .ZN(n3704) );
  AOI21_X1 U4233 ( .B1(n3757), .B2(n3723), .A(n3704), .ZN(n4575) );
  AOI22_X1 U4234 ( .A1(n4462), .A2(REG2_REG_16__SCAN_IN), .B1(n3923), .B2(
        n4866), .ZN(n3627) );
  NAND2_X1 U4235 ( .A1(n4430), .A2(n4177), .ZN(n3626) );
  OAI211_X1 U4236 ( .C1(n4433), .C2(n4571), .A(n3627), .B(n3626), .ZN(n3628)
         );
  AOI21_X1 U4237 ( .B1(n4575), .B2(n4870), .A(n3628), .ZN(n3634) );
  OAI211_X1 U4238 ( .C1(n3631), .C2(n3630), .A(n3629), .B(n4449), .ZN(n3632)
         );
  OAI21_X1 U4239 ( .B1(n4491), .B2(n3689), .A(n3632), .ZN(n4573) );
  NAND2_X1 U4240 ( .A1(n4573), .A2(n4889), .ZN(n3633) );
  OAI211_X1 U4241 ( .C1(n4577), .C2(n4502), .A(n3634), .B(n3633), .ZN(U3274)
         );
  INV_X1 U4242 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3639) );
  OAI22_X1 U4243 ( .A1(n2927), .A2(n4834), .B1(n3635), .B2(n4833), .ZN(n3636)
         );
  AOI211_X1 U4244 ( .C1(n3638), .C2(n4587), .A(n3637), .B(n3636), .ZN(n3641)
         );
  MUX2_X1 U4245 ( .A(n3639), .B(n3641), .S(n4855), .Z(n3640) );
  OAI21_X1 U4246 ( .B1(n3643), .B2(n4646), .A(n3640), .ZN(U3491) );
  MUX2_X1 U4247 ( .A(n4725), .B(n3641), .S(n4852), .Z(n3642) );
  OAI21_X1 U4248 ( .B1(n3643), .B2(n4591), .A(n3642), .ZN(U3530) );
  INV_X1 U4249 ( .A(n3644), .ZN(n3646) );
  OAI21_X1 U4250 ( .B1(n3646), .B2(n3651), .A(n3645), .ZN(n4882) );
  INV_X1 U4251 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3657) );
  OAI21_X1 U4252 ( .B1(n3648), .B2(n4121), .A(n3647), .ZN(n4881) );
  XNOR2_X1 U4253 ( .A(n3649), .B(n4121), .ZN(n3656) );
  NAND2_X1 U4254 ( .A1(n4881), .A2(n3650), .ZN(n3655) );
  OAI22_X1 U4255 ( .A1(n3652), .A2(n4834), .B1(n3651), .B2(n4833), .ZN(n3653)
         );
  AOI21_X1 U4256 ( .B1(n4838), .B2(n4180), .A(n3653), .ZN(n3654) );
  OAI211_X1 U4257 ( .C1(n4840), .C2(n3656), .A(n3655), .B(n3654), .ZN(n4888)
         );
  AOI21_X1 U4258 ( .B1(n4802), .B2(n4881), .A(n4888), .ZN(n3659) );
  MUX2_X1 U4259 ( .A(n3657), .B(n3659), .S(n4855), .Z(n3658) );
  OAI21_X1 U4260 ( .B1(n4882), .B2(n4646), .A(n3658), .ZN(U3489) );
  INV_X1 U4261 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3660) );
  MUX2_X1 U4262 ( .A(n3660), .B(n3659), .S(n4852), .Z(n3661) );
  OAI21_X1 U4263 ( .B1(n4591), .B2(n4882), .A(n3661), .ZN(U3529) );
  INV_X1 U4264 ( .A(n3662), .ZN(n3663) );
  OR2_X1 U4265 ( .A1(n3664), .A2(n3663), .ZN(n4147) );
  XNOR2_X1 U4266 ( .A(n3665), .B(n4147), .ZN(n3711) );
  INV_X1 U4267 ( .A(n4871), .ZN(n4884) );
  OAI22_X1 U4268 ( .A1(n3666), .A2(n4834), .B1(n3677), .B2(n4833), .ZN(n3674)
         );
  INV_X1 U4269 ( .A(n3667), .ZN(n3668) );
  AOI21_X1 U4270 ( .B1(n3670), .B2(n3669), .A(n3668), .ZN(n3671) );
  XNOR2_X1 U4271 ( .A(n3671), .B(n4147), .ZN(n3672) );
  NOR2_X1 U4272 ( .A1(n3672), .A2(n4840), .ZN(n3673) );
  AOI211_X1 U4273 ( .C1(n4838), .C2(n4178), .A(n3674), .B(n3673), .ZN(n3675)
         );
  OAI21_X1 U4274 ( .B1(n3711), .B2(n4452), .A(n3675), .ZN(n3712) );
  NAND2_X1 U4275 ( .A1(n3712), .A2(n4889), .ZN(n3684) );
  INV_X1 U4276 ( .A(n3691), .ZN(n3676) );
  OAI21_X1 U4277 ( .B1(n3678), .B2(n3677), .A(n3676), .ZN(n3719) );
  INV_X1 U4278 ( .A(n3719), .ZN(n3682) );
  INV_X1 U4279 ( .A(n3679), .ZN(n3680) );
  OAI22_X1 U4280 ( .A1(n4826), .A2(n4734), .B1(n3680), .B2(n4879), .ZN(n3681)
         );
  AOI21_X1 U4281 ( .B1(n3682), .B2(n4870), .A(n3681), .ZN(n3683) );
  OAI211_X1 U4282 ( .C1(n3711), .C2(n4884), .A(n3684), .B(n3683), .ZN(U3277)
         );
  INV_X1 U4283 ( .A(n3685), .ZN(n3687) );
  NAND2_X1 U4284 ( .A1(n3688), .A2(n4139), .ZN(n3721) );
  OAI21_X1 U4285 ( .B1(n3688), .B2(n4139), .A(n3721), .ZN(n4588) );
  INV_X1 U4286 ( .A(n4588), .ZN(n3698) );
  XNOR2_X1 U4287 ( .A(n4032), .B(n4139), .ZN(n3690) );
  OAI22_X1 U4288 ( .A1(n3690), .A2(n4840), .B1(n4572), .B2(n3689), .ZN(n4586)
         );
  OAI21_X1 U4289 ( .B1(n3691), .B2(n4583), .A(n3725), .ZN(n4647) );
  AOI22_X1 U4290 ( .A1(n4462), .A2(REG2_REG_14__SCAN_IN), .B1(n3692), .B2(
        n4866), .ZN(n3693) );
  OAI21_X1 U4291 ( .B1(n4583), .B2(n4433), .A(n3693), .ZN(n3694) );
  AOI21_X1 U4292 ( .B1(n4430), .B2(n4179), .A(n3694), .ZN(n3695) );
  OAI21_X1 U4293 ( .B1(n4647), .B2(n4883), .A(n3695), .ZN(n3696) );
  AOI21_X1 U4294 ( .B1(n4586), .B2(n4889), .A(n3696), .ZN(n3697) );
  OAI21_X1 U4295 ( .B1(n3698), .B2(n4502), .A(n3697), .ZN(U3276) );
  NAND2_X1 U4296 ( .A1(n4466), .A2(n4465), .ZN(n4142) );
  XOR2_X1 U4297 ( .A(n4142), .B(n3699), .Z(n4569) );
  INV_X1 U4298 ( .A(n4569), .ZN(n3710) );
  XNOR2_X1 U4299 ( .A(n4468), .B(n4142), .ZN(n3700) );
  NAND2_X1 U4300 ( .A1(n3700), .A2(n4449), .ZN(n3702) );
  NAND2_X1 U4301 ( .A1(n4174), .A2(n4838), .ZN(n3701) );
  NAND2_X1 U4302 ( .A1(n3702), .A2(n3701), .ZN(n4568) );
  INV_X1 U4303 ( .A(n4489), .ZN(n3703) );
  OAI21_X1 U4304 ( .B1(n4566), .B2(n3704), .A(n3703), .ZN(n4640) );
  NOR2_X1 U4305 ( .A1(n4640), .A2(n4883), .ZN(n3708) );
  AOI22_X1 U4306 ( .A1(n4462), .A2(REG2_REG_17__SCAN_IN), .B1(n3932), .B2(
        n4866), .ZN(n3706) );
  NAND2_X1 U4307 ( .A1(n4430), .A2(n4176), .ZN(n3705) );
  OAI211_X1 U4308 ( .C1(n4566), .C2(n4433), .A(n3706), .B(n3705), .ZN(n3707)
         );
  AOI211_X1 U4309 ( .C1(n4568), .C2(n4826), .A(n3708), .B(n3707), .ZN(n3709)
         );
  OAI21_X1 U4310 ( .B1(n3710), .B2(n4502), .A(n3709), .ZN(U3273) );
  INV_X1 U4311 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3714) );
  INV_X1 U4312 ( .A(n3711), .ZN(n3713) );
  AOI21_X1 U4313 ( .B1(n4802), .B2(n3713), .A(n3712), .ZN(n3716) );
  MUX2_X1 U4314 ( .A(n3714), .B(n3716), .S(n4852), .Z(n3715) );
  OAI21_X1 U4315 ( .B1(n4591), .B2(n3719), .A(n3715), .ZN(U3531) );
  INV_X1 U4316 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3717) );
  MUX2_X1 U4317 ( .A(n3717), .B(n3716), .S(n4855), .Z(n3718) );
  OAI21_X1 U4318 ( .B1(n3719), .B2(n4646), .A(n3718), .ZN(U3493) );
  NAND2_X1 U4319 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  XOR2_X1 U4320 ( .A(n4140), .B(n3722), .Z(n4582) );
  INV_X1 U4321 ( .A(n3723), .ZN(n3724) );
  AOI21_X1 U4322 ( .B1(n3751), .B2(n3725), .A(n3724), .ZN(n4579) );
  INV_X1 U4323 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4217) );
  OAI22_X1 U4324 ( .A1(n4889), .A2(n4217), .B1(n4911), .B2(n4879), .ZN(n3726)
         );
  AOI21_X1 U4325 ( .B1(n4430), .B2(n4178), .A(n3726), .ZN(n3727) );
  OAI21_X1 U4326 ( .B1(n4901), .B2(n4433), .A(n3727), .ZN(n3732) );
  AOI21_X1 U4327 ( .B1(n3728), .B2(n4140), .A(n4840), .ZN(n3730) );
  AOI22_X1 U4328 ( .A1(n3730), .A2(n3729), .B1(n4838), .B2(n4176), .ZN(n4581)
         );
  NOR2_X1 U4329 ( .A1(n4581), .A2(n4462), .ZN(n3731) );
  AOI211_X1 U4330 ( .C1(n4579), .C2(n4870), .A(n3732), .B(n3731), .ZN(n3733)
         );
  OAI21_X1 U4331 ( .B1(n4582), .B2(n4502), .A(n3733), .ZN(U3275) );
  MUX2_X1 U4332 ( .A(n3734), .B(REG2_REG_2__SCAN_IN), .S(n4462), .Z(n3743) );
  NAND2_X1 U4333 ( .A1(n3735), .A2(n4871), .ZN(n3741) );
  AOI22_X1 U4334 ( .A1(n4870), .A2(n3736), .B1(REG3_REG_2__SCAN_IN), .B2(n4866), .ZN(n3740) );
  AOI22_X1 U4335 ( .A1(n3738), .A2(n3737), .B1(n4430), .B2(n3194), .ZN(n3739)
         );
  NAND3_X1 U4336 ( .A1(n3741), .A2(n3740), .A3(n3739), .ZN(n3742) );
  OR2_X1 U4337 ( .A1(n3743), .A2(n3742), .ZN(U3288) );
  NAND2_X1 U4338 ( .A1(n4177), .A2(n2274), .ZN(n3749) );
  NAND2_X1 U4339 ( .A1(n3751), .A2(n2277), .ZN(n3748) );
  NAND2_X1 U4340 ( .A1(n3749), .A2(n3748), .ZN(n3750) );
  XNOR2_X1 U4341 ( .A(n3750), .B(n3835), .ZN(n4905) );
  NAND2_X1 U4342 ( .A1(n4177), .A2(n3854), .ZN(n3753) );
  NAND2_X1 U4343 ( .A1(n3751), .A2(n2280), .ZN(n3752) );
  NAND2_X1 U4344 ( .A1(n4176), .A2(n2274), .ZN(n3755) );
  NAND2_X1 U4345 ( .A1(n3757), .A2(n2277), .ZN(n3754) );
  NAND2_X1 U4346 ( .A1(n3755), .A2(n3754), .ZN(n3756) );
  XNOR2_X1 U4347 ( .A(n3756), .B(n3855), .ZN(n3760) );
  NAND2_X1 U4348 ( .A1(n4176), .A2(n3854), .ZN(n3759) );
  NAND2_X1 U4349 ( .A1(n3757), .A2(n2273), .ZN(n3758) );
  NAND2_X1 U4350 ( .A1(n3759), .A2(n3758), .ZN(n3761) );
  NAND2_X1 U4351 ( .A1(n3760), .A2(n3761), .ZN(n3914) );
  OAI21_X1 U4352 ( .B1(n4905), .B2(n4904), .A(n3914), .ZN(n3765) );
  NAND3_X1 U4353 ( .A1(n3914), .A2(n4904), .A3(n4905), .ZN(n3764) );
  INV_X1 U4354 ( .A(n3760), .ZN(n3763) );
  INV_X1 U4355 ( .A(n3761), .ZN(n3762) );
  NAND2_X1 U4356 ( .A1(n3763), .A2(n3762), .ZN(n3913) );
  NAND2_X1 U4357 ( .A1(n4175), .A2(n2280), .ZN(n3767) );
  NAND2_X1 U4358 ( .A1(n3769), .A2(n2276), .ZN(n3766) );
  NAND2_X1 U4359 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  XNOR2_X1 U4360 ( .A(n3768), .B(n3855), .ZN(n3773) );
  NAND2_X1 U4361 ( .A1(n4175), .A2(n3854), .ZN(n3771) );
  NAND2_X1 U4362 ( .A1(n3769), .A2(n2280), .ZN(n3770) );
  NAND2_X1 U4363 ( .A1(n3771), .A2(n3770), .ZN(n3772) );
  NAND2_X1 U4364 ( .A1(n3773), .A2(n3772), .ZN(n3927) );
  NAND2_X1 U4365 ( .A1(n4174), .A2(n2273), .ZN(n3775) );
  INV_X1 U4366 ( .A(n4490), .ZN(n3777) );
  NAND2_X1 U4367 ( .A1(n3777), .A2(n2277), .ZN(n3774) );
  NAND2_X1 U4368 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  XNOR2_X1 U4369 ( .A(n3776), .B(n3855), .ZN(n3992) );
  NAND2_X1 U4370 ( .A1(n4174), .A2(n3854), .ZN(n3779) );
  NAND2_X1 U4371 ( .A1(n3777), .A2(n2280), .ZN(n3778) );
  NAND2_X1 U4372 ( .A1(n3779), .A2(n3778), .ZN(n3780) );
  INV_X1 U4373 ( .A(n3992), .ZN(n3781) );
  INV_X1 U4374 ( .A(n3780), .ZN(n3991) );
  NAND2_X1 U4375 ( .A1(n4496), .A2(n2273), .ZN(n3785) );
  NAND2_X1 U4376 ( .A1(n3783), .A2(n2277), .ZN(n3784) );
  NAND2_X1 U4377 ( .A1(n3785), .A2(n3784), .ZN(n3786) );
  XNOR2_X1 U4378 ( .A(n3786), .B(n3835), .ZN(n3789) );
  NOR2_X1 U4379 ( .A1(n4480), .A2(n2279), .ZN(n3787) );
  AOI21_X1 U4380 ( .B1(n4496), .B2(n3854), .A(n3787), .ZN(n3788) );
  NAND2_X1 U4381 ( .A1(n3789), .A2(n3788), .ZN(n3894) );
  OAI21_X1 U4382 ( .B1(n3789), .B2(n3788), .A(n3894), .ZN(n3888) );
  NAND2_X1 U4383 ( .A1(n4547), .A2(n2273), .ZN(n3791) );
  NAND2_X1 U4384 ( .A1(n4444), .A2(n2276), .ZN(n3790) );
  NAND2_X1 U4385 ( .A1(n3791), .A2(n3790), .ZN(n3792) );
  XNOR2_X1 U4386 ( .A(n3792), .B(n3855), .ZN(n3804) );
  NAND2_X1 U4387 ( .A1(n4547), .A2(n3854), .ZN(n3794) );
  NAND2_X1 U4388 ( .A1(n4444), .A2(n2274), .ZN(n3793) );
  NAND2_X1 U4389 ( .A1(n3794), .A2(n3793), .ZN(n3805) );
  NAND2_X1 U4390 ( .A1(n3804), .A2(n3805), .ZN(n3970) );
  INV_X1 U4391 ( .A(n3970), .ZN(n3796) );
  OR2_X1 U4392 ( .A1(n3888), .A2(n3796), .ZN(n3795) );
  NOR2_X1 U4393 ( .A1(n3886), .A2(n3795), .ZN(n3798) );
  NOR2_X1 U4394 ( .A1(n3796), .A2(n3894), .ZN(n3797) );
  NOR2_X1 U4395 ( .A1(n3798), .A2(n3797), .ZN(n3810) );
  NOR2_X1 U4396 ( .A1(n3837), .A2(n4548), .ZN(n3799) );
  AOI21_X1 U4397 ( .B1(n4445), .B2(n3854), .A(n3799), .ZN(n3897) );
  NAND2_X1 U4398 ( .A1(n4445), .A2(n2274), .ZN(n3802) );
  NAND2_X1 U4399 ( .A1(n3800), .A2(n2276), .ZN(n3801) );
  NAND2_X1 U4400 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  XNOR2_X1 U4401 ( .A(n3803), .B(n3835), .ZN(n3896) );
  INV_X1 U4402 ( .A(n3804), .ZN(n3807) );
  INV_X1 U4403 ( .A(n3805), .ZN(n3806) );
  AND2_X1 U4404 ( .A1(n3807), .A2(n3806), .ZN(n3969) );
  AOI21_X1 U4405 ( .B1(n3897), .B2(n3896), .A(n3969), .ZN(n3809) );
  NOR2_X1 U4406 ( .A1(n3896), .A2(n3897), .ZN(n3808) );
  AOI21_X1 U4407 ( .B1(n3810), .B2(n3809), .A(n3808), .ZN(n3980) );
  AOI22_X1 U4408 ( .A1(n4425), .A2(n3854), .B1(n2274), .B2(n3811), .ZN(n3816)
         );
  AOI22_X1 U4409 ( .A1(n4425), .A2(n2273), .B1(n2277), .B2(n3811), .ZN(n3812)
         );
  XNOR2_X1 U4410 ( .A(n3812), .B(n3855), .ZN(n3815) );
  XOR2_X1 U4411 ( .A(n3816), .B(n3815), .Z(n3981) );
  NOR2_X1 U4412 ( .A1(n2279), .A2(n4395), .ZN(n3813) );
  AOI21_X1 U4413 ( .B1(n4405), .B2(n3854), .A(n3813), .ZN(n3821) );
  XNOR2_X1 U4414 ( .A(n3814), .B(n3855), .ZN(n3820) );
  XOR2_X1 U4415 ( .A(n3821), .B(n3820), .Z(n3876) );
  INV_X1 U4416 ( .A(n3815), .ZN(n3818) );
  INV_X1 U4417 ( .A(n3816), .ZN(n3817) );
  NOR2_X1 U4418 ( .A1(n3818), .A2(n3817), .ZN(n3877) );
  NOR2_X1 U4419 ( .A1(n3876), .A2(n3877), .ZN(n3819) );
  INV_X1 U4420 ( .A(n3820), .ZN(n3822) );
  NAND2_X1 U4421 ( .A1(n4389), .A2(n2281), .ZN(n3825) );
  NAND2_X1 U4422 ( .A1(n3823), .A2(n2276), .ZN(n3824) );
  NAND2_X1 U4423 ( .A1(n3825), .A2(n3824), .ZN(n3826) );
  XNOR2_X1 U4424 ( .A(n3826), .B(n3835), .ZN(n3829) );
  OAI22_X1 U4425 ( .A1(n4345), .A2(n3827), .B1(n3837), .B2(n4369), .ZN(n3937)
         );
  AOI22_X1 U4426 ( .A1(n4364), .A2(n2280), .B1(n2277), .B2(n3839), .ZN(n3831)
         );
  XNOR2_X1 U4427 ( .A(n3831), .B(n3855), .ZN(n3906) );
  NAND2_X1 U4428 ( .A1(n4347), .A2(n2273), .ZN(n3834) );
  NAND2_X1 U4429 ( .A1(n3832), .A2(n2276), .ZN(n3833) );
  NAND2_X1 U4430 ( .A1(n3834), .A2(n3833), .ZN(n3836) );
  XNOR2_X1 U4431 ( .A(n3836), .B(n3835), .ZN(n3841) );
  NOR2_X1 U4432 ( .A1(n2279), .A2(n4524), .ZN(n3838) );
  AOI21_X1 U4433 ( .B1(n4347), .B2(n3854), .A(n3838), .ZN(n3840) );
  NOR2_X1 U4434 ( .A1(n3841), .A2(n3840), .ZN(n4007) );
  AOI22_X1 U4435 ( .A1(n4364), .A2(n3854), .B1(n2281), .B2(n3839), .ZN(n3905)
         );
  AOI21_X2 U4436 ( .B1(n3904), .B2(n3906), .A(n3905), .ZN(n4004) );
  NAND2_X1 U4437 ( .A1(n3841), .A2(n3840), .ZN(n4005) );
  INV_X1 U4438 ( .A(n3867), .ZN(n3851) );
  NAND2_X1 U4439 ( .A1(n4324), .A2(n2274), .ZN(n3843) );
  NAND2_X1 U4440 ( .A1(n3845), .A2(n2277), .ZN(n3842) );
  NAND2_X1 U4441 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  XNOR2_X1 U4442 ( .A(n3844), .B(n3855), .ZN(n3849) );
  NAND2_X1 U4443 ( .A1(n4324), .A2(n3854), .ZN(n3847) );
  NAND2_X1 U4444 ( .A1(n3845), .A2(n2274), .ZN(n3846) );
  NAND2_X1 U4445 ( .A1(n3847), .A2(n3846), .ZN(n3848) );
  NAND2_X1 U4446 ( .A1(n3849), .A2(n3848), .ZN(n3852) );
  OAI21_X1 U4447 ( .B1(n3849), .B2(n3848), .A(n3852), .ZN(n3868) );
  INV_X1 U4448 ( .A(n3868), .ZN(n3850) );
  NAND2_X1 U4449 ( .A1(n3851), .A2(n3850), .ZN(n3869) );
  NAND2_X1 U4450 ( .A1(n3869), .A2(n3852), .ZN(n3860) );
  AOI22_X1 U4451 ( .A1(n4299), .A2(n2280), .B1(n2276), .B2(n3853), .ZN(n3858)
         );
  AOI22_X1 U4452 ( .A1(n4299), .A2(n3854), .B1(n2273), .B2(n3853), .ZN(n3856)
         );
  XNOR2_X1 U4453 ( .A(n3856), .B(n3855), .ZN(n3857) );
  XOR2_X1 U4454 ( .A(n3858), .B(n3857), .Z(n3859) );
  XNOR2_X1 U4455 ( .A(n3860), .B(n3859), .ZN(n3866) );
  OAI22_X1 U4456 ( .A1(n3996), .A2(n4288), .B1(STATE_REG_SCAN_IN), .B2(n3861), 
        .ZN(n3864) );
  INV_X1 U4457 ( .A(n4292), .ZN(n3862) );
  OAI22_X1 U4458 ( .A1(n3862), .A2(n4897), .B1(n4896), .B2(n4011), .ZN(n3863)
         );
  AOI211_X1 U4459 ( .C1(n4014), .C2(n4283), .A(n3864), .B(n3863), .ZN(n3865)
         );
  OAI21_X1 U4460 ( .B1(n3866), .B2(n4016), .A(n3865), .ZN(U3217) );
  NAND2_X1 U4461 ( .A1(n3870), .A2(n3869), .ZN(n3875) );
  AOI22_X1 U4462 ( .A1(n3994), .A2(n4299), .B1(n3995), .B2(n4347), .ZN(n3874)
         );
  OAI22_X1 U4463 ( .A1(n3996), .A2(n4517), .B1(STATE_REG_SCAN_IN), .B2(n3871), 
        .ZN(n3872) );
  AOI21_X1 U4464 ( .B1(n4014), .B2(n4302), .A(n3872), .ZN(n3873) );
  NAND3_X1 U4465 ( .A1(n3875), .A2(n3874), .A3(n3873), .ZN(U3211) );
  INV_X1 U4466 ( .A(n3979), .ZN(n3878) );
  OAI21_X1 U4467 ( .B1(n3878), .B2(n3877), .A(n3876), .ZN(n3880) );
  NAND3_X1 U4468 ( .A1(n3880), .A2(n4907), .A3(n3879), .ZN(n3885) );
  AOI22_X1 U4469 ( .A1(n3994), .A2(n4389), .B1(n3995), .B2(n4425), .ZN(n3884)
         );
  OAI22_X1 U4470 ( .A1(n3996), .A2(n4395), .B1(STATE_REG_SCAN_IN), .B2(n3881), 
        .ZN(n3882) );
  AOI21_X1 U4471 ( .B1(n4014), .B2(n4396), .A(n3882), .ZN(n3883) );
  NAND3_X1 U4472 ( .A1(n3885), .A2(n3884), .A3(n3883), .ZN(U3213) );
  INV_X1 U4473 ( .A(n3895), .ZN(n3887) );
  AOI21_X1 U4474 ( .B1(n3886), .B2(n3888), .A(n3887), .ZN(n3893) );
  AOI22_X1 U4475 ( .A1(n3995), .A2(n4174), .B1(n3994), .B2(n4547), .ZN(n3892)
         );
  NOR2_X1 U4476 ( .A1(STATE_REG_SCAN_IN), .A2(n3889), .ZN(n4763) );
  NOR2_X1 U4477 ( .A1(n3996), .A2(n4480), .ZN(n3890) );
  AOI211_X1 U4478 ( .C1(n4014), .C2(n4482), .A(n4763), .B(n3890), .ZN(n3891)
         );
  OAI211_X1 U4479 ( .C1(n3893), .C2(n4016), .A(n3892), .B(n3891), .ZN(U3216)
         );
  NAND2_X1 U4480 ( .A1(n3895), .A2(n3894), .ZN(n3973) );
  OAI21_X1 U4481 ( .B1(n3973), .B2(n3969), .A(n3970), .ZN(n3899) );
  XOR2_X1 U4482 ( .A(n3897), .B(n3896), .Z(n3898) );
  XNOR2_X1 U4483 ( .A(n3899), .B(n3898), .ZN(n3903) );
  AOI22_X1 U4484 ( .A1(n3995), .A2(n4547), .B1(n3994), .B2(n4425), .ZN(n3902)
         );
  OAI22_X1 U4485 ( .A1(n3996), .A2(n4548), .B1(STATE_REG_SCAN_IN), .B2(n2805), 
        .ZN(n3900) );
  AOI21_X1 U4486 ( .B1(n4014), .B2(n4429), .A(n3900), .ZN(n3901) );
  OAI211_X1 U4487 ( .C1(n3903), .C2(n4016), .A(n3902), .B(n3901), .ZN(U3220)
         );
  XNOR2_X1 U4488 ( .A(n3906), .B(n3905), .ZN(n3907) );
  XNOR2_X1 U4489 ( .A(n3904), .B(n3907), .ZN(n3912) );
  OAI22_X1 U4490 ( .A1(n3996), .A2(n4350), .B1(STATE_REG_SCAN_IN), .B2(n3908), 
        .ZN(n3910) );
  OAI22_X1 U4491 ( .A1(n4345), .A2(n4896), .B1(n4897), .B2(n4518), .ZN(n3909)
         );
  AOI211_X1 U4492 ( .C1(n4014), .C2(n4352), .A(n3910), .B(n3909), .ZN(n3911)
         );
  OAI21_X1 U4493 ( .B1(n3912), .B2(n4016), .A(n3911), .ZN(U3222) );
  NAND2_X1 U4494 ( .A1(n3914), .A2(n3913), .ZN(n3920) );
  INV_X1 U4495 ( .A(n4904), .ZN(n3916) );
  NOR2_X1 U4496 ( .A1(n3915), .A2(n3916), .ZN(n3918) );
  INV_X1 U4497 ( .A(n3915), .ZN(n3917) );
  OAI22_X1 U4498 ( .A1(n3918), .A2(n4905), .B1(n3917), .B2(n4904), .ZN(n3919)
         );
  XOR2_X1 U4499 ( .A(n3920), .B(n3919), .Z(n3926) );
  AOI22_X1 U4500 ( .A1(n3995), .A2(n4177), .B1(n3994), .B2(n4175), .ZN(n3925)
         );
  NOR2_X1 U4501 ( .A1(STATE_REG_SCAN_IN), .A2(n3921), .ZN(n4752) );
  NOR2_X1 U4502 ( .A1(n3996), .A2(n4571), .ZN(n3922) );
  AOI211_X1 U4503 ( .C1(n4014), .C2(n3923), .A(n4752), .B(n3922), .ZN(n3924)
         );
  OAI211_X1 U4504 ( .C1(n3926), .C2(n4016), .A(n3925), .B(n3924), .ZN(U3223)
         );
  NAND2_X1 U4505 ( .A1(n2310), .A2(n3927), .ZN(n3928) );
  XNOR2_X1 U4506 ( .A(n3929), .B(n3928), .ZN(n3935) );
  AOI22_X1 U4507 ( .A1(n3995), .A2(n4176), .B1(n3994), .B2(n4174), .ZN(n3934)
         );
  NOR2_X1 U4508 ( .A1(STATE_REG_SCAN_IN), .A2(n3930), .ZN(n4249) );
  NOR2_X1 U4509 ( .A1(n3996), .A2(n4566), .ZN(n3931) );
  AOI211_X1 U4510 ( .C1(n4014), .C2(n3932), .A(n4249), .B(n3931), .ZN(n3933)
         );
  OAI211_X1 U4511 ( .C1(n3935), .C2(n4016), .A(n3934), .B(n3933), .ZN(U3225)
         );
  NOR2_X1 U4512 ( .A1(n2291), .A2(n3936), .ZN(n3938) );
  XNOR2_X1 U4513 ( .A(n3938), .B(n3937), .ZN(n3944) );
  OAI22_X1 U4514 ( .A1(n3996), .A2(n4369), .B1(STATE_REG_SCAN_IN), .B2(n3939), 
        .ZN(n3941) );
  INV_X1 U4515 ( .A(n4364), .ZN(n4525) );
  OAI22_X1 U4516 ( .A1(n4362), .A2(n4896), .B1(n4897), .B2(n4525), .ZN(n3940)
         );
  AOI211_X1 U4517 ( .C1(n4014), .C2(n3942), .A(n3941), .B(n3940), .ZN(n3943)
         );
  OAI21_X1 U4518 ( .B1(n3944), .B2(n4016), .A(n3943), .ZN(U3226) );
  INV_X1 U4519 ( .A(n3945), .ZN(n3950) );
  OAI21_X1 U4520 ( .B1(n3948), .B2(n3947), .A(n3946), .ZN(n3949) );
  NAND3_X1 U4521 ( .A1(n3950), .A2(n4907), .A3(n3949), .ZN(n3957) );
  AOI22_X1 U4522 ( .A1(n3995), .A2(n2433), .B1(n3994), .B2(n4186), .ZN(n3956)
         );
  NOR2_X1 U4523 ( .A1(n3996), .A2(n3951), .ZN(n3953) );
  AOI211_X1 U4524 ( .C1(n4014), .C2(n3954), .A(n3953), .B(n3952), .ZN(n3955)
         );
  NAND3_X1 U4525 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(U3227) );
  OAI21_X1 U4526 ( .B1(n3960), .B2(n3959), .A(n3958), .ZN(n3961) );
  NAND2_X1 U4527 ( .A1(n3961), .A2(n4907), .ZN(n3968) );
  AOI22_X1 U4528 ( .A1(n3995), .A2(n4837), .B1(n3994), .B2(n4182), .ZN(n3967)
         );
  NOR2_X1 U4529 ( .A1(n3996), .A2(n3962), .ZN(n3964) );
  AOI211_X1 U4530 ( .C1(n4014), .C2(n3965), .A(n3964), .B(n3963), .ZN(n3966)
         );
  NAND3_X1 U4531 ( .A1(n3968), .A2(n3967), .A3(n3966), .ZN(U3228) );
  INV_X1 U4532 ( .A(n3969), .ZN(n3971) );
  NAND2_X1 U4533 ( .A1(n3971), .A2(n3970), .ZN(n3972) );
  XNOR2_X1 U4534 ( .A(n3973), .B(n3972), .ZN(n3978) );
  OAI22_X1 U4535 ( .A1(n3996), .A2(n4456), .B1(STATE_REG_SCAN_IN), .B2(n3974), 
        .ZN(n3976) );
  OAI22_X1 U4536 ( .A1(n3984), .A2(n4897), .B1(n4896), .B2(n4447), .ZN(n3975)
         );
  AOI211_X1 U4537 ( .C1(n4014), .C2(n4458), .A(n3976), .B(n3975), .ZN(n3977)
         );
  OAI21_X1 U4538 ( .B1(n3978), .B2(n4016), .A(n3977), .ZN(U3230) );
  OAI21_X1 U4539 ( .B1(n3981), .B2(n3980), .A(n3979), .ZN(n3982) );
  NAND2_X1 U4540 ( .A1(n3982), .A2(n4907), .ZN(n3989) );
  OAI22_X1 U4541 ( .A1(n3996), .A2(n4415), .B1(STATE_REG_SCAN_IN), .B2(n3983), 
        .ZN(n3986) );
  OAI22_X1 U4542 ( .A1(n4362), .A2(n4897), .B1(n4896), .B2(n3984), .ZN(n3985)
         );
  AOI211_X1 U4543 ( .C1(n4014), .C2(n3987), .A(n3986), .B(n3985), .ZN(n3988)
         );
  NAND2_X1 U4544 ( .A1(n3989), .A2(n3988), .ZN(U3232) );
  XNOR2_X1 U4545 ( .A(n3992), .B(n3991), .ZN(n3993) );
  XNOR2_X1 U4546 ( .A(n3990), .B(n3993), .ZN(n4002) );
  AOI22_X1 U4547 ( .A1(n3995), .A2(n4175), .B1(n3994), .B2(n4496), .ZN(n4001)
         );
  NOR2_X1 U4548 ( .A1(n3996), .A2(n4490), .ZN(n3998) );
  INV_X1 U4549 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3997) );
  NOR2_X1 U4550 ( .A1(STATE_REG_SCAN_IN), .A2(n3997), .ZN(n4258) );
  AOI211_X1 U4551 ( .C1(n4014), .C2(n3999), .A(n3998), .B(n4258), .ZN(n4000)
         );
  OAI211_X1 U4552 ( .C1(n4002), .C2(n4016), .A(n4001), .B(n4000), .ZN(U3235)
         );
  OR2_X1 U4553 ( .A1(n4004), .A2(n4003), .ZN(n4009) );
  INV_X1 U4554 ( .A(n4005), .ZN(n4006) );
  NOR2_X1 U4555 ( .A1(n4007), .A2(n4006), .ZN(n4008) );
  XNOR2_X1 U4556 ( .A(n4009), .B(n4008), .ZN(n4017) );
  INV_X1 U4557 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4010) );
  OAI22_X1 U4558 ( .A1(n3996), .A2(n4524), .B1(STATE_REG_SCAN_IN), .B2(n4010), 
        .ZN(n4013) );
  OAI22_X1 U4559 ( .A1(n4525), .A2(n4896), .B1(n4897), .B2(n4011), .ZN(n4012)
         );
  AOI211_X1 U4560 ( .C1(n4014), .C2(n4330), .A(n4013), .B(n4012), .ZN(n4015)
         );
  OAI21_X1 U4561 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(U3237) );
  NAND2_X1 U4562 ( .A1(n2270), .A2(DATAI_31_), .ZN(n4269) );
  INV_X1 U4563 ( .A(n4269), .ZN(n4272) );
  OAI22_X1 U4564 ( .A1(n4022), .A2(n4047), .B1(n4173), .B2(n4269), .ZN(n4148)
         );
  NAND2_X1 U4565 ( .A1(n4019), .A2(n4018), .ZN(n4042) );
  INV_X1 U4566 ( .A(n4020), .ZN(n4021) );
  AOI21_X1 U4567 ( .B1(n4292), .B2(n4280), .A(n4021), .ZN(n4114) );
  NAND2_X1 U4568 ( .A1(n4022), .A2(n4047), .ZN(n4023) );
  NAND2_X1 U4569 ( .A1(n4173), .A2(n4269), .ZN(n4117) );
  NAND2_X1 U4570 ( .A1(n4023), .A2(n4117), .ZN(n4146) );
  NOR2_X1 U4571 ( .A1(n4292), .A2(n4280), .ZN(n4024) );
  OR2_X1 U4572 ( .A1(n4146), .A2(n4024), .ZN(n4040) );
  AOI21_X1 U4573 ( .B1(n4042), .B2(n4114), .A(n4040), .ZN(n4116) );
  NAND3_X1 U4574 ( .A1(n4114), .A2(n4297), .A3(n2359), .ZN(n4045) );
  INV_X1 U4575 ( .A(n4025), .ZN(n4026) );
  NOR2_X1 U4576 ( .A1(n4130), .A2(n4026), .ZN(n4105) );
  NAND2_X1 U4577 ( .A1(n4027), .A2(n4030), .ZN(n4062) );
  NAND2_X1 U4578 ( .A1(n4029), .A2(n4028), .ZN(n4090) );
  AND2_X1 U4579 ( .A1(n4090), .A2(n4030), .ZN(n4095) );
  INV_X1 U4580 ( .A(n4095), .ZN(n4031) );
  OAI211_X1 U4581 ( .C1(n4032), .C2(n4062), .A(n4099), .B(n4031), .ZN(n4033)
         );
  AND2_X1 U4582 ( .A1(n4033), .A2(n4096), .ZN(n4036) );
  OR2_X1 U4583 ( .A1(n4035), .A2(n4034), .ZN(n4101) );
  OAI21_X1 U4584 ( .B1(n4036), .B2(n4101), .A(n4100), .ZN(n4038) );
  OAI21_X1 U4585 ( .B1(n4103), .B2(n4038), .A(n4037), .ZN(n4039) );
  AOI21_X1 U4586 ( .B1(n4105), .B2(n4039), .A(n2358), .ZN(n4043) );
  NOR4_X1 U4587 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  AOI21_X1 U4588 ( .B1(n4116), .B2(n4045), .A(n4044), .ZN(n4046) );
  AOI21_X1 U4589 ( .B1(n4048), .B2(n4047), .A(n4046), .ZN(n4049) );
  AOI21_X1 U4590 ( .B1(n4272), .B2(n4148), .A(n4049), .ZN(n4050) );
  XNOR2_X1 U4591 ( .A(n4050), .B(n4766), .ZN(n4165) );
  INV_X1 U4592 ( .A(n4051), .ZN(n4164) );
  NAND2_X1 U4593 ( .A1(n4053), .A2(n4052), .ZN(n4054) );
  NOR2_X1 U4594 ( .A1(n4054), .A2(n4084), .ZN(n4088) );
  INV_X1 U4595 ( .A(n4079), .ZN(n4056) );
  NOR2_X1 U4596 ( .A1(n4056), .A2(n4055), .ZN(n4059) );
  INV_X1 U4597 ( .A(n4057), .ZN(n4058) );
  AOI21_X1 U4598 ( .B1(n4088), .B2(n4059), .A(n4058), .ZN(n4065) );
  NAND2_X1 U4599 ( .A1(n4061), .A2(n4060), .ZN(n4092) );
  INV_X1 U4600 ( .A(n4062), .ZN(n4064) );
  OAI211_X1 U4601 ( .C1(n4065), .C2(n4092), .A(n4064), .B(n4063), .ZN(n4066)
         );
  INV_X1 U4602 ( .A(n4066), .ZN(n4094) );
  OAI211_X1 U4603 ( .C1(n4069), .C2(n4157), .A(n4068), .B(n4067), .ZN(n4072)
         );
  NAND3_X1 U4604 ( .A1(n4072), .A2(n4071), .A3(n4070), .ZN(n4075) );
  NAND3_X1 U4605 ( .A1(n4075), .A2(n4074), .A3(n4073), .ZN(n4077) );
  NAND2_X1 U4606 ( .A1(n4077), .A2(n4076), .ZN(n4080) );
  NAND4_X1 U4607 ( .A1(n4080), .A2(n4079), .A3(n2304), .A4(n4078), .ZN(n4083)
         );
  NAND3_X1 U4608 ( .A1(n4083), .A2(n4082), .A3(n4081), .ZN(n4089) );
  AOI21_X1 U4609 ( .B1(n4086), .B2(n4085), .A(n4084), .ZN(n4087) );
  AOI21_X1 U4610 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4091) );
  OR2_X1 U4611 ( .A1(n4091), .A2(n4090), .ZN(n4093) );
  OAI22_X1 U4612 ( .A1(n4095), .A2(n4094), .B1(n4093), .B2(n4092), .ZN(n4098)
         );
  INV_X1 U4613 ( .A(n4096), .ZN(n4097) );
  AOI21_X1 U4614 ( .B1(n4099), .B2(n4098), .A(n4097), .ZN(n4102) );
  OAI21_X1 U4615 ( .B1(n4102), .B2(n4101), .A(n4100), .ZN(n4104) );
  AOI21_X1 U4616 ( .B1(n4384), .B2(n4104), .A(n4103), .ZN(n4106) );
  OAI21_X1 U4617 ( .B1(n4107), .B2(n4106), .A(n4105), .ZN(n4109) );
  NAND2_X1 U4618 ( .A1(n4109), .A2(n4108), .ZN(n4111) );
  AOI211_X1 U4619 ( .C1(n4112), .C2(n4111), .A(n4110), .B(n4148), .ZN(n4115)
         );
  AND3_X1 U4620 ( .A1(n4115), .A2(n4114), .A3(n4113), .ZN(n4119) );
  AOI21_X1 U4621 ( .B1(n4148), .B2(n4117), .A(n4116), .ZN(n4118) );
  OAI21_X1 U4622 ( .B1(n4119), .B2(n4118), .A(n3046), .ZN(n4160) );
  NOR4_X1 U4623 ( .A1(n4122), .A2(n4121), .A3(n4830), .A4(n4120), .ZN(n4137)
         );
  NAND2_X1 U4624 ( .A1(n4124), .A2(n4123), .ZN(n4442) );
  NOR4_X1 U4625 ( .A1(n4127), .A2(n4442), .A3(n4126), .A4(n4125), .ZN(n4136)
         );
  NOR4_X1 U4626 ( .A1(n4289), .A2(n4128), .A3(n4403), .A4(n4781), .ZN(n4135)
         );
  INV_X1 U4627 ( .A(n4341), .ZN(n4129) );
  OR2_X1 U4628 ( .A1(n4130), .A2(n4129), .ZN(n4360) );
  NAND2_X1 U4629 ( .A1(n4319), .A2(n4131), .ZN(n4344) );
  NOR4_X1 U4630 ( .A1(n4360), .A2(n4133), .A3(n4132), .A4(n4344), .ZN(n4134)
         );
  NAND4_X1 U4631 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4154)
         );
  NOR4_X1 U4632 ( .A1(n4141), .A2(n4140), .A3(n4139), .A4(n4138), .ZN(n4144)
         );
  NAND2_X1 U4633 ( .A1(n4382), .A2(n4384), .ZN(n4421) );
  XNOR2_X1 U4634 ( .A(n4496), .B(n4480), .ZN(n4473) );
  NOR4_X1 U4635 ( .A1(n4499), .A2(n4421), .A3(n4473), .A4(n4142), .ZN(n4143)
         );
  NAND2_X1 U4636 ( .A1(n4144), .A2(n4143), .ZN(n4145) );
  NOR4_X1 U4637 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4151)
         );
  NAND2_X1 U4638 ( .A1(n2359), .A2(n4149), .ZN(n4317) );
  INV_X1 U4639 ( .A(n4317), .ZN(n4321) );
  NAND4_X1 U4640 ( .A1(n4151), .A2(n4150), .A3(n4297), .A4(n4321), .ZN(n4153)
         );
  XNOR2_X1 U4641 ( .A(n4405), .B(n4388), .ZN(n4380) );
  INV_X1 U4642 ( .A(n4380), .ZN(n4386) );
  NAND3_X1 U4643 ( .A1(n4158), .A2(n4652), .A3(n4155), .ZN(n4156) );
  NAND2_X1 U4644 ( .A1(n4160), .A2(n4156), .ZN(n4162) );
  OAI21_X1 U4645 ( .B1(n4158), .B2(n4157), .A(n4652), .ZN(n4159) );
  AND2_X1 U4646 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  MUX2_X1 U4647 ( .A(n4162), .B(n4161), .S(n4829), .Z(n4163) );
  AOI21_X1 U4648 ( .B1(n4165), .B2(n4164), .A(n4163), .ZN(n4172) );
  NOR4_X1 U4649 ( .A1(n4916), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4169)
         );
  NAND2_X1 U4650 ( .A1(n4169), .A2(n2273), .ZN(n4170) );
  OAI211_X1 U4651 ( .C1(n4651), .C2(n4656), .A(n4170), .B(B_REG_SCAN_IN), .ZN(
        n4171) );
  OAI21_X1 U4652 ( .B1(n4172), .B2(n4656), .A(n4171), .ZN(U3239) );
  MUX2_X1 U4653 ( .A(n4173), .B(DATAO_REG_31__SCAN_IN), .S(n4189), .Z(U3581)
         );
  MUX2_X1 U4654 ( .A(n4292), .B(DATAO_REG_29__SCAN_IN), .S(n4189), .Z(U3579)
         );
  MUX2_X1 U4655 ( .A(n4299), .B(DATAO_REG_28__SCAN_IN), .S(n4189), .Z(U3578)
         );
  MUX2_X1 U4656 ( .A(n4324), .B(DATAO_REG_27__SCAN_IN), .S(n4189), .Z(U3577)
         );
  MUX2_X1 U4657 ( .A(n4347), .B(DATAO_REG_26__SCAN_IN), .S(n4189), .Z(U3576)
         );
  MUX2_X1 U4658 ( .A(n4364), .B(DATAO_REG_25__SCAN_IN), .S(n4189), .Z(U3575)
         );
  MUX2_X1 U4659 ( .A(n4389), .B(DATAO_REG_24__SCAN_IN), .S(n4189), .Z(U3574)
         );
  MUX2_X1 U4660 ( .A(n4405), .B(DATAO_REG_23__SCAN_IN), .S(n4189), .Z(U3573)
         );
  MUX2_X1 U4661 ( .A(n4425), .B(DATAO_REG_22__SCAN_IN), .S(n4189), .Z(U3572)
         );
  MUX2_X1 U4662 ( .A(n4445), .B(DATAO_REG_21__SCAN_IN), .S(n4189), .Z(U3571)
         );
  MUX2_X1 U4663 ( .A(n4547), .B(DATAO_REG_20__SCAN_IN), .S(n4189), .Z(U3570)
         );
  MUX2_X1 U4664 ( .A(n4496), .B(DATAO_REG_19__SCAN_IN), .S(n4189), .Z(U3569)
         );
  MUX2_X1 U4665 ( .A(n4174), .B(DATAO_REG_18__SCAN_IN), .S(n4189), .Z(U3568)
         );
  MUX2_X1 U4666 ( .A(n4175), .B(DATAO_REG_17__SCAN_IN), .S(n4189), .Z(U3567)
         );
  MUX2_X1 U4667 ( .A(n4176), .B(DATAO_REG_16__SCAN_IN), .S(n4189), .Z(U3566)
         );
  MUX2_X1 U4668 ( .A(n4177), .B(DATAO_REG_15__SCAN_IN), .S(n4189), .Z(U3565)
         );
  MUX2_X1 U4669 ( .A(n4178), .B(DATAO_REG_14__SCAN_IN), .S(n4189), .Z(U3564)
         );
  MUX2_X1 U4670 ( .A(n4179), .B(DATAO_REG_13__SCAN_IN), .S(n4189), .Z(U3563)
         );
  MUX2_X1 U4671 ( .A(DATAO_REG_12__SCAN_IN), .B(n4180), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4672 ( .A(n4181), .B(DATAO_REG_11__SCAN_IN), .S(n4189), .Z(U3561)
         );
  MUX2_X1 U4673 ( .A(DATAO_REG_10__SCAN_IN), .B(n4182), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4674 ( .A(DATAO_REG_9__SCAN_IN), .B(n4183), .S(U4043), .Z(U3559) );
  MUX2_X1 U4675 ( .A(DATAO_REG_8__SCAN_IN), .B(n4837), .S(U4043), .Z(U3558) );
  MUX2_X1 U4676 ( .A(n4184), .B(DATAO_REG_7__SCAN_IN), .S(n4189), .Z(U3557) );
  MUX2_X1 U4677 ( .A(n4185), .B(DATAO_REG_6__SCAN_IN), .S(n4189), .Z(U3556) );
  MUX2_X1 U4678 ( .A(n4186), .B(DATAO_REG_5__SCAN_IN), .S(n4189), .Z(U3555) );
  MUX2_X1 U4679 ( .A(n4187), .B(DATAO_REG_4__SCAN_IN), .S(n4189), .Z(U3554) );
  MUX2_X1 U4680 ( .A(DATAO_REG_3__SCAN_IN), .B(n2433), .S(U4043), .Z(U3553) );
  MUX2_X1 U4681 ( .A(n4188), .B(DATAO_REG_2__SCAN_IN), .S(n4189), .Z(U3552) );
  MUX2_X1 U4682 ( .A(n3194), .B(DATAO_REG_1__SCAN_IN), .S(n4189), .Z(U3551) );
  MUX2_X1 U4683 ( .A(n4190), .B(DATAO_REG_0__SCAN_IN), .S(n4189), .Z(U3550) );
  OAI211_X1 U4684 ( .C1(n4193), .C2(n4192), .A(n4729), .B(n4191), .ZN(n4202)
         );
  MUX2_X1 U4685 ( .A(REG1_REG_1__SCAN_IN), .B(n4790), .S(n4194), .Z(n4196) );
  NAND2_X1 U4686 ( .A1(n4196), .A2(n4195), .ZN(n4197) );
  NAND3_X1 U4687 ( .A1(n4769), .A2(n4198), .A3(n4197), .ZN(n4201) );
  NAND2_X1 U4688 ( .A1(n4682), .A2(n2524), .ZN(n4200) );
  AOI22_X1 U4689 ( .A1(n4764), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4199) );
  NAND4_X1 U4690 ( .A1(n4202), .A2(n4201), .A3(n4200), .A4(n4199), .ZN(U3241)
         );
  AOI22_X1 U4691 ( .A1(n4764), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4213) );
  OAI211_X1 U4692 ( .C1(n4205), .C2(n4204), .A(n4729), .B(n4203), .ZN(n4210)
         );
  XNOR2_X1 U4693 ( .A(n4207), .B(n4206), .ZN(n4208) );
  NAND2_X1 U4694 ( .A1(n4769), .A2(n4208), .ZN(n4209) );
  AND2_X1 U4695 ( .A1(n4210), .A2(n4209), .ZN(n4212) );
  NAND2_X1 U4696 ( .A1(n4682), .A2(n2527), .ZN(n4211) );
  NAND4_X1 U4697 ( .A1(n4214), .A2(n4213), .A3(n4212), .A4(n4211), .ZN(U3242)
         );
  AND2_X1 U4698 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4899) );
  NOR2_X1 U4699 ( .A1(n4216), .A2(n4215), .ZN(n4221) );
  NAND2_X1 U4700 ( .A1(n4223), .A2(REG2_REG_15__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U4701 ( .A1(n4232), .A2(n4217), .ZN(n4218) );
  NAND2_X1 U4702 ( .A1(n4242), .A2(n4218), .ZN(n4220) );
  INV_X1 U4703 ( .A(n4243), .ZN(n4219) );
  AOI211_X1 U4704 ( .C1(n4221), .C2(n4220), .A(n4219), .B(n4771), .ZN(n4222)
         );
  AOI211_X1 U4705 ( .C1(n4764), .C2(ADDR_REG_15__SCAN_IN), .A(n4899), .B(n4222), .ZN(n4230) );
  XNOR2_X1 U4706 ( .A(n4223), .B(REG1_REG_15__SCAN_IN), .ZN(n4233) );
  INV_X1 U4707 ( .A(n4224), .ZN(n4654) );
  NAND2_X1 U4708 ( .A1(n4654), .A2(n4225), .ZN(n4227) );
  XNOR2_X1 U4709 ( .A(n4233), .B(n4231), .ZN(n4228) );
  NAND2_X1 U4710 ( .A1(n4769), .A2(n4228), .ZN(n4229) );
  OAI211_X1 U4711 ( .C1(n4767), .C2(n4232), .A(n4230), .B(n4229), .ZN(U3255)
         );
  NOR2_X1 U4712 ( .A1(n4234), .A2(n4235), .ZN(n4236) );
  XNOR2_X1 U4713 ( .A(n4235), .B(n4234), .ZN(n4753) );
  NOR2_X1 U4714 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4753), .ZN(n4754) );
  INV_X1 U4715 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4238) );
  INV_X1 U4716 ( .A(n4241), .ZN(n4653) );
  NOR2_X1 U4717 ( .A1(n4653), .A2(REG1_REG_17__SCAN_IN), .ZN(n4264) );
  INV_X1 U4718 ( .A(n4264), .ZN(n4237) );
  OAI21_X1 U4719 ( .B1(n4241), .B2(n4238), .A(n4237), .ZN(n4239) );
  NOR2_X1 U4720 ( .A1(n4240), .A2(n4239), .ZN(n4263) );
  AOI21_X1 U4721 ( .B1(n4240), .B2(n4239), .A(n4263), .ZN(n4252) );
  INV_X1 U4722 ( .A(n4769), .ZN(n4743) );
  XNOR2_X1 U4723 ( .A(n4241), .B(REG2_REG_17__SCAN_IN), .ZN(n4247) );
  AND2_X2 U4724 ( .A1(n4243), .A2(n4242), .ZN(n4244) );
  NAND2_X1 U4725 ( .A1(n4244), .A2(n4914), .ZN(n4245) );
  XNOR2_X2 U4726 ( .A(n4244), .B(n4234), .ZN(n4750) );
  INV_X1 U4727 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4748) );
  NAND2_X2 U4728 ( .A1(n4750), .A2(n4748), .ZN(n4749) );
  NAND2_X1 U4729 ( .A1(n4245), .A2(n4749), .ZN(n4246) );
  AOI221_X1 U4730 ( .B1(n4247), .B2(n4253), .C1(n4246), .C2(n4253), .A(n4771), 
        .ZN(n4248) );
  AOI211_X1 U4731 ( .C1(n4764), .C2(ADDR_REG_17__SCAN_IN), .A(n4249), .B(n4248), .ZN(n4251) );
  NAND2_X1 U4732 ( .A1(n4682), .A2(n4653), .ZN(n4250) );
  OAI211_X1 U4733 ( .C1(n4252), .C2(n4743), .A(n4251), .B(n4250), .ZN(U3257)
         );
  INV_X1 U4734 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4255) );
  INV_X1 U4735 ( .A(n4268), .ZN(n4759) );
  NOR2_X1 U4736 ( .A1(n4759), .A2(n4255), .ZN(n4254) );
  AOI21_X1 U4737 ( .B1(n4255), .B2(n4759), .A(n4254), .ZN(n4256) );
  NAND2_X1 U4738 ( .A1(n4764), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4260) );
  INV_X1 U4739 ( .A(n4258), .ZN(n4259) );
  NAND2_X1 U4740 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  XNOR2_X1 U4741 ( .A(n4268), .B(REG1_REG_18__SCAN_IN), .ZN(n4761) );
  XOR2_X1 U4742 ( .A(n4760), .B(n4761), .Z(n4265) );
  NAND2_X1 U4743 ( .A1(n4769), .A2(n4265), .ZN(n4266) );
  OAI211_X1 U4744 ( .C1(n4767), .C2(n4268), .A(n4267), .B(n4266), .ZN(U3258)
         );
  XNOR2_X1 U4745 ( .A(n4270), .B(n4269), .ZN(n4595) );
  AOI21_X1 U4746 ( .B1(n4272), .B2(n4443), .A(n4271), .ZN(n4592) );
  NOR2_X1 U4747 ( .A1(n4592), .A2(n4462), .ZN(n4273) );
  AOI21_X1 U4748 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4462), .A(n4273), .ZN(n4274) );
  OAI21_X1 U4749 ( .B1(n4595), .B2(n4883), .A(n4274), .ZN(U3260) );
  OAI22_X1 U4750 ( .A1(n4276), .A2(n4883), .B1(n4275), .B2(n4879), .ZN(n4277)
         );
  AOI22_X1 U4751 ( .A1(n4430), .A2(n4299), .B1(n4462), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n4279) );
  XNOR2_X1 U4752 ( .A(n4282), .B(n4289), .ZN(n4516) );
  AOI22_X1 U4753 ( .A1(n4462), .A2(REG2_REG_28__SCAN_IN), .B1(n4283), .B2(
        n4866), .ZN(n4295) );
  INV_X1 U4754 ( .A(n4306), .ZN(n4286) );
  INV_X1 U4755 ( .A(n4284), .ZN(n4285) );
  OAI211_X1 U4756 ( .C1(n4286), .C2(n4288), .A(n4285), .B(n3093), .ZN(n4514)
         );
  NAND2_X1 U4757 ( .A1(n4324), .A2(n4406), .ZN(n4287) );
  OAI21_X1 U4758 ( .B1(n4833), .B2(n4288), .A(n4287), .ZN(n4291) );
  OAI21_X1 U4759 ( .B1(n4829), .B2(n4514), .A(n4515), .ZN(n4293) );
  NAND2_X1 U4760 ( .A1(n4293), .A2(n4889), .ZN(n4294) );
  OAI211_X1 U4761 ( .C1(n4516), .C2(n4502), .A(n4295), .B(n4294), .ZN(U3262)
         );
  OAI21_X1 U4762 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n4300) );
  AOI22_X1 U4763 ( .A1(n4300), .A2(n4449), .B1(n4838), .B2(n4299), .ZN(n4301)
         );
  INV_X1 U4764 ( .A(n4301), .ZN(n4520) );
  AOI21_X1 U4765 ( .B1(n4302), .B2(n4866), .A(n4520), .ZN(n4313) );
  XNOR2_X1 U4766 ( .A(n4304), .B(n4303), .ZN(n4521) );
  NAND2_X1 U4767 ( .A1(n4521), .A2(n4305), .ZN(n4312) );
  INV_X1 U4768 ( .A(n4328), .ZN(n4307) );
  OAI21_X1 U4769 ( .B1(n4307), .B2(n4517), .A(n4306), .ZN(n4606) );
  INV_X1 U4770 ( .A(n4606), .ZN(n4310) );
  AOI22_X1 U4771 ( .A1(n4430), .A2(n4347), .B1(n4462), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4308) );
  OAI21_X1 U4772 ( .B1(n4517), .B2(n4433), .A(n4308), .ZN(n4309) );
  AOI21_X1 U4773 ( .B1(n4310), .B2(n4870), .A(n4309), .ZN(n4311) );
  OAI211_X1 U4774 ( .C1(n4462), .C2(n4313), .A(n4312), .B(n4311), .ZN(U3263)
         );
  OR2_X1 U4775 ( .A1(n4358), .A2(n4314), .ZN(n4316) );
  INV_X1 U4776 ( .A(n4528), .ZN(n4336) );
  NAND2_X1 U4777 ( .A1(n4320), .A2(n4319), .ZN(n4322) );
  XNOR2_X1 U4778 ( .A(n4322), .B(n4321), .ZN(n4323) );
  NAND2_X1 U4779 ( .A1(n4323), .A2(n4449), .ZN(n4326) );
  NAND2_X1 U4780 ( .A1(n4324), .A2(n4838), .ZN(n4325) );
  NAND2_X1 U4781 ( .A1(n4326), .A2(n4325), .ZN(n4527) );
  INV_X1 U4782 ( .A(n4327), .ZN(n4329) );
  OAI21_X1 U4783 ( .B1(n4329), .B2(n4524), .A(n4328), .ZN(n4610) );
  NOR2_X1 U4784 ( .A1(n4610), .A2(n4883), .ZN(n4334) );
  AOI22_X1 U4785 ( .A1(n4462), .A2(REG2_REG_26__SCAN_IN), .B1(n4330), .B2(
        n4866), .ZN(n4332) );
  NAND2_X1 U4786 ( .A1(n4430), .A2(n4364), .ZN(n4331) );
  OAI211_X1 U4787 ( .C1(n4433), .C2(n4524), .A(n4332), .B(n4331), .ZN(n4333)
         );
  AOI211_X1 U4788 ( .C1(n4527), .C2(n4826), .A(n4334), .B(n4333), .ZN(n4335)
         );
  OAI21_X1 U4789 ( .B1(n4336), .B2(n4502), .A(n4335), .ZN(U3264) );
  OR2_X1 U4790 ( .A1(n4358), .A2(n4337), .ZN(n4339) );
  NAND2_X1 U4791 ( .A1(n4339), .A2(n4338), .ZN(n4340) );
  XNOR2_X1 U4792 ( .A(n4340), .B(n4344), .ZN(n4532) );
  INV_X1 U4793 ( .A(n4532), .ZN(n4356) );
  NAND2_X1 U4794 ( .A1(n4342), .A2(n4341), .ZN(n4343) );
  XOR2_X1 U4795 ( .A(n4344), .B(n4343), .Z(n4349) );
  OAI22_X1 U4796 ( .A1(n4345), .A2(n4834), .B1(n4350), .B2(n4833), .ZN(n4346)
         );
  AOI21_X1 U4797 ( .B1(n4838), .B2(n4347), .A(n4346), .ZN(n4348) );
  OAI21_X1 U4798 ( .B1(n4349), .B2(n4840), .A(n4348), .ZN(n4531) );
  OR2_X1 U4799 ( .A1(n4367), .A2(n4350), .ZN(n4351) );
  NAND2_X1 U4800 ( .A1(n4327), .A2(n4351), .ZN(n4614) );
  AOI22_X1 U4801 ( .A1(n4462), .A2(REG2_REG_25__SCAN_IN), .B1(n4352), .B2(
        n4866), .ZN(n4353) );
  OAI21_X1 U4802 ( .B1(n4614), .B2(n4883), .A(n4353), .ZN(n4354) );
  AOI21_X1 U4803 ( .B1(n4531), .B2(n4826), .A(n4354), .ZN(n4355) );
  OAI21_X1 U4804 ( .B1(n4356), .B2(n4502), .A(n4355), .ZN(U3265) );
  OR2_X1 U4805 ( .A1(n4358), .A2(n4357), .ZN(n4359) );
  XOR2_X1 U4806 ( .A(n4360), .B(n4359), .Z(n4536) );
  INV_X1 U4807 ( .A(n4536), .ZN(n4375) );
  XNOR2_X1 U4808 ( .A(n4361), .B(n4360), .ZN(n4366) );
  OAI22_X1 U4809 ( .A1(n4362), .A2(n4834), .B1(n4833), .B2(n4369), .ZN(n4363)
         );
  AOI21_X1 U4810 ( .B1(n4838), .B2(n4364), .A(n4363), .ZN(n4365) );
  OAI21_X1 U4811 ( .B1(n4366), .B2(n4840), .A(n4365), .ZN(n4535) );
  INV_X1 U4812 ( .A(n4367), .ZN(n4368) );
  OAI21_X1 U4813 ( .B1(n2339), .B2(n4369), .A(n4368), .ZN(n4618) );
  NOR2_X1 U4814 ( .A1(n4618), .A2(n4883), .ZN(n4373) );
  INV_X1 U4815 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4371) );
  OAI22_X1 U4816 ( .A1(n4826), .A2(n4371), .B1(n4370), .B2(n4879), .ZN(n4372)
         );
  AOI211_X1 U4817 ( .C1(n4535), .C2(n4826), .A(n4373), .B(n4372), .ZN(n4374)
         );
  OAI21_X1 U4818 ( .B1(n4375), .B2(n4502), .A(n4374), .ZN(U3266) );
  AOI21_X1 U4819 ( .B1(n4420), .B2(n4377), .A(n4376), .ZN(n4378) );
  INV_X1 U4820 ( .A(n4378), .ZN(n4402) );
  NAND2_X1 U4821 ( .A1(n4402), .A2(n4403), .ZN(n4401) );
  NAND2_X1 U4822 ( .A1(n4401), .A2(n4379), .ZN(n4381) );
  XNOR2_X1 U4823 ( .A(n4381), .B(n4380), .ZN(n4540) );
  INV_X1 U4824 ( .A(n4540), .ZN(n4400) );
  INV_X1 U4825 ( .A(n4382), .ZN(n4383) );
  AOI21_X1 U4826 ( .B1(n4423), .B2(n4384), .A(n4383), .ZN(n4404) );
  OAI21_X1 U4827 ( .B1(n4404), .B2(n4403), .A(n4385), .ZN(n4387) );
  XNOR2_X1 U4828 ( .A(n4387), .B(n4386), .ZN(n4392) );
  AOI22_X1 U4829 ( .A1(n4425), .A2(n4406), .B1(n4443), .B2(n4388), .ZN(n4391)
         );
  NAND2_X1 U4830 ( .A1(n4389), .A2(n4838), .ZN(n4390) );
  OAI211_X1 U4831 ( .C1(n4392), .C2(n4840), .A(n4391), .B(n4390), .ZN(n4539)
         );
  OAI21_X1 U4832 ( .B1(n2336), .B2(n4395), .A(n4394), .ZN(n4622) );
  AOI22_X1 U4833 ( .A1(n4462), .A2(REG2_REG_23__SCAN_IN), .B1(n4396), .B2(
        n4866), .ZN(n4397) );
  OAI21_X1 U4834 ( .B1(n4622), .B2(n4883), .A(n4397), .ZN(n4398) );
  AOI21_X1 U4835 ( .B1(n4539), .B2(n4826), .A(n4398), .ZN(n4399) );
  OAI21_X1 U4836 ( .B1(n4400), .B2(n4502), .A(n4399), .ZN(U3267) );
  OAI21_X1 U4837 ( .B1(n4402), .B2(n4403), .A(n4401), .ZN(n4546) );
  XNOR2_X1 U4838 ( .A(n4404), .B(n4403), .ZN(n4410) );
  NAND2_X1 U4839 ( .A1(n4405), .A2(n4838), .ZN(n4408) );
  NAND2_X1 U4840 ( .A1(n4445), .A2(n4406), .ZN(n4407) );
  OAI211_X1 U4841 ( .C1(n4833), .C2(n4415), .A(n4408), .B(n4407), .ZN(n4409)
         );
  AOI21_X1 U4842 ( .B1(n4410), .B2(n4449), .A(n4409), .ZN(n4545) );
  INV_X1 U4843 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4412) );
  OAI22_X1 U4844 ( .A1(n4826), .A2(n4412), .B1(n4411), .B2(n4879), .ZN(n4413)
         );
  INV_X1 U4845 ( .A(n4413), .ZN(n4417) );
  OR2_X1 U4846 ( .A1(n4414), .A2(n4415), .ZN(n4543) );
  NAND3_X1 U4847 ( .A1(n4543), .A2(n4393), .A3(n4870), .ZN(n4416) );
  OAI211_X1 U4848 ( .C1(n4545), .C2(n4462), .A(n4417), .B(n4416), .ZN(n4418)
         );
  INV_X1 U4849 ( .A(n4418), .ZN(n4419) );
  OAI21_X1 U4850 ( .B1(n4546), .B2(n4502), .A(n4419), .ZN(U3268) );
  XOR2_X1 U4851 ( .A(n4421), .B(n4420), .Z(n4552) );
  INV_X1 U4852 ( .A(n4552), .ZN(n4437) );
  INV_X1 U4853 ( .A(n4421), .ZN(n4422) );
  XNOR2_X1 U4854 ( .A(n4423), .B(n4422), .ZN(n4424) );
  NAND2_X1 U4855 ( .A1(n4424), .A2(n4449), .ZN(n4427) );
  NAND2_X1 U4856 ( .A1(n4425), .A2(n4838), .ZN(n4426) );
  NAND2_X1 U4857 ( .A1(n4427), .A2(n4426), .ZN(n4551) );
  INV_X1 U4858 ( .A(n4414), .ZN(n4428) );
  OAI21_X1 U4859 ( .B1(n4454), .B2(n4548), .A(n4428), .ZN(n4627) );
  NOR2_X1 U4860 ( .A1(n4627), .A2(n4883), .ZN(n4435) );
  AOI22_X1 U4861 ( .A1(n4462), .A2(REG2_REG_21__SCAN_IN), .B1(n4429), .B2(
        n4866), .ZN(n4432) );
  NAND2_X1 U4862 ( .A1(n4430), .A2(n4547), .ZN(n4431) );
  OAI211_X1 U4863 ( .C1(n4433), .C2(n4548), .A(n4432), .B(n4431), .ZN(n4434)
         );
  AOI211_X1 U4864 ( .C1(n4551), .C2(n4826), .A(n4435), .B(n4434), .ZN(n4436)
         );
  OAI21_X1 U4865 ( .B1(n4437), .B2(n4502), .A(n4436), .ZN(U3269) );
  XNOR2_X1 U4866 ( .A(n4438), .B(n4442), .ZN(n4453) );
  NAND2_X1 U4867 ( .A1(n4440), .A2(n4439), .ZN(n4441) );
  XOR2_X1 U4868 ( .A(n4442), .B(n4441), .Z(n4450) );
  AOI22_X1 U4869 ( .A1(n4445), .A2(n4838), .B1(n4444), .B2(n4443), .ZN(n4446)
         );
  OAI21_X1 U4870 ( .B1(n4447), .B2(n4834), .A(n4446), .ZN(n4448) );
  AOI21_X1 U4871 ( .B1(n4450), .B2(n4449), .A(n4448), .ZN(n4451) );
  OAI21_X1 U4872 ( .B1(n4453), .B2(n4452), .A(n4451), .ZN(n4555) );
  INV_X1 U4873 ( .A(n4555), .ZN(n4463) );
  INV_X1 U4874 ( .A(n4453), .ZN(n4556) );
  INV_X1 U4875 ( .A(n4479), .ZN(n4457) );
  INV_X1 U4876 ( .A(n4454), .ZN(n4455) );
  OAI21_X1 U4877 ( .B1(n4457), .B2(n4456), .A(n4455), .ZN(n4631) );
  AOI22_X1 U4878 ( .A1(n4462), .A2(REG2_REG_20__SCAN_IN), .B1(n4458), .B2(
        n4866), .ZN(n4459) );
  OAI21_X1 U4879 ( .B1(n4631), .B2(n4883), .A(n4459), .ZN(n4460) );
  AOI21_X1 U4880 ( .B1(n4556), .B2(n4871), .A(n4460), .ZN(n4461) );
  OAI21_X1 U4881 ( .B1(n4463), .B2(n4462), .A(n4461), .ZN(U3270) );
  XNOR2_X1 U4882 ( .A(n4464), .B(n4473), .ZN(n4560) );
  INV_X1 U4883 ( .A(n4560), .ZN(n4488) );
  INV_X1 U4884 ( .A(n4465), .ZN(n4467) );
  OAI21_X1 U4885 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n4492) );
  INV_X1 U4886 ( .A(n4469), .ZN(n4471) );
  OAI21_X1 U4887 ( .B1(n4492), .B2(n4471), .A(n4470), .ZN(n4472) );
  XOR2_X1 U4888 ( .A(n4473), .B(n4472), .Z(n4477) );
  OAI22_X1 U4889 ( .A1(n4474), .A2(n4834), .B1(n4480), .B2(n4833), .ZN(n4475)
         );
  AOI21_X1 U4890 ( .B1(n4838), .B2(n4547), .A(n4475), .ZN(n4476) );
  OAI21_X1 U4891 ( .B1(n4477), .B2(n4840), .A(n4476), .ZN(n4559) );
  INV_X1 U4892 ( .A(n4478), .ZN(n4481) );
  OAI21_X1 U4893 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n4635) );
  NOR2_X1 U4894 ( .A1(n4635), .A2(n4883), .ZN(n4486) );
  INV_X1 U4895 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4484) );
  INV_X1 U4896 ( .A(n4482), .ZN(n4483) );
  OAI22_X1 U4897 ( .A1(n4826), .A2(n4484), .B1(n4483), .B2(n4879), .ZN(n4485)
         );
  AOI211_X1 U4898 ( .C1(n4559), .C2(n4826), .A(n4486), .B(n4485), .ZN(n4487)
         );
  OAI21_X1 U4899 ( .B1(n4488), .B2(n4502), .A(n4487), .ZN(U3271) );
  OAI211_X1 U4900 ( .C1(n4489), .C2(n4490), .A(n4478), .B(n3093), .ZN(n4563)
         );
  OAI22_X1 U4901 ( .A1(n4491), .A2(n4834), .B1(n4490), .B2(n4833), .ZN(n4495)
         );
  XNOR2_X1 U4902 ( .A(n4492), .B(n4499), .ZN(n4493) );
  NOR2_X1 U4903 ( .A1(n4493), .A2(n4840), .ZN(n4494) );
  AOI211_X1 U4904 ( .C1(n4838), .C2(n4496), .A(n4495), .B(n4494), .ZN(n4564)
         );
  OAI21_X1 U4905 ( .B1(n4829), .B2(n4563), .A(n4564), .ZN(n4505) );
  OAI22_X1 U4906 ( .A1(n4826), .A2(n4255), .B1(n4497), .B2(n4879), .ZN(n4504)
         );
  OAI21_X1 U4907 ( .B1(n4500), .B2(n4499), .A(n4498), .ZN(n4501) );
  INV_X1 U4908 ( .A(n4501), .ZN(n4565) );
  NOR2_X1 U4909 ( .A1(n4565), .A2(n4502), .ZN(n4503) );
  AOI211_X1 U4910 ( .C1(n4826), .C2(n4505), .A(n4504), .B(n4503), .ZN(n4506)
         );
  INV_X1 U4911 ( .A(n4506), .ZN(U3272) );
  NOR2_X1 U4912 ( .A1(n4592), .A2(n3091), .ZN(n4507) );
  AOI21_X1 U4913 ( .B1(REG1_REG_31__SCAN_IN), .B2(n3091), .A(n4507), .ZN(n4508) );
  OAI21_X1 U4914 ( .B1(n4595), .B2(n4591), .A(n4508), .ZN(U3549) );
  INV_X1 U4915 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4513) );
  INV_X1 U4916 ( .A(n4509), .ZN(n4597) );
  NAND2_X1 U4917 ( .A1(n4597), .A2(n4510), .ZN(n4512) );
  NAND2_X1 U4918 ( .A1(n4598), .A2(n4852), .ZN(n4511) );
  OAI211_X1 U4919 ( .C1(n4852), .C2(n4513), .A(n4512), .B(n4511), .ZN(U3548)
         );
  INV_X1 U4920 ( .A(n4587), .ZN(n4845) );
  MUX2_X1 U4921 ( .A(REG1_REG_28__SCAN_IN), .B(n4602), .S(n4852), .Z(U3546) );
  INV_X1 U4922 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4522) );
  OAI22_X1 U4923 ( .A1(n4518), .A2(n4834), .B1(n4517), .B2(n4833), .ZN(n4519)
         );
  AOI211_X1 U4924 ( .C1(n4521), .C2(n4587), .A(n4520), .B(n4519), .ZN(n4603)
         );
  MUX2_X1 U4925 ( .A(n4522), .B(n4603), .S(n4852), .Z(n4523) );
  OAI21_X1 U4926 ( .B1(n4591), .B2(n4606), .A(n4523), .ZN(U3545) );
  INV_X1 U4927 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4529) );
  OAI22_X1 U4928 ( .A1(n4525), .A2(n4834), .B1(n4524), .B2(n4833), .ZN(n4526)
         );
  AOI211_X1 U4929 ( .C1(n4528), .C2(n4587), .A(n4527), .B(n4526), .ZN(n4607)
         );
  MUX2_X1 U4930 ( .A(n4529), .B(n4607), .S(n4852), .Z(n4530) );
  OAI21_X1 U4931 ( .B1(n4591), .B2(n4610), .A(n4530), .ZN(U3544) );
  INV_X1 U4932 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4533) );
  AOI21_X1 U4933 ( .B1(n4532), .B2(n4587), .A(n4531), .ZN(n4611) );
  MUX2_X1 U4934 ( .A(n4533), .B(n4611), .S(n4852), .Z(n4534) );
  OAI21_X1 U4935 ( .B1(n4591), .B2(n4614), .A(n4534), .ZN(U3543) );
  INV_X1 U4936 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4537) );
  AOI21_X1 U4937 ( .B1(n4536), .B2(n4587), .A(n4535), .ZN(n4615) );
  MUX2_X1 U4938 ( .A(n4537), .B(n4615), .S(n4852), .Z(n4538) );
  OAI21_X1 U4939 ( .B1(n4591), .B2(n4618), .A(n4538), .ZN(U3542) );
  INV_X1 U4940 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4541) );
  AOI21_X1 U4941 ( .B1(n4540), .B2(n4587), .A(n4539), .ZN(n4619) );
  MUX2_X1 U4942 ( .A(n4541), .B(n4619), .S(n4852), .Z(n4542) );
  OAI21_X1 U4943 ( .B1(n4591), .B2(n4622), .A(n4542), .ZN(U3541) );
  NAND3_X1 U4944 ( .A1(n4543), .A2(n3093), .A3(n4393), .ZN(n4544) );
  OAI211_X1 U4945 ( .C1(n4546), .C2(n4845), .A(n4545), .B(n4544), .ZN(n4623)
         );
  MUX2_X1 U4946 ( .A(REG1_REG_22__SCAN_IN), .B(n4623), .S(n4852), .Z(U3540) );
  INV_X1 U4947 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4553) );
  INV_X1 U4948 ( .A(n4547), .ZN(n4549) );
  OAI22_X1 U4949 ( .A1(n4549), .A2(n4834), .B1(n4833), .B2(n4548), .ZN(n4550)
         );
  AOI211_X1 U4950 ( .C1(n4552), .C2(n4587), .A(n4551), .B(n4550), .ZN(n4624)
         );
  MUX2_X1 U4951 ( .A(n4553), .B(n4624), .S(n4852), .Z(n4554) );
  OAI21_X1 U4952 ( .B1(n4591), .B2(n4627), .A(n4554), .ZN(U3539) );
  INV_X1 U4953 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4557) );
  AOI21_X1 U4954 ( .B1(n4802), .B2(n4556), .A(n4555), .ZN(n4628) );
  MUX2_X1 U4955 ( .A(n4557), .B(n4628), .S(n4852), .Z(n4558) );
  OAI21_X1 U4956 ( .B1(n4591), .B2(n4631), .A(n4558), .ZN(U3538) );
  INV_X1 U4957 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4561) );
  AOI21_X1 U4958 ( .B1(n4560), .B2(n4587), .A(n4559), .ZN(n4632) );
  MUX2_X1 U4959 ( .A(n4561), .B(n4632), .S(n4852), .Z(n4562) );
  OAI21_X1 U4960 ( .B1(n4591), .B2(n4635), .A(n4562), .ZN(U3537) );
  OAI211_X1 U4961 ( .C1(n4565), .C2(n4845), .A(n4564), .B(n4563), .ZN(n4636)
         );
  MUX2_X1 U4962 ( .A(REG1_REG_18__SCAN_IN), .B(n4636), .S(n4852), .Z(U3536) );
  OAI22_X1 U4963 ( .A1(n4898), .A2(n4834), .B1(n4566), .B2(n4833), .ZN(n4567)
         );
  AOI211_X1 U4964 ( .C1(n4569), .C2(n4587), .A(n4568), .B(n4567), .ZN(n4637)
         );
  MUX2_X1 U4965 ( .A(n4238), .B(n4637), .S(n4852), .Z(n4570) );
  OAI21_X1 U4966 ( .B1(n4591), .B2(n4640), .A(n4570), .ZN(U3535) );
  OAI22_X1 U4967 ( .A1(n4572), .A2(n4834), .B1(n4571), .B2(n4833), .ZN(n4574)
         );
  AOI211_X1 U4968 ( .C1(n3093), .C2(n4575), .A(n4574), .B(n4573), .ZN(n4576)
         );
  OAI21_X1 U4969 ( .B1(n4577), .B2(n4845), .A(n4576), .ZN(n4641) );
  MUX2_X1 U4970 ( .A(REG1_REG_16__SCAN_IN), .B(n4641), .S(n4852), .Z(U3534) );
  OAI22_X1 U4971 ( .A1(n4895), .A2(n4834), .B1(n4833), .B2(n4901), .ZN(n4578)
         );
  AOI21_X1 U4972 ( .B1(n4579), .B2(n3093), .A(n4578), .ZN(n4580) );
  OAI211_X1 U4973 ( .C1(n4582), .C2(n4845), .A(n4581), .B(n4580), .ZN(n4642)
         );
  MUX2_X1 U4974 ( .A(REG1_REG_15__SCAN_IN), .B(n4642), .S(n4852), .Z(U3533) );
  INV_X1 U4975 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4589) );
  OAI22_X1 U4976 ( .A1(n4584), .A2(n4834), .B1(n4833), .B2(n4583), .ZN(n4585)
         );
  AOI211_X1 U4977 ( .C1(n4588), .C2(n4587), .A(n4586), .B(n4585), .ZN(n4643)
         );
  MUX2_X1 U4978 ( .A(n4589), .B(n4643), .S(n4852), .Z(n4590) );
  OAI21_X1 U4979 ( .B1(n4591), .B2(n4647), .A(n4590), .ZN(U3532) );
  NOR2_X1 U4980 ( .A1(n4592), .A2(n3099), .ZN(n4593) );
  AOI21_X1 U4981 ( .B1(REG0_REG_31__SCAN_IN), .B2(n3099), .A(n4593), .ZN(n4594) );
  OAI21_X1 U4982 ( .B1(n4595), .B2(n4646), .A(n4594), .ZN(U3517) );
  INV_X1 U4983 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U4984 ( .A1(n4597), .A2(n4596), .ZN(n4600) );
  NAND2_X1 U4985 ( .A1(n4598), .A2(n4855), .ZN(n4599) );
  OAI211_X1 U4986 ( .C1(n4855), .C2(n4601), .A(n4600), .B(n4599), .ZN(U3516)
         );
  MUX2_X1 U4987 ( .A(REG0_REG_28__SCAN_IN), .B(n4602), .S(n4855), .Z(U3514) );
  INV_X1 U4988 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4604) );
  MUX2_X1 U4989 ( .A(n4604), .B(n4603), .S(n4855), .Z(n4605) );
  OAI21_X1 U4990 ( .B1(n4606), .B2(n4646), .A(n4605), .ZN(U3513) );
  INV_X1 U4991 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4608) );
  MUX2_X1 U4992 ( .A(n4608), .B(n4607), .S(n4855), .Z(n4609) );
  OAI21_X1 U4993 ( .B1(n4610), .B2(n4646), .A(n4609), .ZN(U3512) );
  INV_X1 U4994 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4612) );
  MUX2_X1 U4995 ( .A(n4612), .B(n4611), .S(n4855), .Z(n4613) );
  OAI21_X1 U4996 ( .B1(n4614), .B2(n4646), .A(n4613), .ZN(U3511) );
  INV_X1 U4997 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4616) );
  MUX2_X1 U4998 ( .A(n4616), .B(n4615), .S(n4855), .Z(n4617) );
  OAI21_X1 U4999 ( .B1(n4618), .B2(n4646), .A(n4617), .ZN(U3510) );
  INV_X1 U5000 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4620) );
  MUX2_X1 U5001 ( .A(n4620), .B(n4619), .S(n4855), .Z(n4621) );
  OAI21_X1 U5002 ( .B1(n4622), .B2(n4646), .A(n4621), .ZN(U3509) );
  MUX2_X1 U5003 ( .A(REG0_REG_22__SCAN_IN), .B(n4623), .S(n4855), .Z(U3508) );
  INV_X1 U5004 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4625) );
  MUX2_X1 U5005 ( .A(n4625), .B(n4624), .S(n4855), .Z(n4626) );
  OAI21_X1 U5006 ( .B1(n4627), .B2(n4646), .A(n4626), .ZN(U3507) );
  INV_X1 U5007 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4629) );
  MUX2_X1 U5008 ( .A(n4629), .B(n4628), .S(n4855), .Z(n4630) );
  OAI21_X1 U5009 ( .B1(n4631), .B2(n4646), .A(n4630), .ZN(U3506) );
  INV_X1 U5010 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4633) );
  MUX2_X1 U5011 ( .A(n4633), .B(n4632), .S(n4855), .Z(n4634) );
  OAI21_X1 U5012 ( .B1(n4635), .B2(n4646), .A(n4634), .ZN(U3505) );
  MUX2_X1 U5013 ( .A(REG0_REG_18__SCAN_IN), .B(n4636), .S(n4855), .Z(U3503) );
  INV_X1 U5014 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4638) );
  MUX2_X1 U5015 ( .A(n4638), .B(n4637), .S(n4855), .Z(n4639) );
  OAI21_X1 U5016 ( .B1(n4640), .B2(n4646), .A(n4639), .ZN(U3501) );
  MUX2_X1 U5017 ( .A(REG0_REG_16__SCAN_IN), .B(n4641), .S(n4855), .Z(U3499) );
  MUX2_X1 U5018 ( .A(REG0_REG_15__SCAN_IN), .B(n4642), .S(n4855), .Z(U3497) );
  INV_X1 U5019 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4644) );
  MUX2_X1 U5020 ( .A(n4644), .B(n4643), .S(n4855), .Z(n4645) );
  OAI21_X1 U5021 ( .B1(n4647), .B2(n4646), .A(n4645), .ZN(U3495) );
  MUX2_X1 U5022 ( .A(n4648), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5023 ( .A(n4649), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5024 ( .A(n4650), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5025 ( .A(DATAI_22_), .B(n4651), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5026 ( .A(DATAI_20_), .B(n4652), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5027 ( .A(n4829), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5028 ( .A(DATAI_18_), .B(n4759), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5029 ( .A(DATAI_17_), .B(n4653), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U5030 ( .A(DATAI_14_), .B(n4654), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5031 ( .A(n2403), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5032 ( .A(DATAI_4_), .B(n4655), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5033 ( .A(DATAI_3_), .B(n3144), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5034 ( .A(n2527), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5035 ( .A(n2524), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5036 ( .A(DATAI_23_), .ZN(n4657) );
  OAI21_X1 U5037 ( .B1(STATE_REG_SCAN_IN), .B2(n4657), .A(n4656), .ZN(U3329)
         );
  AND2_X1 U5038 ( .A1(D_REG_2__SCAN_IN), .A2(n4658), .ZN(U3320) );
  AND2_X1 U5039 ( .A1(D_REG_3__SCAN_IN), .A2(n4658), .ZN(U3319) );
  AND2_X1 U5040 ( .A1(D_REG_4__SCAN_IN), .A2(n4658), .ZN(U3318) );
  AND2_X1 U5041 ( .A1(D_REG_5__SCAN_IN), .A2(n4658), .ZN(U3317) );
  AND2_X1 U5042 ( .A1(D_REG_6__SCAN_IN), .A2(n4658), .ZN(U3316) );
  AND2_X1 U5043 ( .A1(D_REG_7__SCAN_IN), .A2(n4658), .ZN(U3315) );
  AND2_X1 U5044 ( .A1(D_REG_8__SCAN_IN), .A2(n4658), .ZN(U3314) );
  AND2_X1 U5045 ( .A1(D_REG_9__SCAN_IN), .A2(n4658), .ZN(U3313) );
  AND2_X1 U5046 ( .A1(D_REG_10__SCAN_IN), .A2(n4658), .ZN(U3312) );
  AND2_X1 U5047 ( .A1(D_REG_11__SCAN_IN), .A2(n4658), .ZN(U3311) );
  AND2_X1 U5048 ( .A1(D_REG_12__SCAN_IN), .A2(n4658), .ZN(U3310) );
  AND2_X1 U5049 ( .A1(D_REG_13__SCAN_IN), .A2(n4658), .ZN(U3309) );
  AND2_X1 U5050 ( .A1(D_REG_14__SCAN_IN), .A2(n4658), .ZN(U3308) );
  AND2_X1 U5051 ( .A1(D_REG_15__SCAN_IN), .A2(n4658), .ZN(U3307) );
  AND2_X1 U5052 ( .A1(D_REG_16__SCAN_IN), .A2(n4658), .ZN(U3306) );
  AND2_X1 U5053 ( .A1(D_REG_17__SCAN_IN), .A2(n4658), .ZN(U3305) );
  AND2_X1 U5054 ( .A1(D_REG_18__SCAN_IN), .A2(n4658), .ZN(U3304) );
  AND2_X1 U5055 ( .A1(D_REG_19__SCAN_IN), .A2(n4658), .ZN(U3303) );
  AND2_X1 U5056 ( .A1(D_REG_20__SCAN_IN), .A2(n4658), .ZN(U3302) );
  AND2_X1 U5057 ( .A1(D_REG_21__SCAN_IN), .A2(n4658), .ZN(U3301) );
  AND2_X1 U5058 ( .A1(D_REG_22__SCAN_IN), .A2(n4658), .ZN(U3300) );
  AND2_X1 U5059 ( .A1(D_REG_23__SCAN_IN), .A2(n4658), .ZN(U3299) );
  AND2_X1 U5060 ( .A1(D_REG_24__SCAN_IN), .A2(n4658), .ZN(U3298) );
  AND2_X1 U5061 ( .A1(D_REG_25__SCAN_IN), .A2(n4658), .ZN(U3297) );
  AND2_X1 U5062 ( .A1(D_REG_26__SCAN_IN), .A2(n4658), .ZN(U3296) );
  AND2_X1 U5063 ( .A1(D_REG_27__SCAN_IN), .A2(n4658), .ZN(U3295) );
  AND2_X1 U5064 ( .A1(D_REG_28__SCAN_IN), .A2(n4658), .ZN(U3294) );
  AND2_X1 U5065 ( .A1(D_REG_29__SCAN_IN), .A2(n4658), .ZN(U3293) );
  AND2_X1 U5066 ( .A1(D_REG_30__SCAN_IN), .A2(n4658), .ZN(U3292) );
  AND2_X1 U5067 ( .A1(D_REG_31__SCAN_IN), .A2(n4658), .ZN(U3291) );
  AOI211_X1 U5068 ( .C1(n4661), .C2(n4660), .A(n4659), .B(n4771), .ZN(n4663)
         );
  AOI211_X1 U5069 ( .C1(n4764), .C2(ADDR_REG_5__SCAN_IN), .A(n4663), .B(n4662), 
        .ZN(n4668) );
  OAI211_X1 U5070 ( .C1(n4666), .C2(n4665), .A(n4769), .B(n4664), .ZN(n4667)
         );
  OAI211_X1 U5071 ( .C1(n4767), .C2(n4807), .A(n4668), .B(n4667), .ZN(U3245)
         );
  AOI211_X1 U5072 ( .C1(n4671), .C2(n4670), .A(n4669), .B(n4771), .ZN(n4673)
         );
  AOI211_X1 U5073 ( .C1(n4764), .C2(ADDR_REG_6__SCAN_IN), .A(n4673), .B(n4672), 
        .ZN(n4677) );
  OAI211_X1 U5074 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4675), .A(n4769), .B(n4674), 
        .ZN(n4676) );
  OAI211_X1 U5075 ( .C1(n4767), .C2(n3275), .A(n4677), .B(n4676), .ZN(U3246)
         );
  INV_X1 U5076 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5077 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4680), .B1(n4679), .B2(n4678), .ZN(n4681) );
  XNOR2_X1 U5078 ( .A(n4817), .B(n4681), .ZN(n4685) );
  NOR2_X1 U5079 ( .A1(n4851), .A2(n4743), .ZN(n4683) );
  AOI21_X1 U5080 ( .B1(n4683), .B2(n4689), .A(n4682), .ZN(n4684) );
  OAI22_X1 U5081 ( .A1(n4771), .A2(n4685), .B1(n4817), .B2(n4684), .ZN(n4686)
         );
  AOI211_X1 U5082 ( .C1(n4764), .C2(ADDR_REG_7__SCAN_IN), .A(n4687), .B(n4686), 
        .ZN(n4692) );
  OAI211_X1 U5083 ( .C1(n4690), .C2(n4689), .A(n4769), .B(n4688), .ZN(n4691)
         );
  NAND2_X1 U5084 ( .A1(n4692), .A2(n4691), .ZN(U3247) );
  AOI211_X1 U5085 ( .C1(n4695), .C2(n4694), .A(n4693), .B(n4743), .ZN(n4697)
         );
  AOI211_X1 U5086 ( .C1(n4764), .C2(ADDR_REG_8__SCAN_IN), .A(n4697), .B(n4696), 
        .ZN(n4701) );
  OAI211_X1 U5087 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4699), .A(n4729), .B(n4698), 
        .ZN(n4700) );
  OAI211_X1 U5088 ( .C1(n4767), .C2(n4702), .A(n4701), .B(n4700), .ZN(U3248)
         );
  OAI211_X1 U5089 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4704), .A(n4769), .B(n4703), .ZN(n4708) );
  OAI211_X1 U5090 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4706), .A(n4729), .B(n4705), .ZN(n4707) );
  OAI211_X1 U5091 ( .C1(n4767), .C2(n4865), .A(n4708), .B(n4707), .ZN(n4709)
         );
  AOI211_X1 U5092 ( .C1(n4764), .C2(ADDR_REG_10__SCAN_IN), .A(n4710), .B(n4709), .ZN(n4711) );
  INV_X1 U5093 ( .A(n4711), .ZN(U3250) );
  AOI22_X1 U5094 ( .A1(n4712), .A2(REG1_REG_11__SCAN_IN), .B1(n3660), .B2(
        n4877), .ZN(n4715) );
  OAI21_X1 U5095 ( .B1(n4715), .B2(n4714), .A(n4769), .ZN(n4713) );
  AOI21_X1 U5096 ( .B1(n4715), .B2(n4714), .A(n4713), .ZN(n4717) );
  AOI211_X1 U5097 ( .C1(n4764), .C2(ADDR_REG_11__SCAN_IN), .A(n4717), .B(n4716), .ZN(n4722) );
  OAI211_X1 U5098 ( .C1(n4720), .C2(n4719), .A(n4729), .B(n4718), .ZN(n4721)
         );
  OAI211_X1 U5099 ( .C1(n4767), .C2(n4877), .A(n4722), .B(n4721), .ZN(U3251)
         );
  AOI211_X1 U5100 ( .C1(n4725), .C2(n4724), .A(n4723), .B(n4743), .ZN(n4727)
         );
  AOI211_X1 U5101 ( .C1(n4764), .C2(ADDR_REG_12__SCAN_IN), .A(n4727), .B(n4726), .ZN(n4732) );
  OAI211_X1 U5102 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4730), .A(n4729), .B(n4728), .ZN(n4731) );
  OAI211_X1 U5103 ( .C1(n4767), .C2(n4892), .A(n4732), .B(n4731), .ZN(U3252)
         );
  AOI21_X1 U5104 ( .B1(n4894), .B2(n4734), .A(n4733), .ZN(n4735) );
  XNOR2_X1 U5105 ( .A(n4736), .B(n4735), .ZN(n4747) );
  INV_X1 U5106 ( .A(n4737), .ZN(n4738) );
  NAND2_X1 U5107 ( .A1(n4739), .A2(n4738), .ZN(n4740) );
  XNOR2_X1 U5108 ( .A(n4741), .B(n4740), .ZN(n4742) );
  OAI22_X1 U5109 ( .A1(n4894), .A2(n4767), .B1(n4743), .B2(n4742), .ZN(n4744)
         );
  AOI211_X1 U5110 ( .C1(n4764), .C2(ADDR_REG_13__SCAN_IN), .A(n4745), .B(n4744), .ZN(n4746) );
  OAI21_X1 U5111 ( .B1(n4747), .B2(n4771), .A(n4746), .ZN(U3253) );
  AOI221_X1 U5112 ( .B1(n4750), .B2(n4749), .C1(n4748), .C2(n4749), .A(n4771), 
        .ZN(n4751) );
  AOI211_X1 U5113 ( .C1(n4764), .C2(ADDR_REG_16__SCAN_IN), .A(n4752), .B(n4751), .ZN(n4756) );
  OAI221_X1 U5114 ( .B1(n4754), .B2(REG1_REG_16__SCAN_IN), .C1(n4754), .C2(
        n4753), .A(n4769), .ZN(n4755) );
  OAI211_X1 U5115 ( .C1(n4767), .C2(n4914), .A(n4756), .B(n4755), .ZN(U3256)
         );
  MUX2_X1 U5116 ( .A(REG2_REG_19__SCAN_IN), .B(n4484), .S(n4766), .Z(n4757) );
  XNOR2_X1 U5117 ( .A(n4758), .B(n4757), .ZN(n4772) );
  MUX2_X1 U5118 ( .A(REG1_REG_19__SCAN_IN), .B(n4561), .S(n4766), .Z(n4762) );
  AOI21_X1 U5119 ( .B1(n4764), .B2(ADDR_REG_19__SCAN_IN), .A(n4763), .ZN(n4765) );
  OAI21_X1 U5120 ( .B1(n4767), .B2(n4766), .A(n4765), .ZN(n4768) );
  OAI21_X1 U5121 ( .B1(n4772), .B2(n4771), .A(n4770), .ZN(U3259) );
  AOI22_X1 U5122 ( .A1(STATE_REG_SCAN_IN), .A2(n4774), .B1(n4773), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5123 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4775) );
  AOI22_X1 U5124 ( .A1(n4855), .A2(n4776), .B1(n4775), .B2(n3099), .ZN(U3467)
         );
  INV_X1 U5125 ( .A(n4777), .ZN(n4779) );
  AOI21_X1 U5126 ( .B1(n4780), .B2(n4779), .A(n4778), .ZN(n4784) );
  INV_X1 U5127 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5128 ( .A1(n4781), .A2(n4871), .B1(REG3_REG_0__SCAN_IN), .B2(n4866), .ZN(n4782) );
  OAI221_X1 U5129 ( .B1(n4462), .B2(n4784), .C1(n4889), .C2(n4783), .A(n4782), 
        .ZN(U3290) );
  INV_X1 U5130 ( .A(n3093), .ZN(n4818) );
  OAI22_X1 U5131 ( .A1(n4787), .A2(n4786), .B1(n4818), .B2(n4785), .ZN(n4788)
         );
  NOR2_X1 U5132 ( .A1(n4789), .A2(n4788), .ZN(n4792) );
  AOI22_X1 U5133 ( .A1(n4852), .A2(n4792), .B1(n4790), .B2(n3091), .ZN(U3519)
         );
  INV_X1 U5134 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5135 ( .A1(n4855), .A2(n4792), .B1(n4791), .B2(n3099), .ZN(U3469)
         );
  AOI22_X1 U5136 ( .A1(n4462), .A2(REG2_REG_3__SCAN_IN), .B1(n4866), .B2(n4793), .ZN(n4797) );
  AOI22_X1 U5137 ( .A1(n4795), .A2(n4871), .B1(n4870), .B2(n4794), .ZN(n4796)
         );
  OAI211_X1 U5138 ( .C1(n4462), .C2(n4798), .A(n4797), .B(n4796), .ZN(U3287)
         );
  INV_X1 U5139 ( .A(n4799), .ZN(n4801) );
  AOI211_X1 U5140 ( .C1(n4803), .C2(n4802), .A(n4801), .B(n4800), .ZN(n4805)
         );
  AOI22_X1 U5141 ( .A1(n4852), .A2(n4805), .B1(n3272), .B2(n3091), .ZN(U3522)
         );
  INV_X1 U5142 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5143 ( .A1(n4855), .A2(n4805), .B1(n4804), .B2(n3099), .ZN(U3475)
         );
  AOI22_X1 U5144 ( .A1(STATE_REG_SCAN_IN), .A2(n4807), .B1(n4806), .B2(U3149), 
        .ZN(U3347) );
  AOI22_X1 U5145 ( .A1(STATE_REG_SCAN_IN), .A2(n3275), .B1(n4808), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5146 ( .A1(n4809), .A2(n4866), .B1(REG2_REG_6__SCAN_IN), .B2(n4462), .ZN(n4814) );
  INV_X1 U5147 ( .A(n4810), .ZN(n4811) );
  AOI22_X1 U5148 ( .A1(n4812), .A2(n4871), .B1(n4870), .B2(n4811), .ZN(n4813)
         );
  OAI211_X1 U5149 ( .C1(n4462), .C2(n4815), .A(n4814), .B(n4813), .ZN(U3284)
         );
  AOI22_X1 U5150 ( .A1(STATE_REG_SCAN_IN), .A2(n4817), .B1(n4816), .B2(U3149), 
        .ZN(U3345) );
  AOI21_X1 U5151 ( .B1(n4820), .B2(n4819), .A(n4818), .ZN(n4822) );
  AND2_X1 U5152 ( .A1(n4822), .A2(n4821), .ZN(n4848) );
  INV_X1 U5153 ( .A(n4848), .ZN(n4828) );
  NOR2_X1 U5154 ( .A1(n4823), .A2(n4830), .ZN(n4846) );
  INV_X1 U5155 ( .A(n4846), .ZN(n4825) );
  NAND3_X1 U5156 ( .A1(n4825), .A2(n4849), .A3(n4824), .ZN(n4827) );
  OAI211_X1 U5157 ( .C1(n4829), .C2(n4828), .A(n4827), .B(n4826), .ZN(n4842)
         );
  XNOR2_X1 U5158 ( .A(n4831), .B(n4830), .ZN(n4841) );
  OAI22_X1 U5159 ( .A1(n4835), .A2(n4834), .B1(n4833), .B2(n4832), .ZN(n4836)
         );
  AOI21_X1 U5160 ( .B1(n4838), .B2(n4837), .A(n4836), .ZN(n4839) );
  OAI21_X1 U5161 ( .B1(n4841), .B2(n4840), .A(n4839), .ZN(n4847) );
  OAI22_X1 U5162 ( .A1(n4842), .A2(n4847), .B1(REG2_REG_7__SCAN_IN), .B2(n4889), .ZN(n4843) );
  OAI21_X1 U5163 ( .B1(n4844), .B2(n4879), .A(n4843), .ZN(U3283) );
  NOR2_X1 U5164 ( .A1(n4846), .A2(n4845), .ZN(n4850) );
  AOI211_X1 U5165 ( .C1(n4850), .C2(n4849), .A(n4848), .B(n4847), .ZN(n4854)
         );
  AOI22_X1 U5166 ( .A1(n4852), .A2(n4854), .B1(n4851), .B2(n3091), .ZN(U3525)
         );
  INV_X1 U5167 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4853) );
  AOI22_X1 U5168 ( .A1(n4855), .A2(n4854), .B1(n4853), .B2(n3099), .ZN(U3481)
         );
  OAI22_X1 U5169 ( .A1(U3149), .A2(n4856), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4857) );
  INV_X1 U5170 ( .A(n4857), .ZN(U3344) );
  AOI22_X1 U5171 ( .A1(n4858), .A2(n4866), .B1(REG2_REG_8__SCAN_IN), .B2(n4462), .ZN(n4862) );
  AOI22_X1 U5172 ( .A1(n4860), .A2(n4871), .B1(n4870), .B2(n4859), .ZN(n4861)
         );
  OAI211_X1 U5173 ( .C1(n4462), .C2(n4863), .A(n4862), .B(n4861), .ZN(U3282)
         );
  AOI22_X1 U5174 ( .A1(STATE_REG_SCAN_IN), .A2(n4865), .B1(n4864), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5175 ( .A1(n4867), .A2(n4866), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4462), .ZN(n4874) );
  INV_X1 U5176 ( .A(n4868), .ZN(n4869) );
  AOI22_X1 U5177 ( .A1(n4872), .A2(n4871), .B1(n4870), .B2(n4869), .ZN(n4873)
         );
  OAI211_X1 U5178 ( .C1(n4462), .C2(n4875), .A(n4874), .B(n4873), .ZN(U3280)
         );
  AOI22_X1 U5179 ( .A1(STATE_REG_SCAN_IN), .A2(n4877), .B1(n4876), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5180 ( .A1(n4880), .A2(n4879), .B1(n4878), .B2(n4889), .ZN(n4887)
         );
  INV_X1 U5181 ( .A(n4881), .ZN(n4885) );
  OAI22_X1 U5182 ( .A1(n4885), .A2(n4884), .B1(n4883), .B2(n4882), .ZN(n4886)
         );
  AOI211_X1 U5183 ( .C1(n4889), .C2(n4888), .A(n4887), .B(n4886), .ZN(n4890)
         );
  INV_X1 U5184 ( .A(n4890), .ZN(U3279) );
  AOI22_X1 U5185 ( .A1(STATE_REG_SCAN_IN), .A2(n4892), .B1(n4891), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5186 ( .A1(STATE_REG_SCAN_IN), .A2(n4894), .B1(n4893), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5187 ( .A1(n4898), .A2(n4897), .B1(n4896), .B2(n4895), .ZN(n4903)
         );
  INV_X1 U5188 ( .A(n4899), .ZN(n4900) );
  OAI21_X1 U5189 ( .B1(n3996), .B2(n4901), .A(n4900), .ZN(n4902) );
  NOR2_X1 U5190 ( .A1(n4903), .A2(n4902), .ZN(n4910) );
  XNOR2_X1 U5191 ( .A(n4905), .B(n4904), .ZN(n4906) );
  XNOR2_X1 U5192 ( .A(n3915), .B(n4906), .ZN(n4908) );
  NAND2_X1 U5193 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  OAI211_X1 U5194 ( .C1(n4912), .C2(n4911), .A(n4910), .B(n4909), .ZN(U3238)
         );
  AOI22_X1 U5195 ( .A1(STATE_REG_SCAN_IN), .A2(n4914), .B1(n4913), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n4916), .B1(n4915), .B2(U3149), 
        .ZN(U3324) );
  CLKBUF_X2 U2307 ( .A(n3302), .Z(n2274) );
  CLKBUF_X3 U2311 ( .A(n3302), .Z(n2273) );
  CLKBUF_X1 U2420 ( .A(n2874), .Z(n2998) );
endmodule

