

module b22_C_gen_AntiSAT_k_256_5 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777;

  OR2_X1 U7416 ( .A1(n9087), .A2(n6707), .ZN(n7109) );
  INV_X2 U7417 ( .A(n14636), .ZN(n15074) );
  NAND2_X1 U7418 ( .A1(n8148), .A2(n8147), .ZN(n14039) );
  OAI22_X1 U7419 ( .A1(n12513), .A2(n7577), .B1(n12511), .B2(n12512), .ZN(
        n12518) );
  CLKBUF_X1 U7420 ( .A(n14700), .Z(n6677) );
  OAI21_X1 U7421 ( .B1(n15046), .B2(n10969), .A(n10971), .ZN(n11100) );
  OR2_X2 U7422 ( .A1(n10476), .A2(n11911), .ZN(n14630) );
  INV_X2 U7423 ( .A(n12560), .ZN(n12575) );
  OAI21_X1 U7424 ( .B1(n7386), .B2(n7119), .A(n7117), .ZN(n7928) );
  NAND2_X1 U7425 ( .A1(n7845), .A2(n7387), .ZN(n7386) );
  INV_X1 U7426 ( .A(n12387), .ZN(n15363) );
  BUF_X2 U7427 ( .A(n11935), .Z(n11967) );
  BUF_X2 U7428 ( .A(n7728), .Z(n8203) );
  INV_X1 U7429 ( .A(n10120), .ZN(n11884) );
  INV_X2 U7430 ( .A(n6675), .ZN(n10273) );
  NAND4_X2 U7431 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n14320)
         );
  NAND2_X1 U7432 ( .A1(n6670), .A2(n10090), .ZN(n11817) );
  BUF_X1 U7433 ( .A(n11896), .Z(n6674) );
  CLKBUF_X1 U7434 ( .A(n15665), .Z(n6668) );
  NOR2_X1 U7435 ( .A1(n10794), .A2(n10793), .ZN(n15665) );
  NAND2_X2 U7436 ( .A1(n6928), .A2(n7605), .ZN(n13851) );
  AOI21_X1 U7437 ( .B1(n13822), .B2(n15293), .A(n13821), .ZN(n14030) );
  OAI22_X1 U7438 ( .A1(n7576), .A2(n12461), .B1(n12466), .B2(n12467), .ZN(
        n12475) );
  AOI21_X1 U7439 ( .B1(n12463), .B2(n12462), .A(n12460), .ZN(n12461) );
  INV_X2 U7441 ( .A(n12292), .ZN(n12320) );
  NAND2_X1 U7442 ( .A1(n14141), .A2(n8293), .ZN(n7705) );
  INV_X2 U7443 ( .A(n7705), .ZN(n9740) );
  INV_X1 U7444 ( .A(n13703), .ZN(n6878) );
  INV_X2 U7445 ( .A(n12824), .ZN(n12807) );
  INV_X1 U7446 ( .A(n6686), .ZN(n11309) );
  CLKBUF_X3 U7447 ( .A(n9448), .Z(n10389) );
  CLKBUF_X2 U7448 ( .A(n8454), .Z(n8951) );
  CLKBUF_X2 U7449 ( .A(n13078), .Z(n6678) );
  OR2_X1 U7450 ( .A1(n14881), .A2(n14880), .ZN(n7289) );
  INV_X1 U7451 ( .A(n9868), .ZN(n8725) );
  NAND2_X1 U7452 ( .A1(n8835), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8836) );
  CLKBUF_X2 U7453 ( .A(n11893), .Z(n6676) );
  INV_X1 U7454 ( .A(n12817), .ZN(n12826) );
  CLKBUF_X3 U7455 ( .A(n11896), .Z(n6675) );
  NAND2_X1 U7456 ( .A1(n13624), .A2(n13623), .ZN(n13622) );
  XNOR2_X1 U7457 ( .A(n13508), .B(n13507), .ZN(n13642) );
  XNOR2_X1 U7458 ( .A(n13476), .B(n13474), .ZN(n11669) );
  NOR2_X1 U7459 ( .A1(n13766), .A2(n10446), .ZN(n14009) );
  INV_X1 U7460 ( .A(n14479), .ZN(n14674) );
  NAND2_X1 U7461 ( .A1(n9591), .A2(n9590), .ZN(n10092) );
  NAND2_X1 U7462 ( .A1(n7099), .A2(n9050), .ZN(n9052) );
  XNOR2_X1 U7463 ( .A(n9052), .B(n7562), .ZN(n15770) );
  OR2_X1 U7464 ( .A1(n6684), .A2(n9095), .ZN(n6669) );
  XNOR2_X1 U7465 ( .A(n10621), .B(n10636), .ZN(n15473) );
  NOR2_X2 U7466 ( .A1(n14787), .A2(n14788), .ZN(n14786) );
  NAND2_X2 U7467 ( .A1(n15240), .A2(n15239), .ZN(n15238) );
  MUX2_X1 U7468 ( .A(n11912), .B(n11911), .S(n12091), .Z(n11935) );
  INV_X2 U7469 ( .A(n11935), .ZN(n12017) );
  AND2_X1 U7470 ( .A1(n12083), .A2(n12082), .ZN(n6732) );
  AND2_X2 U7471 ( .A1(n6844), .A2(n6842), .ZN(n8247) );
  INV_X2 U7472 ( .A(n14317), .ZN(n10219) );
  NAND2_X1 U7473 ( .A1(n9591), .A2(n9590), .ZN(n6670) );
  OAI21_X2 U7474 ( .B1(n13096), .B2(n14895), .A(n15541), .ZN(n13097) );
  XNOR2_X2 U7475 ( .A(n7820), .B(n7818), .ZN(n10904) );
  NAND2_X1 U7476 ( .A1(n7803), .A2(n7802), .ZN(n7820) );
  NOR2_X2 U7477 ( .A1(n9056), .A2(n9057), .ZN(n9060) );
  INV_X1 U7478 ( .A(n11936), .ZN(n10266) );
  INV_X1 U7479 ( .A(n6676), .ZN(n6671) );
  NAND2_X1 U7480 ( .A1(n14141), .A2(n8293), .ZN(n6672) );
  NOR2_X4 U7481 ( .A1(n6940), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7675) );
  AOI21_X2 U7482 ( .B1(n13513), .B2(n13643), .A(n6799), .ZN(n13624) );
  CLKBUF_X3 U7483 ( .A(n12368), .Z(n12655) );
  INV_X2 U7484 ( .A(n12368), .ZN(n12383) );
  NAND2_X2 U7485 ( .A1(n7791), .A2(n7790), .ZN(n12411) );
  NOR2_X2 U7486 ( .A1(n15557), .A2(n13051), .ZN(n15576) );
  NOR2_X2 U7487 ( .A1(n15558), .A2(n15559), .ZN(n15557) );
  NAND3_X2 U7488 ( .A1(n6939), .A2(n6941), .A3(n6942), .ZN(n6940) );
  XNOR2_X2 U7489 ( .A(n9771), .B(P1_IR_REG_20__SCAN_IN), .ZN(n11911) );
  BUF_X2 U7490 ( .A(n7908), .Z(n7909) );
  XNOR2_X2 U7491 ( .A(n7088), .B(n9055), .ZN(n14783) );
  NAND2_X2 U7492 ( .A1(n9054), .A2(n9053), .ZN(n7088) );
  XNOR2_X2 U7493 ( .A(n8834), .B(n8833), .ZN(n10344) );
  OAI21_X2 U7494 ( .B1(n10067), .B2(n15749), .A(n10066), .ZN(n10631) );
  NAND2_X1 U7495 ( .A1(n13575), .A2(n9456), .ZN(n13574) );
  NAND4_X2 U7496 ( .A1(n7734), .A2(n7733), .A3(n7732), .A4(n7731), .ZN(n13702)
         );
  NAND2_X1 U7497 ( .A1(n7292), .A2(n7293), .ZN(n7295) );
  AND2_X4 U7498 ( .A1(n13461), .A2(n8443), .ZN(n10766) );
  OAI22_X2 U7499 ( .A1(n13801), .A2(n13789), .B1(n8246), .B2(n8300), .ZN(n8244) );
  OAI21_X2 U7500 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n8991), .A(n8990), .ZN(
        n9029) );
  XNOR2_X2 U7501 ( .A(n9578), .B(n9577), .ZN(n11912) );
  OAI21_X2 U7502 ( .B1(n9770), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9578) );
  NAND4_X4 U7503 ( .A1(n7697), .A2(n7696), .A3(n7695), .A4(n7694), .ZN(n13705)
         );
  INV_X2 U7504 ( .A(n11911), .ZN(n12089) );
  AND2_X1 U7505 ( .A1(n9784), .A2(n9782), .ZN(n11896) );
  NAND2_X1 U7506 ( .A1(n6670), .A2(n11804), .ZN(n11893) );
  OAI21_X1 U7507 ( .B1(n11790), .B2(n11817), .A(n11792), .ZN(n14700) );
  NAND2_X1 U7508 ( .A1(n8419), .A2(n8420), .ZN(n13078) );
  NOR2_X2 U7509 ( .A1(n15620), .A2(n10055), .ZN(n10619) );
  XNOR2_X2 U7510 ( .A(n7297), .B(n10646), .ZN(n10055) );
  XNOR2_X2 U7511 ( .A(n10635), .B(n10636), .ZN(n15469) );
  NAND2_X2 U7512 ( .A1(n10634), .A2(n6865), .ZN(n10635) );
  OAI211_X4 U7513 ( .C1(n7715), .C2(n10091), .A(n7192), .B(n7191), .ZN(n12363)
         );
  OR2_X2 U7514 ( .A1(n7704), .A2(n9501), .ZN(n7192) );
  NAND2_X1 U7515 ( .A1(n10968), .A2(n10967), .ZN(n15046) );
  BUF_X4 U7516 ( .A(n10426), .Z(n6686) );
  NAND4_X2 U7517 ( .A1(n7753), .A2(n7752), .A3(n7751), .A4(n7750), .ZN(n13701)
         );
  AOI21_X2 U7518 ( .B1(n7602), .B2(n7600), .A(n6744), .ZN(n6943) );
  NOR2_X2 U7519 ( .A1(n15455), .A2(n15454), .ZN(n15453) );
  NOR2_X2 U7520 ( .A1(n10619), .A2(n10620), .ZN(n15455) );
  XNOR2_X2 U7521 ( .A(n8836), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12171) );
  OAI222_X1 U7522 ( .A1(n11724), .A2(P2_U3088), .B1(n14150), .B2(n14763), .C1(
        n12144), .C2(n14152), .ZN(P2_U3297) );
  AND2_X1 U7523 ( .A1(n6681), .A2(n11724), .ZN(n7729) );
  AOI21_X2 U7524 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9925), .A(n10025), .ZN(
        n9936) );
  NOR2_X2 U7525 ( .A1(n15453), .A2(n7300), .ZN(n10621) );
  OAI222_X1 U7526 ( .A1(P3_U3151), .A2(n9886), .B1(n11518), .B2(n7383), .C1(
        n13468), .C2(n6816), .ZN(P3_U3293) );
  NOR2_X2 U7527 ( .A1(n15473), .A2(n15474), .ZN(n15472) );
  CLKBUF_X1 U7528 ( .A(n9590), .Z(n6679) );
  XNOR2_X1 U7529 ( .A(n9585), .B(n9584), .ZN(n9590) );
  BUF_X2 U7530 ( .A(n10019), .Z(n6680) );
  OAI211_X1 U7531 ( .C1(n8460), .C2(n8459), .A(n8462), .B(n7296), .ZN(n10019)
         );
  NOR2_X2 U7532 ( .A1(n15001), .A2(n9066), .ZN(n15004) );
  NOR2_X2 U7533 ( .A1(n9065), .A2(n9064), .ZN(n15001) );
  OAI21_X1 U7534 ( .B1(n12533), .B2(n12532), .A(n12531), .ZN(n12538) );
  NAND2_X1 U7535 ( .A1(n8287), .A2(n8286), .ZN(n13833) );
  XNOR2_X1 U7536 ( .A(n13055), .B(n13054), .ZN(n14853) );
  OR2_X1 U7537 ( .A1(n14569), .A2(n14557), .ZN(n14556) );
  NAND2_X1 U7538 ( .A1(n7333), .A2(n7331), .ZN(n14972) );
  OR2_X1 U7539 ( .A1(n11509), .A2(n11510), .ZN(n11583) );
  NAND2_X1 U7540 ( .A1(n7886), .A2(n7885), .ZN(n11032) );
  XNOR2_X1 U7541 ( .A(n7295), .B(n15528), .ZN(n15522) );
  OR2_X1 U7542 ( .A1(n14929), .A2(n11394), .ZN(n11466) );
  NAND2_X1 U7543 ( .A1(n6966), .A2(n10492), .ZN(n10502) );
  NAND2_X1 U7544 ( .A1(n10559), .A2(n15298), .ZN(n15303) );
  NAND2_X1 U7545 ( .A1(n10265), .A2(n10264), .ZN(n11941) );
  INV_X4 U7546 ( .A(n13044), .ZN(P3_U3897) );
  NOR2_X1 U7547 ( .A1(n6713), .A2(n6839), .ZN(n6838) );
  INV_X4 U7551 ( .A(n11160), .ZN(n13922) );
  INV_X2 U7552 ( .A(n8749), .ZN(n7160) );
  INV_X4 U7553 ( .A(n7809), .ZN(n12554) );
  NOR2_X2 U7554 ( .A1(n7652), .A2(n7651), .ZN(n12656) );
  BUF_X1 U7555 ( .A(n9591), .Z(n6688) );
  INV_X2 U7557 ( .A(n11912), .ZN(n12092) );
  XNOR2_X1 U7558 ( .A(n9436), .B(n9441), .ZN(n12838) );
  XNOR2_X1 U7559 ( .A(n9582), .B(n9581), .ZN(n9591) );
  INV_X1 U7560 ( .A(n12682), .ZN(n6681) );
  INV_X1 U7561 ( .A(n9782), .ZN(n9786) );
  BUF_X4 U7562 ( .A(n7692), .Z(n11804) );
  AND2_X1 U7563 ( .A1(n7761), .A2(n7662), .ZN(n6942) );
  OR2_X1 U7564 ( .A1(n7256), .A2(n12124), .ZN(n7255) );
  AOI21_X1 U7565 ( .B1(n13133), .B2(n15732), .A(n13129), .ZN(n13397) );
  AOI211_X1 U7566 ( .C1(n14018), .C2(n15390), .A(n14017), .B(n14016), .ZN(
        n14102) );
  OAI21_X1 U7567 ( .B1(n8962), .B2(n15641), .A(n8961), .ZN(n13121) );
  AOI21_X1 U7568 ( .B1(n14488), .B2(n14792), .A(n14487), .ZN(n14683) );
  AND2_X1 U7569 ( .A1(n12645), .A2(n12644), .ZN(n12647) );
  NAND2_X1 U7570 ( .A1(n12311), .A2(n12310), .ZN(n12313) );
  NAND2_X1 U7571 ( .A1(n11739), .A2(n11738), .ZN(n14397) );
  NAND2_X1 U7572 ( .A1(n14163), .A2(n14164), .ZN(n12784) );
  XNOR2_X1 U7573 ( .A(n13148), .B(n13158), .ZN(n13141) );
  NAND2_X1 U7574 ( .A1(n12774), .A2(n14256), .ZN(n14163) );
  AOI21_X1 U7575 ( .B1(n14495), .B2(n14426), .A(n14447), .ZN(n14485) );
  NAND2_X1 U7576 ( .A1(n13642), .A2(n13510), .ZN(n13643) );
  NAND2_X1 U7577 ( .A1(n7102), .A2(n7108), .ZN(n7105) );
  NAND2_X1 U7578 ( .A1(n13205), .A2(n13204), .ZN(n13207) );
  NAND2_X1 U7579 ( .A1(n8220), .A2(n8219), .ZN(n13797) );
  NAND2_X1 U7580 ( .A1(n12766), .A2(n12765), .ZN(n14186) );
  NAND2_X1 U7581 ( .A1(n11772), .A2(n11771), .ZN(n14688) );
  NAND2_X1 U7582 ( .A1(n7596), .A2(n7595), .ZN(n13882) );
  XNOR2_X1 U7583 ( .A(n8196), .B(n8195), .ZN(n12133) );
  OAI21_X1 U7584 ( .B1(n14268), .B2(n7084), .A(n7413), .ZN(n7083) );
  AND2_X1 U7585 ( .A1(n8161), .A2(n8160), .ZN(n13842) );
  OR2_X1 U7586 ( .A1(n8193), .A2(n8192), .ZN(n8218) );
  NAND2_X1 U7587 ( .A1(n13941), .A2(n8279), .ZN(n13918) );
  AND2_X1 U7588 ( .A1(n6929), .A2(n8277), .ZN(n13942) );
  NAND2_X1 U7589 ( .A1(n8159), .A2(n8146), .ZN(n11790) );
  OR2_X1 U7590 ( .A1(n13949), .A2(n8275), .ZN(n6929) );
  XNOR2_X1 U7591 ( .A(n12728), .B(n12725), .ZN(n14291) );
  NAND2_X1 U7592 ( .A1(n7095), .A2(n7094), .ZN(n7096) );
  XNOR2_X1 U7593 ( .A(n14557), .B(n14566), .ZN(n14548) );
  NAND2_X1 U7594 ( .A1(n6841), .A2(n12631), .ZN(n11632) );
  NAND2_X1 U7595 ( .A1(n11583), .A2(n6965), .ZN(n11667) );
  NAND2_X1 U7596 ( .A1(n8088), .A2(n8087), .ZN(n14120) );
  NAND2_X1 U7597 ( .A1(n11821), .A2(n11820), .ZN(n14590) );
  NAND2_X1 U7598 ( .A1(n14793), .A2(n11291), .ZN(n11292) );
  NAND2_X1 U7599 ( .A1(n11833), .A2(n11832), .ZN(n14728) );
  NAND2_X1 U7600 ( .A1(n8041), .A2(n8040), .ZN(n13934) );
  OAI21_X1 U7601 ( .B1(n11491), .B2(n11490), .A(n11489), .ZN(n11567) );
  NAND2_X1 U7602 ( .A1(n10750), .A2(n8261), .ZN(n10562) );
  OAI21_X1 U7603 ( .B1(n8852), .B2(n7221), .A(n7220), .ZN(n11444) );
  AOI21_X1 U7604 ( .B1(n11278), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11169), .ZN(
        n14356) );
  NAND2_X1 U7605 ( .A1(n10502), .A2(n7366), .ZN(n10610) );
  NAND2_X1 U7606 ( .A1(n7194), .A2(n7193), .ZN(n10839) );
  INV_X1 U7607 ( .A(n10757), .ZN(n7194) );
  NAND2_X1 U7608 ( .A1(n15610), .A2(n15609), .ZN(n15608) );
  NAND2_X1 U7609 ( .A1(n7875), .A2(n7874), .ZN(n15393) );
  NAND2_X1 U7610 ( .A1(n10465), .A2(n10464), .ZN(n10962) );
  INV_X2 U7611 ( .A(n15682), .ZN(n15649) );
  NAND2_X1 U7612 ( .A1(n10912), .A2(n10911), .ZN(n15107) );
  NAND2_X1 U7613 ( .A1(n7841), .A2(n7840), .ZN(n7845) );
  AND2_X1 U7614 ( .A1(n10422), .A2(n10421), .ZN(n11947) );
  NAND2_X1 U7615 ( .A1(n7717), .A2(n7716), .ZN(n15282) );
  BUF_X2 U7616 ( .A(n13493), .Z(n13505) );
  NAND2_X1 U7617 ( .A1(n7299), .A2(n7298), .ZN(n7297) );
  NAND4_X1 U7618 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n15652)
         );
  AND4_X1 U7619 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n15636)
         );
  NAND2_X2 U7620 ( .A1(n6973), .A2(n7652), .ZN(n13493) );
  OR2_X1 U7621 ( .A1(n15718), .A2(n15663), .ZN(n10793) );
  NAND4_X2 U7622 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n14316) );
  INV_X2 U7623 ( .A(n11817), .ZN(n11892) );
  OR2_X1 U7624 ( .A1(n15440), .A2(n15439), .ZN(n7299) );
  AND2_X2 U7625 ( .A1(n12804), .A2(n14630), .ZN(n12817) );
  NAND2_X1 U7626 ( .A1(n7738), .A2(n7739), .ZN(n7741) );
  CLKBUF_X1 U7627 ( .A(n9792), .Z(n9813) );
  NAND4_X2 U7628 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n14317) );
  NAND2_X2 U7629 ( .A1(n11016), .A2(n10086), .ZN(n12824) );
  INV_X4 U7630 ( .A(n7853), .ZN(n8204) );
  NOR2_X1 U7631 ( .A1(n10052), .A2(n10053), .ZN(n15440) );
  NOR2_X1 U7632 ( .A1(n9889), .A2(n9890), .ZN(n10052) );
  OR2_X1 U7633 ( .A1(n15292), .A2(n12610), .ZN(n10446) );
  NAND2_X1 U7634 ( .A1(n7079), .A2(n6724), .ZN(n9792) );
  NAND2_X1 U7635 ( .A1(n8996), .A2(n8997), .ZN(n8998) );
  INV_X1 U7636 ( .A(n11928), .ZN(n11016) );
  AND2_X4 U7637 ( .A1(n8444), .A2(n8443), .ZN(n8465) );
  AND2_X1 U7638 ( .A1(n12092), .A2(n12089), .ZN(n11928) );
  INV_X2 U7639 ( .A(n7704), .ZN(n7760) );
  XNOR2_X1 U7640 ( .A(n8995), .B(n15450), .ZN(n9023) );
  AND2_X1 U7641 ( .A1(n11724), .A2(n12682), .ZN(n7730) );
  AOI21_X1 U7642 ( .B1(n7756), .B2(n7378), .A(n7377), .ZN(n7376) );
  XNOR2_X1 U7643 ( .A(n9438), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U7644 ( .A1(n14762), .A2(n9782), .ZN(n10120) );
  NAND2_X1 U7645 ( .A1(n8417), .A2(n8441), .ZN(n13469) );
  OAI21_X1 U7646 ( .B1(n9035), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n8994), .ZN(
        n8995) );
  OAI21_X1 U7647 ( .B1(n7713), .B2(n7712), .A(n7711), .ZN(n7714) );
  CLKBUF_X1 U7648 ( .A(n8247), .Z(n12646) );
  NAND2_X2 U7649 ( .A1(n12140), .A2(n7668), .ZN(n12682) );
  XNOR2_X1 U7650 ( .A(n9773), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U7651 ( .A1(n9778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9582) );
  OAI21_X1 U7652 ( .B1(n9437), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9436) );
  XNOR2_X1 U7653 ( .A(n9576), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14773) );
  NAND2_X1 U7654 ( .A1(n7669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7670) );
  XNOR2_X1 U7655 ( .A(n9781), .B(n9780), .ZN(n9782) );
  AND2_X1 U7656 ( .A1(n7725), .A2(n7743), .ZN(n9853) );
  MUX2_X1 U7657 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8418), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8420) );
  NAND2_X1 U7658 ( .A1(n7283), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U7659 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U7661 ( .A1(n7465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U7662 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7674), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n7677) );
  AND2_X1 U7663 ( .A1(n10389), .A2(n7085), .ZN(n9450) );
  AND2_X1 U7664 ( .A1(n8693), .A2(n8722), .ZN(n8829) );
  AND3_X1 U7665 ( .A1(n6895), .A2(n8616), .A3(n6894), .ZN(n8904) );
  NOR2_X1 U7666 ( .A1(n9447), .A2(n9446), .ZN(n7405) );
  CLKBUF_X1 U7667 ( .A(n7761), .Z(n7910) );
  AND2_X1 U7668 ( .A1(n7639), .A2(n7664), .ZN(n6941) );
  NAND2_X1 U7669 ( .A1(n7682), .A2(n7707), .ZN(n13711) );
  NAND2_X2 U7670 ( .A1(n7689), .A2(n7688), .ZN(n10090) );
  AND2_X1 U7671 ( .A1(n7636), .A2(n7635), .ZN(n7639) );
  AND3_X1 U7672 ( .A1(n8409), .A2(n8408), .A3(n8407), .ZN(n8616) );
  NAND2_X1 U7673 ( .A1(n7665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7666) );
  AND2_X1 U7674 ( .A1(n7100), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9026) );
  AND2_X1 U7675 ( .A1(n7302), .A2(n7062), .ZN(n7061) );
  NAND2_X1 U7676 ( .A1(n8415), .A2(n7540), .ZN(n7539) );
  INV_X2 U7677 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7302) );
  INV_X1 U7678 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9432) );
  NOR2_X1 U7679 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7064) );
  INV_X1 U7680 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9341) );
  NOR2_X1 U7681 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9819) );
  INV_X4 U7682 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X2 U7683 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10149) );
  INV_X1 U7684 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9822) );
  INV_X1 U7685 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9602) );
  INV_X1 U7686 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9530) );
  INV_X1 U7687 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9431) );
  XNOR2_X1 U7688 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n9025) );
  INV_X4 U7689 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7690 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7100) );
  INV_X1 U7691 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7684) );
  INV_X1 U7692 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10146) );
  NOR2_X1 U7693 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8406) );
  NOR2_X1 U7694 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8405) );
  NOR2_X1 U7695 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7659) );
  NOR2_X1 U7696 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7660) );
  NOR3_X1 U7697 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .A3(
        P2_IR_REG_25__SCAN_IN), .ZN(n7662) );
  INV_X1 U7698 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7640) );
  NOR2_X1 U7699 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7633) );
  NOR2_X1 U7700 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7632) );
  NOR2_X1 U7701 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7638) );
  NOR2_X1 U7702 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7637) );
  INV_X1 U7703 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7763) );
  INV_X1 U7704 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7681) );
  INV_X4 U7705 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7706 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9584) );
  NOR2_X2 U7707 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8461) );
  NOR2_X1 U7708 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7171) );
  BUF_X1 U7709 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n13472) );
  INV_X1 U7710 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9441) );
  NOR2_X1 U7711 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9445) );
  OAI211_X1 U7712 ( .C1(n11567), .C2(n7066), .A(1'b1), .B(n7065), .ZN(n14947)
         );
  NOR2_X2 U7714 ( .A1(n12559), .A2(n13795), .ZN(n13772) );
  NOR2_X2 U7715 ( .A1(n13972), .A2(n13961), .ZN(n7201) );
  NOR2_X1 U7716 ( .A1(n6869), .A2(n6868), .ZN(n6683) );
  AND2_X1 U7717 ( .A1(n7101), .A2(n7105), .ZN(n6684) );
  NOR2_X1 U7718 ( .A1(n6869), .A2(n6868), .ZN(n15000) );
  OR2_X2 U7719 ( .A1(n8340), .A2(n15407), .ZN(n8338) );
  OR2_X2 U7720 ( .A1(n8340), .A2(n15424), .ZN(n8343) );
  INV_X1 U7721 ( .A(n11817), .ZN(n6685) );
  NAND2_X2 U7722 ( .A1(n11292), .A2(n11871), .ZN(n11383) );
  AOI211_X1 U7723 ( .C1(n14320), .C2(n10242), .A(n10241), .B(n10240), .ZN(
        n11126) );
  NAND2_X1 U7724 ( .A1(n11928), .A2(n9792), .ZN(n10426) );
  NOR2_X2 U7725 ( .A1(n15490), .A2(n10624), .ZN(n10626) );
  NOR2_X2 U7726 ( .A1(n15492), .A2(n15491), .ZN(n15490) );
  OR2_X1 U7727 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  AND2_X1 U7728 ( .A1(n12530), .A2(n12529), .ZN(n12533) );
  NAND2_X2 U7729 ( .A1(n10932), .A2(n10931), .ZN(n11349) );
  NAND2_X1 U7730 ( .A1(n14618), .A2(n14617), .ZN(n14616) );
  NAND4_X2 U7731 ( .A1(n7703), .A2(n7702), .A3(n7701), .A4(n7700), .ZN(n13703)
         );
  XNOR2_X2 U7732 ( .A(n9085), .B(n7561), .ZN(n15017) );
  XNOR2_X2 U7733 ( .A(n9518), .B(n9517), .ZN(n10094) );
  NAND2_X2 U7734 ( .A1(n8247), .A2(n11216), .ZN(n7652) );
  NAND2_X1 U7735 ( .A1(n7647), .A2(n7644), .ZN(n11216) );
  AND2_X2 U7736 ( .A1(n8489), .A2(n10069), .ZN(n8502) );
  NOR2_X2 U7737 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8489) );
  NOR2_X2 U7738 ( .A1(n14556), .A2(n6677), .ZN(n7179) );
  AOI22_X2 U7739 ( .A1(n14438), .A2(n14624), .B1(n14735), .B2(n14437), .ZN(
        n14618) );
  XNOR2_X1 U7740 ( .A(n11941), .B(n14316), .ZN(n11936) );
  NAND2_X2 U7741 ( .A1(n14531), .A2(n14543), .ZN(n14535) );
  NOR2_X2 U7742 ( .A1(n14506), .A2(n14425), .ZN(n14491) );
  AOI21_X2 U7743 ( .B1(n12321), .B2(n7529), .A(n12351), .ZN(n12324) );
  NOR2_X2 U7744 ( .A1(n7110), .A2(n15015), .ZN(n9085) );
  NOR2_X2 U7745 ( .A1(n13994), .A2(n14084), .ZN(n13993) );
  OAI22_X2 U7746 ( .A1(n14527), .A2(n14526), .B1(n7178), .B2(n14445), .ZN(
        n14503) );
  INV_X1 U7747 ( .A(n7704), .ZN(n6687) );
  NAND2_X1 U7748 ( .A1(n7705), .A2(n10090), .ZN(n7704) );
  AOI21_X2 U7749 ( .B1(n14519), .B2(n14526), .A(n7130), .ZN(n14508) );
  OAI21_X2 U7750 ( .B1(n11100), .B2(n10973), .A(n10972), .ZN(n11256) );
  CLKBUF_X1 U7751 ( .A(n10120), .Z(n6689) );
  NOR2_X1 U7752 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8409) );
  NOR2_X1 U7753 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8408) );
  NOR2_X1 U7754 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8407) );
  AND2_X1 U7755 ( .A1(n8444), .A2(n13463), .ZN(n8454) );
  NAND2_X1 U7756 ( .A1(n12883), .A2(n13169), .ZN(n7150) );
  OR2_X1 U7757 ( .A1(n13209), .A2(n13217), .ZN(n12291) );
  NOR2_X1 U7758 ( .A1(n8861), .A2(n7236), .ZN(n7235) );
  INV_X1 U7759 ( .A(n8858), .ZN(n7236) );
  AND2_X1 U7760 ( .A1(n8924), .A2(n8910), .ZN(n9429) );
  NOR2_X1 U7761 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n6901) );
  NOR2_X1 U7762 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n6902) );
  AND2_X1 U7763 ( .A1(n8412), .A2(n8413), .ZN(n6898) );
  INV_X1 U7764 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8412) );
  AND2_X1 U7765 ( .A1(n8404), .A2(n8511), .ZN(n6899) );
  NAND2_X1 U7766 ( .A1(n8748), .A2(n7028), .ZN(n7492) );
  NOR2_X1 U7767 ( .A1(n7031), .A2(n7029), .ZN(n7028) );
  INV_X1 U7768 ( .A(n8390), .ZN(n7029) );
  INV_X1 U7769 ( .A(n7495), .ZN(n7031) );
  NOR2_X1 U7770 ( .A1(n7922), .A2(n7520), .ZN(n7519) );
  INV_X1 U7771 ( .A(n7522), .ZN(n7520) );
  NAND2_X1 U7772 ( .A1(n14566), .A2(n7074), .ZN(n12775) );
  NAND2_X1 U7773 ( .A1(n14587), .A2(n14564), .ZN(n7452) );
  NOR2_X1 U7774 ( .A1(n7324), .A2(n14617), .ZN(n7323) );
  INV_X1 U7775 ( .A(n7326), .ZN(n7324) );
  NAND2_X1 U7776 ( .A1(n14735), .A2(n14416), .ZN(n7330) );
  NAND2_X1 U7777 ( .A1(n7149), .A2(n7150), .ZN(n7148) );
  INV_X1 U7778 ( .A(n13019), .ZN(n7149) );
  AND2_X1 U7779 ( .A1(n13461), .A2(n13463), .ZN(n8488) );
  OR2_X1 U7780 ( .A1(n13278), .A2(n13256), .ZN(n12264) );
  AND4_X1 U7781 ( .A1(n8494), .A2(n8493), .A3(n8492), .A4(n8491), .ZN(n15623)
         );
  AND2_X1 U7782 ( .A1(n8904), .A2(n6773), .ZN(n8439) );
  INV_X1 U7783 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U7784 ( .A1(n8904), .A2(n7538), .ZN(n8419) );
  NAND2_X1 U7785 ( .A1(n11667), .A2(n11666), .ZN(n13476) );
  AOI21_X1 U7786 ( .B1(n6933), .B2(n6934), .A(n13800), .ZN(n6932) );
  NAND2_X1 U7787 ( .A1(n14773), .A2(n11166), .ZN(n10086) );
  OR2_X1 U7788 ( .A1(n14773), .A2(n12092), .ZN(n10476) );
  NAND2_X1 U7789 ( .A1(n12365), .A2(n12364), .ZN(n12376) );
  AOI22_X1 U7790 ( .A1(n12383), .A2(n13704), .B1(n12368), .B2(n12363), .ZN(
        n12375) );
  OAI21_X1 U7791 ( .B1(n6691), .B2(n6702), .A(n6753), .ZN(n12055) );
  NAND2_X1 U7792 ( .A1(n12085), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U7793 ( .A1(n7266), .A2(n12088), .ZN(n7265) );
  INV_X1 U7794 ( .A(n7269), .ZN(n7266) );
  OAI21_X1 U7795 ( .B1(n7866), .B2(SI_10_), .A(n7890), .ZN(n7887) );
  AOI21_X1 U7796 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n9090), .A(n9089), .ZN(
        n9091) );
  NAND2_X1 U7797 ( .A1(n13215), .A2(n8875), .ZN(n7208) );
  OR2_X1 U7798 ( .A1(n13220), .A2(n13199), .ZN(n12285) );
  OR2_X1 U7799 ( .A1(n12933), .A2(n13238), .ZN(n12281) );
  INV_X1 U7800 ( .A(n8851), .ZN(n7227) );
  NAND2_X1 U7801 ( .A1(n12191), .A2(n12190), .ZN(n8847) );
  NAND2_X1 U7802 ( .A1(n12183), .A2(n12184), .ZN(n8844) );
  AND2_X1 U7803 ( .A1(n10344), .A2(n13089), .ZN(n10194) );
  INV_X1 U7804 ( .A(n12359), .ZN(n8843) );
  NOR2_X1 U7805 ( .A1(n7539), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7538) );
  AOI21_X1 U7806 ( .B1(n7495), .B2(n7494), .A(n6810), .ZN(n7493) );
  INV_X1 U7807 ( .A(n8391), .ZN(n7494) );
  NAND2_X1 U7808 ( .A1(n8615), .A2(n8370), .ZN(n8371) );
  NAND2_X1 U7809 ( .A1(n7022), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7021) );
  OAI21_X1 U7810 ( .B1(n7482), .B2(n7481), .A(n8557), .ZN(n7480) );
  NAND2_X1 U7811 ( .A1(n9546), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8355) );
  AOI21_X1 U7812 ( .B1(n13490), .B2(n13654), .A(n6760), .ZN(n7354) );
  AND2_X1 U7813 ( .A1(n8282), .A2(n7598), .ZN(n7597) );
  OR2_X1 U7814 ( .A1(n13917), .A2(n7599), .ZN(n7598) );
  NAND2_X1 U7815 ( .A1(n13942), .A2(n13943), .ZN(n13941) );
  AOI21_X1 U7816 ( .B1(n12624), .B2(n7587), .A(n7586), .ZN(n7585) );
  NAND2_X1 U7817 ( .A1(n10562), .A2(n7584), .ZN(n7583) );
  INV_X1 U7818 ( .A(n8263), .ZN(n7586) );
  XNOR2_X1 U7819 ( .A(n15363), .B(n13702), .ZN(n12613) );
  NAND2_X1 U7820 ( .A1(n7370), .A2(n7369), .ZN(n7368) );
  NOR2_X1 U7821 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7369) );
  INV_X1 U7822 ( .A(n12101), .ZN(n7259) );
  AOI21_X1 U7823 ( .B1(n12104), .B2(n12103), .A(n12102), .ZN(n7258) );
  NAND2_X1 U7824 ( .A1(n14583), .A2(n14419), .ZN(n6891) );
  OR2_X1 U7825 ( .A1(n12721), .A2(n12726), .ZN(n12013) );
  AND2_X1 U7826 ( .A1(n9518), .A2(n9432), .ZN(n7063) );
  AND2_X1 U7827 ( .A1(n7172), .A2(n7171), .ZN(n7407) );
  NOR2_X1 U7828 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7172) );
  NAND2_X1 U7829 ( .A1(n8060), .A2(n8059), .ZN(n8080) );
  NAND2_X1 U7830 ( .A1(n8037), .A2(n8023), .ZN(n8038) );
  NAND2_X1 U7831 ( .A1(n7986), .A2(n7985), .ZN(n8003) );
  XNOR2_X1 U7832 ( .A(n7925), .B(n9541), .ZN(n7923) );
  XNOR2_X1 U7833 ( .A(n7903), .B(SI_11_), .ZN(n7906) );
  NAND2_X1 U7834 ( .A1(n9604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U7835 ( .A1(n7379), .A2(n7381), .ZN(n7739) );
  NAND2_X1 U7836 ( .A1(n7382), .A2(n7720), .ZN(n7379) );
  AOI21_X1 U7837 ( .B1(n7145), .B2(n7143), .A(n6751), .ZN(n7142) );
  INV_X1 U7838 ( .A(n6709), .ZN(n7143) );
  AOI211_X1 U7839 ( .C1(n12900), .C2(n13229), .A(n12874), .B(n12901), .ZN(
        n12880) );
  OR2_X1 U7840 ( .A1(n13010), .A2(n13011), .ZN(n13008) );
  OAI21_X1 U7841 ( .B1(n13141), .B2(n13140), .A(n13139), .ZN(n13142) );
  NAND2_X1 U7842 ( .A1(n7219), .A2(n7218), .ZN(n13139) );
  AND2_X1 U7843 ( .A1(n7219), .A2(n6721), .ZN(n13140) );
  NAND2_X1 U7844 ( .A1(n13154), .A2(n8882), .ZN(n7219) );
  AOI21_X1 U7845 ( .B1(n13141), .B2(n13138), .A(n6913), .ZN(n13147) );
  OAI21_X1 U7846 ( .B1(n13156), .B2(n12301), .A(n12299), .ZN(n13136) );
  NAND2_X1 U7847 ( .A1(n13198), .A2(n7629), .ZN(n13185) );
  OR2_X1 U7848 ( .A1(n13343), .A2(n13217), .ZN(n7629) );
  AND2_X1 U7849 ( .A1(n12291), .A2(n8779), .ZN(n13204) );
  NAND2_X1 U7850 ( .A1(n8432), .A2(n9388), .ZN(n8761) );
  INV_X1 U7851 ( .A(n8752), .ZN(n8432) );
  NAND2_X1 U7852 ( .A1(n8733), .A2(n7525), .ZN(n13244) );
  NOR2_X1 U7853 ( .A1(n13241), .A2(n7526), .ZN(n7525) );
  INV_X1 U7854 ( .A(n12276), .ZN(n7526) );
  AND4_X1 U7855 ( .A1(n8716), .A2(n8715), .A3(n8714), .A4(n8713), .ZN(n13256)
         );
  OR2_X1 U7856 ( .A1(n13448), .A2(n12992), .ZN(n12246) );
  NAND2_X1 U7857 ( .A1(n8859), .A2(n7235), .ZN(n7234) );
  AND4_X1 U7858 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n12849)
         );
  NAND2_X1 U7859 ( .A1(n7224), .A2(n7228), .ZN(n11247) );
  INV_X1 U7860 ( .A(n15655), .ZN(n15624) );
  NAND2_X1 U7861 ( .A1(n7054), .A2(n8474), .ZN(n15646) );
  AND2_X1 U7862 ( .A1(n8473), .A2(n7055), .ZN(n7054) );
  NAND2_X1 U7863 ( .A1(n7160), .A2(n6816), .ZN(n8474) );
  NAND2_X1 U7864 ( .A1(n13469), .A2(n6717), .ZN(n8473) );
  INV_X1 U7865 ( .A(n15673), .ZN(n15654) );
  INV_X1 U7866 ( .A(n15641), .ZN(n15671) );
  AND2_X1 U7867 ( .A1(n8932), .A2(n8931), .ZN(n10792) );
  INV_X1 U7868 ( .A(n12152), .ZN(n8947) );
  NAND2_X1 U7869 ( .A1(n8924), .A2(n8912), .ZN(n9547) );
  INV_X1 U7870 ( .A(n9547), .ZN(n8928) );
  XNOR2_X1 U7871 ( .A(n8440), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U7872 ( .A1(n13453), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8440) );
  XNOR2_X1 U7873 ( .A(n8442), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U7874 ( .A1(n8441), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8442) );
  AND2_X1 U7875 ( .A1(n7135), .A2(n6899), .ZN(n6894) );
  NOR2_X1 U7876 ( .A1(n6897), .A2(n6896), .ZN(n6895) );
  OAI21_X1 U7877 ( .B1(n8780), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8394), .ZN(
        n8792) );
  NAND2_X1 U7878 ( .A1(n7030), .A2(n7475), .ZN(n8748) );
  AOI21_X1 U7879 ( .B1(n8388), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n7476), .ZN(
        n7475) );
  INV_X1 U7880 ( .A(n8745), .ZN(n7476) );
  INV_X1 U7881 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U7882 ( .A1(n8358), .A2(n7482), .ZN(n8542) );
  NAND2_X1 U7883 ( .A1(n8351), .A2(n8350), .ZN(n8496) );
  NAND2_X1 U7884 ( .A1(n6969), .A2(n6968), .ZN(n11509) );
  AOI21_X1 U7885 ( .B1(n6970), .B2(n6692), .A(n6754), .ZN(n6968) );
  NAND2_X1 U7886 ( .A1(n13851), .A2(n13850), .ZN(n8287) );
  NAND2_X1 U7887 ( .A1(n8138), .A2(n13881), .ZN(n7508) );
  NAND2_X1 U7888 ( .A1(n7509), .A2(n8138), .ZN(n7507) );
  INV_X1 U7889 ( .A(n12633), .ZN(n13943) );
  NAND2_X1 U7890 ( .A1(n7582), .A2(n14912), .ZN(n7580) );
  AOI21_X1 U7891 ( .B1(n7519), .B2(n7902), .A(n6716), .ZN(n7518) );
  OR2_X1 U7892 ( .A1(n12459), .A2(n13693), .ZN(n7522) );
  NAND2_X1 U7893 ( .A1(n6940), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U7894 ( .A1(n8104), .A2(SI_22_), .ZN(n8119) );
  INV_X1 U7895 ( .A(n7370), .ZN(n7367) );
  AOI21_X1 U7896 ( .B1(n7415), .B2(n7416), .A(n7414), .ZN(n7413) );
  INV_X1 U7897 ( .A(n14237), .ZN(n7414) );
  NAND2_X1 U7898 ( .A1(n7422), .A2(n14231), .ZN(n7421) );
  INV_X1 U7899 ( .A(n14165), .ZN(n7422) );
  NAND2_X1 U7900 ( .A1(n9793), .A2(n7614), .ZN(n9794) );
  NAND2_X1 U7901 ( .A1(n9791), .A2(n14775), .ZN(n9793) );
  NAND2_X1 U7902 ( .A1(n14927), .A2(n12720), .ZN(n12728) );
  NOR4_X1 U7903 ( .A1(n12122), .A2(n11909), .A3(n14450), .A4(n11908), .ZN(
        n11910) );
  NOR2_X1 U7904 ( .A1(n7338), .A2(n7344), .ZN(n7337) );
  NOR2_X1 U7905 ( .A1(n14421), .A2(n14444), .ZN(n7344) );
  NAND2_X1 U7906 ( .A1(n7448), .A2(n7452), .ZN(n7446) );
  NAND2_X1 U7907 ( .A1(n14442), .A2(n7449), .ZN(n7448) );
  NAND2_X1 U7908 ( .A1(n14595), .A2(n7451), .ZN(n7449) );
  NAND2_X1 U7909 ( .A1(n6770), .A2(n7330), .ZN(n7326) );
  XNOR2_X1 U7910 ( .A(n14638), .B(n14416), .ZN(n14629) );
  AND2_X1 U7911 ( .A1(n12013), .A2(n12014), .ZN(n11876) );
  INV_X1 U7912 ( .A(n7460), .ZN(n7459) );
  INV_X1 U7913 ( .A(n10976), .ZN(n7461) );
  NAND2_X1 U7914 ( .A1(n7348), .A2(n10248), .ZN(n10234) );
  INV_X1 U7915 ( .A(n14667), .ZN(n6858) );
  NAND2_X1 U7916 ( .A1(n11722), .A2(n11721), .ZN(n11734) );
  NAND2_X1 U7917 ( .A1(n10389), .A2(n7284), .ZN(n11025) );
  NAND2_X1 U7918 ( .A1(n7845), .A2(n7844), .ZN(n7865) );
  OR2_X1 U7919 ( .A1(n7690), .A2(SI_1_), .ZN(n7691) );
  NAND2_X1 U7920 ( .A1(n6821), .A2(n9063), .ZN(n6871) );
  NAND2_X1 U7921 ( .A1(n7101), .A2(n7105), .ZN(n7554) );
  INV_X1 U7922 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U7923 ( .A1(n10703), .A2(n10702), .ZN(n10822) );
  OAI21_X1 U7924 ( .B1(n6926), .B2(n12357), .A(n6734), .ZN(n7034) );
  XNOR2_X1 U7925 ( .A(n6927), .B(n13058), .ZN(n6926) );
  AOI21_X1 U7926 ( .B1(n7531), .B2(n7530), .A(n7527), .ZN(n6927) );
  NAND2_X1 U7927 ( .A1(n14871), .A2(n6862), .ZN(n13107) );
  OR2_X1 U7928 ( .A1(n14869), .A2(n13371), .ZN(n6862) );
  NAND2_X1 U7929 ( .A1(n8738), .A2(n8737), .ZN(n13247) );
  INV_X1 U7930 ( .A(n13604), .ZN(n7350) );
  NAND2_X1 U7931 ( .A1(n9481), .A2(n15298), .ZN(n13668) );
  NAND2_X1 U7932 ( .A1(n14947), .A2(n12696), .ZN(n14200) );
  NAND2_X1 U7933 ( .A1(n14450), .A2(n6708), .ZN(n7372) );
  NAND2_X1 U7934 ( .A1(n7121), .A2(n6741), .ZN(n7305) );
  XNOR2_X1 U7935 ( .A(n14451), .B(n14428), .ZN(n14669) );
  NAND2_X1 U7936 ( .A1(n6840), .A2(n6740), .ZN(n14451) );
  INV_X1 U7937 ( .A(n9086), .ZN(n7561) );
  INV_X1 U7938 ( .A(n12386), .ZN(n6829) );
  NAND2_X1 U7939 ( .A1(n7180), .A2(n10219), .ZN(n7245) );
  OAI21_X1 U7940 ( .B1(n11966), .B2(n7281), .A(n7280), .ZN(n11970) );
  NAND2_X1 U7941 ( .A1(n7282), .A2(n11964), .ZN(n7280) );
  NOR2_X1 U7942 ( .A1(n7282), .A2(n11964), .ZN(n7281) );
  INV_X1 U7943 ( .A(n11970), .ZN(n11973) );
  AOI21_X1 U7944 ( .B1(n12012), .B2(n7276), .A(n7275), .ZN(n7274) );
  INV_X1 U7945 ( .A(n12015), .ZN(n7275) );
  NAND2_X1 U7946 ( .A1(n7279), .A2(n6736), .ZN(n7276) );
  AND2_X1 U7947 ( .A1(n12500), .A2(n7544), .ZN(n7542) );
  NAND2_X1 U7948 ( .A1(n12494), .A2(n12493), .ZN(n7544) );
  NAND2_X1 U7949 ( .A1(n6768), .A2(n12500), .ZN(n7543) );
  NAND2_X1 U7950 ( .A1(n7550), .A2(n7549), .ZN(n7548) );
  NAND2_X1 U7951 ( .A1(n7547), .A2(n7546), .ZN(n7545) );
  NAND2_X1 U7952 ( .A1(n12057), .A2(n12056), .ZN(n12060) );
  AND2_X1 U7953 ( .A1(n12511), .A2(n12512), .ZN(n7577) );
  OAI21_X1 U7954 ( .B1(n12524), .B2(n7568), .A(n7565), .ZN(n12530) );
  AND2_X1 U7955 ( .A1(n12522), .A2(n12523), .ZN(n7568) );
  NAND2_X1 U7956 ( .A1(n7567), .A2(n7566), .ZN(n7565) );
  INV_X1 U7957 ( .A(n13155), .ZN(n7012) );
  AND2_X1 U7958 ( .A1(n12084), .A2(n7270), .ZN(n7269) );
  AOI21_X1 U7959 ( .B1(n12088), .B2(n7264), .A(n7263), .ZN(n7262) );
  INV_X1 U7960 ( .A(n7267), .ZN(n7264) );
  INV_X1 U7961 ( .A(n12086), .ZN(n7263) );
  NAND2_X1 U7962 ( .A1(n8021), .A2(n9840), .ZN(n7394) );
  NAND2_X1 U7963 ( .A1(n7491), .A2(n12316), .ZN(n12319) );
  AND2_X1 U7964 ( .A1(n12305), .A2(n12304), .ZN(n7491) );
  OR2_X1 U7965 ( .A1(n13335), .A2(n13157), .ZN(n12162) );
  AND2_X1 U7966 ( .A1(n7042), .A2(n13316), .ZN(n7041) );
  OR2_X1 U7967 ( .A1(n7532), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U7968 ( .A1(n15431), .A2(n15650), .ZN(n12180) );
  INV_X1 U7969 ( .A(n13480), .ZN(n6987) );
  INV_X1 U7970 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6845) );
  OAI21_X1 U7971 ( .B1(n11099), .B2(n7319), .A(n11865), .ZN(n7318) );
  INV_X1 U7972 ( .A(n10908), .ZN(n7319) );
  NAND2_X1 U7973 ( .A1(n7968), .A2(n9638), .ZN(n7985) );
  OAI21_X1 U7974 ( .B1(n11804), .B2(n9508), .A(n6875), .ZN(n7722) );
  NAND2_X1 U7975 ( .A1(n7692), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U7976 ( .A1(n10652), .A2(n7301), .ZN(n7300) );
  NAND2_X1 U7977 ( .A1(n6697), .A2(n12163), .ZN(n6912) );
  NAND2_X1 U7978 ( .A1(n6909), .A2(n8965), .ZN(n6908) );
  NAND2_X1 U7979 ( .A1(n6697), .A2(n6910), .ZN(n6909) );
  NOR2_X1 U7980 ( .A1(n8803), .A2(n13173), .ZN(n6910) );
  NAND2_X1 U7981 ( .A1(n8826), .A2(n6916), .ZN(n6915) );
  NAND2_X1 U7982 ( .A1(n12301), .A2(n12299), .ZN(n6916) );
  NOR2_X1 U7983 ( .A1(n13025), .A2(n13169), .ZN(n12301) );
  NAND2_X1 U7984 ( .A1(n8434), .A2(n8433), .ZN(n8795) );
  INV_X1 U7985 ( .A(n8783), .ZN(n8434) );
  INV_X1 U7986 ( .A(n7038), .ZN(n6918) );
  AOI21_X1 U7987 ( .B1(n7041), .B2(n7043), .A(n7039), .ZN(n7038) );
  INV_X1 U7988 ( .A(n12243), .ZN(n7039) );
  AND2_X1 U7989 ( .A1(n7041), .A2(n6921), .ZN(n6920) );
  NAND2_X1 U7990 ( .A1(n12337), .A2(n7534), .ZN(n6921) );
  NOR2_X1 U7991 ( .A1(n12249), .A2(n7535), .ZN(n7534) );
  INV_X1 U7992 ( .A(n12240), .ZN(n7535) );
  NOR2_X1 U7993 ( .A1(n7052), .A2(n12223), .ZN(n7051) );
  INV_X1 U7994 ( .A(n8563), .ZN(n7052) );
  OR2_X1 U7995 ( .A1(n12218), .A2(n12216), .ZN(n7228) );
  AND3_X1 U7996 ( .A1(n8486), .A2(n8485), .A3(n8484), .ZN(n10366) );
  OR2_X1 U7997 ( .A1(n12171), .A2(n10344), .ZN(n12353) );
  INV_X1 U7998 ( .A(n7008), .ZN(n7007) );
  INV_X1 U7999 ( .A(n7470), .ZN(n7004) );
  AOI21_X1 U8000 ( .B1(n7472), .B2(n7474), .A(n7471), .ZN(n7470) );
  INV_X1 U8001 ( .A(n8366), .ZN(n7471) );
  AOI21_X1 U8002 ( .B1(n7479), .B2(n7481), .A(n7009), .ZN(n7008) );
  INV_X1 U8003 ( .A(n8362), .ZN(n7009) );
  AND2_X1 U8004 ( .A1(n7483), .A2(n8357), .ZN(n7482) );
  INV_X1 U8005 ( .A(n8539), .ZN(n7483) );
  NOR2_X1 U8006 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6900) );
  NAND2_X1 U8007 ( .A1(n7552), .A2(n12550), .ZN(n7551) );
  AND2_X1 U8008 ( .A1(n12645), .A2(n12567), .ZN(n12600) );
  OR2_X1 U8009 ( .A1(n6938), .A2(n6718), .ZN(n6934) );
  INV_X1 U8010 ( .A(n7506), .ZN(n7502) );
  NOR2_X1 U8011 ( .A1(n8190), .A2(n7505), .ZN(n7504) );
  INV_X1 U8012 ( .A(n8170), .ZN(n7505) );
  OR2_X1 U8013 ( .A1(n14111), .A2(n13808), .ZN(n12637) );
  AND2_X1 U8014 ( .A1(n12638), .A2(n8157), .ZN(n7506) );
  INV_X1 U8015 ( .A(n6961), .ZN(n6960) );
  NAND2_X1 U8016 ( .A1(n7876), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U8017 ( .A1(n10562), .A2(n10563), .ZN(n10561) );
  INV_X1 U8018 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U8019 ( .A1(n14420), .A2(n7074), .ZN(n12767) );
  NOR2_X1 U8020 ( .A1(n14728), .A2(n7189), .ZN(n7188) );
  INV_X1 U8021 ( .A(n7190), .ZN(n7189) );
  NOR2_X1 U8022 ( .A1(n7312), .A2(n11869), .ZN(n7311) );
  NOR2_X1 U8023 ( .A1(n11866), .A2(n7313), .ZN(n7312) );
  INV_X1 U8024 ( .A(n10947), .ZN(n7313) );
  AND2_X1 U8025 ( .A1(n11357), .A2(n10975), .ZN(n7464) );
  OAI21_X1 U8026 ( .B1(n8235), .B2(n8234), .A(n8233), .ZN(n11718) );
  OAI21_X1 U8027 ( .B1(n8172), .B2(n8171), .A(n8175), .ZN(n8193) );
  AND2_X1 U8028 ( .A1(n7086), .A2(n6774), .ZN(n7085) );
  INV_X1 U8029 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U8030 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U8031 ( .A1(n8141), .A2(SI_24_), .ZN(n8158) );
  INV_X1 U8032 ( .A(n10090), .ZN(n7692) );
  AND2_X1 U8033 ( .A1(n7625), .A2(n7087), .ZN(n7086) );
  INV_X1 U8034 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U8035 ( .A1(n7987), .A2(n9711), .ZN(n8004) );
  AND2_X1 U8036 ( .A1(n9439), .A2(n9440), .ZN(n7286) );
  INV_X1 U8037 ( .A(n7906), .ZN(n7120) );
  AOI21_X1 U8038 ( .B1(n7888), .B2(n7390), .A(n7389), .ZN(n7388) );
  INV_X1 U8039 ( .A(n7890), .ZN(n7389) );
  INV_X1 U8040 ( .A(n7864), .ZN(n7390) );
  NOR2_X1 U8041 ( .A1(n7391), .A2(n7843), .ZN(n7387) );
  INV_X1 U8042 ( .A(n7888), .ZN(n7391) );
  AND2_X1 U8043 ( .A1(n7124), .A2(n7802), .ZN(n7123) );
  AND2_X1 U8044 ( .A1(n7821), .A2(n7780), .ZN(n7124) );
  NAND2_X1 U8045 ( .A1(n7384), .A2(n7821), .ZN(n7125) );
  OAI21_X1 U8046 ( .B1(n7785), .B2(n7385), .A(n7819), .ZN(n7384) );
  OR2_X1 U8047 ( .A1(n9555), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9596) );
  INV_X1 U8048 ( .A(n10090), .ZN(n7239) );
  INV_X1 U8049 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n8991) );
  INV_X1 U8050 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9024) );
  AOI22_X1 U8051 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9047), .B1(n9049), .B2(
        n9001), .ZN(n9002) );
  OAI21_X1 U8052 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n9632), .A(n9005), .ZN(
        n9058) );
  OAI21_X1 U8053 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14359), .A(n9076), .ZN(
        n9082) );
  NOR2_X1 U8054 ( .A1(n9094), .A2(n9093), .ZN(n9097) );
  AND2_X1 U8055 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9092), .ZN(n9093) );
  NAND2_X1 U8056 ( .A1(n11535), .A2(n7168), .ZN(n11649) );
  NOR2_X1 U8057 ( .A1(n11538), .A2(n7169), .ZN(n7168) );
  INV_X1 U8058 ( .A(n11534), .ZN(n7169) );
  NAND2_X1 U8059 ( .A1(n12879), .A2(n7140), .ZN(n7139) );
  INV_X1 U8060 ( .A(n12919), .ZN(n7146) );
  INV_X1 U8061 ( .A(n12942), .ZN(n7140) );
  INV_X1 U8062 ( .A(n6680), .ZN(n7241) );
  NOR2_X1 U8063 ( .A1(n11804), .A2(n9527), .ZN(n7238) );
  NOR2_X1 U8064 ( .A1(n15652), .A2(n12170), .ZN(n15651) );
  AND2_X1 U8065 ( .A1(n10300), .A2(n10177), .ZN(n10184) );
  NOR2_X1 U8066 ( .A1(n7159), .A2(n7155), .ZN(n7154) );
  INV_X1 U8067 ( .A(n12890), .ZN(n7155) );
  INV_X1 U8068 ( .A(n13031), .ZN(n7159) );
  NAND2_X1 U8069 ( .A1(n13031), .A2(n7158), .ZN(n7157) );
  INV_X1 U8070 ( .A(n12854), .ZN(n7158) );
  AND3_X1 U8071 ( .A1(n8580), .A2(n8579), .A3(n8578), .ZN(n11434) );
  OR2_X1 U8072 ( .A1(n11432), .A2(n11433), .ZN(n11535) );
  NAND2_X1 U8073 ( .A1(n12934), .A2(n12873), .ZN(n12901) );
  NAND2_X1 U8074 ( .A1(n12159), .A2(n12311), .ZN(n7531) );
  NOR2_X1 U8075 ( .A1(n12351), .A2(n12158), .ZN(n7530) );
  AND4_X1 U8076 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n11228)
         );
  INV_X1 U8077 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9885) );
  INV_X1 U8078 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U8079 ( .A1(n15437), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7298) );
  XNOR2_X1 U8080 ( .A(n10640), .B(n10625), .ZN(n15509) );
  AOI21_X1 U8081 ( .B1(n10627), .B2(n7294), .A(n13045), .ZN(n7293) );
  AND2_X1 U8082 ( .A1(n15552), .A2(n13067), .ZN(n15569) );
  NOR2_X1 U8083 ( .A1(n15538), .A2(n6889), .ZN(n13050) );
  NOR2_X1 U8084 ( .A1(n13096), .A2(n11525), .ZN(n6889) );
  NOR2_X1 U8085 ( .A1(n15574), .A2(n7291), .ZN(n13052) );
  AND2_X1 U8086 ( .A1(n15583), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U8087 ( .A1(n14872), .A2(n14873), .ZN(n14871) );
  OR2_X1 U8088 ( .A1(n8885), .A2(n12922), .ZN(n8887) );
  NAND2_X1 U8089 ( .A1(n7210), .A2(n7215), .ZN(n8885) );
  OAI21_X1 U8090 ( .B1(n13154), .B2(n7214), .A(n7211), .ZN(n8942) );
  AOI21_X1 U8091 ( .B1(n7215), .B2(n7213), .A(n7212), .ZN(n7211) );
  INV_X1 U8092 ( .A(n7215), .ZN(n7214) );
  INV_X1 U8093 ( .A(n7217), .ZN(n7213) );
  XNOR2_X1 U8094 ( .A(n12976), .B(n13200), .ZN(n13184) );
  NAND2_X1 U8095 ( .A1(n7035), .A2(n12285), .ZN(n13205) );
  NAND2_X1 U8096 ( .A1(n7208), .A2(n6737), .ZN(n13198) );
  INV_X1 U8097 ( .A(n13254), .ZN(n13261) );
  NAND2_X1 U8098 ( .A1(n8431), .A2(n8430), .ZN(n8739) );
  INV_X1 U8099 ( .A(n8728), .ZN(n8431) );
  INV_X1 U8100 ( .A(n7232), .ZN(n7231) );
  AOI21_X1 U8101 ( .B1(n7232), .B2(n7230), .A(n6746), .ZN(n7229) );
  AND2_X1 U8102 ( .A1(n12340), .A2(n11620), .ZN(n7532) );
  AND2_X1 U8103 ( .A1(n12257), .A2(n12243), .ZN(n13316) );
  NAND2_X1 U8104 ( .A1(n8629), .A2(n7534), .ZN(n7533) );
  NOR2_X1 U8105 ( .A1(n12340), .A2(n7233), .ZN(n7232) );
  INV_X1 U8106 ( .A(n8860), .ZN(n7233) );
  NAND2_X1 U8107 ( .A1(n7234), .A2(n8860), .ZN(n11678) );
  NAND2_X1 U8108 ( .A1(n11528), .A2(n11527), .ZN(n8629) );
  AND4_X1 U8109 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n12994)
         );
  AOI21_X1 U8110 ( .B1(n7049), .B2(n7051), .A(n7048), .ZN(n7047) );
  INV_X1 U8111 ( .A(n12225), .ZN(n7048) );
  INV_X1 U8112 ( .A(n15601), .ZN(n7049) );
  INV_X1 U8113 ( .A(n7051), .ZN(n7050) );
  NOR2_X1 U8114 ( .A1(n12332), .A2(n7223), .ZN(n7222) );
  INV_X1 U8115 ( .A(n7228), .ZN(n7223) );
  NAND2_X1 U8116 ( .A1(n8852), .A2(n7225), .ZN(n7224) );
  NAND2_X1 U8117 ( .A1(n10998), .A2(n8850), .ZN(n11044) );
  AND2_X1 U8118 ( .A1(n10797), .A2(n10783), .ZN(n7631) );
  AND4_X1 U8119 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n15611)
         );
  AND3_X1 U8120 ( .A1(n8518), .A2(n8517), .A3(n8516), .ZN(n15617) );
  AND2_X1 U8121 ( .A1(n8847), .A2(n8846), .ZN(n7209) );
  INV_X1 U8122 ( .A(n8847), .ZN(n15628) );
  NAND3_X1 U8123 ( .A1(n9880), .A2(n12320), .A3(n9868), .ZN(n15637) );
  OR2_X1 U8124 ( .A1(n9509), .A2(n9429), .ZN(n10794) );
  INV_X1 U8125 ( .A(n15637), .ZN(n15653) );
  NAND2_X1 U8126 ( .A1(n8895), .A2(n12320), .ZN(n15673) );
  NAND2_X1 U8127 ( .A1(n10792), .A2(n10791), .ZN(n10795) );
  NAND2_X1 U8128 ( .A1(n8751), .A2(n8750), .ZN(n12933) );
  NAND2_X1 U8129 ( .A1(n8930), .A2(n8929), .ZN(n8968) );
  OR2_X1 U8130 ( .A1(n8805), .A2(n8398), .ZN(n8400) );
  NOR2_X1 U8131 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7135) );
  AND2_X1 U8132 ( .A1(n7537), .A2(n8908), .ZN(n7058) );
  INV_X1 U8133 ( .A(n7539), .ZN(n7537) );
  XNOR2_X1 U8134 ( .A(n8903), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8924) );
  INV_X1 U8135 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8908) );
  AND3_X1 U8136 ( .A1(n6898), .A2(n6902), .A3(n6901), .ZN(n8414) );
  AND2_X1 U8137 ( .A1(n6893), .A2(n6899), .ZN(n8410) );
  AND2_X1 U8138 ( .A1(n8406), .A2(n8405), .ZN(n6893) );
  AND3_X1 U8139 ( .A1(n8616), .A2(n7135), .A3(n8512), .ZN(n7134) );
  NAND2_X1 U8140 ( .A1(n7032), .A2(n8394), .ZN(n8780) );
  NAND2_X1 U8141 ( .A1(n8393), .A2(n11630), .ZN(n7032) );
  XNOR2_X1 U8142 ( .A(n8901), .B(n8900), .ZN(n10160) );
  NAND2_X1 U8143 ( .A1(n8748), .A2(n8390), .ZN(n8758) );
  AND2_X1 U8144 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  INV_X1 U8145 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8833) );
  OR2_X1 U8146 ( .A1(n8386), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8387) );
  OAI21_X1 U8147 ( .B1(n8706), .B2(n7001), .A(n6998), .ZN(n8386) );
  AOI21_X1 U8148 ( .B1(n6998), .B2(n7001), .A(n6996), .ZN(n6995) );
  NAND2_X1 U8149 ( .A1(n8706), .A2(n6998), .ZN(n6997) );
  NAND2_X1 U8150 ( .A1(n7477), .A2(n8387), .ZN(n8736) );
  AND2_X1 U8151 ( .A1(n8388), .A2(n7478), .ZN(n7477) );
  AND2_X1 U8152 ( .A1(n8385), .A2(n8384), .ZN(n8718) );
  NAND2_X1 U8153 ( .A1(n7023), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8154 ( .A1(n8371), .A2(n10152), .ZN(n7024) );
  INV_X1 U8155 ( .A(n7021), .ZN(n7020) );
  INV_X1 U8156 ( .A(n8364), .ZN(n7474) );
  AND2_X1 U8157 ( .A1(n8366), .A2(n8365), .ZN(n8587) );
  NAND2_X1 U8158 ( .A1(n7005), .A2(n7008), .ZN(n8571) );
  NAND2_X1 U8159 ( .A1(n8358), .A2(n7479), .ZN(n7005) );
  NAND2_X1 U8160 ( .A1(n8571), .A2(n8570), .ZN(n8573) );
  OR2_X1 U8161 ( .A1(n8574), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8576) );
  AND2_X1 U8162 ( .A1(n8362), .A2(n8361), .ZN(n8557) );
  AOI21_X1 U8163 ( .B1(n7017), .B2(n7019), .A(n7015), .ZN(n7014) );
  INV_X1 U8164 ( .A(n8355), .ZN(n7015) );
  AND2_X1 U8165 ( .A1(n8355), .A2(n8354), .ZN(n8509) );
  AND2_X1 U8166 ( .A1(n8353), .A2(n8352), .ZN(n8495) );
  AND2_X1 U8167 ( .A1(n6900), .A2(n8461), .ZN(n8512) );
  NAND2_X1 U8168 ( .A1(n7466), .A2(n8348), .ZN(n8481) );
  NOR2_X1 U8169 ( .A1(n7361), .A2(n7364), .ZN(n7360) );
  AND2_X1 U8170 ( .A1(n13524), .A2(n13523), .ZN(n7364) );
  NAND2_X1 U8171 ( .A1(n10449), .A2(n6967), .ZN(n10487) );
  AND2_X1 U8172 ( .A1(n10448), .A2(n10447), .ZN(n6967) );
  OR2_X1 U8173 ( .A1(n9474), .A2(n9473), .ZN(n10449) );
  AOI21_X1 U8174 ( .B1(n7354), .B2(n7352), .A(n6794), .ZN(n7351) );
  INV_X1 U8175 ( .A(n13490), .ZN(n7352) );
  INV_X1 U8176 ( .A(n6985), .ZN(n6981) );
  INV_X1 U8177 ( .A(n7354), .ZN(n7353) );
  NAND2_X1 U8178 ( .A1(n13585), .A2(n13504), .ZN(n13508) );
  AND2_X1 U8179 ( .A1(n10507), .A2(n10501), .ZN(n7366) );
  NOR2_X1 U8180 ( .A1(n7365), .A2(n7362), .ZN(n7361) );
  INV_X1 U8181 ( .A(n13594), .ZN(n7362) );
  NAND2_X1 U8182 ( .A1(n13622), .A2(n7363), .ZN(n7358) );
  NOR2_X1 U8183 ( .A1(n7365), .A2(n13515), .ZN(n7363) );
  AND2_X1 U8184 ( .A1(n8169), .A2(n8168), .ZN(n13664) );
  NOR2_X1 U8185 ( .A1(n6681), .A2(n11724), .ZN(n7699) );
  NOR2_X1 U8186 ( .A1(n11724), .A2(n12682), .ZN(n7728) );
  NAND2_X1 U8187 ( .A1(n7699), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7694) );
  XNOR2_X1 U8188 ( .A(n13726), .B(n13735), .ZN(n15246) );
  XNOR2_X1 U8189 ( .A(n8291), .B(n6950), .ZN(n6949) );
  INV_X1 U8190 ( .A(n12641), .ZN(n6950) );
  OR2_X1 U8191 ( .A1(n13833), .A2(n6934), .ZN(n6930) );
  OR2_X1 U8192 ( .A1(n6936), .A2(n6718), .ZN(n6933) );
  OAI21_X1 U8193 ( .B1(n7589), .B2(n6938), .A(n13811), .ZN(n6937) );
  INV_X1 U8194 ( .A(n8221), .ZN(n8223) );
  NAND2_X1 U8195 ( .A1(n13833), .A2(n13846), .ZN(n7594) );
  NAND2_X1 U8196 ( .A1(n13859), .A2(n7506), .ZN(n13843) );
  INV_X1 U8197 ( .A(n7628), .ZN(n7511) );
  INV_X1 U8198 ( .A(n8285), .ZN(n7607) );
  AOI21_X1 U8199 ( .B1(n7597), .B2(n7599), .A(n6720), .ZN(n7595) );
  NAND2_X1 U8200 ( .A1(n13918), .A2(n7597), .ZN(n7596) );
  NAND2_X1 U8201 ( .A1(n8284), .A2(n8283), .ZN(n13884) );
  INV_X1 U8202 ( .A(n13882), .ZN(n8284) );
  NAND2_X1 U8203 ( .A1(n13918), .A2(n13917), .ZN(n13916) );
  AOI21_X1 U8204 ( .B1(n7499), .B2(n13956), .A(n6762), .ZN(n7498) );
  NAND2_X1 U8205 ( .A1(n11030), .A2(n6963), .ZN(n6962) );
  NAND2_X1 U8206 ( .A1(n11032), .A2(n7519), .ZN(n7517) );
  OR2_X1 U8207 ( .A1(n7896), .A2(n7895), .ZN(n7916) );
  NAND2_X1 U8208 ( .A1(n7894), .A2(n7893), .ZN(n12459) );
  NAND2_X1 U8209 ( .A1(n7727), .A2(n7726), .ZN(n12387) );
  OR2_X1 U8210 ( .A1(n7653), .A2(n12656), .ZN(n7657) );
  NAND2_X1 U8211 ( .A1(n12553), .A2(n12552), .ZN(n13765) );
  INV_X1 U8212 ( .A(n11790), .ZN(n6956) );
  OR2_X1 U8213 ( .A1(n15292), .A2(n9482), .ZN(n15403) );
  OAI21_X1 U8214 ( .B1(n8303), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8319) );
  INV_X1 U8215 ( .A(n8107), .ZN(n7396) );
  AND4_X1 U8216 ( .A1(n6777), .A2(n7761), .A3(n7909), .A4(n7639), .ZN(n7654)
         );
  INV_X1 U8217 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6989) );
  INV_X1 U8218 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7641) );
  AND2_X1 U8219 ( .A1(n7640), .A2(n6992), .ZN(n6991) );
  AND3_X1 U8220 ( .A1(n7909), .A2(n7639), .A3(n7761), .ZN(n7603) );
  INV_X1 U8221 ( .A(n7430), .ZN(n7428) );
  NAND2_X1 U8222 ( .A1(n7076), .A2(n7075), .ZN(n11489) );
  AOI21_X1 U8223 ( .B1(n6694), .B2(n7078), .A(n6767), .ZN(n7075) );
  AOI21_X1 U8224 ( .B1(n7419), .B2(n7423), .A(n7418), .ZN(n7417) );
  INV_X1 U8225 ( .A(n14210), .ZN(n7418) );
  AND2_X1 U8226 ( .A1(n12803), .A2(n12802), .ZN(n14208) );
  INV_X1 U8227 ( .A(n14231), .ZN(n7423) );
  AND2_X1 U8228 ( .A1(n14210), .A2(n12793), .ZN(n14229) );
  NAND2_X1 U8229 ( .A1(n10417), .A2(n6723), .ZN(n10576) );
  INV_X1 U8230 ( .A(n14310), .ZN(n11492) );
  INV_X1 U8231 ( .A(n12750), .ZN(n7416) );
  AOI21_X1 U8232 ( .B1(n14271), .B2(n12750), .A(n6763), .ZN(n7415) );
  NAND2_X1 U8233 ( .A1(n6764), .A2(n7068), .ZN(n7067) );
  INV_X1 U8234 ( .A(n6710), .ZN(n7068) );
  INV_X1 U8235 ( .A(n11568), .ZN(n7069) );
  AND2_X1 U8236 ( .A1(n7612), .A2(n12736), .ZN(n7412) );
  NAND2_X1 U8237 ( .A1(n7074), .A2(n14304), .ZN(n12722) );
  INV_X1 U8238 ( .A(n12120), .ZN(n12124) );
  NAND2_X1 U8239 ( .A1(n7257), .A2(n6739), .ZN(n7256) );
  NAND2_X1 U8240 ( .A1(n7259), .A2(n7258), .ZN(n7257) );
  AND2_X1 U8241 ( .A1(n11299), .A2(n11298), .ZN(n12713) );
  AND2_X1 U8242 ( .A1(n9518), .A2(n7302), .ZN(n9513) );
  AND2_X1 U8243 ( .A1(n14694), .A2(n14445), .ZN(n7130) );
  INV_X1 U8244 ( .A(n14532), .ZN(n14543) );
  INV_X1 U8245 ( .A(n7345), .ZN(n7341) );
  NOR2_X1 U8246 ( .A1(n7335), .A2(n14543), .ZN(n7334) );
  INV_X1 U8247 ( .A(n7337), .ZN(n7335) );
  XNOR2_X1 U8248 ( .A(n14700), .B(n7399), .ZN(n14532) );
  NAND2_X1 U8249 ( .A1(n7444), .A2(n7450), .ZN(n7439) );
  OR2_X1 U8250 ( .A1(n11793), .A2(n11817), .ZN(n11796) );
  NAND2_X1 U8251 ( .A1(n7346), .A2(n14443), .ZN(n7345) );
  INV_X1 U8252 ( .A(n6891), .ZN(n14574) );
  AND2_X1 U8253 ( .A1(n7452), .A2(n7451), .ZN(n7443) );
  AND2_X1 U8254 ( .A1(n14440), .A2(n14418), .ZN(n6826) );
  NAND2_X1 U8255 ( .A1(n14722), .A2(n14418), .ZN(n7451) );
  OR2_X1 U8256 ( .A1(n14596), .A2(n14595), .ZN(n7447) );
  AND2_X1 U8257 ( .A1(n14419), .A2(n11830), .ZN(n14584) );
  AOI21_X1 U8258 ( .B1(n7323), .B2(n7328), .A(n6752), .ZN(n7321) );
  XNOR2_X1 U8259 ( .A(n14728), .B(n14417), .ZN(n14617) );
  OR2_X1 U8260 ( .A1(n14652), .A2(n14435), .ZN(n14415) );
  NAND2_X1 U8261 ( .A1(n7453), .A2(n7456), .ZN(n11595) );
  INV_X1 U8262 ( .A(n7457), .ZN(n7456) );
  OAI21_X1 U8263 ( .B1(n12006), .B2(n7458), .A(n11876), .ZN(n7457) );
  OR2_X1 U8264 ( .A1(n14929), .A2(n12713), .ZN(n12008) );
  INV_X1 U8265 ( .A(n11876), .ZN(n11459) );
  NAND2_X1 U8266 ( .A1(n11383), .A2(n11382), .ZN(n11387) );
  NAND2_X1 U8267 ( .A1(n11387), .A2(n12006), .ZN(n11463) );
  NAND2_X1 U8268 ( .A1(n11009), .A2(n7464), .ZN(n11359) );
  INV_X1 U8269 ( .A(n14630), .ZN(n15055) );
  AND2_X1 U8270 ( .A1(n11855), .A2(n11854), .ZN(n14961) );
  OR2_X1 U8271 ( .A1(n10476), .A2(n9774), .ZN(n15126) );
  INV_X1 U8272 ( .A(n15126), .ZN(n15116) );
  NAND2_X1 U8273 ( .A1(n10248), .A2(n10247), .ZN(n15066) );
  NAND2_X1 U8274 ( .A1(n14756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9779) );
  XNOR2_X1 U8275 ( .A(n11734), .B(n11723), .ZN(n12577) );
  XNOR2_X1 U8276 ( .A(n11718), .B(n11717), .ZN(n12681) );
  INV_X1 U8277 ( .A(n9447), .ZN(n7173) );
  AND2_X1 U8278 ( .A1(n7401), .A2(n7175), .ZN(n7174) );
  INV_X1 U8279 ( .A(n9446), .ZN(n7175) );
  AND2_X1 U8280 ( .A1(n8083), .A2(n7624), .ZN(n8084) );
  NAND2_X1 U8281 ( .A1(n9432), .A2(n9513), .ZN(n9503) );
  NAND2_X1 U8282 ( .A1(n7400), .A2(n9433), .ZN(n9529) );
  INV_X1 U8283 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9433) );
  INV_X1 U8284 ( .A(n9503), .ZN(n7400) );
  NAND2_X1 U8285 ( .A1(n14782), .A2(n14781), .ZN(n7099) );
  AOI21_X1 U8286 ( .B1(n9012), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9011), .ZN(
        n9071) );
  AND2_X1 U8287 ( .A1(n9067), .A2(n9068), .ZN(n9011) );
  NAND2_X1 U8288 ( .A1(n8817), .A2(n8816), .ZN(n13148) );
  NAND2_X1 U8289 ( .A1(n12852), .A2(n12988), .ZN(n12891) );
  AND3_X1 U8290 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(n11541) );
  NAND2_X1 U8291 ( .A1(n13008), .A2(n12865), .ZN(n12911) );
  NAND2_X1 U8292 ( .A1(n10529), .A2(n6728), .ZN(n10703) );
  NAND2_X1 U8293 ( .A1(n7166), .A2(n7165), .ZN(n12981) );
  AOI21_X1 U8294 ( .B1(n6693), .B2(n13011), .A(n6757), .ZN(n7165) );
  AND4_X1 U8295 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(n11658)
         );
  NAND2_X1 U8296 ( .A1(n8710), .A2(n8709), .ZN(n13278) );
  AND2_X1 U8297 ( .A1(n10771), .A2(n8894), .ZN(n12928) );
  INV_X1 U8298 ( .A(n12849), .ZN(n12893) );
  NAND4_X1 U8299 ( .A1(n8569), .A2(n8568), .A3(n8567), .A4(n8566), .ZN(n15598)
         );
  INV_X1 U8300 ( .A(n11228), .ZN(n15597) );
  NAND3_X1 U8301 ( .A1(n7524), .A2(n8467), .A3(n7523), .ZN(n15655) );
  NAND2_X1 U8302 ( .A1(n8454), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7523) );
  AND2_X1 U8303 ( .A1(n8466), .A2(n8468), .ZN(n7524) );
  NOR2_X1 U8304 ( .A1(n15522), .A2(n15523), .ZN(n15521) );
  NOR2_X1 U8305 ( .A1(n15540), .A2(n15539), .ZN(n15538) );
  NOR2_X1 U8306 ( .A1(n15576), .A2(n15575), .ZN(n15574) );
  AND2_X1 U8307 ( .A1(n9882), .A2(n9881), .ZN(n14879) );
  INV_X1 U8308 ( .A(n15488), .ZN(n15586) );
  NAND2_X1 U8309 ( .A1(n13090), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7288) );
  NAND2_X1 U8310 ( .A1(n13146), .A2(n6846), .ZN(n13327) );
  INV_X1 U8311 ( .A(n6847), .ZN(n6846) );
  OAI21_X1 U8312 ( .B1(n13147), .B2(n15662), .A(n13145), .ZN(n6847) );
  NAND2_X1 U8313 ( .A1(n8771), .A2(n8770), .ZN(n13209) );
  NAND2_X1 U8314 ( .A1(n8733), .A2(n12276), .ZN(n13242) );
  AND3_X1 U8315 ( .A1(n8546), .A2(n8545), .A3(n8544), .ZN(n11051) );
  MUX2_X1 U8316 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8416), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8417) );
  XNOR2_X1 U8317 ( .A(n8830), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12359) );
  XNOR2_X1 U8318 ( .A(n8724), .B(n8828), .ZN(n13089) );
  NAND2_X1 U8319 ( .A1(n8127), .A2(n8126), .ZN(n14045) );
  NAND2_X1 U8320 ( .A1(n6955), .A2(n12576), .ZN(n8127) );
  INV_X1 U8321 ( .A(n11793), .ZN(n6955) );
  OR2_X1 U8322 ( .A1(n7705), .A2(n13711), .ZN(n7191) );
  AND2_X1 U8323 ( .A1(n11201), .A2(n11195), .ZN(n7357) );
  AND2_X1 U8324 ( .A1(n6971), .A2(n11343), .ZN(n6970) );
  OR2_X1 U8325 ( .A1(n11203), .A2(n6692), .ZN(n6971) );
  NAND2_X1 U8326 ( .A1(n7913), .A2(n7912), .ZN(n14912) );
  NAND2_X1 U8327 ( .A1(n7994), .A2(n7993), .ZN(n14084) );
  NAND2_X1 U8328 ( .A1(n13618), .A2(n13480), .ZN(n6984) );
  NAND2_X1 U8329 ( .A1(n8011), .A2(n8010), .ZN(n14079) );
  NAND2_X1 U8330 ( .A1(n8063), .A2(n8062), .ZN(n14063) );
  OR2_X1 U8331 ( .A1(n9484), .A2(n9483), .ZN(n13646) );
  NAND2_X1 U8332 ( .A1(n7358), .A2(n7359), .ZN(n6994) );
  INV_X1 U8333 ( .A(n7361), .ZN(n7359) );
  AOI21_X1 U8334 ( .B1(n13622), .B2(n13520), .A(n13594), .ZN(n13595) );
  NAND2_X1 U8335 ( .A1(n11669), .A2(n11668), .ZN(n13478) );
  INV_X1 U8336 ( .A(n13653), .ZN(n13676) );
  OR2_X1 U8337 ( .A1(n13787), .A2(n8238), .ZN(n8229) );
  INV_X1 U8338 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7685) );
  AND2_X1 U8339 ( .A1(n9745), .A2(n12668), .ZN(n15274) );
  NAND2_X1 U8340 ( .A1(n13957), .A2(n8036), .ZN(n13931) );
  NAND2_X1 U8341 ( .A1(n15343), .A2(n9480), .ZN(n15298) );
  NAND2_X1 U8342 ( .A1(n8110), .A2(n8109), .ZN(n14118) );
  NAND2_X1 U8343 ( .A1(n6954), .A2(n12576), .ZN(n8110) );
  INV_X1 U8344 ( .A(n11714), .ZN(n6954) );
  INV_X1 U8345 ( .A(n12660), .ZN(n13759) );
  XNOR2_X1 U8346 ( .A(n7060), .B(n14155), .ZN(n7059) );
  NOR2_X1 U8347 ( .A1(n10089), .A2(n10088), .ZN(n10207) );
  AND2_X1 U8348 ( .A1(n10087), .A2(n12824), .ZN(n10088) );
  NAND2_X1 U8349 ( .A1(n10922), .A2(n10921), .ZN(n15115) );
  NAND2_X1 U8350 ( .A1(n7408), .A2(n7409), .ZN(n14923) );
  AND2_X1 U8351 ( .A1(n14247), .A2(n6779), .ZN(n7409) );
  NAND2_X1 U8352 ( .A1(n10951), .A2(n10950), .ZN(n14986) );
  NAND2_X1 U8353 ( .A1(n11842), .A2(n11841), .ZN(n14638) );
  INV_X1 U8354 ( .A(n14277), .ZN(n14951) );
  AND2_X1 U8355 ( .A1(n10119), .A2(n10118), .ZN(n14563) );
  XNOR2_X1 U8356 ( .A(n10339), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14361) );
  NAND2_X1 U8357 ( .A1(n10389), .A2(n7625), .ZN(n9772) );
  OAI21_X1 U8358 ( .B1(n14484), .B2(n14447), .A(n7436), .ZN(n14468) );
  OR2_X1 U8359 ( .A1(n10091), .A2(n11817), .ZN(n10097) );
  OR2_X1 U8360 ( .A1(n11893), .A2(n10093), .ZN(n10096) );
  NAND2_X1 U8361 ( .A1(n6836), .A2(n14670), .ZN(n14741) );
  AOI21_X1 U8362 ( .B1(n14669), .B2(n14792), .A(n6857), .ZN(n14670) );
  NAND2_X1 U8363 ( .A1(n6859), .A2(n6858), .ZN(n6857) );
  XNOR2_X1 U8364 ( .A(n9060), .B(n7564), .ZN(n14785) );
  INV_X1 U8365 ( .A(n9061), .ZN(n7564) );
  INV_X1 U8366 ( .A(n9065), .ZN(n6868) );
  NAND2_X1 U8367 ( .A1(n7091), .A2(n7089), .ZN(n15012) );
  NAND2_X1 U8368 ( .A1(n7095), .A2(n7090), .ZN(n7089) );
  NOR2_X1 U8369 ( .A1(n9073), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U8370 ( .A1(n15017), .A2(n7106), .ZN(n7104) );
  NOR2_X1 U8371 ( .A1(n6707), .A2(n7107), .ZN(n7106) );
  INV_X1 U8372 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7107) );
  AND2_X1 U8373 ( .A1(n9087), .A2(n6707), .ZN(n7108) );
  INV_X1 U8374 ( .A(n12385), .ZN(n6828) );
  NAND2_X1 U8375 ( .A1(n7248), .A2(n7243), .ZN(n7242) );
  NAND2_X1 U8376 ( .A1(n7245), .A2(n7244), .ZN(n7243) );
  NAND2_X1 U8377 ( .A1(n11934), .A2(n14317), .ZN(n7244) );
  NAND2_X1 U8378 ( .A1(n12017), .A2(n7247), .ZN(n7246) );
  AND2_X1 U8379 ( .A1(n7180), .A2(n14317), .ZN(n7247) );
  OAI21_X1 U8380 ( .B1(n7574), .B2(n7571), .A(n6759), .ZN(n12416) );
  NAND2_X1 U8381 ( .A1(n6748), .A2(n7575), .ZN(n6880) );
  NAND2_X1 U8382 ( .A1(n11975), .A2(n11974), .ZN(n11978) );
  OAI21_X1 U8383 ( .B1(n12463), .B2(n12462), .A(n6761), .ZN(n7576) );
  NAND2_X1 U8384 ( .A1(n7251), .A2(n7250), .ZN(n11990) );
  NAND2_X1 U8385 ( .A1(n11985), .A2(n11987), .ZN(n7250) );
  OAI21_X1 U8386 ( .B1(n12472), .B2(n12655), .A(n12471), .ZN(n12473) );
  NAND2_X1 U8387 ( .A1(n11999), .A2(n12000), .ZN(n7278) );
  INV_X1 U8388 ( .A(n12497), .ZN(n7547) );
  INV_X1 U8389 ( .A(n12498), .ZN(n7546) );
  INV_X1 U8390 ( .A(n12494), .ZN(n7549) );
  NAND2_X1 U8391 ( .A1(n7277), .A2(n7274), .ZN(n12025) );
  NAND2_X1 U8392 ( .A1(n12048), .A2(n12049), .ZN(n7249) );
  OR2_X1 U8393 ( .A1(n6831), .A2(n12485), .ZN(n7541) );
  AND2_X1 U8394 ( .A1(n12508), .A2(n12507), .ZN(n6849) );
  INV_X1 U8395 ( .A(n12523), .ZN(n7567) );
  INV_X1 U8396 ( .A(n12522), .ZN(n7566) );
  NAND2_X1 U8397 ( .A1(n7272), .A2(n7271), .ZN(n12070) );
  OR2_X1 U8398 ( .A1(n12067), .A2(n7273), .ZN(n7271) );
  OAI21_X1 U8399 ( .B1(n12314), .B2(n12313), .A(n12312), .ZN(n12315) );
  NAND2_X1 U8400 ( .A1(n12347), .A2(n7010), .ZN(n12304) );
  AOI21_X1 U8401 ( .B1(n12303), .B2(n7011), .A(n13141), .ZN(n7010) );
  NAND2_X1 U8402 ( .A1(n8883), .A2(n13158), .ZN(n8884) );
  INV_X1 U8403 ( .A(n12246), .ZN(n7043) );
  INV_X1 U8404 ( .A(n8768), .ZN(n7496) );
  NOR2_X1 U8405 ( .A1(n7588), .A2(n12622), .ZN(n7584) );
  INV_X1 U8406 ( .A(n8262), .ZN(n7587) );
  XNOR2_X1 U8407 ( .A(n14773), .B(n14390), .ZN(n12091) );
  NOR2_X1 U8408 ( .A1(n7262), .A2(n6696), .ZN(n7261) );
  AOI22_X1 U8409 ( .A1(n7262), .A2(n7265), .B1(n6696), .B2(n7269), .ZN(n7260)
         );
  OR2_X1 U8410 ( .A1(n14318), .A2(n11129), .ZN(n11929) );
  INV_X1 U8411 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7062) );
  NOR2_X1 U8412 ( .A1(n8050), .A2(SI_18_), .ZN(n8055) );
  NAND2_X1 U8413 ( .A1(n7393), .A2(n7392), .ZN(n8056) );
  NAND2_X1 U8414 ( .A1(n6801), .A2(n6703), .ZN(n7392) );
  NAND2_X1 U8415 ( .A1(n7866), .A2(SI_10_), .ZN(n7890) );
  INV_X1 U8416 ( .A(n11226), .ZN(n7164) );
  OR2_X1 U8417 ( .A1(n10652), .A2(n15753), .ZN(n6865) );
  INV_X1 U8418 ( .A(n10629), .ZN(n7294) );
  INV_X1 U8419 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13033) );
  NAND2_X1 U8420 ( .A1(n14835), .A2(n6863), .ZN(n13104) );
  OR2_X1 U8421 ( .A1(n13103), .A2(n13379), .ZN(n6863) );
  OR2_X1 U8422 ( .A1(n8820), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13117) );
  AND2_X1 U8423 ( .A1(n8884), .A2(n8882), .ZN(n7217) );
  OR2_X1 U8424 ( .A1(n7218), .A2(n7216), .ZN(n7215) );
  INV_X1 U8425 ( .A(n8884), .ZN(n7216) );
  INV_X1 U8426 ( .A(n12922), .ZN(n7212) );
  AND2_X1 U8427 ( .A1(n13141), .A2(n6721), .ZN(n7218) );
  NAND2_X1 U8428 ( .A1(n8435), .A2(n12943), .ZN(n8807) );
  INV_X1 U8429 ( .A(n8795), .ZN(n8435) );
  OR2_X1 U8430 ( .A1(n8761), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8772) );
  INV_X1 U8431 ( .A(n7235), .ZN(n7230) );
  OR2_X1 U8432 ( .A1(n8581), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8596) );
  AND2_X1 U8433 ( .A1(n8502), .A2(n8423), .ZN(n8520) );
  XNOR2_X1 U8434 ( .A(n12199), .B(n15617), .ZN(n15607) );
  NAND2_X1 U8435 ( .A1(n9868), .A2(n6730), .ZN(n7055) );
  NAND2_X1 U8436 ( .A1(n15608), .A2(n8849), .ZN(n10996) );
  NOR2_X1 U8437 ( .A1(n12326), .A2(n7207), .ZN(n7206) );
  INV_X1 U8438 ( .A(n8849), .ZN(n7207) );
  INV_X1 U8439 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7540) );
  INV_X1 U8440 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U8441 ( .A1(n7492), .A2(n6704), .ZN(n8394) );
  AOI21_X1 U8442 ( .B1(n8718), .B2(n7000), .A(n6999), .ZN(n6998) );
  INV_X1 U8443 ( .A(n8385), .ZN(n6999) );
  INV_X1 U8444 ( .A(n8383), .ZN(n7000) );
  INV_X1 U8445 ( .A(n8718), .ZN(n7001) );
  AND2_X1 U8446 ( .A1(n7134), .A2(n8410), .ZN(n8693) );
  INV_X1 U8447 ( .A(n7018), .ZN(n7017) );
  OAI21_X1 U8448 ( .B1(n8495), .B2(n7019), .A(n8509), .ZN(n7018) );
  INV_X1 U8449 ( .A(n8353), .ZN(n7019) );
  AND2_X1 U8450 ( .A1(n6986), .A2(n13484), .ZN(n6985) );
  NAND2_X1 U8451 ( .A1(n13614), .A2(n6987), .ZN(n6986) );
  OR2_X1 U8452 ( .A1(n13667), .A2(n13522), .ZN(n7365) );
  AOI21_X1 U8453 ( .B1(n12637), .B2(n7592), .A(n7591), .ZN(n7590) );
  INV_X1 U8454 ( .A(n8288), .ZN(n7592) );
  INV_X1 U8455 ( .A(n12636), .ZN(n7591) );
  NOR2_X1 U8456 ( .A1(n7593), .A2(n12638), .ZN(n7589) );
  INV_X1 U8457 ( .A(n12637), .ZN(n7593) );
  NOR2_X1 U8458 ( .A1(n7198), .A2(n14107), .ZN(n7197) );
  INV_X1 U8459 ( .A(n7199), .ZN(n7198) );
  NOR2_X1 U8460 ( .A1(n14111), .A2(n14034), .ZN(n7199) );
  INV_X1 U8461 ( .A(n8281), .ZN(n7599) );
  NOR2_X1 U8462 ( .A1(n8049), .A2(n7500), .ZN(n7499) );
  INV_X1 U8463 ( .A(n8036), .ZN(n7500) );
  NAND2_X1 U8464 ( .A1(n7995), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8014) );
  INV_X1 U8465 ( .A(n7956), .ZN(n7954) );
  NOR2_X1 U8466 ( .A1(n8266), .A2(n7579), .ZN(n6961) );
  INV_X1 U8467 ( .A(n7518), .ZN(n7516) );
  NAND2_X1 U8468 ( .A1(n11030), .A2(n12625), .ZN(n11029) );
  AND2_X1 U8469 ( .A1(n12621), .A2(n12620), .ZN(n7484) );
  INV_X1 U8470 ( .A(n7817), .ZN(n7487) );
  INV_X1 U8471 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7854) );
  OR2_X1 U8472 ( .A1(n7855), .A2(n7854), .ZN(n7878) );
  INV_X1 U8473 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7829) );
  OR2_X1 U8474 ( .A1(n7830), .A2(n7829), .ZN(n7855) );
  NOR2_X1 U8475 ( .A1(n6749), .A2(n7601), .ZN(n7600) );
  INV_X1 U8476 ( .A(n8259), .ZN(n7601) );
  NAND2_X1 U8477 ( .A1(n6943), .A2(n6944), .ZN(n10750) );
  INV_X1 U8478 ( .A(n12621), .ZN(n6944) );
  NOR2_X1 U8479 ( .A1(n10395), .A2(n12424), .ZN(n10758) );
  NOR2_X1 U8480 ( .A1(n7649), .A2(n6843), .ZN(n6842) );
  OR2_X1 U8481 ( .A1(n7643), .A2(n6845), .ZN(n6844) );
  NOR2_X1 U8482 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6843) );
  AND2_X1 U8483 ( .A1(n7641), .A2(n7642), .ZN(n7370) );
  INV_X1 U8484 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6992) );
  OR2_X1 U8485 ( .A1(n7805), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7823) );
  INV_X1 U8486 ( .A(n11315), .ZN(n7432) );
  NAND2_X1 U8487 ( .A1(n14445), .A2(n7074), .ZN(n12794) );
  NAND2_X1 U8488 ( .A1(n14303), .A2(n7074), .ZN(n12785) );
  NAND2_X1 U8489 ( .A1(n7074), .A2(n14314), .ZN(n10584) );
  NAND2_X1 U8490 ( .A1(n14424), .A2(n7074), .ZN(n12805) );
  INV_X1 U8491 ( .A(n12110), .ZN(n12115) );
  NOR2_X1 U8492 ( .A1(n14674), .A2(n14492), .ZN(n14452) );
  NOR2_X1 U8493 ( .A1(n14638), .A2(n14652), .ZN(n7190) );
  INV_X1 U8494 ( .A(n12008), .ZN(n7458) );
  NOR2_X1 U8495 ( .A1(n7458), .A2(n7455), .ZN(n7454) );
  INV_X1 U8496 ( .A(n11382), .ZN(n7455) );
  NOR2_X1 U8497 ( .A1(n11984), .A2(n14986), .ZN(n7186) );
  NAND2_X1 U8498 ( .A1(n7179), .A2(n7178), .ZN(n14510) );
  AOI21_X1 U8499 ( .B1(n7317), .B2(n7319), .A(n6743), .ZN(n7315) );
  NOR2_X1 U8500 ( .A1(n11893), .A2(n9515), .ZN(n6839) );
  AOI21_X1 U8501 ( .B1(n8218), .B2(n8217), .A(n7615), .ZN(n8235) );
  NOR2_X1 U8502 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9574) );
  OR2_X1 U8503 ( .A1(n8056), .A2(n10082), .ZN(n8037) );
  AOI21_X1 U8504 ( .B1(n6690), .B2(n7119), .A(n7397), .ZN(n7115) );
  AND2_X1 U8505 ( .A1(n9607), .A2(n7946), .ZN(n7945) );
  NAND2_X1 U8506 ( .A1(n7786), .A2(n7785), .ZN(n7803) );
  INV_X1 U8507 ( .A(n7758), .ZN(n7377) );
  INV_X1 U8508 ( .A(n7740), .ZN(n7378) );
  NAND2_X1 U8509 ( .A1(n8992), .A2(n7569), .ZN(n8993) );
  NAND2_X1 U8510 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7570), .ZN(n7569) );
  INV_X1 U8511 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U8512 ( .A1(n9004), .A2(n9003), .ZN(n9022) );
  AOI21_X1 U8513 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9704), .A(n9006), .ZN(
        n9007) );
  AOI21_X1 U8514 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15028), .A(n9083), .ZN(
        n9088) );
  OR2_X1 U8515 ( .A1(n12880), .A2(n12879), .ZN(n7141) );
  NOR2_X1 U8516 ( .A1(n7164), .A2(n11223), .ZN(n7162) );
  OR2_X1 U8517 ( .A1(n11224), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U8518 ( .A1(n8426), .A2(n11693), .ZN(n8639) );
  INV_X1 U8519 ( .A(n8623), .ZN(n8426) );
  NAND2_X1 U8520 ( .A1(n11649), .A2(n6731), .ZN(n11689) );
  INV_X1 U8521 ( .A(n11651), .ZN(n7170) );
  NAND2_X1 U8522 ( .A1(n10184), .A2(n10180), .ZN(n10301) );
  NAND2_X1 U8523 ( .A1(n12881), .A2(n13157), .ZN(n7151) );
  NAND2_X1 U8524 ( .A1(n7141), .A2(n7140), .ZN(n7152) );
  NAND2_X1 U8525 ( .A1(n8428), .A2(n13033), .ZN(n8680) );
  INV_X1 U8526 ( .A(n8666), .ZN(n8428) );
  NAND2_X1 U8527 ( .A1(n7529), .A2(n7528), .ZN(n7527) );
  NAND2_X1 U8528 ( .A1(n12161), .A2(n12160), .ZN(n7528) );
  OR2_X1 U8529 ( .A1(n12354), .A2(n12353), .ZN(n12355) );
  OR2_X1 U8530 ( .A1(n12324), .A2(n12322), .ZN(n7469) );
  OR2_X1 U8531 ( .A1(n10013), .A2(n10012), .ZN(n10015) );
  INV_X1 U8532 ( .A(n7297), .ZN(n10617) );
  NAND2_X1 U8533 ( .A1(n10639), .A2(n6864), .ZN(n10640) );
  OR2_X1 U8534 ( .A1(n10654), .A2(n15757), .ZN(n6864) );
  CLKBUF_X1 U8535 ( .A(n15504), .Z(n6874) );
  XNOR2_X1 U8536 ( .A(n13097), .B(n13069), .ZN(n15561) );
  NAND2_X1 U8537 ( .A1(n15561), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15560) );
  NOR2_X1 U8538 ( .A1(n13103), .A2(n13053), .ZN(n6888) );
  XNOR2_X1 U8539 ( .A(n13104), .B(n13054), .ZN(n14856) );
  AND2_X1 U8540 ( .A1(n6911), .A2(n6907), .ZN(n12159) );
  NOR2_X1 U8541 ( .A1(n6914), .A2(n6908), .ZN(n6907) );
  AND2_X1 U8542 ( .A1(n6915), .A2(n12307), .ZN(n6914) );
  OR2_X1 U8543 ( .A1(n12301), .A2(n12300), .ZN(n13155) );
  INV_X1 U8544 ( .A(n8880), .ZN(n13173) );
  NAND2_X1 U8545 ( .A1(n13207), .A2(n12291), .ZN(n13182) );
  NAND2_X1 U8546 ( .A1(n7208), .A2(n8876), .ZN(n13196) );
  AND2_X1 U8547 ( .A1(n12285), .A2(n12286), .ZN(n13214) );
  NAND2_X1 U8548 ( .A1(n7036), .A2(n12281), .ZN(n13219) );
  NAND2_X1 U8549 ( .A1(n13227), .A2(n13231), .ZN(n13226) );
  OR2_X1 U8550 ( .A1(n8739), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8752) );
  NOR2_X1 U8551 ( .A1(n6925), .A2(n6924), .ZN(n6923) );
  INV_X1 U8552 ( .A(n12264), .ZN(n6924) );
  INV_X1 U8553 ( .A(n12275), .ZN(n6925) );
  OR2_X1 U8554 ( .A1(n8711), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8728) );
  AND3_X1 U8555 ( .A1(n8732), .A2(n8731), .A3(n8730), .ZN(n13274) );
  AND2_X1 U8556 ( .A1(n12264), .A2(n12268), .ZN(n13276) );
  OR2_X1 U8557 ( .A1(n8680), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U8558 ( .A1(n8429), .A2(n9234), .ZN(n8711) );
  INV_X1 U8559 ( .A(n8697), .ZN(n8429) );
  INV_X1 U8560 ( .A(n8868), .ZN(n13291) );
  NAND2_X1 U8561 ( .A1(n6919), .A2(n6917), .ZN(n13305) );
  AOI21_X1 U8562 ( .B1(n6920), .B2(n6922), .A(n6918), .ZN(n6917) );
  INV_X1 U8563 ( .A(n7534), .ZN(n6922) );
  NAND2_X1 U8564 ( .A1(n8427), .A2(n12991), .ZN(n8654) );
  INV_X1 U8565 ( .A(n8639), .ZN(n8427) );
  OR2_X1 U8566 ( .A1(n8654), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U8567 ( .A1(n8859), .A2(n8858), .ZN(n11621) );
  NAND2_X1 U8568 ( .A1(n6905), .A2(n6903), .ZN(n11558) );
  AOI21_X1 U8569 ( .B1(n6698), .B2(n7050), .A(n6904), .ZN(n6903) );
  INV_X1 U8570 ( .A(n12229), .ZN(n6904) );
  AND2_X1 U8571 ( .A1(n12232), .A2(n12236), .ZN(n12335) );
  AOI21_X1 U8572 ( .B1(n7222), .B2(n7226), .A(n6699), .ZN(n7220) );
  INV_X1 U8573 ( .A(n7222), .ZN(n7221) );
  NAND2_X1 U8574 ( .A1(n8425), .A2(n8424), .ZN(n8581) );
  INV_X1 U8575 ( .A(n8564), .ZN(n8425) );
  NAND2_X1 U8576 ( .A1(n8520), .A2(n9327), .ZN(n8548) );
  OR2_X1 U8577 ( .A1(n8548), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8564) );
  AND3_X1 U8578 ( .A1(n8500), .A2(n8499), .A3(n8498), .ZN(n10525) );
  NAND2_X1 U8579 ( .A1(n15634), .A2(n12184), .ZN(n15629) );
  INV_X1 U8580 ( .A(n10366), .ZN(n15630) );
  NAND2_X1 U8581 ( .A1(n15640), .A2(n15635), .ZN(n15634) );
  AND2_X1 U8582 ( .A1(n8842), .A2(n8933), .ZN(n15662) );
  CLKBUF_X1 U8583 ( .A(n10181), .Z(n15658) );
  AND4_X2 U8584 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n15674)
         );
  NAND2_X1 U8585 ( .A1(n12146), .A2(n12145), .ZN(n12156) );
  NOR2_X1 U8586 ( .A1(n8401), .A2(n7514), .ZN(n7513) );
  INV_X1 U8587 ( .A(n8399), .ZN(n7514) );
  OR2_X1 U8588 ( .A1(n8835), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8899) );
  AND2_X1 U8589 ( .A1(n8381), .A2(n8380), .ZN(n8686) );
  AND2_X1 U8590 ( .A1(n8379), .A2(n8378), .ZN(n8672) );
  NAND2_X1 U8591 ( .A1(n7021), .A2(n7024), .ZN(n8646) );
  OR2_X1 U8592 ( .A1(n8649), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8662) );
  AND2_X1 U8593 ( .A1(n8370), .A2(n8369), .ZN(n8612) );
  NAND2_X1 U8594 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  AOI21_X1 U8595 ( .B1(n7006), .B2(n7007), .A(n7004), .ZN(n7003) );
  AOI21_X1 U8596 ( .B1(n7008), .B2(n7480), .A(n7473), .ZN(n7006) );
  NOR2_X1 U8597 ( .A1(n8618), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8555) );
  INV_X1 U8598 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8554) );
  OR2_X1 U8599 ( .A1(n8514), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8618) );
  INV_X1 U8600 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8511) );
  AND2_X1 U8601 ( .A1(n8350), .A2(n8349), .ZN(n8480) );
  NAND2_X1 U8602 ( .A1(n7467), .A2(n8346), .ZN(n8470) );
  AND2_X1 U8603 ( .A1(n8348), .A2(n8347), .ZN(n8469) );
  XNOR2_X1 U8604 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8464) );
  NAND2_X1 U8605 ( .A1(n8344), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8463) );
  INV_X1 U8606 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7810) );
  OR2_X1 U8607 ( .A1(n7811), .A2(n7810), .ZN(n7830) );
  NAND2_X1 U8608 ( .A1(n8012), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8028) );
  INV_X1 U8609 ( .A(n8014), .ZN(n8012) );
  NAND2_X1 U8610 ( .A1(n6982), .A2(n6985), .ZN(n13655) );
  NAND2_X1 U8611 ( .A1(n6983), .A2(n13614), .ZN(n6982) );
  AND2_X1 U8612 ( .A1(n12600), .A2(n12572), .ZN(n12573) );
  INV_X1 U8613 ( .A(n8203), .ZN(n8238) );
  NAND3_X1 U8614 ( .A1(n7608), .A2(n7673), .A3(n7610), .ZN(n13704) );
  NAND2_X1 U8615 ( .A1(n7699), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7610) );
  AND2_X1 U8616 ( .A1(n7672), .A2(n7609), .ZN(n7608) );
  AND3_X1 U8617 ( .A1(n13706), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n13708) );
  AOI21_X1 U8618 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n13710), .A(n13708), .ZN(
        n15159) );
  AOI21_X1 U8619 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n9853), .A(n15168), .ZN(
        n10040) );
  NOR2_X1 U8620 ( .A1(n10038), .A2(n6860), .ZN(n15185) );
  AND2_X1 U8621 ( .A1(n9854), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6860) );
  AOI21_X1 U8622 ( .B1(n9922), .B2(P2_REG2_REG_6__SCAN_IN), .A(n9918), .ZN(
        n15205) );
  AOI21_X1 U8623 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10380), .A(n10379), .ZN(
        n10382) );
  NAND2_X1 U8624 ( .A1(n13724), .A2(n13725), .ZN(n13726) );
  NAND2_X1 U8625 ( .A1(n15259), .A2(n6820), .ZN(n15275) );
  OR2_X1 U8626 ( .A1(n15264), .A2(n13728), .ZN(n6820) );
  NAND2_X1 U8627 ( .A1(n15275), .A2(n15276), .ZN(n15273) );
  NOR2_X1 U8628 ( .A1(n13730), .A2(n13750), .ZN(n13748) );
  NAND2_X1 U8629 ( .A1(n13855), .A2(n7195), .ZN(n13795) );
  NOR2_X1 U8630 ( .A1(n13797), .A2(n7196), .ZN(n7195) );
  INV_X1 U8631 ( .A(n7197), .ZN(n7196) );
  INV_X1 U8632 ( .A(n7504), .ZN(n7503) );
  NAND2_X1 U8633 ( .A1(n7502), .A2(n7504), .ZN(n7501) );
  NAND2_X1 U8634 ( .A1(n13855), .A2(n7199), .ZN(n13825) );
  NAND2_X1 U8635 ( .A1(n13855), .A2(n13842), .ZN(n13837) );
  AOI21_X1 U8636 ( .B1(n7606), .B2(n13881), .A(n6729), .ZN(n7605) );
  NAND2_X1 U8637 ( .A1(n13882), .A2(n7606), .ZN(n6928) );
  NAND2_X1 U8638 ( .A1(n8089), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8111) );
  OR2_X1 U8639 ( .A1(n8028), .A2(n8027), .ZN(n8043) );
  NAND2_X1 U8640 ( .A1(n7201), .A2(n7200), .ZN(n13932) );
  AND2_X1 U8641 ( .A1(n7622), .A2(n8272), .ZN(n6951) );
  OR2_X1 U8642 ( .A1(n13955), .A2(n13956), .ZN(n13957) );
  NAND2_X1 U8643 ( .A1(n7203), .A2(n7202), .ZN(n13994) );
  INV_X1 U8644 ( .A(n7203), .ZN(n11640) );
  NAND2_X1 U8645 ( .A1(n6959), .A2(n6957), .ZN(n11405) );
  AOI21_X1 U8646 ( .B1(n6961), .B2(n6964), .A(n6958), .ZN(n6957) );
  OR2_X1 U8647 ( .A1(n11030), .A2(n6960), .ZN(n6959) );
  INV_X1 U8648 ( .A(n11236), .ZN(n6958) );
  NAND2_X1 U8649 ( .A1(n7914), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7934) );
  INV_X1 U8650 ( .A(n7205), .ZN(n11241) );
  NAND2_X1 U8651 ( .A1(n11029), .A2(n8265), .ZN(n11153) );
  NOR2_X2 U8652 ( .A1(n10839), .A2(n15393), .ZN(n11036) );
  NAND2_X1 U8653 ( .A1(n10561), .A2(n8262), .ZN(n10835) );
  NAND2_X1 U8654 ( .A1(n10835), .A2(n12624), .ZN(n10834) );
  NAND2_X1 U8655 ( .A1(n10758), .A2(n15385), .ZN(n10757) );
  INV_X1 U8656 ( .A(n6943), .ZN(n10752) );
  NAND2_X1 U8657 ( .A1(n10325), .A2(n12618), .ZN(n7602) );
  NOR2_X2 U8658 ( .A1(n10852), .A2(n15377), .ZN(n10855) );
  XNOR2_X1 U8659 ( .A(n13704), .B(n12363), .ZN(n12612) );
  NAND2_X1 U8660 ( .A1(n12579), .A2(n12578), .ZN(n13764) );
  NAND2_X1 U8661 ( .A1(n8026), .A2(n8025), .ZN(n13961) );
  INV_X1 U8662 ( .A(n15403), .ZN(n15392) );
  NAND2_X1 U8663 ( .A1(n8333), .A2(n15339), .ZN(n10556) );
  NAND2_X1 U8664 ( .A1(n7909), .A2(n7910), .ZN(n6993) );
  NAND2_X1 U8665 ( .A1(n7639), .A2(n7640), .ZN(n6990) );
  NAND2_X1 U8666 ( .A1(n13713), .A2(n7681), .ZN(n7707) );
  INV_X1 U8667 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8344) );
  OR2_X1 U8668 ( .A1(n10718), .A2(n7078), .ZN(n7077) );
  INV_X1 U8669 ( .A(n11058), .ZN(n7078) );
  OR2_X1 U8670 ( .A1(n11282), .A2(n11281), .ZN(n11294) );
  AND2_X1 U8671 ( .A1(n14231), .A2(n12783), .ZN(n14165) );
  AND2_X1 U8672 ( .A1(n7073), .A2(n7072), .ZN(n10419) );
  NAND2_X1 U8673 ( .A1(n12817), .A2(n14316), .ZN(n7072) );
  NAND2_X1 U8674 ( .A1(n7074), .A2(n11941), .ZN(n7073) );
  NAND2_X1 U8675 ( .A1(n12784), .A2(n14165), .ZN(n14232) );
  INV_X1 U8676 ( .A(n11798), .ZN(n11784) );
  INV_X1 U8677 ( .A(n12804), .ZN(n12823) );
  INV_X1 U8678 ( .A(n14270), .ZN(n12745) );
  NAND2_X1 U8679 ( .A1(n7411), .A2(n12702), .ZN(n14198) );
  INV_X1 U8680 ( .A(n14200), .ZN(n7411) );
  INV_X1 U8681 ( .A(n14307), .ZN(n12697) );
  AND2_X1 U8682 ( .A1(n14164), .A2(n12773), .ZN(n14256) );
  OR2_X1 U8683 ( .A1(n10939), .A2(n10938), .ZN(n10953) );
  NAND2_X1 U8684 ( .A1(n7074), .A2(n14308), .ZN(n12684) );
  AND2_X1 U8685 ( .A1(n11388), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11468) );
  AND4_X1 U8686 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n14461) );
  INV_X1 U8687 ( .A(n11902), .ZN(n11807) );
  INV_X1 U8688 ( .A(n11900), .ZN(n11889) );
  NAND2_X1 U8689 ( .A1(n9623), .A2(n9622), .ZN(n14326) );
  AOI21_X1 U8690 ( .B1(n10713), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9672), .ZN(
        n9648) );
  OR2_X1 U8691 ( .A1(n9596), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9597) );
  INV_X1 U8692 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U8693 ( .A1(n7436), .A2(n14447), .ZN(n7435) );
  NAND2_X1 U8694 ( .A1(n14484), .A2(n7436), .ZN(n6840) );
  NAND2_X1 U8695 ( .A1(n14495), .A2(n12830), .ZN(n7122) );
  INV_X1 U8696 ( .A(n7437), .ZN(n7436) );
  OAI21_X1 U8697 ( .B1(n14485), .B2(n14447), .A(n14472), .ZN(n7437) );
  AND2_X1 U8698 ( .A1(n14449), .A2(n11770), .ZN(n14472) );
  OR2_X1 U8699 ( .A1(n14674), .A2(n14461), .ZN(n11770) );
  NOR2_X1 U8700 ( .A1(n14510), .A2(n14688), .ZN(n14513) );
  NAND2_X1 U8701 ( .A1(n14513), .A2(n14495), .ZN(n14492) );
  INV_X1 U8702 ( .A(n14423), .ZN(n14507) );
  NAND2_X1 U8703 ( .A1(n7334), .A2(n7339), .ZN(n7132) );
  NOR2_X1 U8704 ( .A1(n11822), .A2(n14261), .ZN(n11809) );
  NAND2_X1 U8705 ( .A1(n7439), .A2(n14548), .ZN(n7438) );
  OR2_X1 U8706 ( .A1(n11818), .A2(n11817), .ZN(n11821) );
  AND2_X1 U8707 ( .A1(n11881), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U8708 ( .A1(n11883), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11822) );
  NAND2_X1 U8709 ( .A1(n14585), .A2(n14584), .ZN(n14583) );
  NAND2_X1 U8710 ( .A1(n14651), .A2(n7187), .ZN(n14600) );
  AND2_X1 U8711 ( .A1(n14722), .A2(n7188), .ZN(n7187) );
  INV_X1 U8712 ( .A(n7323), .ZN(n7322) );
  NAND2_X1 U8713 ( .A1(n14651), .A2(n7190), .ZN(n14631) );
  NAND2_X1 U8714 ( .A1(n14651), .A2(n14961), .ZN(n14650) );
  NAND2_X1 U8715 ( .A1(n11350), .A2(n7182), .ZN(n11394) );
  NOR2_X1 U8716 ( .A1(n14245), .A2(n7184), .ZN(n7182) );
  NOR2_X1 U8717 ( .A1(n10953), .A2(n10952), .ZN(n10978) );
  NAND2_X1 U8718 ( .A1(n14795), .A2(n14794), .ZN(n14793) );
  AOI21_X1 U8719 ( .B1(n7311), .B2(n7313), .A(n6742), .ZN(n7309) );
  NAND2_X1 U8720 ( .A1(n11350), .A2(n7186), .ZN(n14802) );
  NAND2_X1 U8721 ( .A1(n11350), .A2(n15127), .ZN(n11352) );
  OR2_X1 U8722 ( .A1(n10924), .A2(n10923), .ZN(n10939) );
  AND2_X1 U8723 ( .A1(n11485), .A2(n11258), .ZN(n11350) );
  NOR2_X1 U8724 ( .A1(n15107), .A2(n11259), .ZN(n11258) );
  NAND2_X1 U8725 ( .A1(n7177), .A2(n7176), .ZN(n11259) );
  INV_X1 U8726 ( .A(n15054), .ZN(n7177) );
  NAND2_X1 U8727 ( .A1(n15056), .A2(n15092), .ZN(n15054) );
  NAND2_X1 U8728 ( .A1(n10964), .A2(n10963), .ZN(n11144) );
  NAND2_X1 U8729 ( .A1(n7307), .A2(n11947), .ZN(n7306) );
  NAND2_X1 U8730 ( .A1(n7181), .A2(n7180), .ZN(n10270) );
  INV_X1 U8731 ( .A(n10237), .ZN(n7181) );
  INV_X1 U8732 ( .A(n7348), .ZN(n11856) );
  OR2_X1 U8733 ( .A1(n11915), .A2(n10118), .ZN(n14401) );
  OR2_X1 U8734 ( .A1(n10471), .A2(n10470), .ZN(n14459) );
  INV_X1 U8735 ( .A(n14668), .ZN(n6859) );
  INV_X1 U8736 ( .A(n15056), .ZN(n11139) );
  INV_X1 U8737 ( .A(n11129), .ZN(n10244) );
  AND2_X1 U8738 ( .A1(n9449), .A2(n9583), .ZN(n9567) );
  NAND2_X1 U8739 ( .A1(n9437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9438) );
  INV_X1 U8740 ( .A(n8144), .ZN(n8142) );
  AND2_X1 U8741 ( .A1(n7286), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U8742 ( .A1(n8075), .A2(n8061), .ZN(n8078) );
  XNOR2_X1 U8743 ( .A(n8078), .B(n8082), .ZN(n11878) );
  XNOR2_X1 U8744 ( .A(n8038), .B(n8050), .ZN(n11840) );
  NAND2_X1 U8745 ( .A1(n7395), .A2(n8004), .ZN(n8022) );
  NAND2_X1 U8746 ( .A1(n8003), .A2(n7626), .ZN(n7395) );
  AND2_X1 U8747 ( .A1(n10389), .A2(n9439), .ZN(n10405) );
  NAND2_X1 U8748 ( .A1(n10389), .A2(n7286), .ZN(n10551) );
  AND2_X1 U8749 ( .A1(n10338), .A2(n10151), .ZN(n11278) );
  NAND2_X1 U8750 ( .A1(n7116), .A2(n7905), .ZN(n7924) );
  NAND2_X1 U8751 ( .A1(n7386), .A2(n6711), .ZN(n7116) );
  NAND2_X1 U8752 ( .A1(n7386), .A2(n7388), .ZN(n7907) );
  NAND2_X1 U8753 ( .A1(n7865), .A2(n7864), .ZN(n7889) );
  AND2_X1 U8754 ( .A1(n7125), .A2(n7126), .ZN(n7839) );
  NAND2_X1 U8755 ( .A1(n7741), .A2(n7740), .ZN(n7757) );
  NAND2_X1 U8756 ( .A1(n7382), .A2(n7381), .ZN(n7721) );
  INV_X1 U8757 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7687) );
  INV_X1 U8758 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9231) );
  XNOR2_X1 U8759 ( .A(n8993), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n9035) );
  NOR2_X1 U8760 ( .A1(n9044), .A2(n9045), .ZN(n9046) );
  INV_X1 U8761 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U8762 ( .A1(n9000), .A2(n8999), .ZN(n9049) );
  OAI21_X1 U8763 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n9830), .A(n9010), .ZN(
        n9068) );
  NOR2_X1 U8764 ( .A1(n9073), .A2(n15009), .ZN(n7090) );
  NAND2_X1 U8765 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  NAND2_X1 U8766 ( .A1(n11112), .A2(n11222), .ZN(n11225) );
  NAND2_X1 U8767 ( .A1(n7147), .A2(n7148), .ZN(n12920) );
  NAND2_X1 U8768 ( .A1(n7152), .A2(n6709), .ZN(n7147) );
  NAND2_X1 U8769 ( .A1(n12891), .A2(n12890), .ZN(n12889) );
  NAND2_X1 U8770 ( .A1(n11535), .A2(n11534), .ZN(n11537) );
  NAND2_X1 U8771 ( .A1(n6823), .A2(n6822), .ZN(n10529) );
  INV_X1 U8772 ( .A(n10367), .ZN(n6822) );
  INV_X1 U8773 ( .A(n10368), .ZN(n6823) );
  NAND2_X1 U8774 ( .A1(n13008), .A2(n6693), .ZN(n12912) );
  INV_X1 U8775 ( .A(n7138), .ZN(n7137) );
  OAI21_X1 U8776 ( .B1(n7144), .B2(n7139), .A(n7142), .ZN(n7138) );
  NAND2_X1 U8777 ( .A1(n8422), .A2(n8421), .ZN(n12930) );
  NAND2_X1 U8778 ( .A1(n11225), .A2(n11224), .ZN(n11227) );
  NAND2_X1 U8779 ( .A1(n11227), .A2(n11226), .ZN(n11430) );
  NAND2_X1 U8780 ( .A1(n6678), .A2(n6725), .ZN(n7240) );
  OAI21_X1 U8781 ( .B1(n6701), .B2(n7238), .A(n9868), .ZN(n7237) );
  INV_X1 U8782 ( .A(n13229), .ZN(n13199) );
  AND2_X1 U8783 ( .A1(n8813), .A2(n8812), .ZN(n13169) );
  INV_X1 U8784 ( .A(n7141), .ZN(n12941) );
  INV_X1 U8785 ( .A(n13042), .ZN(n13302) );
  NAND2_X1 U8786 ( .A1(n7153), .A2(n7156), .ZN(n12952) );
  AND2_X1 U8787 ( .A1(n7157), .A2(n12857), .ZN(n7156) );
  AND4_X1 U8788 ( .A1(n8685), .A2(n8684), .A3(n8683), .A4(n8682), .ZN(n13315)
         );
  NAND2_X1 U8789 ( .A1(n8782), .A2(n8781), .ZN(n12976) );
  AND2_X1 U8790 ( .A1(n10529), .A2(n10528), .ZN(n10530) );
  AND3_X1 U8791 ( .A1(n8756), .A2(n8755), .A3(n8754), .ZN(n13238) );
  AND2_X1 U8792 ( .A1(n8778), .A2(n8777), .ZN(n13217) );
  NAND2_X1 U8793 ( .A1(n8760), .A2(n8759), .ZN(n13220) );
  AND4_X1 U8794 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n11696)
         );
  NAND2_X1 U8795 ( .A1(n12959), .A2(n12863), .ZN(n13010) );
  AOI21_X1 U8796 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(n10825) );
  NAND2_X1 U8797 ( .A1(n10189), .A2(n10195), .ZN(n13027) );
  AND2_X1 U8798 ( .A1(n10193), .A2(n10192), .ZN(n15429) );
  NAND2_X1 U8799 ( .A1(n7152), .A2(n7151), .ZN(n13018) );
  NAND2_X1 U8800 ( .A1(n7033), .A2(n8806), .ZN(n13025) );
  NAND2_X1 U8801 ( .A1(n13032), .A2(n13031), .ZN(n13030) );
  NAND2_X1 U8802 ( .A1(n12889), .A2(n12854), .ZN(n13032) );
  NAND2_X1 U8803 ( .A1(n10170), .A2(n10169), .ZN(n13037) );
  INV_X1 U8804 ( .A(n12362), .ZN(n7046) );
  INV_X1 U8805 ( .A(n13169), .ZN(n13143) );
  AND2_X1 U8806 ( .A1(n8789), .A2(n8788), .ZN(n13200) );
  INV_X1 U8807 ( .A(n13238), .ZN(n13002) );
  INV_X1 U8808 ( .A(n13301), .ZN(n12954) );
  INV_X1 U8809 ( .A(n11696), .ZN(n11688) );
  INV_X1 U8810 ( .A(n11658), .ZN(n11647) );
  INV_X1 U8811 ( .A(n15611), .ZN(n11109) );
  INV_X1 U8812 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15450) );
  INV_X1 U8813 ( .A(n7299), .ZN(n15438) );
  INV_X1 U8814 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15499) );
  INV_X1 U8815 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15520) );
  NOR2_X1 U8816 ( .A1(n6874), .A2(n10627), .ZN(n10630) );
  NOR2_X1 U8817 ( .A1(n10630), .A2(n10629), .ZN(n13046) );
  NOR2_X1 U8818 ( .A1(n15521), .A2(n13049), .ZN(n15540) );
  OR2_X1 U8819 ( .A1(n15551), .A2(n15550), .ZN(n15552) );
  AND2_X1 U8820 ( .A1(n15567), .A2(n13071), .ZN(n15591) );
  INV_X1 U8821 ( .A(n7290), .ZN(n14815) );
  NOR2_X1 U8822 ( .A1(n7620), .A2(n8896), .ZN(n8897) );
  NAND2_X1 U8823 ( .A1(n8794), .A2(n8793), .ZN(n13335) );
  NAND2_X1 U8824 ( .A1(n7037), .A2(n12264), .ZN(n13262) );
  NAND2_X1 U8825 ( .A1(n7040), .A2(n12246), .ZN(n13317) );
  NAND2_X1 U8826 ( .A1(n7533), .A2(n7532), .ZN(n7040) );
  NAND2_X1 U8827 ( .A1(n7533), .A2(n11620), .ZN(n11684) );
  NAND2_X1 U8828 ( .A1(n7234), .A2(n7232), .ZN(n11680) );
  NAND2_X1 U8829 ( .A1(n8629), .A2(n12240), .ZN(n11627) );
  NAND2_X1 U8830 ( .A1(n6906), .A2(n7047), .ZN(n11442) );
  OR2_X1 U8831 ( .A1(n15602), .A2(n7050), .ZN(n6906) );
  NAND2_X1 U8832 ( .A1(n7224), .A2(n7222), .ZN(n11249) );
  NAND2_X1 U8833 ( .A1(n7053), .A2(n8563), .ZN(n11251) );
  NAND2_X1 U8834 ( .A1(n15602), .A2(n15601), .ZN(n7053) );
  NAND2_X1 U8835 ( .A1(n8852), .A2(n8851), .ZN(n15596) );
  NAND2_X1 U8836 ( .A1(n15638), .A2(n8846), .ZN(n15622) );
  NAND2_X1 U8837 ( .A1(n11453), .A2(n11003), .ZN(n15631) );
  NOR2_X1 U8838 ( .A1(n10795), .A2(n12323), .ZN(n15679) );
  NAND2_X1 U8839 ( .A1(n10795), .A2(n15676), .ZN(n15682) );
  AOI21_X1 U8840 ( .B1(n13456), .B2(n7160), .A(n12153), .ZN(n13393) );
  NOR2_X1 U8841 ( .A1(n13327), .A2(n6733), .ZN(n13401) );
  INV_X1 U8842 ( .A(n13148), .ZN(n8883) );
  OR2_X1 U8843 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  NAND2_X1 U8844 ( .A1(n8653), .A2(n8652), .ZN(n13448) );
  AND2_X1 U8845 ( .A1(n8926), .A2(n8925), .ZN(n10788) );
  INV_X1 U8846 ( .A(n8968), .ZN(n10172) );
  INV_X1 U8847 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8438) );
  INV_X1 U8848 ( .A(n8444), .ZN(n13461) );
  NAND2_X1 U8849 ( .A1(n8400), .A2(n8399), .ZN(n8815) );
  OAI21_X1 U8850 ( .B1(n7056), .B2(n7057), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8418) );
  NAND2_X1 U8851 ( .A1(n8512), .A2(n7135), .ZN(n7057) );
  AND2_X1 U8852 ( .A1(n8414), .A2(n8410), .ZN(n7133) );
  OAI21_X1 U8853 ( .B1(n8758), .B2(n8757), .A(n8391), .ZN(n8769) );
  NAND2_X1 U8854 ( .A1(n8736), .A2(n8388), .ZN(n8746) );
  NAND2_X1 U8855 ( .A1(n8387), .A2(n8388), .ZN(n8734) );
  NAND2_X1 U8856 ( .A1(n8719), .A2(n8718), .ZN(n8721) );
  NAND2_X1 U8857 ( .A1(n8706), .A2(n8383), .ZN(n8719) );
  INV_X1 U8858 ( .A(SI_19_), .ZN(n10156) );
  INV_X1 U8859 ( .A(SI_17_), .ZN(n9840) );
  INV_X1 U8860 ( .A(SI_16_), .ZN(n9711) );
  INV_X1 U8861 ( .A(SI_15_), .ZN(n9638) );
  NAND2_X1 U8862 ( .A1(n7020), .A2(n7024), .ZN(n8632) );
  NAND2_X1 U8863 ( .A1(n7022), .A2(n7024), .ZN(n8630) );
  INV_X1 U8864 ( .A(SI_12_), .ZN(n9541) );
  INV_X1 U8865 ( .A(SI_11_), .ZN(n9536) );
  OAI21_X1 U8866 ( .B1(n8571), .B2(n7474), .A(n7472), .ZN(n8590) );
  NAND2_X1 U8867 ( .A1(n8573), .A2(n8364), .ZN(n8588) );
  XNOR2_X1 U8868 ( .A(n8592), .B(n8591), .ZN(n13091) );
  OAI21_X1 U8869 ( .B1(n8358), .B2(n7481), .A(n7479), .ZN(n8560) );
  NAND2_X1 U8870 ( .A1(n8542), .A2(n8360), .ZN(n8558) );
  NAND2_X1 U8871 ( .A1(n8358), .A2(n8357), .ZN(n8540) );
  NAND2_X1 U8872 ( .A1(n7016), .A2(n8353), .ZN(n8510) );
  NAND2_X1 U8873 ( .A1(n8496), .A2(n8495), .ZN(n7016) );
  XNOR2_X1 U8874 ( .A(n8483), .B(n8482), .ZN(n10062) );
  NAND2_X1 U8875 ( .A1(n8462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U8876 ( .A1(n8459), .A2(n8619), .ZN(n7296) );
  AND2_X1 U8877 ( .A1(n7358), .A2(n7360), .ZN(n13529) );
  AND2_X1 U8878 ( .A1(n11590), .A2(n11582), .ZN(n6965) );
  NAND2_X1 U8879 ( .A1(n7953), .A2(n7952), .ZN(n12483) );
  NAND2_X1 U8880 ( .A1(n11196), .A2(n11195), .ZN(n11332) );
  INV_X1 U8881 ( .A(n13992), .ZN(n13605) );
  NAND2_X1 U8882 ( .A1(n13478), .A2(n13477), .ZN(n13603) );
  NAND2_X1 U8883 ( .A1(n10487), .A2(n10486), .ZN(n6966) );
  NAND2_X1 U8884 ( .A1(n6976), .A2(n6977), .ZN(n13640) );
  INV_X1 U8885 ( .A(n6978), .ZN(n6977) );
  OAI21_X1 U8886 ( .B1(n6979), .B2(n13614), .A(n7351), .ZN(n6978) );
  NAND2_X1 U8887 ( .A1(n13547), .A2(n13490), .ZN(n13637) );
  NAND2_X1 U8888 ( .A1(n11330), .A2(n11203), .ZN(n11341) );
  NOR2_X1 U8889 ( .A1(n13646), .A2(n13953), .ZN(n13659) );
  NAND2_X1 U8890 ( .A1(n7356), .A2(n7355), .ZN(n13547) );
  INV_X1 U8891 ( .A(n13654), .ZN(n7355) );
  INV_X1 U8892 ( .A(n13655), .ZN(n7356) );
  NAND2_X1 U8893 ( .A1(n10502), .A2(n10501), .ZN(n10612) );
  INV_X1 U8894 ( .A(n13674), .ZN(n13649) );
  NAND2_X1 U8895 ( .A1(n8210), .A2(n8209), .ZN(n13683) );
  NAND2_X1 U8896 ( .A1(n8203), .A2(n7747), .ZN(n7734) );
  CLKBUF_X1 U8897 ( .A(n13704), .Z(n6854) );
  NAND2_X1 U8898 ( .A1(n7728), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7697) );
  OR2_X1 U8899 ( .A1(n15185), .A2(n15184), .ZN(n15187) );
  XNOR2_X1 U8900 ( .A(n13722), .B(n13733), .ZN(n11078) );
  NAND2_X1 U8901 ( .A1(n11078), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13724) );
  NAND2_X1 U8902 ( .A1(n6948), .A2(n8302), .ZN(n13776) );
  NAND2_X1 U8903 ( .A1(n6949), .A2(n15293), .ZN(n6948) );
  OAI22_X1 U8904 ( .A1(n8300), .A2(n13953), .B1(n13768), .B2(n8299), .ZN(n8301) );
  NAND2_X1 U8905 ( .A1(n6930), .A2(n6933), .ZN(n13790) );
  NAND2_X1 U8906 ( .A1(n13843), .A2(n8170), .ZN(n13824) );
  NAND2_X1 U8907 ( .A1(n7594), .A2(n8288), .ZN(n13819) );
  NAND2_X1 U8908 ( .A1(n13859), .A2(n8157), .ZN(n13845) );
  NOR2_X1 U8909 ( .A1(n13887), .A2(n7628), .ZN(n13871) );
  NAND2_X1 U8910 ( .A1(n13890), .A2(n7510), .ZN(n13869) );
  NAND2_X1 U8911 ( .A1(n13884), .A2(n7606), .ZN(n13865) );
  AND2_X1 U8912 ( .A1(n13886), .A2(n13885), .ZN(n14050) );
  NAND2_X1 U8913 ( .A1(n13916), .A2(n8281), .ZN(n13899) );
  NAND3_X1 U8914 ( .A1(n13945), .A2(n6974), .A3(n13946), .ZN(n14068) );
  NAND2_X1 U8915 ( .A1(n6952), .A2(n8272), .ZN(n13969) );
  NAND2_X1 U8916 ( .A1(n6962), .A2(n7578), .ZN(n11237) );
  NAND2_X1 U8917 ( .A1(n7517), .A2(n7518), .ZN(n11239) );
  NAND2_X1 U8918 ( .A1(n7521), .A2(n7522), .ZN(n11157) );
  OR2_X1 U8919 ( .A1(n11032), .A2(n7902), .ZN(n7521) );
  NAND2_X1 U8920 ( .A1(n10566), .A2(n6972), .ZN(n10890) );
  NAND2_X1 U8921 ( .A1(n7488), .A2(n7817), .ZN(n10749) );
  INV_X1 U8922 ( .A(n15285), .ZN(n13907) );
  INV_X1 U8923 ( .A(n15298), .ZN(n15283) );
  INV_X1 U8924 ( .A(n13998), .ZN(n15281) );
  AND2_X1 U8925 ( .A1(n15303), .A2(n13759), .ZN(n15285) );
  INV_X2 U8926 ( .A(n15303), .ZN(n15305) );
  INV_X1 U8927 ( .A(n13765), .ZN(n14097) );
  INV_X1 U8928 ( .A(n13764), .ZN(n14101) );
  NAND2_X1 U8929 ( .A1(n6953), .A2(n12576), .ZN(n8088) );
  INV_X1 U8930 ( .A(n11818), .ZN(n6953) );
  OR2_X1 U8931 ( .A1(n10919), .A2(n7715), .ZN(n7852) );
  NOR2_X1 U8932 ( .A1(n15358), .A2(n14093), .ZN(n15365) );
  AND2_X1 U8933 ( .A1(n9475), .A2(n8320), .ZN(n15343) );
  CLKBUF_X1 U8934 ( .A(n15321), .Z(n15338) );
  NAND2_X1 U8935 ( .A1(n8313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7679) );
  INV_X1 U8936 ( .A(n7663), .ZN(n8307) );
  XNOR2_X1 U8937 ( .A(n8306), .B(n8305), .ZN(n11631) );
  INV_X1 U8938 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U8939 ( .A1(n8304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8306) );
  INV_X1 U8940 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11716) );
  NAND2_X1 U8941 ( .A1(n8119), .A2(n7127), .ZN(n8120) );
  INV_X1 U8942 ( .A(n7128), .ZN(n7127) );
  INV_X1 U8943 ( .A(n12646), .ZN(n12659) );
  NAND2_X1 U8944 ( .A1(n7654), .A2(n7641), .ZN(n7645) );
  INV_X1 U8945 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10411) );
  INV_X1 U8946 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10077) );
  INV_X1 U8947 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9739) );
  INV_X1 U8948 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9645) );
  INV_X1 U8949 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9601) );
  INV_X1 U8950 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9600) );
  INV_X1 U8951 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9559) );
  INV_X1 U8952 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9550) );
  INV_X1 U8953 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9546) );
  INV_X1 U8954 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9535) );
  INV_X1 U8955 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9502) );
  INV_X1 U8956 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U8957 ( .A1(n11059), .A2(n11058), .ZN(n11063) );
  NAND2_X1 U8958 ( .A1(n10104), .A2(n6695), .ZN(n7434) );
  NAND2_X1 U8959 ( .A1(n10116), .A2(n6695), .ZN(n7433) );
  NAND2_X1 U8960 ( .A1(n14176), .A2(n12750), .ZN(n14179) );
  OAI22_X1 U8961 ( .A1(n7428), .A2(n7427), .B1(n12829), .B2(n7430), .ZN(n7426)
         );
  NAND2_X1 U8962 ( .A1(n11316), .A2(n11315), .ZN(n11318) );
  NAND2_X1 U8963 ( .A1(n7083), .A2(n12758), .ZN(n14188) );
  INV_X1 U8964 ( .A(n7415), .ZN(n7084) );
  INV_X1 U8965 ( .A(n7417), .ZN(n7082) );
  AND2_X1 U8966 ( .A1(n7081), .A2(n14208), .ZN(n7080) );
  NAND2_X1 U8967 ( .A1(n7417), .A2(n7420), .ZN(n7081) );
  NAND2_X1 U8968 ( .A1(n11599), .A2(n11598), .ZN(n14940) );
  NAND2_X1 U8969 ( .A1(n14289), .A2(n12733), .ZN(n14938) );
  AOI21_X1 U8970 ( .B1(n10579), .B2(n10578), .A(n10577), .ZN(n10711) );
  AND2_X1 U8971 ( .A1(n10576), .A2(n10575), .ZN(n10577) );
  OAI21_X1 U8972 ( .B1(n12784), .B2(n7423), .A(n7419), .ZN(n14207) );
  OAI21_X1 U8973 ( .B1(n12745), .B2(n7416), .A(n7415), .ZN(n14238) );
  NAND2_X1 U8974 ( .A1(n14198), .A2(n12706), .ZN(n14246) );
  NAND2_X1 U8975 ( .A1(n6769), .A2(n7067), .ZN(n7065) );
  NOR2_X1 U8976 ( .A1(n7067), .A2(n6712), .ZN(n7066) );
  NOR2_X1 U8977 ( .A1(n10205), .A2(n10105), .ZN(n10117) );
  OR2_X1 U8978 ( .A1(n9801), .A2(n9800), .ZN(n14277) );
  NAND2_X1 U8979 ( .A1(n10292), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14958) );
  OAI21_X2 U8980 ( .B1(n10711), .B2(n10710), .A(n10709), .ZN(n10719) );
  NAND2_X1 U8981 ( .A1(n10719), .A2(n10718), .ZN(n11059) );
  NAND2_X1 U8982 ( .A1(n7256), .A2(n12123), .ZN(n7253) );
  INV_X1 U8983 ( .A(n12132), .ZN(n6818) );
  OR3_X1 U8984 ( .A1(n11730), .A2(n11729), .A3(n11728), .ZN(n14402) );
  OR2_X1 U8985 ( .A1(n11900), .A2(n9783), .ZN(n9789) );
  OR2_X1 U8986 ( .A1(n11902), .A2(n9797), .ZN(n9787) );
  AOI21_X1 U8987 ( .B1(n14344), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14345), .ZN(
        n9725) );
  AOI21_X1 U8988 ( .B1(n9695), .B2(n9693), .A(n9694), .ZN(n9697) );
  NOR2_X1 U8989 ( .A1(n9828), .A2(n9829), .ZN(n10140) );
  NOR2_X1 U8990 ( .A1(n15018), .A2(n6856), .ZN(n11175) );
  XNOR2_X1 U8991 ( .A(n6855), .B(n11837), .ZN(n14385) );
  NAND2_X1 U8992 ( .A1(n15029), .A2(n14375), .ZN(n6855) );
  AOI21_X1 U8993 ( .B1(n12577), .B2(n11892), .A(n6811), .ZN(n14663) );
  AOI21_X1 U8994 ( .B1(n12681), .B2(n11892), .A(n11743), .ZN(n14666) );
  AND2_X1 U8995 ( .A1(n7336), .A2(n7334), .ZN(n14541) );
  NAND2_X1 U8996 ( .A1(n7337), .A2(n7336), .ZN(n14542) );
  NAND2_X1 U8997 ( .A1(n14574), .A2(n7340), .ZN(n7336) );
  NAND2_X1 U8998 ( .A1(n7343), .A2(n7347), .ZN(n7342) );
  INV_X1 U8999 ( .A(n14574), .ZN(n7343) );
  NAND2_X1 U9000 ( .A1(n14596), .A2(n7443), .ZN(n7441) );
  NAND2_X1 U9001 ( .A1(n7447), .A2(n7451), .ZN(n14579) );
  NAND2_X1 U9002 ( .A1(n7325), .A2(n7326), .ZN(n14610) );
  NAND2_X1 U9003 ( .A1(n14649), .A2(n7327), .ZN(n7325) );
  AND2_X1 U9004 ( .A1(n7329), .A2(n14413), .ZN(n14628) );
  NAND2_X1 U9005 ( .A1(n14649), .A2(n14415), .ZN(n7329) );
  NAND2_X1 U9006 ( .A1(n11457), .A2(n11456), .ZN(n12721) );
  NAND2_X1 U9007 ( .A1(n11463), .A2(n12008), .ZN(n11464) );
  NOR2_X1 U9008 ( .A1(n12006), .A2(n7332), .ZN(n7331) );
  INV_X1 U9009 ( .A(n11400), .ZN(n7332) );
  NAND2_X1 U9010 ( .A1(n7333), .A2(n11400), .ZN(n11401) );
  NAND2_X1 U9011 ( .A1(n11386), .A2(n11385), .ZN(n14929) );
  NAND2_X1 U9012 ( .A1(n11349), .A2(n11866), .ZN(n7310) );
  NAND2_X1 U9013 ( .A1(n11359), .A2(n10976), .ZN(n10977) );
  NOR2_X1 U9014 ( .A1(n7463), .A2(n7462), .ZN(n11358) );
  INV_X1 U9015 ( .A(n10975), .ZN(n7462) );
  INV_X1 U9016 ( .A(n11009), .ZN(n7463) );
  NAND2_X1 U9017 ( .A1(n11094), .A2(n11099), .ZN(n7316) );
  INV_X1 U9018 ( .A(n15067), .ZN(n14656) );
  INV_X1 U9019 ( .A(n15058), .ZN(n14654) );
  NAND2_X1 U9020 ( .A1(n10461), .A2(n14161), .ZN(n14633) );
  INV_X1 U9021 ( .A(n6833), .ZN(n6832) );
  OAI21_X1 U9022 ( .B1(n14678), .B2(n14677), .A(n14675), .ZN(n6833) );
  XNOR2_X1 U9023 ( .A(n11737), .B(n11736), .ZN(n14759) );
  OAI22_X1 U9024 ( .A1(n11734), .A2(n11733), .B1(n11732), .B2(n13460), .ZN(
        n11737) );
  INV_X1 U9025 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9577) );
  INV_X1 U9026 ( .A(n14390), .ZN(n11166) );
  INV_X1 U9027 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10410) );
  INV_X1 U9028 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10391) );
  INV_X1 U9029 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10341) );
  INV_X1 U9030 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9825) );
  INV_X1 U9031 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9643) );
  INV_X1 U9032 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9605) );
  INV_X1 U9033 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9598) );
  INV_X1 U9034 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9562) );
  INV_X1 U9035 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9558) );
  INV_X1 U9036 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9533) );
  AND2_X1 U9037 ( .A1(n9505), .A2(n9529), .ZN(n14324) );
  CLKBUF_X1 U9038 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14775) );
  INV_X1 U9039 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7113) );
  XNOR2_X1 U9040 ( .A(n9031), .B(n7111), .ZN(n14780) );
  INV_X1 U9041 ( .A(n9032), .ZN(n7111) );
  INV_X1 U9042 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6866) );
  XNOR2_X1 U9043 ( .A(n9046), .B(n7563), .ZN(n14782) );
  INV_X1 U9044 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7563) );
  INV_X1 U9045 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U9046 ( .A1(n7114), .A2(n9062), .ZN(n14787) );
  NAND2_X1 U9047 ( .A1(n14785), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7114) );
  INV_X1 U9048 ( .A(n9095), .ZN(n7553) );
  NAND2_X1 U9049 ( .A1(n7045), .A2(n7044), .ZN(P3_U3296) );
  OR2_X1 U9050 ( .A1(n12361), .A2(n12360), .ZN(n7044) );
  NAND2_X1 U9051 ( .A1(n7034), .A2(n7046), .ZN(n7045) );
  AND2_X1 U9052 ( .A1(n14885), .A2(n14883), .ZN(n6890) );
  OAI21_X1 U9053 ( .B1(n14882), .B2(n6873), .A(n14879), .ZN(n6872) );
  AOI211_X1 U9054 ( .C1(n15588), .C2(n13111), .A(n13110), .B(n13109), .ZN(
        n13112) );
  OAI21_X1 U9055 ( .B1(n11330), .B2(n6692), .A(n6970), .ZN(n11508) );
  NAND2_X1 U9056 ( .A1(n6984), .A2(n13614), .ZN(n13621) );
  AOI21_X1 U9057 ( .B1(n6994), .B2(n13676), .A(n13675), .ZN(n13677) );
  MUX2_X1 U9058 ( .A(n13761), .B(n13760), .S(n13759), .Z(n13763) );
  NAND2_X1 U9059 ( .A1(n7059), .A2(n14951), .ZN(n14160) );
  INV_X1 U9060 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6834) );
  INV_X1 U9061 ( .A(n7096), .ZN(n15007) );
  INV_X1 U9062 ( .A(n7558), .ZN(n15011) );
  NAND2_X1 U9063 ( .A1(n7105), .A2(n6738), .ZN(n14814) );
  AND2_X1 U9064 ( .A1(n7117), .A2(n7946), .ZN(n6690) );
  AND3_X1 U9065 ( .A1(n12040), .A2(n14617), .A3(n12039), .ZN(n6691) );
  INV_X1 U9066 ( .A(n13842), .ZN(n14034) );
  INV_X1 U9067 ( .A(n7346), .ZN(n14711) );
  NAND2_X1 U9068 ( .A1(n14772), .A2(n10092), .ZN(n7346) );
  AND2_X1 U9069 ( .A1(n11338), .A2(n11337), .ZN(n6692) );
  AND2_X1 U9070 ( .A1(n7167), .A2(n12865), .ZN(n6693) );
  AND2_X1 U9071 ( .A1(n7077), .A2(n11062), .ZN(n6694) );
  NAND2_X1 U9072 ( .A1(n10288), .A2(n10287), .ZN(n6695) );
  AND2_X1 U9073 ( .A1(n12087), .A2(n7267), .ZN(n6696) );
  AND2_X1 U9074 ( .A1(n12307), .A2(n12299), .ZN(n6697) );
  INV_X1 U9075 ( .A(n12425), .ZN(n7575) );
  INV_X1 U9076 ( .A(n14067), .ZN(n6975) );
  AND2_X1 U9077 ( .A1(n7047), .A2(n12230), .ZN(n6698) );
  INV_X1 U9078 ( .A(n13881), .ZN(n8283) );
  NOR2_X1 U9079 ( .A1(n13888), .A2(n8283), .ZN(n13887) );
  AND2_X1 U9080 ( .A1(n15598), .A2(n11434), .ZN(n6699) );
  NAND2_X1 U9081 ( .A1(n11280), .A2(n11279), .ZN(n14245) );
  INV_X1 U9082 ( .A(n7480), .ZN(n7479) );
  INV_X1 U9083 ( .A(n12493), .ZN(n7550) );
  AND2_X1 U9084 ( .A1(n8263), .A2(n7884), .ZN(n12624) );
  INV_X1 U9085 ( .A(n12624), .ZN(n7588) );
  AND2_X1 U9086 ( .A1(n9584), .A2(n9581), .ZN(n6700) );
  INV_X1 U9087 ( .A(n7328), .ZN(n7327) );
  NAND2_X1 U9088 ( .A1(n7330), .A2(n14415), .ZN(n7328) );
  INV_X1 U9089 ( .A(n7905), .ZN(n7119) );
  NAND2_X1 U9090 ( .A1(n11273), .A2(n11272), .ZN(n14801) );
  INV_X1 U9091 ( .A(n14801), .ZN(n7185) );
  AND2_X1 U9092 ( .A1(n11804), .A2(SI_1_), .ZN(n6701) );
  NAND2_X1 U9093 ( .A1(n6765), .A2(n7249), .ZN(n6702) );
  INV_X1 U9094 ( .A(n10446), .ZN(n9715) );
  OR2_X1 U9095 ( .A1(n8021), .A2(n9840), .ZN(n6703) );
  AND2_X1 U9096 ( .A1(n8802), .A2(n8801), .ZN(n13157) );
  AND2_X1 U9097 ( .A1(n7493), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6704) );
  CLKBUF_X1 U9098 ( .A(n12368), .Z(n12580) );
  INV_X1 U9099 ( .A(n7729), .ZN(n7853) );
  NOR2_X1 U9100 ( .A1(n12249), .A2(n12248), .ZN(n6705) );
  OR2_X1 U9101 ( .A1(n13932), .A2(n14063), .ZN(n6706) );
  INV_X1 U9102 ( .A(n14303), .ZN(n7399) );
  NAND2_X1 U9103 ( .A1(n8904), .A2(n8415), .ZN(n8902) );
  XNOR2_X1 U9104 ( .A(n14861), .B(n9092), .ZN(n6707) );
  NAND2_X1 U9105 ( .A1(n12745), .A2(n12744), .ZN(n14176) );
  NAND2_X1 U9106 ( .A1(n8237), .A2(n8236), .ZN(n12559) );
  INV_X1 U9107 ( .A(n8360), .ZN(n7481) );
  AND2_X1 U9108 ( .A1(n14674), .A2(n14427), .ZN(n6708) );
  AND2_X1 U9109 ( .A1(n7150), .A2(n7151), .ZN(n6709) );
  NOR2_X1 U9110 ( .A1(n14548), .A2(n7341), .ZN(n7340) );
  NAND2_X1 U9111 ( .A1(n14948), .A2(n14946), .ZN(n6710) );
  INV_X1 U9112 ( .A(n7579), .ZN(n7578) );
  OAI21_X1 U9113 ( .B1(n7581), .B2(n13692), .A(n7580), .ZN(n7579) );
  INV_X1 U9114 ( .A(n6913), .ZN(n13137) );
  AOI21_X1 U9115 ( .B1(n13156), .B2(n12299), .A(n6915), .ZN(n6913) );
  AND2_X1 U9116 ( .A1(n7388), .A2(n7120), .ZN(n6711) );
  AND2_X1 U9117 ( .A1(n11575), .A2(n11494), .ZN(n6712) );
  AND2_X1 U9118 ( .A1(n11852), .A2(n10113), .ZN(n6713) );
  AND2_X1 U9119 ( .A1(n7927), .A2(n7943), .ZN(n6714) );
  NAND2_X1 U9120 ( .A1(n7928), .A2(n7927), .ZN(n6715) );
  INV_X1 U9121 ( .A(n13934), .ZN(n7200) );
  XNOR2_X1 U9122 ( .A(n8527), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U9123 ( .A1(n11895), .A2(n11894), .ZN(n14694) );
  INV_X1 U9124 ( .A(n14694), .ZN(n7178) );
  INV_X1 U9125 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9325) );
  AND2_X1 U9126 ( .A1(n14912), .A2(n13692), .ZN(n6716) );
  AND2_X1 U9127 ( .A1(n6678), .A2(n9886), .ZN(n6717) );
  INV_X1 U9128 ( .A(n14961), .ZN(n14652) );
  NAND2_X1 U9129 ( .A1(n14291), .A2(n14290), .ZN(n14289) );
  AND2_X1 U9130 ( .A1(n14107), .A2(n8289), .ZN(n6718) );
  INV_X1 U9131 ( .A(n15009), .ZN(n7094) );
  OR3_X1 U9132 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        n13472), .ZN(n6719) );
  AND2_X1 U9133 ( .A1(n14120), .A2(n13632), .ZN(n6720) );
  NAND2_X1 U9134 ( .A1(n13025), .A2(n13143), .ZN(n6721) );
  AND2_X1 U9135 ( .A1(n9575), .A2(n9574), .ZN(n6722) );
  OR2_X1 U9136 ( .A1(n10419), .A2(n10418), .ZN(n6723) );
  NAND2_X1 U9137 ( .A1(n10936), .A2(n10935), .ZN(n11984) );
  AND2_X1 U9138 ( .A1(n9568), .A2(n9567), .ZN(n6724) );
  INV_X1 U9139 ( .A(n11965), .ZN(n7282) );
  AND2_X1 U9140 ( .A1(n13469), .A2(n7241), .ZN(n6725) );
  NAND2_X1 U9141 ( .A1(n13855), .A2(n7197), .ZN(n6726) );
  AND2_X1 U9142 ( .A1(n14638), .A2(n14437), .ZN(n6727) );
  AND2_X1 U9143 ( .A1(n10528), .A2(n10531), .ZN(n6728) );
  NOR2_X1 U9144 ( .A1(n13870), .A2(n7607), .ZN(n7606) );
  AND2_X1 U9145 ( .A1(n12008), .A2(n12001), .ZN(n12006) );
  INV_X1 U9146 ( .A(n6964), .ZN(n6963) );
  NAND2_X1 U9147 ( .A1(n6745), .A2(n12625), .ZN(n6964) );
  AND2_X1 U9148 ( .A1(n14045), .A2(n13540), .ZN(n6729) );
  AND2_X1 U9149 ( .A1(n11804), .A2(n7383), .ZN(n6730) );
  AND2_X1 U9150 ( .A1(n11648), .A2(n7170), .ZN(n6731) );
  AND2_X1 U9151 ( .A1(n13328), .A2(n15739), .ZN(n6733) );
  AND3_X1 U9152 ( .A1(n7469), .A2(n12355), .A3(n12356), .ZN(n6734) );
  NOR2_X1 U9153 ( .A1(n8008), .A2(n7368), .ZN(n7649) );
  OR2_X1 U9154 ( .A1(n13101), .A2(n13052), .ZN(n6735) );
  OR2_X1 U9155 ( .A1(n11999), .A2(n12000), .ZN(n6736) );
  AND2_X1 U9156 ( .A1(n8877), .A2(n8876), .ZN(n6737) );
  INV_X1 U9157 ( .A(n7226), .ZN(n7225) );
  OR2_X1 U9158 ( .A1(n8853), .A2(n7227), .ZN(n7226) );
  AND2_X1 U9159 ( .A1(n7104), .A2(n7109), .ZN(n6738) );
  AND2_X1 U9160 ( .A1(n12210), .A2(n12205), .ZN(n12326) );
  AND2_X1 U9161 ( .A1(n12115), .A2(n12114), .ZN(n6739) );
  AND2_X1 U9162 ( .A1(n7435), .A2(n14449), .ZN(n6740) );
  NOR2_X1 U9163 ( .A1(n14450), .A2(n6708), .ZN(n6741) );
  INV_X1 U9164 ( .A(n7420), .ZN(n7419) );
  NAND2_X1 U9165 ( .A1(n14229), .A2(n7421), .ZN(n7420) );
  NOR2_X1 U9166 ( .A1(n14986), .A2(n14308), .ZN(n6742) );
  NOR2_X1 U9167 ( .A1(n15107), .A2(n14311), .ZN(n6743) );
  NOR2_X1 U9168 ( .A1(n12424), .A2(n8260), .ZN(n6744) );
  OR2_X1 U9169 ( .A1(n14912), .A2(n11151), .ZN(n6745) );
  NOR2_X1 U9170 ( .A1(n13448), .A2(n13314), .ZN(n6746) );
  XOR2_X1 U9171 ( .A(n7611), .B(n9428), .Z(n6747) );
  INV_X1 U9172 ( .A(n7340), .ZN(n7339) );
  AND2_X1 U9173 ( .A1(n12423), .A2(n12422), .ZN(n6748) );
  AND2_X1 U9174 ( .A1(n12424), .A2(n8260), .ZN(n6749) );
  OR2_X1 U9175 ( .A1(n12930), .A2(n13041), .ZN(n8965) );
  OR2_X1 U9176 ( .A1(n8189), .A2(n13808), .ZN(n6750) );
  AND4_X1 U9177 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n11946) );
  NOR2_X1 U9178 ( .A1(n12918), .A2(n12925), .ZN(n6751) );
  NOR2_X1 U9179 ( .A1(n14728), .A2(n14417), .ZN(n6752) );
  OR2_X1 U9180 ( .A1(n12048), .A2(n12049), .ZN(n6753) );
  INV_X1 U9181 ( .A(n14155), .ZN(n7431) );
  AND2_X1 U9182 ( .A1(n11507), .A2(n11506), .ZN(n6754) );
  NAND2_X1 U9183 ( .A1(n13730), .A2(n13750), .ZN(n6755) );
  NAND2_X1 U9184 ( .A1(n7133), .A2(n7134), .ZN(n6756) );
  AND2_X1 U9185 ( .A1(n12867), .A2(n12982), .ZN(n6757) );
  INV_X1 U9186 ( .A(n7184), .ZN(n7183) );
  NAND2_X1 U9187 ( .A1(n7186), .A2(n7185), .ZN(n7184) );
  AND2_X1 U9188 ( .A1(n12428), .A2(n13697), .ZN(n6758) );
  OR2_X1 U9189 ( .A1(n12407), .A2(n12408), .ZN(n6759) );
  OR2_X1 U9190 ( .A1(n14473), .A2(n14472), .ZN(n7121) );
  INV_X1 U9191 ( .A(n12337), .ZN(n11527) );
  INV_X1 U9192 ( .A(n7473), .ZN(n7472) );
  OAI21_X1 U9193 ( .B1(n8570), .B2(n7474), .A(n8587), .ZN(n7473) );
  AND2_X1 U9194 ( .A1(n13635), .A2(n13492), .ZN(n6760) );
  INV_X1 U9195 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9508) );
  INV_X1 U9196 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U9197 ( .A1(n12466), .A2(n12467), .ZN(n6761) );
  NOR2_X1 U9198 ( .A1(n7200), .A2(n13954), .ZN(n6762) );
  AND2_X1 U9199 ( .A1(n12754), .A2(n12753), .ZN(n6763) );
  OAI21_X1 U9200 ( .B1(n6714), .B2(n7398), .A(SI_14_), .ZN(n7397) );
  NAND2_X1 U9201 ( .A1(n7069), .A2(n11575), .ZN(n6764) );
  AND2_X1 U9202 ( .A1(n12160), .A2(n12155), .ZN(n12350) );
  INV_X1 U9203 ( .A(n12350), .ZN(n7529) );
  AND2_X1 U9204 ( .A1(n12046), .A2(n12047), .ZN(n6765) );
  OR2_X1 U9205 ( .A1(n7431), .A2(n7429), .ZN(n6766) );
  OR2_X1 U9206 ( .A1(n11319), .A2(n7432), .ZN(n6767) );
  NAND2_X1 U9207 ( .A1(n7545), .A2(n7548), .ZN(n6768) );
  OR2_X1 U9208 ( .A1(n6710), .A2(n11494), .ZN(n6769) );
  OR2_X1 U9209 ( .A1(n14414), .A2(n6727), .ZN(n6770) );
  AND2_X1 U9210 ( .A1(n14557), .A2(n14444), .ZN(n6771) );
  INV_X1 U9211 ( .A(n12629), .ZN(n11410) );
  NAND2_X2 U9212 ( .A1(n10114), .A2(n6838), .ZN(n11934) );
  AND2_X1 U9213 ( .A1(n7321), .A2(n14595), .ZN(n6772) );
  AND2_X1 U9214 ( .A1(n7538), .A2(n7536), .ZN(n6773) );
  NOR2_X1 U9215 ( .A1(n9435), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6774) );
  AND2_X1 U9216 ( .A1(n7360), .A2(n13528), .ZN(n6775) );
  INV_X1 U9217 ( .A(n7802), .ZN(n7385) );
  AND2_X1 U9218 ( .A1(n12012), .A2(n7278), .ZN(n6776) );
  AND3_X1 U9219 ( .A1(n7640), .A2(n6992), .A3(n6989), .ZN(n6777) );
  AND2_X1 U9220 ( .A1(n11880), .A2(n11879), .ZN(n14722) );
  INV_X1 U9221 ( .A(n14722), .ZN(n14440) );
  INV_X1 U9222 ( .A(n12706), .ZN(n7410) );
  AND2_X1 U9223 ( .A1(n13884), .A2(n8285), .ZN(n6778) );
  OR2_X1 U9224 ( .A1(n12702), .A2(n7410), .ZN(n6779) );
  INV_X1 U9225 ( .A(n7946), .ZN(n7398) );
  INV_X1 U9226 ( .A(n12084), .ZN(n7268) );
  AND2_X1 U9227 ( .A1(n7163), .A2(n11429), .ZN(n6780) );
  OR2_X1 U9228 ( .A1(n7552), .A2(n12550), .ZN(n6781) );
  NAND2_X1 U9229 ( .A1(n6997), .A2(n6995), .ZN(n8388) );
  OR2_X1 U9230 ( .A1(n7560), .A2(n12456), .ZN(n6782) );
  INV_X1 U9231 ( .A(n6980), .ZN(n6979) );
  NOR2_X1 U9232 ( .A1(n7353), .A2(n6981), .ZN(n6980) );
  AND2_X1 U9233 ( .A1(n7284), .A2(n6722), .ZN(n6783) );
  AND2_X1 U9234 ( .A1(n8790), .A2(n12291), .ZN(n6784) );
  AND2_X1 U9235 ( .A1(n14315), .A2(n10472), .ZN(n6785) );
  AND2_X1 U9236 ( .A1(n7543), .A2(n12503), .ZN(n6786) );
  NAND2_X1 U9237 ( .A1(n12456), .A2(n7560), .ZN(n6787) );
  NAND2_X1 U9238 ( .A1(n11986), .A2(n7252), .ZN(n6788) );
  AND2_X1 U9239 ( .A1(n12470), .A2(n13691), .ZN(n6789) );
  INV_X1 U9240 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9780) );
  OR2_X1 U9241 ( .A1(n6677), .A2(n14303), .ZN(n6790) );
  INV_X1 U9242 ( .A(n7145), .ZN(n7144) );
  AND2_X1 U9243 ( .A1(n7146), .A2(n7148), .ZN(n7145) );
  OR2_X1 U9244 ( .A1(n7575), .A2(n6748), .ZN(n6791) );
  NAND2_X1 U9245 ( .A1(n12067), .A2(n7273), .ZN(n6792) );
  INV_X1 U9246 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7285) );
  CLKBUF_X3 U9247 ( .A(n7730), .Z(n8030) );
  NAND2_X1 U9248 ( .A1(n7583), .A2(n7585), .ZN(n11030) );
  AND2_X1 U9249 ( .A1(n14651), .A2(n7188), .ZN(n6793) );
  NAND2_X1 U9250 ( .A1(n11567), .A2(n11566), .ZN(n7071) );
  INV_X1 U9251 ( .A(SI_2_), .ZN(n7383) );
  INV_X1 U9252 ( .A(n10654), .ZN(n15487) );
  NAND2_X1 U9253 ( .A1(n14938), .A2(n12736), .ZN(n14216) );
  XOR2_X1 U9254 ( .A(n13494), .B(n13495), .Z(n6794) );
  OR2_X1 U9255 ( .A1(n13400), .A2(n13390), .ZN(n6795) );
  NAND3_X1 U9256 ( .A1(n13478), .A2(n7350), .A3(n13477), .ZN(n13618) );
  INV_X1 U9257 ( .A(n13618), .ZN(n6983) );
  AND2_X1 U9258 ( .A1(n7985), .A2(n7970), .ZN(n6796) );
  NAND2_X1 U9259 ( .A1(n14923), .A2(n12717), .ZN(n14927) );
  OR2_X1 U9260 ( .A1(n6993), .A2(n6990), .ZN(n8006) );
  INV_X1 U9261 ( .A(n7201), .ZN(n13960) );
  INV_X1 U9262 ( .A(n12830), .ZN(n14426) );
  AND4_X1 U9263 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n12830) );
  OR2_X1 U9264 ( .A1(n8883), .A2(n13390), .ZN(n6797) );
  OR2_X1 U9265 ( .A1(n8883), .A2(n13449), .ZN(n6798) );
  INV_X1 U9266 ( .A(n7510), .ZN(n7509) );
  AND2_X1 U9267 ( .A1(n13870), .A2(n7511), .ZN(n7510) );
  INV_X1 U9268 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10152) );
  INV_X1 U9269 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10154) );
  INV_X1 U9270 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9515) );
  INV_X1 U9271 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n7301) );
  AND2_X1 U9272 ( .A1(n13538), .A2(n13543), .ZN(n6799) );
  AND2_X1 U9273 ( .A1(n7071), .A2(n11575), .ZN(n6800) );
  NAND2_X1 U9274 ( .A1(n7394), .A2(n8004), .ZN(n6801) );
  OR2_X1 U9275 ( .A1(n8246), .A2(n14132), .ZN(n6802) );
  AND2_X1 U9276 ( .A1(n8102), .A2(n7129), .ZN(n6803) );
  AND2_X1 U9277 ( .A1(n6703), .A2(n7626), .ZN(n6804) );
  AND2_X1 U9278 ( .A1(n7070), .A2(n7071), .ZN(n6805) );
  INV_X1 U9279 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8411) );
  INV_X1 U9280 ( .A(n13614), .ZN(n6988) );
  NAND2_X1 U9281 ( .A1(n7603), .A2(n7604), .ZN(n8309) );
  NAND2_X1 U9282 ( .A1(n11350), .A2(n7183), .ZN(n6806) );
  INV_X1 U9283 ( .A(n13096), .ZN(n15546) );
  NAND2_X1 U9284 ( .A1(n7602), .A2(n8259), .ZN(n10398) );
  NAND2_X1 U9285 ( .A1(n7974), .A2(n7973), .ZN(n14089) );
  INV_X1 U9286 ( .A(n14089), .ZN(n7202) );
  NAND2_X1 U9287 ( .A1(n7310), .A2(n10947), .ZN(n11269) );
  NAND2_X1 U9288 ( .A1(n7316), .A2(n10908), .ZN(n11257) );
  OR2_X1 U9289 ( .A1(n15150), .A2(n6834), .ZN(n6807) );
  OR2_X1 U9290 ( .A1(n15113), .A2(n11748), .ZN(n6808) );
  NAND2_X1 U9291 ( .A1(n8845), .A2(n8844), .ZN(n15638) );
  NOR2_X1 U9292 ( .A1(n6676), .A2(n11762), .ZN(n6809) );
  AOI21_X1 U9293 ( .B1(n8757), .B2(n8391), .A(n7496), .ZN(n7495) );
  AND2_X1 U9294 ( .A1(n8392), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6810) );
  INV_X1 U9295 ( .A(n6973), .ZN(n15376) );
  INV_X1 U9296 ( .A(SI_22_), .ZN(n7129) );
  NAND2_X1 U9297 ( .A1(n7933), .A2(n7932), .ZN(n12470) );
  INV_X1 U9298 ( .A(n12470), .ZN(n7204) );
  INV_X1 U9299 ( .A(n14732), .ZN(n15134) );
  NAND2_X1 U9300 ( .A1(n10907), .A2(n10906), .ZN(n11963) );
  INV_X1 U9301 ( .A(n11963), .ZN(n7176) );
  AND2_X2 U9302 ( .A1(n10792), .A2(n8939), .ZN(n15764) );
  NOR2_X1 U9303 ( .A1(n6676), .A2(n14761), .ZN(n6811) );
  NAND2_X1 U9304 ( .A1(n6973), .A2(n15359), .ZN(n15390) );
  NAND2_X1 U9305 ( .A1(n7852), .A2(n7851), .ZN(n12441) );
  INV_X1 U9306 ( .A(n12441), .ZN(n7193) );
  NOR2_X1 U9307 ( .A1(n10117), .A2(n10116), .ZN(n6812) );
  NAND2_X1 U9308 ( .A1(n11762), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6813) );
  AND2_X1 U9309 ( .A1(n6813), .A2(n8402), .ZN(n6814) );
  XOR2_X1 U9310 ( .A(n13058), .B(P3_REG2_REG_19__SCAN_IN), .Z(n6815) );
  AND2_X1 U9311 ( .A1(n8292), .A2(n12650), .ZN(n13950) );
  XOR2_X1 U9312 ( .A(n8470), .B(n8469), .Z(n6816) );
  INV_X1 U9313 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7686) );
  INV_X1 U9314 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6996) );
  INV_X1 U9315 ( .A(n9803), .ZN(n14161) );
  AOI21_X2 U9316 ( .B1(n10669), .B2(n6973), .A(n15305), .ZN(n15287) );
  AOI21_X2 U9317 ( .B1(n13810), .B2(n15293), .A(n13809), .ZN(n14023) );
  NAND2_X1 U9318 ( .A1(n10011), .A2(n9883), .ZN(n9908) );
  NAND2_X1 U9319 ( .A1(n8268), .A2(n8269), .ZN(n11636) );
  NAND2_X1 U9320 ( .A1(n6935), .A2(n7590), .ZN(n13805) );
  NAND2_X1 U9321 ( .A1(n13987), .A2(n14000), .ZN(n6952) );
  NAND2_X1 U9322 ( .A1(n7559), .A2(n6782), .ZN(n12463) );
  NAND2_X1 U9323 ( .A1(n12438), .A2(n12437), .ZN(n12445) );
  NAND2_X1 U9324 ( .A1(n6830), .A2(n6827), .ZN(n12393) );
  OR2_X1 U9325 ( .A1(n12508), .A2(n12507), .ZN(n6848) );
  NOR2_X1 U9326 ( .A1(n12540), .A2(n12539), .ZN(n12544) );
  NAND2_X1 U9327 ( .A1(n12416), .A2(n12417), .ZN(n12415) );
  NOR2_X1 U9328 ( .A1(n14550), .A2(n6771), .ZN(n14531) );
  NAND2_X1 U9329 ( .A1(n6817), .A2(n12131), .ZN(P1_U3242) );
  NAND2_X1 U9330 ( .A1(n6819), .A2(n6818), .ZN(n6817) );
  NAND3_X1 U9331 ( .A1(n7254), .A2(n7255), .A3(n7253), .ZN(n6819) );
  NAND2_X1 U9332 ( .A1(n7741), .A2(n7376), .ZN(n7375) );
  AOI21_X2 U9333 ( .B1(n11761), .B2(n11892), .A(n6809), .ZN(n14479) );
  NAND2_X1 U9334 ( .A1(n8143), .A2(n8142), .ZN(n8159) );
  NAND2_X1 U9335 ( .A1(n14676), .A2(n6832), .ZN(n14742) );
  NAND2_X1 U9336 ( .A1(n8103), .A2(n6803), .ZN(n8105) );
  OAI21_X1 U9337 ( .B1(n8141), .B2(SI_24_), .A(n8158), .ZN(n8145) );
  NAND2_X2 U9338 ( .A1(n13982), .A2(n8019), .ZN(n13955) );
  OAI21_X2 U9339 ( .B1(n10848), .B2(n7775), .A(n7776), .ZN(n10322) );
  AOI22_X1 U9340 ( .A1(n13812), .A2(n8211), .B1(n13683), .B2(n14107), .ZN(
        n13801) );
  NAND2_X1 U9341 ( .A1(n6877), .A2(n12629), .ZN(n11407) );
  NAND2_X1 U9342 ( .A1(n7801), .A2(n7800), .ZN(n10394) );
  NAND2_X1 U9343 ( .A1(n7486), .A2(n7485), .ZN(n10555) );
  NAND2_X1 U9344 ( .A1(n8073), .A2(n8072), .ZN(n13911) );
  NAND2_X2 U9345 ( .A1(n8101), .A2(n8100), .ZN(n13888) );
  XNOR2_X1 U9346 ( .A(n10576), .B(n10425), .ZN(n10579) );
  NAND2_X1 U9347 ( .A1(n14279), .A2(n12815), .ZN(n7060) );
  NAND2_X1 U9348 ( .A1(n14212), .A2(n12803), .ZN(n14280) );
  AOI21_X1 U9349 ( .B1(n12549), .B2(n12548), .A(n12547), .ZN(n6825) );
  OAI21_X1 U9350 ( .B1(n6824), .B2(n6825), .A(n7551), .ZN(n12574) );
  NOR2_X1 U9351 ( .A1(n15159), .A2(n15158), .ZN(n15157) );
  XOR2_X2 U9352 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9041), .Z(n9042) );
  NAND2_X1 U9353 ( .A1(n6871), .A2(n6870), .ZN(n6869) );
  NAND2_X1 U9354 ( .A1(n9025), .A2(n9026), .ZN(n8990) );
  INV_X1 U9355 ( .A(n6869), .ZN(n9064) );
  XNOR2_X1 U9356 ( .A(n9038), .B(n6866), .ZN(n15765) );
  NAND2_X1 U9357 ( .A1(n14787), .A2(n14788), .ZN(n6821) );
  NOR2_X1 U9358 ( .A1(n15767), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n9044) );
  XNOR2_X1 U9359 ( .A(n9042), .B(n9043), .ZN(n15767) );
  XNOR2_X2 U9360 ( .A(n8998), .B(n9264), .ZN(n9041) );
  NAND2_X1 U9361 ( .A1(n9069), .A2(n15229), .ZN(n7097) );
  NOR2_X1 U9362 ( .A1(n15014), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U9363 ( .A1(n7289), .A2(n7288), .ZN(n7287) );
  NAND2_X1 U9364 ( .A1(n8831), .A2(n8833), .ZN(n8835) );
  AND2_X4 U9365 ( .A1(n10174), .A2(n10173), .ZN(n12848) );
  NAND2_X1 U9366 ( .A1(n7541), .A2(n6786), .ZN(n12508) );
  OAI21_X1 U9367 ( .B1(n12549), .B2(n12548), .A(n6781), .ZN(n6824) );
  OAI22_X1 U9368 ( .A1(n12373), .A2(n12372), .B1(n12371), .B2(n12370), .ZN(
        n6879) );
  NAND2_X1 U9369 ( .A1(n12398), .A2(n12397), .ZN(n12404) );
  NAND2_X1 U9370 ( .A1(n12480), .A2(n12479), .ZN(n12487) );
  INV_X1 U9371 ( .A(n12384), .ZN(n6885) );
  NAND2_X1 U9372 ( .A1(n6829), .A2(n6828), .ZN(n6827) );
  NAND2_X1 U9373 ( .A1(n6886), .A2(n6885), .ZN(n6830) );
  NAND2_X1 U9374 ( .A1(n12380), .A2(n12379), .ZN(n12386) );
  OAI21_X2 U9375 ( .B1(n13888), .B2(n7508), .A(n7507), .ZN(n13861) );
  NAND2_X1 U9376 ( .A1(n7468), .A2(n7754), .ZN(n10848) );
  INV_X1 U9377 ( .A(n11634), .ZN(n6841) );
  NAND2_X1 U9378 ( .A1(n11399), .A2(n11398), .ZN(n7333) );
  INV_X1 U9379 ( .A(n7121), .ZN(n14678) );
  NOR2_X2 U9380 ( .A1(n14597), .A2(n6826), .ZN(n14585) );
  NAND2_X1 U9381 ( .A1(n14741), .A2(n15150), .ZN(n6835) );
  NAND2_X1 U9382 ( .A1(n6837), .A2(n15134), .ZN(n6836) );
  NOR2_X1 U9383 ( .A1(n14508), .A2(n14507), .ZN(n14506) );
  NAND2_X1 U9384 ( .A1(n14104), .A2(n6802), .ZN(P2_U3495) );
  INV_X1 U9385 ( .A(n8145), .ZN(n8143) );
  INV_X1 U9386 ( .A(n7590), .ZN(n6938) );
  NAND2_X1 U9387 ( .A1(n8124), .A2(n8123), .ZN(n8140) );
  NAND2_X1 U9388 ( .A1(n6932), .A2(n6931), .ZN(n13788) );
  INV_X1 U9389 ( .A(n6937), .ZN(n6936) );
  NAND2_X1 U9390 ( .A1(n7928), .A2(n6714), .ZN(n7947) );
  INV_X1 U9391 ( .A(n12516), .ZN(n6851) );
  OAI21_X1 U9392 ( .B1(n12487), .B2(n12486), .A(n7542), .ZN(n6831) );
  AOI21_X1 U9393 ( .B1(n12487), .B2(n12486), .A(n12484), .ZN(n12485) );
  NAND2_X1 U9394 ( .A1(n12376), .A2(n12375), .ZN(n12374) );
  NAND2_X1 U9395 ( .A1(n7947), .A2(n7945), .ZN(n7966) );
  INV_X1 U9396 ( .A(n14575), .ZN(n7347) );
  NAND2_X1 U9397 ( .A1(n14489), .A2(n7122), .ZN(n14473) );
  NAND2_X1 U9398 ( .A1(n6835), .A2(n6807), .ZN(P1_U3557) );
  INV_X1 U9399 ( .A(n14671), .ZN(n6837) );
  AOI21_X2 U9400 ( .B1(n14471), .B2(n14792), .A(n14470), .ZN(n14676) );
  NAND2_X1 U9401 ( .A1(n10226), .A2(n11857), .ZN(n10272) );
  NOR2_X1 U9402 ( .A1(n14320), .A2(n10238), .ZN(n11925) );
  NAND2_X1 U9403 ( .A1(n11290), .A2(n11289), .ZN(n14795) );
  INV_X1 U9404 ( .A(n9583), .ZN(n9580) );
  NAND3_X1 U9405 ( .A1(n7174), .A2(n7402), .A3(n7173), .ZN(n9583) );
  OR2_X2 U9406 ( .A1(n11008), .A2(n11867), .ZN(n11009) );
  OR2_X2 U9407 ( .A1(n13911), .A2(n8099), .ZN(n8101) );
  NAND2_X1 U9408 ( .A1(n9712), .A2(n9713), .ZN(n7719) );
  XNOR2_X2 U9409 ( .A(n6878), .B(n15282), .ZN(n9712) );
  NAND2_X1 U9410 ( .A1(n7863), .A2(n7862), .ZN(n10833) );
  NAND2_X1 U9411 ( .A1(n10737), .A2(n10735), .ZN(n7468) );
  NOR2_X1 U9412 ( .A1(n6789), .A2(n7516), .ZN(n7515) );
  INV_X1 U9413 ( .A(n13777), .ZN(n6946) );
  NAND2_X1 U9414 ( .A1(n6876), .A2(n13986), .ZN(n14003) );
  NAND2_X1 U9415 ( .A1(n13403), .A2(n6798), .ZN(P3_U3454) );
  NAND2_X1 U9416 ( .A1(n13330), .A2(n6797), .ZN(P3_U3486) );
  NAND2_X1 U9417 ( .A1(n7209), .A2(n15638), .ZN(n15626) );
  OAI21_X2 U9418 ( .B1(n8881), .B2(n13157), .A(n13171), .ZN(n13154) );
  NAND2_X1 U9419 ( .A1(n7205), .A2(n7204), .ZN(n11240) );
  NOR2_X4 U9420 ( .A1(n14039), .A2(n13872), .ZN(n13855) );
  NAND4_X1 U9421 ( .A1(n7909), .A2(n6941), .A3(n6942), .A4(n7663), .ZN(n8313)
         );
  NAND2_X1 U9422 ( .A1(n12545), .A2(n12546), .ZN(n12549) );
  AND3_X2 U9423 ( .A1(n7663), .A2(n7908), .A3(n7678), .ZN(n6939) );
  AND4_X2 U9424 ( .A1(n7661), .A2(n7659), .A3(n7660), .A4(n7658), .ZN(n7663)
         );
  OAI21_X1 U9425 ( .B1(n12544), .B2(n12543), .A(n12542), .ZN(n12545) );
  INV_X1 U9426 ( .A(n12519), .ZN(n6853) );
  OAI21_X1 U9427 ( .B1(n6849), .B2(n12506), .A(n6848), .ZN(n12513) );
  NAND2_X1 U9428 ( .A1(n6853), .A2(n6850), .ZN(n12524) );
  NAND2_X1 U9429 ( .A1(n6852), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U9430 ( .A1(n12518), .A2(n12517), .ZN(n6852) );
  INV_X1 U9431 ( .A(n12402), .ZN(n6883) );
  NAND2_X1 U9432 ( .A1(n7675), .A2(n7665), .ZN(n7669) );
  NAND2_X1 U9433 ( .A1(n11175), .A2(n11174), .ZN(n11364) );
  AND2_X1 U9434 ( .A1(n11170), .A2(n15024), .ZN(n6856) );
  NAND2_X2 U9435 ( .A1(n14502), .A2(n14446), .ZN(n14484) );
  NAND2_X1 U9436 ( .A1(n14483), .A2(n14448), .ZN(n14469) );
  OAI22_X1 U9437 ( .A1(n11256), .A2(n11865), .B1(n10974), .B2(n15107), .ZN(
        n11008) );
  NAND2_X1 U9438 ( .A1(n7440), .A2(n7438), .ZN(n14550) );
  NAND2_X1 U9439 ( .A1(n7710), .A2(n7724), .ZN(n15152) );
  NOR2_X1 U9440 ( .A1(n13731), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U9441 ( .A1(n6755), .A2(n6861), .ZN(n13731) );
  INV_X1 U9442 ( .A(n13748), .ZN(n6861) );
  INV_X1 U9443 ( .A(n14786), .ZN(n6870) );
  NAND2_X1 U9444 ( .A1(n15766), .A2(n15765), .ZN(n9040) );
  XNOR2_X1 U9445 ( .A(n9027), .B(n7113), .ZN(n15776) );
  NAND2_X1 U9446 ( .A1(n15776), .A2(n15777), .ZN(n7112) );
  OAI21_X2 U9447 ( .B1(n14777), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6669), .ZN(
        n6867) );
  NAND2_X1 U9448 ( .A1(n11407), .A2(n7962), .ZN(n11634) );
  INV_X1 U9449 ( .A(n11409), .ZN(n6877) );
  INV_X1 U9450 ( .A(n14001), .ZN(n6876) );
  NAND2_X1 U9451 ( .A1(n6947), .A2(n6946), .ZN(n6945) );
  NAND2_X1 U9452 ( .A1(n7517), .A2(n7515), .ZN(n7941) );
  XNOR2_X1 U9453 ( .A(n10063), .B(n9897), .ZN(n9875) );
  NAND2_X1 U9454 ( .A1(n9904), .A2(n9903), .ZN(n9902) );
  NAND2_X1 U9455 ( .A1(n8125), .A2(n8140), .ZN(n11793) );
  NAND2_X1 U9456 ( .A1(n8105), .A2(n7396), .ZN(n7128) );
  NAND2_X1 U9457 ( .A1(n7115), .A2(n6887), .ZN(n7965) );
  NOR2_X1 U9458 ( .A1(n7347), .A2(n7339), .ZN(n7338) );
  NAND2_X1 U9459 ( .A1(n7373), .A2(n6808), .ZN(P1_U3525) );
  INV_X1 U9460 ( .A(n7118), .ZN(n7117) );
  AND2_X2 U9461 ( .A1(n7556), .A2(n7555), .ZN(n9078) );
  XNOR2_X1 U9462 ( .A(n6867), .B(n6747), .ZN(SUB_1596_U4) );
  INV_X1 U9463 ( .A(n15008), .ZN(n7095) );
  NAND3_X1 U9464 ( .A1(n7093), .A2(n9073), .A3(n7096), .ZN(n7558) );
  NAND2_X1 U9465 ( .A1(n9907), .A2(n9887), .ZN(n9888) );
  NOR2_X1 U9466 ( .A1(n15506), .A2(n15505), .ZN(n15504) );
  NAND3_X1 U9467 ( .A1(n6872), .A2(n6890), .A3(n14884), .ZN(P3_U3200) );
  AND2_X1 U9468 ( .A1(n14881), .A2(n14880), .ZN(n6873) );
  NOR2_X1 U9469 ( .A1(n14852), .A2(n13056), .ZN(n14881) );
  NAND2_X1 U9470 ( .A1(n9888), .A2(n10062), .ZN(n10051) );
  XNOR2_X1 U9471 ( .A(n13052), .B(n13101), .ZN(n14816) );
  XNOR2_X1 U9472 ( .A(n7287), .B(n6815), .ZN(n13113) );
  INV_X1 U9473 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8619) );
  OAI21_X1 U9474 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9909) );
  NAND2_X1 U9475 ( .A1(n8085), .A2(n8084), .ZN(n8103) );
  NAND2_X1 U9476 ( .A1(n10222), .A2(n10221), .ZN(n7303) );
  NAND2_X1 U9477 ( .A1(n14491), .A2(n14490), .ZN(n14489) );
  NAND2_X1 U9478 ( .A1(n7334), .A2(n6891), .ZN(n7131) );
  NAND2_X1 U9479 ( .A1(n14741), .A2(n15113), .ZN(n7373) );
  AOI21_X2 U9480 ( .B1(n14412), .B2(n14429), .A(n14411), .ZN(n14649) );
  XNOR2_X1 U9481 ( .A(n11129), .B(n14318), .ZN(n7348) );
  AND3_X2 U9482 ( .A1(n10096), .A2(n10097), .A3(n10095), .ZN(n11129) );
  NAND2_X2 U9483 ( .A1(n13861), .A2(n13860), .ZN(n13859) );
  NAND2_X1 U9484 ( .A1(n13784), .A2(n15390), .ZN(n6947) );
  INV_X1 U9485 ( .A(n9712), .ZN(n12611) );
  NOR2_X1 U9486 ( .A1(n13776), .A2(n6945), .ZN(n8340) );
  NAND2_X1 U9487 ( .A1(n13915), .A2(n13914), .ZN(n8073) );
  NAND2_X1 U9488 ( .A1(n6881), .A2(n6880), .ZN(n12433) );
  NAND2_X1 U9489 ( .A1(n6879), .A2(n12374), .ZN(n12380) );
  NAND3_X1 U9490 ( .A1(n12421), .A2(n12420), .A3(n6791), .ZN(n6881) );
  OAI21_X1 U9491 ( .B1(n12404), .B2(n12403), .A(n6882), .ZN(n7574) );
  NAND2_X1 U9492 ( .A1(n6884), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U9493 ( .A1(n12404), .A2(n12403), .ZN(n6884) );
  NAND2_X1 U9494 ( .A1(n12386), .A2(n12385), .ZN(n6886) );
  NAND2_X1 U9495 ( .A1(n6690), .A2(n7386), .ZN(n6887) );
  OAI21_X1 U9496 ( .B1(n6711), .B2(n7119), .A(n7923), .ZN(n7118) );
  NAND2_X1 U9497 ( .A1(n8080), .A2(n8079), .ZN(n8085) );
  AOI21_X1 U9498 ( .B1(n12127), .B2(n12126), .A(n12125), .ZN(n7254) );
  NOR2_X2 U9499 ( .A1(n14832), .A2(n6888), .ZN(n13055) );
  NOR2_X2 U9500 ( .A1(n14834), .A2(n14833), .ZN(n14832) );
  INV_X1 U9501 ( .A(n7289), .ZN(n14882) );
  AND2_X1 U9502 ( .A1(n9442), .A2(n9441), .ZN(n7406) );
  NAND2_X1 U9503 ( .A1(n7781), .A2(n7780), .ZN(n7786) );
  NAND2_X1 U9504 ( .A1(n14678), .A2(n14450), .ZN(n7304) );
  INV_X1 U9505 ( .A(n7318), .ZN(n7317) );
  NAND2_X2 U9506 ( .A1(n14616), .A2(n14439), .ZN(n14596) );
  INV_X4 U9507 ( .A(n10092), .ZN(n11852) );
  XNOR2_X1 U9508 ( .A(n6892), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13758) );
  OR2_X1 U9509 ( .A1(n13749), .A2(n13748), .ZN(n6892) );
  NAND4_X1 U9510 ( .A1(n6902), .A2(n6901), .A3(n8405), .A4(n8908), .ZN(n6896)
         );
  NAND4_X1 U9511 ( .A1(n8461), .A2(n8406), .A3(n6898), .A4(n6900), .ZN(n6897)
         );
  NAND2_X1 U9512 ( .A1(n15602), .A2(n6698), .ZN(n6905) );
  AOI21_X1 U9513 ( .B1(n13174), .B2(n13173), .A(n8803), .ZN(n13156) );
  OR2_X1 U9514 ( .A1(n13174), .A2(n6912), .ZN(n6911) );
  NAND2_X1 U9515 ( .A1(n11528), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U9516 ( .A1(n7037), .A2(n6923), .ZN(n8733) );
  NAND2_X1 U9517 ( .A1(n10306), .A2(n15624), .ZN(n12184) );
  INV_X1 U9518 ( .A(n15646), .ZN(n10306) );
  NAND2_X1 U9519 ( .A1(n13833), .A2(n6933), .ZN(n6931) );
  NAND2_X1 U9520 ( .A1(n13833), .A2(n7589), .ZN(n6935) );
  AND4_X2 U9521 ( .A1(n7634), .A2(n7633), .A3(n7632), .A4(n7763), .ZN(n7908)
         );
  NAND2_X1 U9522 ( .A1(n6952), .A2(n6951), .ZN(n8274) );
  INV_X4 U9523 ( .A(n7715), .ZN(n12576) );
  NAND2_X1 U9524 ( .A1(n6956), .A2(n12576), .ZN(n8148) );
  NAND2_X2 U9525 ( .A1(n12656), .A2(n12660), .ZN(n12368) );
  NAND2_X1 U9526 ( .A1(n11330), .A2(n6970), .ZN(n6969) );
  NAND2_X2 U9527 ( .A1(n7657), .A2(n13759), .ZN(n6973) );
  OR2_X1 U9528 ( .A1(n10889), .A2(n6973), .ZN(n6972) );
  NAND2_X1 U9529 ( .A1(n6975), .A2(n15376), .ZN(n6974) );
  NAND2_X1 U9530 ( .A1(n13618), .A2(n6980), .ZN(n6976) );
  NAND4_X1 U9531 ( .A1(n6991), .A2(n7908), .A3(n7639), .A4(n7761), .ZN(n8008)
         );
  NAND2_X1 U9532 ( .A1(n8358), .A2(n7006), .ZN(n7002) );
  NAND2_X1 U9533 ( .A1(n7003), .A2(n7002), .ZN(n8603) );
  NAND3_X1 U9534 ( .A1(n7012), .A2(n12298), .A3(n12164), .ZN(n7011) );
  NAND2_X1 U9535 ( .A1(n8496), .A2(n7017), .ZN(n7013) );
  NAND2_X1 U9536 ( .A1(n7013), .A2(n7014), .ZN(n8529) );
  INV_X1 U9537 ( .A(n8371), .ZN(n7023) );
  NAND2_X1 U9538 ( .A1(n7489), .A2(n7025), .ZN(n12321) );
  NAND2_X1 U9539 ( .A1(n7026), .A2(n12292), .ZN(n7025) );
  NAND2_X1 U9540 ( .A1(n12319), .A2(n12317), .ZN(n7026) );
  INV_X1 U9541 ( .A(n8387), .ZN(n7027) );
  NAND2_X1 U9542 ( .A1(n8388), .A2(n7027), .ZN(n7030) );
  INV_X1 U9543 ( .A(n13025), .ZN(n13407) );
  NAND2_X1 U9544 ( .A1(n11481), .A2(n7160), .ZN(n7033) );
  XNOR2_X1 U9545 ( .A(n8805), .B(n8804), .ZN(n11481) );
  NAND2_X1 U9546 ( .A1(n13219), .A2(n12286), .ZN(n7035) );
  NAND2_X1 U9547 ( .A1(n13232), .A2(n12282), .ZN(n7036) );
  NAND2_X1 U9548 ( .A1(n13290), .A2(n8717), .ZN(n7037) );
  INV_X1 U9549 ( .A(n8844), .ZN(n15640) );
  NAND2_X2 U9550 ( .A1(n9868), .A2(n11804), .ZN(n12152) );
  NAND4_X1 U9551 ( .A1(n8410), .A2(n7058), .A3(n8414), .A4(n8616), .ZN(n7056)
         );
  AND4_X2 U9552 ( .A1(n7063), .A2(n7061), .A3(n7064), .A4(n9819), .ZN(n7402)
         );
  AND2_X2 U9553 ( .A1(n7402), .A2(n7401), .ZN(n9448) );
  XNOR2_X1 U9554 ( .A(n11567), .B(n11494), .ZN(n11569) );
  NAND2_X1 U9555 ( .A1(n7070), .A2(n6800), .ZN(n12692) );
  NAND2_X1 U9556 ( .A1(n11569), .A2(n11568), .ZN(n7070) );
  INV_X2 U9557 ( .A(n6686), .ZN(n7074) );
  NAND2_X1 U9558 ( .A1(n10719), .A2(n6694), .ZN(n7076) );
  OAI21_X1 U9559 ( .B1(n10719), .B2(n7078), .A(n6694), .ZN(n11316) );
  INV_X1 U9560 ( .A(n12838), .ZN(n7079) );
  OAI21_X2 U9561 ( .B1(n12784), .B2(n7082), .A(n7080), .ZN(n14212) );
  NAND2_X1 U9562 ( .A1(n10389), .A2(n7086), .ZN(n9770) );
  NOR2_X1 U9563 ( .A1(n7088), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U9564 ( .A1(n9072), .A2(n7092), .ZN(n7091) );
  NAND2_X1 U9565 ( .A1(n9072), .A2(n15230), .ZN(n7093) );
  INV_X1 U9566 ( .A(n15003), .ZN(n7098) );
  AND2_X2 U9567 ( .A1(n7098), .A2(n7097), .ZN(n15008) );
  NAND3_X1 U9568 ( .A1(n7104), .A2(n7103), .A3(n7109), .ZN(n7101) );
  NAND2_X1 U9569 ( .A1(n15017), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7102) );
  AND2_X2 U9570 ( .A1(n9078), .A2(n9079), .ZN(n15014) );
  NAND2_X1 U9571 ( .A1(n7112), .A2(n9028), .ZN(n9031) );
  NAND2_X1 U9572 ( .A1(n7781), .A2(n7123), .ZN(n7126) );
  NAND3_X1 U9573 ( .A1(n7126), .A2(n7838), .A3(n7125), .ZN(n7841) );
  NAND2_X1 U9574 ( .A1(n8119), .A2(n7128), .ZN(n8124) );
  NAND2_X1 U9575 ( .A1(n8103), .A2(n8102), .ZN(n8104) );
  AND3_X2 U9576 ( .A1(n7132), .A2(n7131), .A3(n6790), .ZN(n14519) );
  MUX2_X1 U9577 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11804), .Z(n7782) );
  MUX2_X1 U9578 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11804), .Z(n7804) );
  MUX2_X1 U9579 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11804), .Z(n7842) );
  MUX2_X1 U9580 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11804), .Z(n7866) );
  MUX2_X1 U9581 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n11804), .Z(n7925) );
  MUX2_X1 U9582 ( .A(n10410), .B(n10411), .S(n11804), .Z(n7987) );
  MUX2_X1 U9583 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n11804), .Z(n8020) );
  NAND2_X2 U9584 ( .A1(n6672), .A2(n11804), .ZN(n7715) );
  NAND2_X1 U9585 ( .A1(n7136), .A2(n7137), .ZN(n12924) );
  NAND3_X1 U9586 ( .A1(n12880), .A2(n7145), .A3(n7140), .ZN(n7136) );
  NAND2_X1 U9587 ( .A1(n12891), .A2(n7154), .ZN(n7153) );
  NAND2_X2 U9588 ( .A1(n9868), .A2(n10090), .ZN(n8749) );
  NAND2_X1 U9589 ( .A1(n7161), .A2(n6780), .ZN(n11432) );
  NAND2_X1 U9590 ( .A1(n11112), .A2(n7162), .ZN(n7161) );
  XNOR2_X1 U9591 ( .A(n10526), .B(n15636), .ZN(n10367) );
  NAND2_X1 U9592 ( .A1(n10365), .A2(n10364), .ZN(n10368) );
  NAND2_X1 U9593 ( .A1(n13010), .A2(n6693), .ZN(n7166) );
  INV_X1 U9594 ( .A(n12910), .ZN(n7167) );
  NAND2_X1 U9595 ( .A1(n11649), .A2(n11648), .ZN(n11652) );
  NAND2_X1 U9596 ( .A1(n9583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9585) );
  NOR2_X1 U9597 ( .A1(n11137), .A2(n15084), .ZN(n15056) );
  INV_X2 U9598 ( .A(n6676), .ZN(n11853) );
  INV_X2 U9599 ( .A(n11934), .ZN(n7180) );
  NOR2_X2 U9600 ( .A1(n6706), .A2(n14120), .ZN(n13906) );
  NOR2_X2 U9601 ( .A1(n11240), .A2(n12483), .ZN(n7203) );
  NOR2_X2 U9602 ( .A1(n11158), .A2(n14912), .ZN(n7205) );
  NAND2_X1 U9603 ( .A1(n15608), .A2(n7206), .ZN(n10998) );
  NAND2_X1 U9604 ( .A1(n13154), .A2(n7217), .ZN(n7210) );
  OAI21_X1 U9605 ( .B1(n8859), .B2(n7231), .A(n7229), .ZN(n13311) );
  NAND2_X1 U9606 ( .A1(n7240), .A2(n7237), .ZN(n10175) );
  NAND3_X1 U9607 ( .A1(n11939), .A2(n7246), .A3(n7242), .ZN(n11945) );
  OAI21_X1 U9608 ( .B1(n11933), .B2(n11932), .A(n11931), .ZN(n7248) );
  INV_X1 U9609 ( .A(n12055), .ZN(n12052) );
  NAND3_X1 U9610 ( .A1(n11983), .A2(n11982), .A3(n6788), .ZN(n7251) );
  INV_X1 U9611 ( .A(n11985), .ZN(n7252) );
  OAI21_X1 U9612 ( .B1(n6732), .B2(n7261), .A(n7260), .ZN(n12100) );
  INV_X1 U9613 ( .A(n12085), .ZN(n7270) );
  NAND3_X1 U9614 ( .A1(n12065), .A2(n12064), .A3(n6792), .ZN(n7272) );
  INV_X1 U9615 ( .A(n12066), .ZN(n7273) );
  NAND3_X1 U9616 ( .A1(n11995), .A2(n11994), .A3(n6776), .ZN(n7277) );
  AND2_X1 U9617 ( .A1(n12006), .A2(n11998), .ZN(n7279) );
  NAND2_X1 U9618 ( .A1(n10389), .A2(n6783), .ZN(n7283) );
  OAI21_X1 U9619 ( .B1(n11950), .B2(n11949), .A(n11948), .ZN(n11952) );
  NAND2_X1 U9620 ( .A1(n11945), .A2(n11944), .ZN(n11950) );
  AND2_X2 U9621 ( .A1(n7290), .A2(n6735), .ZN(n14834) );
  OR2_X2 U9622 ( .A1(n14816), .A2(n14817), .ZN(n7290) );
  NAND2_X1 U9623 ( .A1(n15504), .A2(n7294), .ZN(n7292) );
  INV_X1 U9624 ( .A(n7295), .ZN(n13048) );
  OR2_X1 U9625 ( .A1(n10009), .A2(n15668), .ZN(n10011) );
  OAI21_X1 U9626 ( .B1(n10019), .B2(n9995), .A(n9883), .ZN(n10009) );
  NOR2_X2 U9627 ( .A1(n15472), .A2(n10622), .ZN(n15492) );
  NAND2_X1 U9628 ( .A1(n7303), .A2(n10262), .ZN(n10267) );
  OAI21_X1 U9629 ( .B1(n10221), .B2(n10222), .A(n7303), .ZN(n10223) );
  NAND3_X1 U9630 ( .A1(n7305), .A2(n7372), .A3(n7304), .ZN(n14671) );
  NAND2_X1 U9631 ( .A1(n10899), .A2(n7306), .ZN(n11136) );
  NAND2_X1 U9632 ( .A1(n10473), .A2(n6785), .ZN(n7307) );
  NAND2_X1 U9633 ( .A1(n10473), .A2(n10472), .ZN(n10898) );
  NAND2_X1 U9634 ( .A1(n11136), .A2(n11135), .ZN(n10901) );
  NAND2_X1 U9635 ( .A1(n11349), .A2(n7311), .ZN(n7308) );
  NAND2_X1 U9636 ( .A1(n7308), .A2(n7309), .ZN(n14790) );
  NAND2_X1 U9637 ( .A1(n11094), .A2(n7317), .ZN(n7314) );
  NAND2_X1 U9638 ( .A1(n7314), .A2(n7315), .ZN(n11015) );
  NAND2_X1 U9639 ( .A1(n7320), .A2(n7321), .ZN(n14598) );
  AND2_X2 U9640 ( .A1(n7320), .A2(n6772), .ZN(n14597) );
  OR2_X2 U9641 ( .A1(n14649), .A2(n7322), .ZN(n7320) );
  NAND2_X1 U9642 ( .A1(n7342), .A2(n7345), .ZN(n14549) );
  NAND2_X2 U9643 ( .A1(n7349), .A2(n9809), .ZN(n14318) );
  AND3_X1 U9644 ( .A1(n9810), .A2(n9807), .A3(n9808), .ZN(n7349) );
  NAND3_X1 U9645 ( .A1(n7405), .A2(n9448), .A3(n6700), .ZN(n7465) );
  NAND4_X1 U9646 ( .A1(n7405), .A2(n9448), .A3(n6700), .A4(n9780), .ZN(n14756)
         );
  NAND2_X1 U9647 ( .A1(n11196), .A2(n7357), .ZN(n11330) );
  NAND2_X1 U9648 ( .A1(n7358), .A2(n6775), .ZN(n13560) );
  NAND2_X1 U9649 ( .A1(n10610), .A2(n10514), .ZN(n10516) );
  OR3_X1 U9650 ( .A1(n8008), .A2(n7367), .A3(P2_IR_REG_18__SCAN_IN), .ZN(n7644) );
  OAI21_X1 U9651 ( .B1(n10090), .B2(n9501), .A(n7371), .ZN(n7690) );
  NAND2_X1 U9652 ( .A1(n10090), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7371) );
  OAI21_X1 U9653 ( .B1(n7741), .B2(n7755), .A(n7376), .ZN(n7779) );
  NAND3_X1 U9654 ( .A1(n7375), .A2(n7778), .A3(n7374), .ZN(n7781) );
  NAND2_X1 U9655 ( .A1(n7376), .A2(n7755), .ZN(n7374) );
  NAND2_X1 U9656 ( .A1(n7714), .A2(SI_2_), .ZN(n7381) );
  NAND2_X1 U9657 ( .A1(n7380), .A2(n7383), .ZN(n7382) );
  INV_X1 U9658 ( .A(n7714), .ZN(n7380) );
  NAND2_X1 U9659 ( .A1(n8003), .A2(n6804), .ZN(n7393) );
  NAND2_X1 U9660 ( .A1(n8105), .A2(n8119), .ZN(n11805) );
  NOR2_X2 U9661 ( .A1(n7404), .A2(n7403), .ZN(n7401) );
  NAND3_X1 U9662 ( .A1(n9430), .A2(n10146), .A3(n9822), .ZN(n7403) );
  NAND4_X1 U9663 ( .A1(n9431), .A2(n10149), .A3(n9530), .A4(n9602), .ZN(n7404)
         );
  NAND3_X1 U9664 ( .A1(n7407), .A2(n7406), .A3(n9575), .ZN(n9447) );
  NAND2_X1 U9665 ( .A1(n14200), .A2(n12706), .ZN(n7408) );
  NAND2_X1 U9666 ( .A1(n14938), .A2(n7412), .ZN(n12742) );
  AOI21_X1 U9667 ( .B1(n14155), .B2(n12814), .A(n12822), .ZN(n7430) );
  OAI211_X1 U9668 ( .C1(n14279), .C2(n6766), .A(n7426), .B(n7424), .ZN(n12835)
         );
  NAND2_X1 U9669 ( .A1(n14279), .A2(n7425), .ZN(n7424) );
  NOR2_X1 U9670 ( .A1(n12829), .A2(n7428), .ZN(n7425) );
  NOR2_X1 U9671 ( .A1(n14155), .A2(n12829), .ZN(n7427) );
  INV_X1 U9672 ( .A(n12829), .ZN(n7429) );
  OAI21_X2 U9673 ( .B1(n10205), .B2(n7434), .A(n7433), .ZN(n10291) );
  NAND2_X1 U9674 ( .A1(n10291), .A2(n10290), .ZN(n10417) );
  NAND2_X1 U9675 ( .A1(n14484), .A2(n14485), .ZN(n14483) );
  NAND3_X1 U9676 ( .A1(n7442), .A2(n14596), .A3(n14548), .ZN(n7440) );
  AOI21_X1 U9677 ( .B1(n7442), .B2(n14596), .A(n7439), .ZN(n14552) );
  NAND2_X1 U9678 ( .A1(n7441), .A2(n7446), .ZN(n14562) );
  AND2_X1 U9679 ( .A1(n14575), .A2(n7443), .ZN(n7442) );
  NAND2_X1 U9680 ( .A1(n7445), .A2(n14575), .ZN(n7444) );
  INV_X1 U9681 ( .A(n7446), .ZN(n7445) );
  NAND2_X1 U9682 ( .A1(n14711), .A2(n14443), .ZN(n7450) );
  NAND2_X1 U9683 ( .A1(n11383), .A2(n7454), .ZN(n7453) );
  OAI21_X2 U9684 ( .B1(n11009), .B2(n7461), .A(n7459), .ZN(n11290) );
  OAI21_X1 U9685 ( .B1(n7464), .B2(n7461), .A(n11869), .ZN(n7460) );
  NAND2_X1 U9686 ( .A1(n9580), .A2(n9584), .ZN(n9778) );
  OAI21_X2 U9687 ( .B1(n14644), .B2(n14434), .A(n14436), .ZN(n14624) );
  OAI21_X2 U9688 ( .B1(n14430), .B2(n14429), .A(n14433), .ZN(n14644) );
  NAND2_X1 U9689 ( .A1(n8605), .A2(n8368), .ZN(n8613) );
  NAND2_X1 U9690 ( .A1(n8470), .A2(n8469), .ZN(n7466) );
  NAND2_X1 U9691 ( .A1(n8345), .A2(n8464), .ZN(n7467) );
  INV_X1 U9692 ( .A(n7603), .ZN(n7990) );
  INV_X1 U9693 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7478) );
  NAND2_X1 U9694 ( .A1(n10394), .A2(n7484), .ZN(n7486) );
  NAND2_X1 U9695 ( .A1(n10394), .A2(n12620), .ZN(n7488) );
  AOI21_X1 U9696 ( .B1(n12621), .B2(n7487), .A(n6758), .ZN(n7485) );
  NAND2_X1 U9697 ( .A1(n12319), .A2(n7490), .ZN(n7489) );
  AND2_X1 U9698 ( .A1(n12318), .A2(n12320), .ZN(n7490) );
  NAND2_X1 U9699 ( .A1(n7492), .A2(n7493), .ZN(n8393) );
  NAND2_X1 U9700 ( .A1(n13955), .A2(n7499), .ZN(n7497) );
  NAND2_X1 U9701 ( .A1(n7497), .A2(n7498), .ZN(n13915) );
  OAI211_X2 U9702 ( .C1(n13859), .C2(n7503), .A(n7501), .B(n6750), .ZN(n13812)
         );
  NAND2_X1 U9703 ( .A1(n8400), .A2(n7513), .ZN(n7512) );
  NAND2_X1 U9704 ( .A1(n7512), .A2(n8402), .ZN(n8943) );
  NAND2_X1 U9705 ( .A1(n7512), .A2(n6814), .ZN(n8946) );
  NAND2_X1 U9706 ( .A1(n15646), .A2(n15655), .ZN(n12183) );
  NAND2_X1 U9707 ( .A1(n13244), .A2(n12165), .ZN(n13232) );
  NAND2_X1 U9708 ( .A1(n13207), .A2(n6784), .ZN(n13180) );
  NAND4_X1 U9709 ( .A1(n8410), .A2(n8616), .A3(n8512), .A4(n8411), .ZN(n8690)
         );
  NAND3_X1 U9710 ( .A1(n8410), .A2(n8512), .A3(n8616), .ZN(n8676) );
  INV_X1 U9711 ( .A(n12551), .ZN(n7552) );
  XNOR2_X2 U9712 ( .A(n7554), .B(n7553), .ZN(n14777) );
  NAND2_X1 U9713 ( .A1(n7558), .A2(n7557), .ZN(n7556) );
  INV_X1 U9714 ( .A(n15012), .ZN(n7555) );
  INV_X1 U9715 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7557) );
  NAND3_X1 U9716 ( .A1(n12450), .A2(n12449), .A3(n6787), .ZN(n7559) );
  INV_X1 U9717 ( .A(n12455), .ZN(n7560) );
  NOR2_X1 U9718 ( .A1(n7573), .A2(n7572), .ZN(n7571) );
  INV_X1 U9719 ( .A(n12408), .ZN(n7572) );
  INV_X1 U9720 ( .A(n12407), .ZN(n7573) );
  NAND2_X1 U9721 ( .A1(n12433), .A2(n12434), .ZN(n12432) );
  NAND2_X1 U9722 ( .A1(n12383), .A2(n12363), .ZN(n12365) );
  NOR2_X1 U9723 ( .A1(n7582), .A2(n14912), .ZN(n7581) );
  INV_X1 U9724 ( .A(n8265), .ZN(n7582) );
  AND2_X1 U9725 ( .A1(n7663), .A2(n7662), .ZN(n7604) );
  NAND3_X1 U9726 ( .A1(n7671), .A2(P2_REG3_REG_1__SCAN_IN), .A3(n6681), .ZN(
        n7609) );
  OAI21_X2 U9727 ( .B1(n11636), .B2(n8270), .A(n8271), .ZN(n13987) );
  NAND2_X1 U9728 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  NAND2_X1 U9729 ( .A1(n12113), .A2(n12112), .ZN(n12114) );
  XNOR2_X1 U9730 ( .A(n12903), .B(n12966), .ZN(n12969) );
  NAND2_X1 U9731 ( .A1(n11718), .A2(n11717), .ZN(n11722) );
  XNOR2_X1 U9732 ( .A(n8235), .B(n8234), .ZN(n11761) );
  CLKBUF_X1 U9733 ( .A(n14268), .Z(n14270) );
  NAND2_X2 U9734 ( .A1(n11612), .A2(n11611), .ZN(n14412) );
  NAND2_X1 U9735 ( .A1(n10219), .A2(n11934), .ZN(n11937) );
  NAND2_X1 U9736 ( .A1(n14320), .A2(n10250), .ZN(n10248) );
  AOI21_X1 U9737 ( .B1(n12817), .B2(n14320), .A(n9794), .ZN(n9799) );
  OR2_X1 U9738 ( .A1(n11902), .A2(n10107), .ZN(n10108) );
  OAI22_X1 U9739 ( .A1(n12107), .A2(n12112), .B1(n12106), .B2(n12105), .ZN(
        n12102) );
  NAND2_X1 U9740 ( .A1(n12180), .A2(n12179), .ZN(n10181) );
  INV_X1 U9741 ( .A(n12475), .ZN(n12478) );
  NAND2_X1 U9742 ( .A1(n8439), .A2(n8438), .ZN(n13453) );
  INV_X1 U9743 ( .A(n8439), .ZN(n8441) );
  INV_X1 U9744 ( .A(n8443), .ZN(n13463) );
  INV_X1 U9745 ( .A(n12433), .ZN(n12436) );
  XNOR2_X1 U9746 ( .A(n10100), .B(n12807), .ZN(n10103) );
  INV_X1 U9747 ( .A(n9450), .ZN(n9451) );
  NAND2_X1 U9748 ( .A1(n9450), .A2(n9452), .ZN(n9437) );
  INV_X1 U9749 ( .A(n12416), .ZN(n12419) );
  OAI22_X1 U9750 ( .A1(n12390), .A2(n12655), .B1(n15363), .B2(n12585), .ZN(
        n12391) );
  NAND2_X1 U9751 ( .A1(n15674), .A2(n10175), .ZN(n12179) );
  INV_X1 U9752 ( .A(n10175), .ZN(n15650) );
  INV_X1 U9753 ( .A(n7699), .ZN(n7809) );
  OR2_X1 U9754 ( .A1(n10255), .A2(n10470), .ZN(n15135) );
  NAND2_X2 U9755 ( .A1(n14459), .A2(n14633), .ZN(n14636) );
  XOR2_X1 U9756 ( .A(n9101), .B(n9100), .Z(n7611) );
  OR2_X1 U9757 ( .A1(n14218), .A2(n14217), .ZN(n7612) );
  OR2_X1 U9758 ( .A1(n15407), .A2(n15403), .ZN(n14132) );
  INV_X1 U9759 ( .A(n14132), .ZN(n8335) );
  INV_X2 U9760 ( .A(n15407), .ZN(n15409) );
  AND2_X1 U9761 ( .A1(n12569), .A2(n12568), .ZN(n7613) );
  OR2_X1 U9762 ( .A1(n6686), .A2(n10238), .ZN(n7614) );
  NOR2_X1 U9763 ( .A1(n8216), .A2(n8215), .ZN(n7615) );
  NOR3_X1 U9764 ( .A1(n12602), .A2(n7613), .A3(n12571), .ZN(n7616) );
  AND2_X1 U9765 ( .A1(n8342), .A2(n7621), .ZN(n7617) );
  AND2_X1 U9766 ( .A1(n8337), .A2(n8336), .ZN(n7618) );
  NAND2_X1 U9767 ( .A1(n12599), .A2(n12598), .ZN(n7619) );
  AND2_X1 U9768 ( .A1(n12925), .A2(n15653), .ZN(n7620) );
  OR2_X1 U9769 ( .A1(n15427), .A2(n8341), .ZN(n7621) );
  OR2_X1 U9770 ( .A1(n14079), .A2(n13952), .ZN(n7622) );
  INV_X1 U9771 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7678) );
  OR2_X1 U9772 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9996), .ZN(n7623) );
  INV_X1 U9773 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n7658) );
  INV_X1 U9774 ( .A(n12976), .ZN(n13412) );
  OR2_X1 U9775 ( .A1(n8082), .A2(SI_20_), .ZN(n7624) );
  INV_X1 U9776 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10407) );
  INV_X1 U9777 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8424) );
  INV_X1 U9778 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8691) );
  INV_X1 U9779 ( .A(n13158), .ZN(n12925) );
  AND3_X1 U9780 ( .A1(n9445), .A2(n9434), .A3(n7285), .ZN(n7625) );
  INV_X1 U9781 ( .A(n14245), .ZN(n11302) );
  AND2_X1 U9782 ( .A1(n8004), .A2(n7989), .ZN(n7626) );
  INV_X1 U9783 ( .A(n13241), .ZN(n8744) );
  NAND2_X1 U9784 ( .A1(n13271), .A2(n13270), .ZN(n7627) );
  AND2_X1 U9785 ( .A1(n14118), .A2(n13688), .ZN(n7628) );
  INV_X1 U9786 ( .A(n14450), .ZN(n14428) );
  INV_X1 U9787 ( .A(n12559), .ZN(n13782) );
  AND2_X1 U9788 ( .A1(n10372), .A2(n10525), .ZN(n7630) );
  INV_X1 U9789 ( .A(n15510), .ZN(n10625) );
  INV_X1 U9790 ( .A(n15291), .ZN(n12367) );
  NOR2_X1 U9791 ( .A1(n12368), .A2(n15291), .ZN(n12372) );
  INV_X1 U9792 ( .A(n12376), .ZN(n12377) );
  INV_X1 U9793 ( .A(n11938), .ZN(n11939) );
  INV_X1 U9794 ( .A(n12417), .ZN(n12418) );
  INV_X1 U9795 ( .A(n12434), .ZN(n12435) );
  INV_X1 U9796 ( .A(n12476), .ZN(n12477) );
  AND2_X1 U9797 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  NAND2_X1 U9798 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  INV_X1 U9799 ( .A(n12315), .ZN(n12316) );
  NAND2_X1 U9800 ( .A1(n12544), .A2(n12543), .ZN(n12546) );
  INV_X1 U9801 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9430) );
  INV_X1 U9802 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8404) );
  INV_X1 U9803 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9444) );
  INV_X1 U9804 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U9805 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  OAI21_X1 U9806 ( .B1(n9888), .B2(n10062), .A(n10051), .ZN(n9890) );
  INV_X1 U9807 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8413) );
  INV_X1 U9808 ( .A(n12601), .ZN(n12571) );
  NAND2_X1 U9809 ( .A1(n7942), .A2(n9564), .ZN(n7943) );
  NOR2_X1 U9810 ( .A1(n10654), .A2(n10623), .ZN(n10624) );
  INV_X1 U9811 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11693) );
  NOR2_X1 U9812 ( .A1(n12154), .A2(n13114), .ZN(n8959) );
  INV_X1 U9813 ( .A(n13588), .ZN(n13498) );
  INV_X1 U9814 ( .A(n8130), .ZN(n8128) );
  INV_X1 U9815 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7895) );
  INV_X1 U9816 ( .A(n8091), .ZN(n8089) );
  AND2_X1 U9817 ( .A1(n7977), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7995) );
  INV_X1 U9818 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10720) );
  NOR2_X1 U9819 ( .A1(n9059), .A2(n9058), .ZN(n9006) );
  INV_X1 U9820 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9327) );
  INV_X1 U9821 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9234) );
  INV_X1 U9822 ( .A(n10766), .ZN(n8955) );
  XNOR2_X1 U9823 ( .A(n10626), .B(n10625), .ZN(n15506) );
  AND2_X1 U9824 ( .A1(n13091), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n13045) );
  NAND2_X1 U9825 ( .A1(n8436), .A2(n9236), .ZN(n8820) );
  NAND2_X1 U9826 ( .A1(n13299), .A2(n13298), .ZN(n13285) );
  AND2_X1 U9827 ( .A1(n12246), .A2(n12244), .ZN(n12340) );
  NOR2_X1 U9828 ( .A1(n8960), .A2(n8959), .ZN(n8961) );
  AND2_X1 U9829 ( .A1(n8364), .A2(n8363), .ZN(n8570) );
  NAND2_X1 U9830 ( .A1(n9535), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8353) );
  INV_X1 U9831 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7683) );
  XNOR2_X1 U9832 ( .A(n13493), .B(n12363), .ZN(n10539) );
  AND2_X1 U9833 ( .A1(n8199), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U9834 ( .A1(n8128), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8149) );
  OR2_X1 U9835 ( .A1(n8064), .A2(n13629), .ZN(n8091) );
  NAND2_X1 U9836 ( .A1(n7954), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7978) );
  INV_X1 U9837 ( .A(n13797), .ZN(n8246) );
  INV_X1 U9838 ( .A(n13806), .ZN(n8300) );
  INV_X1 U9839 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7665) );
  INV_X1 U9840 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U9841 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  INV_X1 U9842 ( .A(n12752), .ZN(n12753) );
  INV_X1 U9843 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10938) );
  INV_X1 U9844 ( .A(n11783), .ZN(n11899) );
  NOR2_X1 U9845 ( .A1(n11844), .A2(n11843), .ZN(n11845) );
  NOR2_X1 U9846 ( .A1(n10721), .A2(n10720), .ZN(n10913) );
  INV_X1 U9847 ( .A(n14663), .ZN(n14396) );
  AND2_X1 U9848 ( .A1(n14688), .A2(n14424), .ZN(n14425) );
  NAND2_X1 U9849 ( .A1(n14568), .A2(n7346), .ZN(n14569) );
  AND3_X1 U9850 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10594) );
  OR2_X1 U9851 ( .A1(n14320), .A2(n10250), .ZN(n10247) );
  INV_X1 U9852 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9440) );
  AND2_X1 U9853 ( .A1(n7802), .A2(n7784), .ZN(n7785) );
  NOR2_X1 U9854 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  NAND2_X1 U9855 ( .A1(n11691), .A2(n11690), .ZN(n12843) );
  INV_X1 U9856 ( .A(n13020), .ZN(n13035) );
  AND2_X1 U9857 ( .A1(n8825), .A2(n8824), .ZN(n13158) );
  INV_X1 U9858 ( .A(n15528), .ZN(n13047) );
  INV_X1 U9859 ( .A(n14862), .ZN(n13054) );
  AND2_X1 U9860 ( .A1(n9877), .A2(n9878), .ZN(n9882) );
  INV_X1 U9861 ( .A(n13089), .ZN(n13058) );
  AOI21_X1 U9862 ( .B1(n13237), .B2(n13241), .A(n8873), .ZN(n13227) );
  AND2_X1 U9863 ( .A1(n12275), .A2(n12276), .ZN(n13254) );
  AND4_X1 U9864 ( .A1(n8702), .A2(n8701), .A3(n8700), .A4(n8699), .ZN(n13301)
         );
  AND2_X1 U9865 ( .A1(n13126), .A2(n15732), .ZN(n8966) );
  AND2_X1 U9866 ( .A1(n8971), .A2(n12357), .ZN(n15641) );
  AND2_X1 U9867 ( .A1(n10162), .A2(n15718), .ZN(n15672) );
  OAI21_X1 U9868 ( .B1(n8899), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8901) );
  AND2_X1 U9869 ( .A1(n8383), .A2(n8382), .ZN(n8703) );
  AND2_X1 U9870 ( .A1(n8373), .A2(n8372), .ZN(n8645) );
  AND2_X1 U9871 ( .A1(n8368), .A2(n8367), .ZN(n8602) );
  INV_X1 U9872 ( .A(n13687), .ZN(n13540) );
  OR2_X1 U9873 ( .A1(n8162), .A2(n13599), .ZN(n8181) );
  OR2_X1 U9874 ( .A1(n8149), .A2(n13625), .ZN(n8162) );
  OR2_X1 U9875 ( .A1(n7934), .A2(n15232), .ZN(n7956) );
  OR2_X1 U9876 ( .A1(n8111), .A2(n13645), .ZN(n8130) );
  OR2_X1 U9877 ( .A1(n9484), .A2(n9478), .ZN(n9481) );
  OR2_X1 U9878 ( .A1(n8043), .A2(n8042), .ZN(n8064) );
  INV_X1 U9879 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15232) );
  AND2_X1 U9880 ( .A1(n9751), .A2(n14137), .ZN(n9745) );
  AND2_X1 U9881 ( .A1(n7651), .A2(n12646), .ZN(n9741) );
  OR2_X1 U9882 ( .A1(n9470), .A2(n15342), .ZN(n10558) );
  NAND2_X1 U9883 ( .A1(n15407), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U9884 ( .A1(n12559), .A2(n8335), .ZN(n8337) );
  INV_X1 U9885 ( .A(n12638), .ZN(n13846) );
  INV_X1 U9886 ( .A(n13691), .ZN(n12472) );
  NAND2_X1 U9887 ( .A1(n11831), .A2(n11892), .ZN(n11833) );
  NAND2_X1 U9888 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  INV_X1 U9889 ( .A(n10575), .ZN(n10425) );
  INV_X1 U9890 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10952) );
  OR2_X1 U9891 ( .A1(n9768), .A2(n9767), .ZN(n9804) );
  AND2_X1 U9892 ( .A1(n11845), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11881) );
  INV_X1 U9893 ( .A(n14389), .ZN(n15034) );
  OR2_X1 U9894 ( .A1(n11601), .A2(n11600), .ZN(n11844) );
  NAND2_X1 U9895 ( .A1(n14636), .A2(n10477), .ZN(n14614) );
  OR2_X1 U9896 ( .A1(n9768), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9755) );
  INV_X1 U9897 ( .A(n14638), .ZN(n14735) );
  INV_X1 U9898 ( .A(n11874), .ZN(n14429) );
  NAND2_X1 U9899 ( .A1(n9813), .A2(n9571), .ZN(n9803) );
  INV_X1 U9900 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U9901 ( .A1(n8159), .A2(n8158), .ZN(n8172) );
  NAND2_X1 U9902 ( .A1(n9041), .A2(n9729), .ZN(n8999) );
  OAI22_X1 U9903 ( .A1(n12969), .A2(n13186), .B1(n12968), .B2(n12967), .ZN(
        n12972) );
  INV_X1 U9904 ( .A(n13023), .ZN(n15430) );
  INV_X1 U9905 ( .A(n13027), .ZN(n15432) );
  AOI21_X1 U9906 ( .B1(n13130), .B2(n8465), .A(n8447), .ZN(n13041) );
  AND3_X1 U9907 ( .A1(n8743), .A2(n8742), .A3(n8741), .ZN(n13257) );
  NAND2_X1 U9908 ( .A1(n8898), .A2(n8897), .ZN(n13129) );
  NAND2_X1 U9909 ( .A1(n8767), .A2(n8766), .ZN(n13229) );
  INV_X1 U9910 ( .A(n13315), .ZN(n13287) );
  INV_X1 U9911 ( .A(n6668), .ZN(n15676) );
  INV_X1 U9912 ( .A(n15718), .ZN(n15677) );
  AND2_X1 U9913 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  AND2_X1 U9914 ( .A1(n13116), .A2(n13115), .ZN(n13391) );
  NAND2_X1 U9915 ( .A1(n8843), .A2(n12176), .ZN(n15718) );
  NAND2_X1 U9916 ( .A1(n15662), .A2(n15719), .ZN(n15732) );
  NAND2_X1 U9917 ( .A1(n10160), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9509) );
  INV_X1 U9918 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8828) );
  OR2_X1 U9919 ( .A1(n8576), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8606) );
  AND2_X1 U9920 ( .A1(n8223), .A2(n8202), .ZN(n13814) );
  NAND2_X1 U9921 ( .A1(n10688), .A2(n10685), .ZN(n10877) );
  OR2_X1 U9922 ( .A1(n10558), .A2(n10556), .ZN(n9484) );
  NAND2_X1 U9923 ( .A1(n12605), .A2(n12606), .ZN(n12607) );
  OR2_X1 U9924 ( .A1(n13827), .A2(n8238), .ZN(n8188) );
  INV_X1 U9925 ( .A(n8030), .ZN(n12557) );
  OR2_X1 U9926 ( .A1(n10349), .A2(n10348), .ZN(n10377) );
  INV_X1 U9927 ( .A(n15214), .ZN(n15270) );
  INV_X1 U9928 ( .A(n15265), .ZN(n15268) );
  INV_X1 U9929 ( .A(n12631), .ZN(n11635) );
  INV_X1 U9930 ( .A(n13950), .ZN(n15293) );
  INV_X1 U9931 ( .A(n14077), .ZN(n14059) );
  INV_X1 U9932 ( .A(n15390), .ZN(n14093) );
  AND2_X1 U9933 ( .A1(n11715), .A2(n12666), .ZN(n15399) );
  AND2_X1 U9934 ( .A1(n8316), .A2(n8315), .ZN(n15306) );
  OR3_X1 U9935 ( .A1(n11631), .A2(n14146), .A3(n14147), .ZN(n9475) );
  AND2_X1 U9936 ( .A1(n7873), .A2(n7891), .ZN(n10380) );
  NOR2_X1 U9937 ( .A1(n11294), .A2(n11293), .ZN(n11388) );
  NAND2_X1 U9938 ( .A1(n11468), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11601) );
  AND2_X1 U9939 ( .A1(n14162), .A2(n9775), .ZN(n14950) );
  AND4_X1 U9940 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n12831) );
  INV_X1 U9941 ( .A(n9629), .ZN(n9631) );
  INV_X1 U9942 ( .A(n15036), .ZN(n14383) );
  AND2_X1 U9943 ( .A1(n9631), .A2(n9616), .ZN(n14389) );
  INV_X1 U9944 ( .A(n14422), .ZN(n14526) );
  INV_X1 U9945 ( .A(n14401), .ZN(n14565) );
  NAND2_X1 U9946 ( .A1(n10228), .A2(n10227), .ZN(n14792) );
  INV_X1 U9947 ( .A(n14614), .ZN(n15052) );
  AND2_X1 U9948 ( .A1(n14636), .A2(n11166), .ZN(n15058) );
  NAND2_X1 U9949 ( .A1(n9755), .A2(n9754), .ZN(n10254) );
  INV_X1 U9950 ( .A(n14397), .ZN(n14660) );
  INV_X1 U9951 ( .A(n14792), .ZN(n15128) );
  AND2_X1 U9952 ( .A1(n11018), .A2(n15119), .ZN(n14732) );
  INV_X1 U9953 ( .A(n10254), .ZN(n10470) );
  OR2_X1 U9954 ( .A1(n9568), .A2(n9567), .ZN(n9754) );
  NAND2_X1 U9955 ( .A1(n9040), .A2(n9039), .ZN(n9043) );
  AND2_X1 U9956 ( .A1(n9879), .A2(n9878), .ZN(n15581) );
  INV_X1 U9957 ( .A(n13037), .ZN(n11233) );
  INV_X1 U9958 ( .A(n15429), .ZN(n13040) );
  INV_X1 U9959 ( .A(n13257), .ZN(n13228) );
  OR2_X1 U9960 ( .A1(n9509), .A2(n10161), .ZN(n13044) );
  INV_X1 U9961 ( .A(n15588), .ZN(n15549) );
  INV_X1 U9962 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15466) );
  INV_X1 U9963 ( .A(n14879), .ZN(n15594) );
  NAND2_X1 U9964 ( .A1(n15679), .A2(n15677), .ZN(n13320) );
  AND2_X1 U9965 ( .A1(n11682), .A2(n11681), .ZN(n13387) );
  AOI21_X1 U9966 ( .B1(n8977), .B2(n8986), .A(n8985), .ZN(n8987) );
  NAND2_X1 U9967 ( .A1(n15764), .A2(n15677), .ZN(n13390) );
  INV_X1 U9968 ( .A(n15764), .ZN(n15761) );
  INV_X1 U9969 ( .A(n12930), .ZN(n13400) );
  OR2_X1 U9970 ( .A1(n15742), .A2(n15718), .ZN(n13449) );
  INV_X2 U9971 ( .A(n15742), .ZN(n15740) );
  AND2_X1 U9972 ( .A1(n8976), .A2(n8975), .ZN(n15742) );
  NAND2_X1 U9973 ( .A1(n9548), .A2(n9547), .ZN(n9549) );
  INV_X1 U9974 ( .A(n12171), .ZN(n12176) );
  INV_X1 U9975 ( .A(SI_18_), .ZN(n10082) );
  INV_X1 U9976 ( .A(SI_13_), .ZN(n9564) );
  INV_X1 U9977 ( .A(n10652), .ZN(n15459) );
  NAND2_X1 U9978 ( .A1(n10878), .A2(n10883), .ZN(n11196) );
  NAND2_X1 U9979 ( .A1(n8229), .A2(n8228), .ZN(n13806) );
  INV_X1 U9980 ( .A(n13664), .ZN(n13685) );
  OR2_X1 U9981 ( .A1(n7982), .A2(n7981), .ZN(n13992) );
  NAND2_X1 U9982 ( .A1(n15151), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15265) );
  INV_X1 U9983 ( .A(n15274), .ZN(n15221) );
  INV_X1 U9984 ( .A(n15287), .ZN(n14004) );
  OR2_X1 U9985 ( .A1(n15424), .A2(n15403), .ZN(n14077) );
  OR2_X1 U9986 ( .A1(n8339), .A2(n10556), .ZN(n15424) );
  INV_X2 U9987 ( .A(n15424), .ZN(n15427) );
  AND2_X1 U9988 ( .A1(n14918), .A2(n14917), .ZN(n14922) );
  OR2_X1 U9989 ( .A1(n8339), .A2(n8334), .ZN(n15407) );
  NOR2_X1 U9990 ( .A1(n15306), .A2(n15340), .ZN(n15321) );
  INV_X1 U9991 ( .A(n15343), .ZN(n15340) );
  INV_X1 U9992 ( .A(n7651), .ZN(n11715) );
  INV_X1 U9993 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10393) );
  INV_X1 U9994 ( .A(n14950), .ZN(n14300) );
  INV_X1 U9995 ( .A(n12831), .ZN(n14302) );
  OR2_X1 U9996 ( .A1(n9629), .A2(n12128), .ZN(n15036) );
  INV_X1 U9997 ( .A(n14387), .ZN(n15038) );
  INV_X1 U9998 ( .A(n14343), .ZN(n15042) );
  OR2_X1 U9999 ( .A1(n10255), .A2(n10254), .ZN(n15148) );
  OR3_X1 U10000 ( .A1(n14738), .A2(n14737), .A3(n14736), .ZN(n14752) );
  AND3_X1 U10001 ( .A1(n15104), .A2(n15103), .A3(n15102), .ZN(n15143) );
  AND2_X1 U10002 ( .A1(n9812), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9571) );
  INV_X1 U10003 ( .A(n9567), .ZN(n14769) );
  OR2_X1 U10004 ( .A1(n10409), .A2(n10408), .ZN(n11372) );
  INV_X1 U10005 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10080) );
  AND2_X1 U10006 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9744), .ZN(P2_U3947) );
  NOR2_X1 U10007 ( .A1(n9813), .A2(n9454), .ZN(P1_U4016) );
  NOR2_X1 U10008 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7634) );
  NOR2_X1 U10009 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n7636) );
  NOR2_X1 U10010 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n7635) );
  AND3_X2 U10011 ( .A1(n7638), .A2(n7637), .A3(n7681), .ZN(n7761) );
  NAND2_X1 U10012 ( .A1(n7644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7643) );
  INV_X1 U10013 ( .A(n7649), .ZN(n8303) );
  NAND2_X1 U10014 ( .A1(n7645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7646) );
  MUX2_X1 U10015 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7646), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n7647) );
  INV_X1 U10016 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7648) );
  OR2_X1 U10017 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  XNOR2_X1 U10018 ( .A(n7650), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7651) );
  AND2_X1 U10019 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  INV_X1 U10020 ( .A(n7654), .ZN(n7655) );
  NAND2_X1 U10021 ( .A1(n7655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7656) );
  XNOR2_X1 U10022 ( .A(n7656), .B(P2_IR_REG_19__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U10023 ( .A1(n11216), .A2(n12660), .ZN(n15297) );
  INV_X1 U10024 ( .A(n15297), .ZN(n12666) );
  INV_X1 U10025 ( .A(n15399), .ZN(n15359) );
  NOR2_X1 U10026 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n7661) );
  OAI21_X1 U10027 ( .B1(n7675), .B2(n7648), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n7667) );
  INV_X1 U10028 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n12135) );
  XNOR2_X2 U10029 ( .A(n7670), .B(n12135), .ZN(n11724) );
  NAND2_X1 U10030 ( .A1(n7729), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7673) );
  INV_X1 U10031 ( .A(n11724), .ZN(n7671) );
  NAND2_X1 U10032 ( .A1(n7730), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7672) );
  INV_X1 U10033 ( .A(n7675), .ZN(n7676) );
  NAND2_X2 U10034 ( .A1(n7677), .A2(n7676), .ZN(n8293) );
  XNOR2_X2 U10035 ( .A(n7679), .B(n7678), .ZN(n14141) );
  NAND2_X1 U10036 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7680) );
  MUX2_X1 U10037 ( .A(n7680), .B(P2_IR_REG_31__SCAN_IN), .S(n7681), .Z(n7682)
         );
  INV_X1 U10038 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13713) );
  NAND4_X1 U10039 ( .A1(n7685), .A2(n7684), .A3(n7683), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7689) );
  NAND4_X1 U10040 ( .A1(n7687), .A2(n7686), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U10041 ( .A1(n7690), .A2(SI_1_), .ZN(n7711) );
  INV_X1 U10042 ( .A(SI_1_), .ZN(n9526) );
  NAND2_X1 U10043 ( .A1(n7711), .A2(n7691), .ZN(n7713) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n7239), .Z(n7693) );
  NAND2_X1 U10045 ( .A1(n7693), .A2(SI_0_), .ZN(n7712) );
  XNOR2_X1 U10046 ( .A(n7713), .B(n7712), .ZN(n10091) );
  NAND2_X1 U10047 ( .A1(n7729), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U10048 ( .A1(n7730), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U10049 ( .A1(n11804), .A2(SI_0_), .ZN(n7698) );
  XNOR2_X1 U10050 ( .A(n7698), .B(n8344), .ZN(n14153) );
  MUX2_X1 U10051 ( .A(n13713), .B(n14153), .S(n6672), .Z(n15291) );
  NAND2_X1 U10052 ( .A1(n13705), .A2(n12367), .ZN(n12609) );
  INV_X1 U10053 ( .A(n12609), .ZN(n13572) );
  OAI22_X1 U10054 ( .A1(n12612), .A2(n13572), .B1(n12363), .B2(n6854), .ZN(
        n9713) );
  NAND2_X1 U10055 ( .A1(n7729), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U10056 ( .A1(n8203), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U10057 ( .A1(n8030), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7701) );
  NAND2_X1 U10058 ( .A1(n7699), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U10059 ( .A1(n7707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7706) );
  MUX2_X1 U10060 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7706), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n7710) );
  INV_X1 U10061 ( .A(n7707), .ZN(n7709) );
  INV_X1 U10062 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U10063 ( .A1(n7709), .A2(n7708), .ZN(n7724) );
  INV_X1 U10064 ( .A(n15152), .ZN(n9852) );
  AOI22_X1 U10065 ( .A1(n6687), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9740), .B2(
        n9852), .ZN(n7717) );
  MUX2_X1 U10066 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n11804), .Z(n7720) );
  XNOR2_X1 U10067 ( .A(n7721), .B(n7720), .ZN(n10112) );
  NAND2_X1 U10068 ( .A1(n10112), .A2(n12576), .ZN(n7716) );
  INV_X1 U10069 ( .A(n15282), .ZN(n10538) );
  NAND2_X1 U10070 ( .A1(n6878), .A2(n10538), .ZN(n7718) );
  NAND2_X1 U10071 ( .A1(n7719), .A2(n7718), .ZN(n10862) );
  NAND2_X1 U10072 ( .A1(n7722), .A2(SI_3_), .ZN(n7740) );
  OAI21_X1 U10073 ( .B1(n7722), .B2(SI_3_), .A(n7740), .ZN(n7737) );
  XNOR2_X1 U10074 ( .A(n7739), .B(n7737), .ZN(n10263) );
  NAND2_X1 U10075 ( .A1(n10263), .A2(n12576), .ZN(n7727) );
  NAND2_X1 U10076 ( .A1(n7724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7723) );
  MUX2_X1 U10077 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7723), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7725) );
  OR2_X1 U10078 ( .A1(n7724), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7743) );
  AOI22_X1 U10079 ( .A1(n7760), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9740), .B2(
        n9853), .ZN(n7726) );
  INV_X1 U10080 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U10081 ( .A1(n8204), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U10082 ( .A1(n8030), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U10083 ( .A1(n12554), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10084 ( .A1(n10862), .A2(n12613), .ZN(n7736) );
  INV_X1 U10085 ( .A(n13702), .ZN(n12390) );
  NAND2_X1 U10086 ( .A1(n12390), .A2(n15363), .ZN(n7735) );
  NAND2_X1 U10087 ( .A1(n7736), .A2(n7735), .ZN(n10735) );
  INV_X1 U10088 ( .A(n7737), .ZN(n7738) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7239), .Z(n7742) );
  NAND2_X1 U10090 ( .A1(n7742), .A2(SI_4_), .ZN(n7758) );
  OAI21_X1 U10091 ( .B1(n7742), .B2(SI_4_), .A(n7758), .ZN(n7755) );
  XNOR2_X1 U10092 ( .A(n7757), .B(n7755), .ZN(n10420) );
  NAND2_X1 U10093 ( .A1(n10420), .A2(n12576), .ZN(n7746) );
  NAND2_X1 U10094 ( .A1(n7743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7744) );
  XNOR2_X1 U10095 ( .A(n7744), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U10096 ( .A1(n7760), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9740), .B2(
        n9854), .ZN(n7745) );
  NAND2_X1 U10097 ( .A1(n7746), .A2(n7745), .ZN(n12401) );
  NAND2_X1 U10098 ( .A1(n8204), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10099 ( .A1(n8030), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7752) );
  INV_X1 U10100 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10101 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  NAND2_X1 U10102 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7769) );
  AND2_X1 U10103 ( .A1(n7749), .A2(n7769), .ZN(n10742) );
  NAND2_X1 U10104 ( .A1(n8203), .A2(n10742), .ZN(n7751) );
  NAND2_X1 U10105 ( .A1(n12554), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7750) );
  XNOR2_X1 U10106 ( .A(n12401), .B(n13701), .ZN(n12615) );
  INV_X1 U10107 ( .A(n12615), .ZN(n10737) );
  OR2_X1 U10108 ( .A1(n13701), .A2(n12401), .ZN(n7754) );
  INV_X1 U10109 ( .A(n7755), .ZN(n7756) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n11804), .Z(n7759) );
  NAND2_X1 U10111 ( .A1(n7759), .A2(SI_5_), .ZN(n7780) );
  OAI21_X1 U10112 ( .B1(n7759), .B2(SI_5_), .A(n7780), .ZN(n7777) );
  XNOR2_X1 U10113 ( .A(n7779), .B(n7777), .ZN(n10580) );
  NAND2_X1 U10114 ( .A1(n10580), .A2(n12576), .ZN(n7766) );
  NOR2_X1 U10115 ( .A1(n7910), .A2(n7648), .ZN(n7762) );
  MUX2_X1 U10116 ( .A(n7648), .B(n7762), .S(P2_IR_REG_5__SCAN_IN), .Z(n7764)
         );
  AND2_X1 U10117 ( .A1(n7910), .A2(n7763), .ZN(n7788) );
  NOR2_X1 U10118 ( .A1(n7764), .A2(n7788), .ZN(n9855) );
  AOI22_X1 U10119 ( .A1(n7760), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9740), .B2(
        n9855), .ZN(n7765) );
  NAND2_X1 U10120 ( .A1(n7766), .A2(n7765), .ZN(n15377) );
  NAND2_X1 U10121 ( .A1(n12554), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10122 ( .A1(n8204), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7773) );
  INV_X1 U10123 ( .A(n7769), .ZN(n7767) );
  NAND2_X1 U10124 ( .A1(n7767), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7794) );
  INV_X1 U10125 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U10126 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  AND2_X1 U10127 ( .A1(n7794), .A2(n7770), .ZN(n10856) );
  NAND2_X1 U10128 ( .A1(n8203), .A2(n10856), .ZN(n7772) );
  NAND2_X1 U10129 ( .A1(n8030), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7771) );
  NAND4_X1 U10130 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .ZN(n13700) );
  NOR2_X1 U10131 ( .A1(n15377), .A2(n13700), .ZN(n7775) );
  NAND2_X1 U10132 ( .A1(n15377), .A2(n13700), .ZN(n7776) );
  INV_X1 U10133 ( .A(n7777), .ZN(n7778) );
  NAND2_X1 U10134 ( .A1(n7782), .A2(SI_6_), .ZN(n7802) );
  INV_X1 U10135 ( .A(n7782), .ZN(n7783) );
  INV_X1 U10136 ( .A(SI_6_), .ZN(n9538) );
  NAND2_X1 U10137 ( .A1(n7783), .A2(n9538), .ZN(n7784) );
  OR2_X1 U10138 ( .A1(n7786), .A2(n7785), .ZN(n7787) );
  AND2_X1 U10139 ( .A1(n7803), .A2(n7787), .ZN(n10712) );
  NAND2_X1 U10140 ( .A1(n10712), .A2(n12576), .ZN(n7791) );
  INV_X1 U10141 ( .A(n7788), .ZN(n7805) );
  NAND2_X1 U10142 ( .A1(n7805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7789) );
  XNOR2_X1 U10143 ( .A(n7789), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U10144 ( .A1(n7760), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9740), .B2(
        n9922), .ZN(n7790) );
  NAND2_X1 U10145 ( .A1(n12554), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10146 ( .A1(n8204), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7798) );
  INV_X1 U10147 ( .A(n7794), .ZN(n7792) );
  NAND2_X1 U10148 ( .A1(n7792), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7811) );
  INV_X1 U10149 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U10150 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  AND2_X1 U10151 ( .A1(n7811), .A2(n7795), .ZN(n10775) );
  NAND2_X1 U10152 ( .A1(n8203), .A2(n10775), .ZN(n7797) );
  NAND2_X1 U10153 ( .A1(n8030), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7796) );
  NAND4_X1 U10154 ( .A1(n7799), .A2(n7798), .A3(n7797), .A4(n7796), .ZN(n13699) );
  XNOR2_X1 U10155 ( .A(n12411), .B(n13699), .ZN(n12618) );
  INV_X1 U10156 ( .A(n12618), .ZN(n10326) );
  NAND2_X1 U10157 ( .A1(n10322), .A2(n10326), .ZN(n7801) );
  NAND2_X1 U10158 ( .A1(n12411), .A2(n13699), .ZN(n7800) );
  NAND2_X1 U10159 ( .A1(n7804), .A2(SI_7_), .ZN(n7821) );
  OAI21_X1 U10160 ( .B1(n7804), .B2(SI_7_), .A(n7821), .ZN(n7818) );
  NAND2_X1 U10161 ( .A1(n10904), .A2(n12576), .ZN(n7808) );
  NAND2_X1 U10162 ( .A1(n7823), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7806) );
  XNOR2_X1 U10163 ( .A(n7806), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9924) );
  AOI22_X1 U10164 ( .A1(n7760), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9740), .B2(
        n9924), .ZN(n7807) );
  NAND2_X1 U10165 ( .A1(n7808), .A2(n7807), .ZN(n12424) );
  NAND2_X1 U10166 ( .A1(n8204), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10167 ( .A1(n12554), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U10168 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  AND2_X1 U10169 ( .A1(n7830), .A2(n7812), .ZN(n10807) );
  NAND2_X1 U10170 ( .A1(n8203), .A2(n10807), .ZN(n7814) );
  NAND2_X1 U10171 ( .A1(n8030), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7813) );
  NAND4_X1 U10172 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n13698) );
  INV_X1 U10173 ( .A(n13698), .ZN(n8260) );
  XNOR2_X1 U10174 ( .A(n12424), .B(n8260), .ZN(n12620) );
  NAND2_X1 U10175 ( .A1(n12424), .A2(n13698), .ZN(n7817) );
  INV_X1 U10176 ( .A(n7818), .ZN(n7819) );
  MUX2_X1 U10177 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11804), .Z(n7822) );
  NAND2_X1 U10178 ( .A1(n7822), .A2(SI_8_), .ZN(n7840) );
  OAI21_X1 U10179 ( .B1(SI_8_), .B2(n7822), .A(n7840), .ZN(n7837) );
  XNOR2_X1 U10180 ( .A(n7839), .B(n7837), .ZN(n10909) );
  NAND2_X1 U10181 ( .A1(n10909), .A2(n12576), .ZN(n7828) );
  INV_X1 U10182 ( .A(n7823), .ZN(n7825) );
  INV_X1 U10183 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10184 ( .A1(n7825), .A2(n7824), .ZN(n7847) );
  NAND2_X1 U10185 ( .A1(n7847), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7826) );
  XNOR2_X1 U10186 ( .A(n7826), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U10187 ( .A1(n7760), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9740), .B2(
        n9925), .ZN(n7827) );
  NAND2_X1 U10188 ( .A1(n7828), .A2(n7827), .ZN(n12428) );
  NAND2_X1 U10189 ( .A1(n8204), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10190 ( .A1(n8030), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10191 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U10192 ( .A1(n7855), .A2(n7831), .ZN(n10756) );
  INV_X1 U10193 ( .A(n10756), .ZN(n10693) );
  NAND2_X1 U10194 ( .A1(n8203), .A2(n10693), .ZN(n7833) );
  NAND2_X1 U10195 ( .A1(n12554), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7832) );
  NAND4_X1 U10196 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n13697) );
  INV_X1 U10197 ( .A(n13697), .ZN(n12430) );
  NAND2_X1 U10198 ( .A1(n12428), .A2(n12430), .ZN(n8261) );
  OR2_X1 U10199 ( .A1(n12428), .A2(n12430), .ZN(n7836) );
  NAND2_X1 U10200 ( .A1(n8261), .A2(n7836), .ZN(n12621) );
  INV_X1 U10201 ( .A(n7837), .ZN(n7838) );
  NAND2_X1 U10202 ( .A1(n7842), .A2(SI_9_), .ZN(n7864) );
  OAI21_X1 U10203 ( .B1(n7842), .B2(SI_9_), .A(n7864), .ZN(n7843) );
  INV_X1 U10204 ( .A(n7843), .ZN(n7844) );
  OR2_X1 U10205 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  NAND2_X1 U10206 ( .A1(n7865), .A2(n7846), .ZN(n10919) );
  INV_X1 U10207 ( .A(n7847), .ZN(n7849) );
  INV_X1 U10208 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10209 ( .A1(n7849), .A2(n7848), .ZN(n7867) );
  NAND2_X1 U10210 ( .A1(n7867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7850) );
  XNOR2_X1 U10211 ( .A(n7850), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U10212 ( .A1(n7760), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9740), .B2(
        n10353), .ZN(n7851) );
  NAND2_X1 U10213 ( .A1(n12554), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10214 ( .A1(n8204), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10215 ( .A1(n7855), .A2(n7854), .ZN(n7856) );
  AND2_X1 U10216 ( .A1(n7878), .A2(n7856), .ZN(n10879) );
  NAND2_X1 U10217 ( .A1(n8203), .A2(n10879), .ZN(n7858) );
  NAND2_X1 U10218 ( .A1(n8030), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7857) );
  NAND4_X1 U10219 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n13695) );
  INV_X1 U10220 ( .A(n13695), .ZN(n11329) );
  NAND2_X1 U10221 ( .A1(n12441), .A2(n11329), .ZN(n8262) );
  OR2_X1 U10222 ( .A1(n12441), .A2(n11329), .ZN(n7861) );
  NAND2_X1 U10223 ( .A1(n8262), .A2(n7861), .ZN(n12622) );
  NAND2_X1 U10224 ( .A1(n10555), .A2(n12622), .ZN(n7863) );
  NAND2_X1 U10225 ( .A1(n12441), .A2(n13695), .ZN(n7862) );
  XNOR2_X1 U10226 ( .A(n7889), .B(n7391), .ZN(n10933) );
  NAND2_X1 U10227 ( .A1(n10933), .A2(n12576), .ZN(n7875) );
  INV_X1 U10228 ( .A(n7867), .ZN(n7869) );
  INV_X1 U10229 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7868) );
  AOI21_X1 U10230 ( .B1(n7869), .B2(n7868), .A(n7648), .ZN(n7870) );
  NAND2_X1 U10231 ( .A1(n7870), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7873) );
  INV_X1 U10232 ( .A(n7870), .ZN(n7872) );
  INV_X1 U10233 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10234 ( .A1(n7872), .A2(n7871), .ZN(n7891) );
  AOI22_X1 U10235 ( .A1(n7760), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9740), 
        .B2(n10380), .ZN(n7874) );
  NAND2_X1 U10236 ( .A1(n12554), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10237 ( .A1(n8204), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7882) );
  INV_X1 U10238 ( .A(n7878), .ZN(n7876) );
  INV_X1 U10239 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10240 ( .A1(n7878), .A2(n7877), .ZN(n7879) );
  AND2_X1 U10241 ( .A1(n7896), .A2(n7879), .ZN(n11326) );
  NAND2_X1 U10242 ( .A1(n8203), .A2(n11326), .ZN(n7881) );
  NAND2_X1 U10243 ( .A1(n8030), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7880) );
  NAND4_X1 U10244 ( .A1(n7883), .A2(n7882), .A3(n7881), .A4(n7880), .ZN(n13694) );
  INV_X1 U10245 ( .A(n13694), .ZN(n12454) );
  NAND2_X1 U10246 ( .A1(n15393), .A2(n12454), .ZN(n8263) );
  OR2_X1 U10247 ( .A1(n15393), .A2(n12454), .ZN(n7884) );
  NAND2_X1 U10248 ( .A1(n10833), .A2(n7588), .ZN(n7886) );
  NAND2_X1 U10249 ( .A1(n15393), .A2(n13694), .ZN(n7885) );
  INV_X1 U10250 ( .A(n7887), .ZN(n7888) );
  MUX2_X1 U10251 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11804), .Z(n7903) );
  XNOR2_X1 U10252 ( .A(n7907), .B(n7906), .ZN(n10948) );
  NAND2_X1 U10253 ( .A1(n10948), .A2(n12576), .ZN(n7894) );
  NAND2_X1 U10254 ( .A1(n7891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7892) );
  XNOR2_X1 U10255 ( .A(n7892), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U10256 ( .A1(n7760), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9740), 
        .B2(n11081), .ZN(n7893) );
  NAND2_X1 U10257 ( .A1(n12554), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10258 ( .A1(n8204), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10259 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  AND2_X1 U10260 ( .A1(n7916), .A2(n7897), .ZN(n11207) );
  NAND2_X1 U10261 ( .A1(n8203), .A2(n11207), .ZN(n7899) );
  NAND2_X1 U10262 ( .A1(n8030), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7898) );
  NAND4_X1 U10263 ( .A1(n7901), .A2(n7900), .A3(n7899), .A4(n7898), .ZN(n13693) );
  AND2_X1 U10264 ( .A1(n12459), .A2(n13693), .ZN(n7902) );
  INV_X1 U10265 ( .A(n7903), .ZN(n7904) );
  NAND2_X1 U10266 ( .A1(n7904), .A2(n9536), .ZN(n7905) );
  XNOR2_X1 U10267 ( .A(n7924), .B(n7923), .ZN(n11270) );
  NAND2_X1 U10268 ( .A1(n11270), .A2(n12576), .ZN(n7913) );
  NAND2_X1 U10269 ( .A1(n7909), .A2(n7910), .ZN(n7930) );
  NAND2_X1 U10270 ( .A1(n7930), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7911) );
  XNOR2_X1 U10271 ( .A(n7911), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15226) );
  AOI22_X1 U10272 ( .A1(n7760), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9740), 
        .B2(n15226), .ZN(n7912) );
  NAND2_X1 U10273 ( .A1(n12554), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10274 ( .A1(n8204), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7920) );
  INV_X1 U10275 ( .A(n7916), .ZN(n7914) );
  INV_X1 U10276 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10277 ( .A1(n7916), .A2(n7915), .ZN(n7917) );
  AND2_X1 U10278 ( .A1(n7934), .A2(n7917), .ZN(n11339) );
  NAND2_X1 U10279 ( .A1(n8203), .A2(n11339), .ZN(n7919) );
  NAND2_X1 U10280 ( .A1(n8030), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7918) );
  NAND4_X1 U10281 ( .A1(n7921), .A2(n7920), .A3(n7919), .A4(n7918), .ZN(n13692) );
  NOR2_X1 U10282 ( .A1(n14912), .A2(n13692), .ZN(n7922) );
  INV_X1 U10283 ( .A(n7925), .ZN(n7926) );
  NAND2_X1 U10284 ( .A1(n7926), .A2(n9541), .ZN(n7927) );
  MUX2_X1 U10285 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n11804), .Z(n7944) );
  XNOR2_X1 U10286 ( .A(n7944), .B(n9564), .ZN(n7929) );
  XNOR2_X1 U10287 ( .A(n6715), .B(n7929), .ZN(n11277) );
  NAND2_X1 U10288 ( .A1(n11277), .A2(n12576), .ZN(n7933) );
  NOR2_X1 U10289 ( .A1(n7930), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7950) );
  OR2_X1 U10290 ( .A1(n7950), .A2(n7648), .ZN(n7931) );
  XNOR2_X1 U10291 ( .A(n7931), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U10292 ( .A1(n7760), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9740), 
        .B2(n15234), .ZN(n7932) );
  NAND2_X1 U10293 ( .A1(n8204), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10294 ( .A1(n7934), .A2(n15232), .ZN(n7935) );
  AND2_X1 U10295 ( .A1(n7956), .A2(n7935), .ZN(n11514) );
  NAND2_X1 U10296 ( .A1(n8203), .A2(n11514), .ZN(n7938) );
  NAND2_X1 U10297 ( .A1(n8030), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U10298 ( .A1(n12554), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7936) );
  NAND4_X1 U10299 ( .A1(n7939), .A2(n7938), .A3(n7937), .A4(n7936), .ZN(n13691) );
  OR2_X1 U10300 ( .A1(n12470), .A2(n13691), .ZN(n7940) );
  NAND2_X1 U10301 ( .A1(n7941), .A2(n7940), .ZN(n11409) );
  INV_X1 U10302 ( .A(n7944), .ZN(n7942) );
  NAND2_X1 U10303 ( .A1(n7944), .A2(SI_13_), .ZN(n7946) );
  NAND2_X1 U10304 ( .A1(n7966), .A2(n7965), .ZN(n7948) );
  MUX2_X1 U10305 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n11804), .Z(n7963) );
  XNOR2_X1 U10306 ( .A(n7948), .B(n7963), .ZN(n11384) );
  NAND2_X1 U10307 ( .A1(n11384), .A2(n12576), .ZN(n7953) );
  INV_X1 U10308 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10309 ( .A1(n7950), .A2(n7949), .ZN(n7971) );
  NAND2_X1 U10310 ( .A1(n7971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7951) );
  XNOR2_X1 U10311 ( .A(n7951), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U10312 ( .A1(n7760), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9740), 
        .B2(n13723), .ZN(n7952) );
  NAND2_X1 U10313 ( .A1(n12554), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10314 ( .A1(n8204), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7960) );
  INV_X1 U10315 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10316 ( .A1(n7956), .A2(n7955), .ZN(n7957) );
  AND2_X1 U10317 ( .A1(n7978), .A2(n7957), .ZN(n11584) );
  NAND2_X1 U10318 ( .A1(n8203), .A2(n11584), .ZN(n7959) );
  NAND2_X1 U10319 ( .A1(n8030), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7958) );
  NAND4_X1 U10320 ( .A1(n7961), .A2(n7960), .A3(n7959), .A4(n7958), .ZN(n13690) );
  INV_X1 U10321 ( .A(n13690), .ZN(n11671) );
  XNOR2_X1 U10322 ( .A(n12483), .B(n11671), .ZN(n12629) );
  NAND2_X1 U10323 ( .A1(n12483), .A2(n13690), .ZN(n7962) );
  INV_X1 U10324 ( .A(n7963), .ZN(n7964) );
  NAND2_X1 U10325 ( .A1(n7965), .A2(n7964), .ZN(n7967) );
  NAND2_X1 U10326 ( .A1(n7967), .A2(n7966), .ZN(n7984) );
  MUX2_X1 U10327 ( .A(n10391), .B(n10393), .S(n11804), .Z(n7968) );
  INV_X1 U10328 ( .A(n7968), .ZN(n7969) );
  NAND2_X1 U10329 ( .A1(n7969), .A2(SI_15_), .ZN(n7970) );
  XNOR2_X1 U10330 ( .A(n7984), .B(n6796), .ZN(n11454) );
  NAND2_X1 U10331 ( .A1(n11454), .A2(n12576), .ZN(n7974) );
  OAI21_X1 U10332 ( .B1(n7971), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7972) );
  XNOR2_X1 U10333 ( .A(n7972), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U10334 ( .A1(n7760), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9740), 
        .B2(n15244), .ZN(n7973) );
  INV_X1 U10335 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7976) );
  INV_X1 U10336 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7975) );
  OAI22_X1 U10337 ( .A1(n7809), .A2(n7976), .B1(n7853), .B2(n7975), .ZN(n7982)
         );
  INV_X1 U10338 ( .A(n7978), .ZN(n7977) );
  INV_X1 U10339 ( .A(n7995), .ZN(n7997) );
  INV_X1 U10340 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11670) );
  NAND2_X1 U10341 ( .A1(n7978), .A2(n11670), .ZN(n7979) );
  NAND2_X1 U10342 ( .A1(n7997), .A2(n7979), .ZN(n11672) );
  INV_X1 U10343 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7980) );
  OAI22_X1 U10344 ( .A1(n11672), .A2(n8238), .B1(n12557), .B2(n7980), .ZN(
        n7981) );
  XNOR2_X1 U10345 ( .A(n14089), .B(n13605), .ZN(n12631) );
  OR2_X1 U10346 ( .A1(n14089), .A2(n13992), .ZN(n7983) );
  NAND2_X1 U10347 ( .A1(n11632), .A2(n7983), .ZN(n14001) );
  NAND2_X1 U10348 ( .A1(n7984), .A2(n6796), .ZN(n7986) );
  INV_X1 U10349 ( .A(n7987), .ZN(n7988) );
  NAND2_X1 U10350 ( .A1(n7988), .A2(SI_16_), .ZN(n7989) );
  XNOR2_X1 U10351 ( .A(n8003), .B(n7626), .ZN(n11596) );
  NAND2_X1 U10352 ( .A1(n11596), .A2(n12576), .ZN(n7994) );
  NAND2_X1 U10353 ( .A1(n7990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7991) );
  XNOR2_X1 U10354 ( .A(n7991), .B(n7640), .ZN(n15264) );
  INV_X1 U10355 ( .A(n15264), .ZN(n7992) );
  AOI22_X1 U10356 ( .A1(n7760), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9740), 
        .B2(n7992), .ZN(n7993) );
  INV_X1 U10357 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8001) );
  INV_X1 U10358 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10359 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  NAND2_X1 U10360 ( .A1(n8014), .A2(n7998), .ZN(n13995) );
  OR2_X1 U10361 ( .A1(n13995), .A2(n8238), .ZN(n8000) );
  AOI22_X1 U10362 ( .A1(n12554), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8204), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n7999) );
  OAI211_X1 U10363 ( .C1(n12557), .C2(n8001), .A(n8000), .B(n7999), .ZN(n13689) );
  INV_X1 U10364 ( .A(n13689), .ZN(n13615) );
  XNOR2_X1 U10365 ( .A(n14084), .B(n13615), .ZN(n13986) );
  INV_X1 U10366 ( .A(n13986), .ZN(n14000) );
  NAND2_X1 U10367 ( .A1(n14084), .A2(n13689), .ZN(n8002) );
  NAND2_X1 U10368 ( .A1(n14003), .A2(n8002), .ZN(n13980) );
  XNOR2_X1 U10369 ( .A(n8020), .B(n9840), .ZN(n8005) );
  XNOR2_X1 U10370 ( .A(n8022), .B(n8005), .ZN(n11851) );
  NAND2_X1 U10371 ( .A1(n11851), .A2(n12576), .ZN(n8011) );
  NAND2_X1 U10372 ( .A1(n8006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8007) );
  MUX2_X1 U10373 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8007), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8009) );
  NAND2_X1 U10374 ( .A1(n8009), .A2(n8008), .ZN(n13739) );
  INV_X1 U10375 ( .A(n13739), .ZN(n15267) );
  AOI22_X1 U10376 ( .A1(n7760), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9740), 
        .B2(n15267), .ZN(n8010) );
  INV_X1 U10377 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8018) );
  INV_X1 U10378 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10379 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  NAND2_X1 U10380 ( .A1(n8028), .A2(n8015), .ZN(n13975) );
  OR2_X1 U10381 ( .A1(n13975), .A2(n8238), .ZN(n8017) );
  AOI22_X1 U10382 ( .A1(n12554), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8204), 
        .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n8016) );
  OAI211_X1 U10383 ( .C1(n12557), .C2(n8018), .A(n8017), .B(n8016), .ZN(n13989) );
  INV_X1 U10384 ( .A(n13989), .ZN(n13952) );
  XNOR2_X1 U10385 ( .A(n14079), .B(n13952), .ZN(n13979) );
  NAND2_X1 U10386 ( .A1(n13980), .A2(n13979), .ZN(n13982) );
  NAND2_X1 U10387 ( .A1(n14079), .A2(n13989), .ZN(n8019) );
  INV_X1 U10388 ( .A(n8020), .ZN(n8021) );
  NAND2_X1 U10389 ( .A1(n8056), .A2(n10082), .ZN(n8023) );
  MUX2_X1 U10390 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n11804), .Z(n8050) );
  NAND2_X1 U10391 ( .A1(n11840), .A2(n12576), .ZN(n8026) );
  NAND2_X1 U10392 ( .A1(n8008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8024) );
  XNOR2_X1 U10393 ( .A(n8024), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U10394 ( .A1(n7760), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9740), 
        .B2(n13750), .ZN(n8025) );
  INV_X1 U10395 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U10396 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  NAND2_X1 U10397 ( .A1(n8043), .A2(n8029), .ZN(n13962) );
  OR2_X1 U10398 ( .A1(n13962), .A2(n8238), .ZN(n8035) );
  INV_X1 U10399 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14075) );
  NAND2_X1 U10400 ( .A1(n12554), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10401 ( .A1(n8030), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8031) );
  OAI211_X1 U10402 ( .C1(n7853), .C2(n14075), .A(n8032), .B(n8031), .ZN(n8033)
         );
  INV_X1 U10403 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U10404 ( .A1(n8035), .A2(n8034), .ZN(n13939) );
  XNOR2_X1 U10405 ( .A(n13961), .B(n13939), .ZN(n13956) );
  OR2_X1 U10406 ( .A1(n13961), .A2(n13939), .ZN(n8036) );
  INV_X1 U10407 ( .A(n8050), .ZN(n8051) );
  OAI21_X1 U10408 ( .B1(n8038), .B2(n8051), .A(n8037), .ZN(n8039) );
  MUX2_X1 U10409 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n11804), .Z(n8057) );
  XNOR2_X1 U10410 ( .A(n8057), .B(SI_19_), .ZN(n8053) );
  XNOR2_X1 U10411 ( .A(n8039), .B(n8053), .ZN(n11831) );
  NAND2_X1 U10412 ( .A1(n11831), .A2(n12576), .ZN(n8041) );
  AOI22_X1 U10413 ( .A1(n7760), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12660), 
        .B2(n9740), .ZN(n8040) );
  INV_X1 U10414 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10415 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  NAND2_X1 U10416 ( .A1(n8064), .A2(n8044), .ZN(n13935) );
  INV_X1 U10417 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13936) );
  NAND2_X1 U10418 ( .A1(n8030), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10419 ( .A1(n8204), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8045) );
  OAI211_X1 U10420 ( .C1(n7809), .C2(n13936), .A(n8046), .B(n8045), .ZN(n8047)
         );
  INV_X1 U10421 ( .A(n8047), .ZN(n8048) );
  OAI21_X1 U10422 ( .B1(n13935), .B2(n8238), .A(n8048), .ZN(n13920) );
  NOR2_X1 U10423 ( .A1(n13934), .A2(n13920), .ZN(n8049) );
  INV_X1 U10424 ( .A(n13920), .ZN(n13954) );
  NOR2_X1 U10425 ( .A1(n8051), .A2(n10082), .ZN(n8052) );
  NOR2_X1 U10426 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  OAI21_X1 U10427 ( .B1(n8056), .B2(n8055), .A(n8054), .ZN(n8060) );
  INV_X1 U10428 ( .A(n8057), .ZN(n8058) );
  NAND2_X1 U10429 ( .A1(n8058), .A2(n10156), .ZN(n8059) );
  INV_X1 U10430 ( .A(SI_20_), .ZN(n10345) );
  OR2_X1 U10431 ( .A1(n8080), .A2(n10345), .ZN(n8075) );
  NAND2_X1 U10432 ( .A1(n8080), .A2(n10345), .ZN(n8061) );
  MUX2_X1 U10433 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n11804), .Z(n8082) );
  NAND2_X1 U10434 ( .A1(n11878), .A2(n12576), .ZN(n8063) );
  NAND2_X1 U10435 ( .A1(n7760), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8062) );
  INV_X1 U10436 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U10437 ( .A1(n8064), .A2(n13629), .ZN(n8065) );
  AND2_X1 U10438 ( .A1(n8091), .A2(n8065), .ZN(n13924) );
  NAND2_X1 U10439 ( .A1(n13924), .A2(n8203), .ZN(n8071) );
  INV_X1 U10440 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10441 ( .A1(n12554), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10442 ( .A1(n8204), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8066) );
  OAI211_X1 U10443 ( .C1(n8068), .C2(n12557), .A(n8067), .B(n8066), .ZN(n8069)
         );
  INV_X1 U10444 ( .A(n8069), .ZN(n8070) );
  NAND2_X1 U10445 ( .A1(n8071), .A2(n8070), .ZN(n13940) );
  XNOR2_X1 U10446 ( .A(n14063), .B(n13940), .ZN(n13917) );
  INV_X1 U10447 ( .A(n13917), .ZN(n13914) );
  NAND2_X1 U10448 ( .A1(n14063), .A2(n13940), .ZN(n8072) );
  INV_X1 U10449 ( .A(n8082), .ZN(n8077) );
  MUX2_X1 U10450 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11804), .Z(n8074) );
  NAND2_X1 U10451 ( .A1(n8074), .A2(SI_21_), .ZN(n8102) );
  OAI21_X1 U10452 ( .B1(SI_21_), .B2(n8074), .A(n8102), .ZN(n8081) );
  AND2_X1 U10453 ( .A1(n8075), .A2(n8081), .ZN(n8076) );
  OAI21_X1 U10454 ( .B1(n8078), .B2(n8077), .A(n8076), .ZN(n8086) );
  NAND2_X1 U10455 ( .A1(n8082), .A2(SI_20_), .ZN(n8079) );
  INV_X1 U10456 ( .A(n8081), .ZN(n8083) );
  NAND2_X1 U10457 ( .A1(n8086), .A2(n8103), .ZN(n11818) );
  NAND2_X1 U10458 ( .A1(n7760), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8087) );
  INV_X1 U10459 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10460 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  NAND2_X1 U10461 ( .A1(n8111), .A2(n8092), .ZN(n13902) );
  OR2_X1 U10462 ( .A1(n13902), .A2(n8238), .ZN(n8098) );
  INV_X1 U10463 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U10464 ( .A1(n8204), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10465 ( .A1(n12554), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8093) );
  OAI211_X1 U10466 ( .C1(n12557), .C2(n8095), .A(n8094), .B(n8093), .ZN(n8096)
         );
  INV_X1 U10467 ( .A(n8096), .ZN(n8097) );
  NAND2_X1 U10468 ( .A1(n8098), .A2(n8097), .ZN(n13919) );
  AND2_X1 U10469 ( .A1(n14120), .A2(n13919), .ZN(n8099) );
  OR2_X1 U10470 ( .A1(n14120), .A2(n13919), .ZN(n8100) );
  INV_X1 U10471 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8106) );
  MUX2_X1 U10472 ( .A(n8106), .B(n11716), .S(n11804), .Z(n8107) );
  NAND2_X1 U10473 ( .A1(n11805), .A2(n8107), .ZN(n8108) );
  NAND2_X1 U10474 ( .A1(n8120), .A2(n8108), .ZN(n11714) );
  NAND2_X1 U10475 ( .A1(n7760), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8109) );
  INV_X1 U10476 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U10477 ( .A1(n8111), .A2(n13645), .ZN(n8112) );
  AND2_X1 U10478 ( .A1(n8130), .A2(n8112), .ZN(n13893) );
  NAND2_X1 U10479 ( .A1(n13893), .A2(n8203), .ZN(n8118) );
  INV_X1 U10480 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10481 ( .A1(n12554), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10482 ( .A1(n8204), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8113) );
  OAI211_X1 U10483 ( .C1(n8115), .C2(n12557), .A(n8114), .B(n8113), .ZN(n8116)
         );
  INV_X1 U10484 ( .A(n8116), .ZN(n8117) );
  NAND2_X1 U10485 ( .A1(n8118), .A2(n8117), .ZN(n13688) );
  INV_X1 U10486 ( .A(n13688), .ZN(n13534) );
  XNOR2_X1 U10487 ( .A(n14118), .B(n13534), .ZN(n13881) );
  MUX2_X1 U10488 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11804), .Z(n8121) );
  NAND2_X1 U10489 ( .A1(n8121), .A2(SI_23_), .ZN(n8139) );
  OAI21_X1 U10490 ( .B1(SI_23_), .B2(n8121), .A(n8139), .ZN(n8122) );
  INV_X1 U10491 ( .A(n8122), .ZN(n8123) );
  OR2_X1 U10492 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U10493 ( .A1(n7760), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8126) );
  INV_X1 U10494 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U10495 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  NAND2_X1 U10496 ( .A1(n8149), .A2(n8131), .ZN(n13874) );
  OR2_X1 U10497 ( .A1(n13874), .A2(n8238), .ZN(n8137) );
  INV_X1 U10498 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10499 ( .A1(n12554), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10500 ( .A1(n8204), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8132) );
  OAI211_X1 U10501 ( .C1(n8134), .C2(n12557), .A(n8133), .B(n8132), .ZN(n8135)
         );
  INV_X1 U10502 ( .A(n8135), .ZN(n8136) );
  NAND2_X1 U10503 ( .A1(n8137), .A2(n8136), .ZN(n13687) );
  XNOR2_X1 U10504 ( .A(n14045), .B(n13540), .ZN(n13870) );
  OR2_X1 U10505 ( .A1(n14045), .A2(n13687), .ZN(n8138) );
  INV_X1 U10506 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11791) );
  INV_X1 U10507 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11630) );
  MUX2_X1 U10508 ( .A(n11791), .B(n11630), .S(n11804), .Z(n8144) );
  NAND2_X1 U10509 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  NAND2_X1 U10510 ( .A1(n7760), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8147) );
  INV_X1 U10511 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U10512 ( .A1(n8149), .A2(n13625), .ZN(n8150) );
  AND2_X1 U10513 ( .A1(n8162), .A2(n8150), .ZN(n13856) );
  NAND2_X1 U10514 ( .A1(n13856), .A2(n8203), .ZN(n8156) );
  INV_X1 U10515 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10516 ( .A1(n8204), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10517 ( .A1(n12554), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8151) );
  OAI211_X1 U10518 ( .C1(n12557), .C2(n8153), .A(n8152), .B(n8151), .ZN(n8154)
         );
  INV_X1 U10519 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10520 ( .A1(n8156), .A2(n8155), .ZN(n13686) );
  INV_X1 U10521 ( .A(n13686), .ZN(n13592) );
  XNOR2_X1 U10522 ( .A(n14039), .B(n13592), .ZN(n13860) );
  NAND2_X1 U10523 ( .A1(n14039), .A2(n13686), .ZN(n8157) );
  MUX2_X1 U10524 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n11804), .Z(n8173) );
  XNOR2_X1 U10525 ( .A(n8173), .B(SI_25_), .ZN(n8171) );
  XNOR2_X1 U10526 ( .A(n8172), .B(n8171), .ZN(n12836) );
  NAND2_X1 U10527 ( .A1(n12836), .A2(n12576), .ZN(n8161) );
  NAND2_X1 U10528 ( .A1(n7760), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8160) );
  INV_X1 U10529 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13599) );
  NAND2_X1 U10530 ( .A1(n8162), .A2(n13599), .ZN(n8163) );
  AND2_X1 U10531 ( .A1(n8181), .A2(n8163), .ZN(n13840) );
  NAND2_X1 U10532 ( .A1(n13840), .A2(n8203), .ZN(n8169) );
  INV_X1 U10533 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10534 ( .A1(n8204), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10535 ( .A1(n12554), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8164) );
  OAI211_X1 U10536 ( .C1(n12557), .C2(n8166), .A(n8165), .B(n8164), .ZN(n8167)
         );
  INV_X1 U10537 ( .A(n8167), .ZN(n8168) );
  XNOR2_X1 U10538 ( .A(n14034), .B(n13664), .ZN(n12638) );
  NAND2_X1 U10539 ( .A1(n13842), .A2(n13664), .ZN(n8170) );
  INV_X1 U10540 ( .A(n8173), .ZN(n8174) );
  INV_X1 U10541 ( .A(SI_25_), .ZN(n11379) );
  NAND2_X1 U10542 ( .A1(n8174), .A2(n11379), .ZN(n8175) );
  INV_X1 U10543 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14770) );
  INV_X1 U10544 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14145) );
  MUX2_X1 U10545 ( .A(n14770), .B(n14145), .S(n11804), .Z(n8191) );
  XNOR2_X1 U10546 ( .A(n8191), .B(SI_26_), .ZN(n8176) );
  XNOR2_X1 U10547 ( .A(n8193), .B(n8176), .ZN(n14144) );
  NAND2_X1 U10548 ( .A1(n14144), .A2(n12576), .ZN(n8178) );
  NAND2_X1 U10549 ( .A1(n7760), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8177) );
  NAND2_X2 U10550 ( .A1(n8178), .A2(n8177), .ZN(n14111) );
  INV_X1 U10551 ( .A(n8181), .ZN(n8179) );
  NAND2_X1 U10552 ( .A1(n8179), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8201) );
  INV_X1 U10553 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10554 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U10555 ( .A1(n8201), .A2(n8182), .ZN(n13827) );
  INV_X1 U10556 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U10557 ( .A1(n8204), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10558 ( .A1(n12554), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8183) );
  OAI211_X1 U10559 ( .C1(n12557), .C2(n8185), .A(n8184), .B(n8183), .ZN(n8186)
         );
  INV_X1 U10560 ( .A(n8186), .ZN(n8187) );
  NAND2_X2 U10561 ( .A1(n8188), .A2(n8187), .ZN(n13684) );
  NOR2_X1 U10562 ( .A1(n14111), .A2(n13684), .ZN(n8190) );
  INV_X1 U10563 ( .A(n14111), .ZN(n8189) );
  INV_X1 U10564 ( .A(n13684), .ZN(n13808) );
  INV_X1 U10565 ( .A(n8191), .ZN(n8194) );
  NOR2_X1 U10566 ( .A1(n8194), .A2(SI_26_), .ZN(n8192) );
  NAND2_X1 U10567 ( .A1(n8194), .A2(SI_26_), .ZN(n8213) );
  NAND2_X1 U10568 ( .A1(n8218), .A2(n8213), .ZN(n8196) );
  MUX2_X1 U10569 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n11804), .Z(n8212) );
  INV_X1 U10570 ( .A(SI_27_), .ZN(n11519) );
  XNOR2_X1 U10571 ( .A(n8212), .B(n11519), .ZN(n8215) );
  INV_X1 U10572 ( .A(n8215), .ZN(n8195) );
  NAND2_X1 U10573 ( .A1(n12133), .A2(n12576), .ZN(n8198) );
  NAND2_X1 U10574 ( .A1(n7760), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8197) );
  NAND2_X2 U10575 ( .A1(n8198), .A2(n8197), .ZN(n14107) );
  INV_X1 U10576 ( .A(n8201), .ZN(n8199) );
  INV_X1 U10577 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10578 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  NAND2_X1 U10579 ( .A1(n13814), .A2(n8203), .ZN(n8210) );
  INV_X1 U10580 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U10581 ( .A1(n12554), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10582 ( .A1(n8204), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8205) );
  OAI211_X1 U10583 ( .C1(n8207), .C2(n12557), .A(n8206), .B(n8205), .ZN(n8208)
         );
  INV_X1 U10584 ( .A(n8208), .ZN(n8209) );
  XNOR2_X1 U10585 ( .A(n14107), .B(n13683), .ZN(n13811) );
  INV_X1 U10586 ( .A(n13811), .ZN(n8211) );
  NAND2_X1 U10587 ( .A1(n8212), .A2(SI_27_), .ZN(n8214) );
  AND2_X1 U10588 ( .A1(n8213), .A2(n8214), .ZN(n8217) );
  INV_X1 U10589 ( .A(n8214), .ZN(n8216) );
  MUX2_X1 U10590 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n11804), .Z(n8231) );
  XNOR2_X1 U10591 ( .A(n8231), .B(SI_28_), .ZN(n8234) );
  NAND2_X1 U10592 ( .A1(n11761), .A2(n12576), .ZN(n8220) );
  NAND2_X1 U10593 ( .A1(n6687), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U10594 ( .A1(n8221), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13778) );
  INV_X1 U10595 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U10596 ( .A1(n8223), .A2(n8222), .ZN(n8224) );
  NAND2_X1 U10597 ( .A1(n13778), .A2(n8224), .ZN(n13787) );
  INV_X1 U10598 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U10599 ( .A1(n12554), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10600 ( .A1(n8204), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8225) );
  OAI211_X1 U10601 ( .C1(n14103), .C2(n12557), .A(n8226), .B(n8225), .ZN(n8227) );
  INV_X1 U10602 ( .A(n8227), .ZN(n8228) );
  OR2_X1 U10603 ( .A1(n13797), .A2(n8300), .ZN(n8290) );
  NAND2_X1 U10604 ( .A1(n13797), .A2(n8300), .ZN(n8230) );
  NAND2_X1 U10605 ( .A1(n8290), .A2(n8230), .ZN(n13800) );
  INV_X1 U10606 ( .A(n13800), .ZN(n13789) );
  INV_X1 U10607 ( .A(n8231), .ZN(n8232) );
  INV_X1 U10608 ( .A(SI_28_), .ZN(n13470) );
  NAND2_X1 U10609 ( .A1(n8232), .A2(n13470), .ZN(n8233) );
  MUX2_X1 U10610 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n11804), .Z(n11719) );
  INV_X1 U10611 ( .A(SI_29_), .ZN(n13465) );
  XNOR2_X1 U10612 ( .A(n11719), .B(n13465), .ZN(n11717) );
  NAND2_X1 U10613 ( .A1(n12681), .A2(n12576), .ZN(n8237) );
  NAND2_X1 U10614 ( .A1(n7760), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8236) );
  OR2_X1 U10615 ( .A1(n13778), .A2(n8238), .ZN(n8243) );
  INV_X1 U10616 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10617 ( .A1(n12554), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10618 ( .A1(n8030), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8239) );
  OAI211_X1 U10619 ( .C1(n8341), .C2(n7853), .A(n8240), .B(n8239), .ZN(n8241)
         );
  INV_X1 U10620 ( .A(n8241), .ZN(n8242) );
  NAND2_X1 U10621 ( .A1(n8243), .A2(n8242), .ZN(n13682) );
  XNOR2_X1 U10622 ( .A(n12559), .B(n13682), .ZN(n12641) );
  XNOR2_X1 U10623 ( .A(n8244), .B(n12641), .ZN(n13784) );
  INV_X1 U10624 ( .A(n14079), .ZN(n13978) );
  INV_X1 U10625 ( .A(n12459), .ZN(n15404) );
  INV_X1 U10626 ( .A(n12428), .ZN(n15385) );
  INV_X1 U10627 ( .A(n12363), .ZN(n8245) );
  NAND2_X1 U10628 ( .A1(n8245), .A2(n15291), .ZN(n10670) );
  NOR2_X1 U10629 ( .A1(n10670), .A2(n15282), .ZN(n10863) );
  NAND2_X1 U10630 ( .A1(n10863), .A2(n15363), .ZN(n10741) );
  OR2_X1 U10631 ( .A1(n10741), .A2(n12401), .ZN(n10852) );
  INV_X1 U10632 ( .A(n12411), .ZN(n10332) );
  NAND2_X1 U10633 ( .A1(n10855), .A2(n10332), .ZN(n10395) );
  NAND2_X1 U10634 ( .A1(n15404), .A2(n11036), .ZN(n11158) );
  NAND2_X1 U10635 ( .A1(n13978), .A2(n13993), .ZN(n13972) );
  INV_X1 U10636 ( .A(n14118), .ZN(n13892) );
  NAND2_X1 U10637 ( .A1(n13906), .A2(n13892), .ZN(n13891) );
  OR2_X2 U10638 ( .A1(n13891), .A2(n14045), .ZN(n13872) );
  NAND2_X1 U10639 ( .A1(n11715), .A2(n12659), .ZN(n15292) );
  INV_X1 U10640 ( .A(n11216), .ZN(n12610) );
  AOI211_X1 U10641 ( .C1(n12559), .C2(n13795), .A(n13922), .B(n13772), .ZN(
        n13777) );
  NOR2_X1 U10642 ( .A1(n13705), .A2(n15291), .ZN(n10673) );
  NAND2_X1 U10643 ( .A1(n12612), .A2(n10673), .ZN(n10672) );
  INV_X1 U10644 ( .A(n6854), .ZN(n15295) );
  NAND2_X1 U10645 ( .A1(n15295), .A2(n12363), .ZN(n8248) );
  NAND2_X1 U10646 ( .A1(n10672), .A2(n8248), .ZN(n9718) );
  NAND2_X1 U10647 ( .A1(n9718), .A2(n12611), .ZN(n8250) );
  NAND2_X1 U10648 ( .A1(n6878), .A2(n15282), .ZN(n8249) );
  NAND2_X1 U10649 ( .A1(n8250), .A2(n8249), .ZN(n10868) );
  INV_X1 U10650 ( .A(n12613), .ZN(n10867) );
  NAND2_X1 U10651 ( .A1(n10868), .A2(n10867), .ZN(n8252) );
  NAND2_X1 U10652 ( .A1(n12390), .A2(n12387), .ZN(n8251) );
  NAND2_X1 U10653 ( .A1(n8252), .A2(n8251), .ZN(n10736) );
  NAND2_X1 U10654 ( .A1(n10736), .A2(n12615), .ZN(n8255) );
  INV_X1 U10655 ( .A(n13701), .ZN(n8253) );
  NAND2_X1 U10656 ( .A1(n12401), .A2(n8253), .ZN(n8254) );
  NAND2_X1 U10657 ( .A1(n8255), .A2(n8254), .ZN(n10849) );
  XNOR2_X1 U10658 ( .A(n15377), .B(n13700), .ZN(n12616) );
  NAND2_X1 U10659 ( .A1(n10849), .A2(n12616), .ZN(n8258) );
  INV_X1 U10660 ( .A(n13700), .ZN(n8256) );
  NAND2_X1 U10661 ( .A1(n15377), .A2(n8256), .ZN(n8257) );
  NAND2_X1 U10662 ( .A1(n8258), .A2(n8257), .ZN(n10325) );
  INV_X1 U10663 ( .A(n13699), .ZN(n12413) );
  NAND2_X1 U10664 ( .A1(n12411), .A2(n12413), .ZN(n8259) );
  INV_X1 U10665 ( .A(n12622), .ZN(n10563) );
  XNOR2_X1 U10666 ( .A(n12459), .B(n13693), .ZN(n12625) );
  INV_X1 U10667 ( .A(n13693), .ZN(n8264) );
  NAND2_X1 U10668 ( .A1(n12459), .A2(n8264), .ZN(n8265) );
  INV_X1 U10669 ( .A(n13692), .ZN(n11151) );
  NAND2_X1 U10670 ( .A1(n12470), .A2(n12472), .ZN(n11235) );
  INV_X1 U10671 ( .A(n11235), .ZN(n8266) );
  OR2_X1 U10672 ( .A1(n12470), .A2(n12472), .ZN(n11236) );
  INV_X1 U10673 ( .A(n12483), .ZN(n14907) );
  NAND2_X1 U10674 ( .A1(n11405), .A2(n14907), .ZN(n8267) );
  NAND2_X1 U10675 ( .A1(n8267), .A2(n11671), .ZN(n8269) );
  OR2_X1 U10676 ( .A1(n11405), .A2(n14907), .ZN(n8268) );
  AND2_X1 U10677 ( .A1(n14089), .A2(n13605), .ZN(n8270) );
  OR2_X1 U10678 ( .A1(n14089), .A2(n13605), .ZN(n8271) );
  OR2_X1 U10679 ( .A1(n14084), .A2(n13615), .ZN(n8272) );
  NAND2_X1 U10680 ( .A1(n14079), .A2(n13952), .ZN(n8273) );
  NAND2_X1 U10681 ( .A1(n8274), .A2(n8273), .ZN(n13949) );
  INV_X1 U10682 ( .A(n13939), .ZN(n8276) );
  AND2_X1 U10683 ( .A1(n13961), .A2(n8276), .ZN(n8275) );
  OR2_X1 U10684 ( .A1(n13961), .A2(n8276), .ZN(n8277) );
  NAND2_X1 U10685 ( .A1(n13934), .A2(n13954), .ZN(n8279) );
  OR2_X1 U10686 ( .A1(n13934), .A2(n13954), .ZN(n8278) );
  NAND2_X1 U10687 ( .A1(n8279), .A2(n8278), .ZN(n12633) );
  INV_X1 U10688 ( .A(n13940), .ZN(n8280) );
  NAND2_X1 U10689 ( .A1(n14063), .A2(n8280), .ZN(n8281) );
  INV_X1 U10690 ( .A(n13919), .ZN(n13632) );
  OR2_X1 U10691 ( .A1(n14120), .A2(n13632), .ZN(n8282) );
  OR2_X1 U10692 ( .A1(n14118), .A2(n13534), .ZN(n8285) );
  INV_X1 U10693 ( .A(n13870), .ZN(n13866) );
  INV_X1 U10694 ( .A(n13860), .ZN(n13850) );
  NAND2_X1 U10695 ( .A1(n14039), .A2(n13592), .ZN(n8286) );
  OR2_X1 U10696 ( .A1(n13842), .A2(n13685), .ZN(n8288) );
  NAND2_X1 U10697 ( .A1(n14111), .A2(n13808), .ZN(n12636) );
  INV_X1 U10698 ( .A(n13683), .ZN(n8289) );
  NAND2_X1 U10699 ( .A1(n13788), .A2(n8290), .ZN(n8291) );
  NAND2_X1 U10700 ( .A1(n7651), .A2(n12660), .ZN(n8292) );
  NAND2_X1 U10701 ( .A1(n12646), .A2(n12610), .ZN(n12650) );
  INV_X1 U10702 ( .A(n8293), .ZN(n8294) );
  AND2_X2 U10703 ( .A1(n9741), .A2(n8294), .ZN(n13991) );
  INV_X1 U10704 ( .A(n13991), .ZN(n13953) );
  AND2_X2 U10705 ( .A1(n9741), .A2(n8293), .ZN(n13988) );
  INV_X1 U10706 ( .A(P2_B_REG_SCAN_IN), .ZN(n8295) );
  OR2_X1 U10707 ( .A1(n14141), .A2(n8295), .ZN(n8296) );
  NAND2_X1 U10708 ( .A1(n13988), .A2(n8296), .ZN(n13768) );
  INV_X1 U10709 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14099) );
  NAND2_X1 U10710 ( .A1(n12554), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10711 ( .A1(n8204), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8297) );
  OAI211_X1 U10712 ( .C1(n12557), .C2(n14099), .A(n8298), .B(n8297), .ZN(
        n13681) );
  INV_X1 U10713 ( .A(n13681), .ZN(n8299) );
  INV_X1 U10714 ( .A(n8301), .ZN(n8302) );
  NAND2_X1 U10715 ( .A1(n8319), .A2(n7658), .ZN(n8304) );
  XNOR2_X1 U10716 ( .A(n11631), .B(P2_B_REG_SCAN_IN), .ZN(n8311) );
  OAI21_X1 U10717 ( .B1(n8008), .B2(n8307), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8308) );
  MUX2_X1 U10718 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8308), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8310) );
  NAND2_X1 U10719 ( .A1(n8310), .A2(n8309), .ZN(n14147) );
  NAND2_X1 U10720 ( .A1(n8311), .A2(n14147), .ZN(n8316) );
  NAND2_X1 U10721 ( .A1(n8309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8312) );
  MUX2_X1 U10722 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8312), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8314) );
  NAND2_X1 U10723 ( .A1(n8314), .A2(n8313), .ZN(n14146) );
  INV_X1 U10724 ( .A(n14146), .ZN(n8315) );
  INV_X1 U10725 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15341) );
  NAND2_X1 U10726 ( .A1(n15306), .A2(n15341), .ZN(n8318) );
  NAND2_X1 U10727 ( .A1(n14147), .A2(n14146), .ZN(n8317) );
  NAND2_X1 U10728 ( .A1(n8318), .A2(n8317), .ZN(n15342) );
  XNOR2_X1 U10729 ( .A(n8319), .B(n7658), .ZN(n9742) );
  AND2_X1 U10730 ( .A1(n9742), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10731 ( .A1(n11216), .A2(n13759), .ZN(n12657) );
  NAND2_X1 U10732 ( .A1(n9741), .A2(n12657), .ZN(n12667) );
  NAND2_X1 U10733 ( .A1(n15399), .A2(n12659), .ZN(n9479) );
  AND3_X1 U10734 ( .A1(n15343), .A2(n12667), .A3(n9479), .ZN(n8331) );
  NOR4_X1 U10735 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8324) );
  NOR4_X1 U10736 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8323) );
  NOR4_X1 U10737 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8322) );
  NOR4_X1 U10738 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8321) );
  NAND4_X1 U10739 ( .A1(n8324), .A2(n8323), .A3(n8322), .A4(n8321), .ZN(n8330)
         );
  NOR2_X1 U10740 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8328) );
  NOR4_X1 U10741 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8327) );
  NOR4_X1 U10742 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8326) );
  NOR4_X1 U10743 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8325) );
  NAND4_X1 U10744 ( .A1(n8328), .A2(n8327), .A3(n8326), .A4(n8325), .ZN(n8329)
         );
  OAI21_X1 U10745 ( .B1(n8330), .B2(n8329), .A(n15306), .ZN(n9469) );
  NAND3_X1 U10746 ( .A1(n15342), .A2(n8331), .A3(n9469), .ZN(n8339) );
  INV_X1 U10747 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10748 ( .A1(n15306), .A2(n8332), .ZN(n8333) );
  NAND2_X1 U10749 ( .A1(n11631), .A2(n14146), .ZN(n15339) );
  INV_X1 U10750 ( .A(n10556), .ZN(n8334) );
  INV_X1 U10751 ( .A(n12657), .ZN(n9482) );
  NAND2_X1 U10752 ( .A1(n8338), .A2(n7618), .ZN(P2_U3496) );
  NAND2_X1 U10753 ( .A1(n12559), .A2(n14059), .ZN(n8342) );
  NAND2_X1 U10754 ( .A1(n8343), .A2(n7617), .ZN(P2_U3528) );
  INV_X1 U10755 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8940) );
  INV_X1 U10756 ( .A(n8463), .ZN(n8345) );
  NAND2_X1 U10757 ( .A1(n9501), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10758 ( .A1(n9488), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10759 ( .A1(n9515), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10760 ( .A1(n9502), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10761 ( .A1(n9508), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10762 ( .A1(n8481), .A2(n8480), .ZN(n8351) );
  NAND2_X1 U10763 ( .A1(n9533), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8352) );
  INV_X1 U10764 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U10765 ( .A1(n9544), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10766 ( .A1(n9558), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U10767 ( .A1(n8529), .A2(n8356), .ZN(n8358) );
  NAND2_X1 U10768 ( .A1(n9550), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U10769 ( .A1(n9562), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10770 ( .A1(n9559), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10771 ( .A1(n8360), .A2(n8359), .ZN(n8539) );
  NAND2_X1 U10772 ( .A1(n9598), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10773 ( .A1(n9600), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10774 ( .A1(n9605), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10775 ( .A1(n9601), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10776 ( .A1(n9643), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10777 ( .A1(n9645), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10778 ( .A1(n9825), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10779 ( .A1(n9739), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10780 ( .A1(n8603), .A2(n8602), .ZN(n8605) );
  NAND2_X1 U10781 ( .A1(n10080), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10782 ( .A1(n10077), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U10783 ( .A1(n10341), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8373) );
  INV_X1 U10784 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U10785 ( .A1(n10337), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10786 ( .A1(n8646), .A2(n8645), .ZN(n8648) );
  NAND2_X1 U10787 ( .A1(n8648), .A2(n8373), .ZN(n8661) );
  NAND2_X1 U10788 ( .A1(n10391), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U10789 ( .A1(n10393), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10790 ( .A1(n8376), .A2(n8374), .ZN(n8660) );
  INV_X1 U10791 ( .A(n8660), .ZN(n8375) );
  NAND2_X1 U10792 ( .A1(n8661), .A2(n8375), .ZN(n8377) );
  NAND2_X1 U10793 ( .A1(n8377), .A2(n8376), .ZN(n8673) );
  NAND2_X1 U10794 ( .A1(n10410), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10795 ( .A1(n10411), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10796 ( .A1(n8673), .A2(n8672), .ZN(n8675) );
  NAND2_X1 U10797 ( .A1(n8675), .A2(n8379), .ZN(n8687) );
  INV_X1 U10798 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10554) );
  NAND2_X1 U10799 ( .A1(n10554), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8381) );
  INV_X1 U10800 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U10801 ( .A1(n10550), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U10802 ( .A1(n8687), .A2(n8686), .ZN(n8689) );
  NAND2_X1 U10803 ( .A1(n8689), .A2(n8381), .ZN(n8704) );
  INV_X1 U10804 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U10805 ( .A1(n11028), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8383) );
  INV_X1 U10806 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U10807 ( .A1(n11024), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10808 ( .A1(n8704), .A2(n8703), .ZN(n8706) );
  INV_X1 U10809 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11168) );
  NAND2_X1 U10810 ( .A1(n11168), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8385) );
  INV_X1 U10811 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U10812 ( .A1(n11165), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8384) );
  INV_X1 U10813 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U10814 ( .A1(n11819), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8390) );
  INV_X1 U10815 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U10816 ( .A1(n11191), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8389) );
  AND2_X1 U10817 ( .A1(n8390), .A2(n8389), .ZN(n8745) );
  XNOR2_X1 U10818 ( .A(n11716), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U10819 ( .A1(n11716), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U10820 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8768) );
  INV_X1 U10821 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8392) );
  INV_X1 U10822 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14151) );
  NAND2_X1 U10823 ( .A1(n14151), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10824 ( .A1(n8792), .A2(n8395), .ZN(n8397) );
  INV_X1 U10825 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12839) );
  NAND2_X1 U10826 ( .A1(n12839), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10827 ( .A1(n8397), .A2(n8396), .ZN(n8805) );
  AND2_X1 U10828 ( .A1(n14770), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10829 ( .A1(n14145), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8399) );
  INV_X1 U10830 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14143) );
  AND2_X1 U10831 ( .A1(n14143), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8401) );
  INV_X1 U10832 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12134) );
  NAND2_X1 U10833 ( .A1(n12134), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8402) );
  INV_X1 U10834 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8944) );
  XNOR2_X1 U10835 ( .A(n8944), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8403) );
  XNOR2_X1 U10836 ( .A(n8943), .B(n8403), .ZN(n13466) );
  NAND2_X1 U10837 ( .A1(n8419), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10838 ( .A1(n13466), .A2(n7160), .ZN(n8422) );
  OR2_X1 U10839 ( .A1(n12152), .A2(n13470), .ZN(n8421) );
  INV_X2 U10840 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10069) );
  INV_X1 U10841 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n8423) );
  OR2_X2 U10842 ( .A1(n8596), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8623) );
  INV_X1 U10843 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8430) );
  OR2_X2 U10844 ( .A1(n8772), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8783) );
  INV_X1 U10845 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8433) );
  INV_X1 U10846 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12943) );
  OR2_X2 U10847 ( .A1(n8807), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8818) );
  INV_X1 U10848 ( .A(n8818), .ZN(n8436) );
  INV_X1 U10849 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U10850 ( .A1(n8820), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10851 ( .A1(n13117), .A2(n8437), .ZN(n13130) );
  NAND2_X1 U10852 ( .A1(n8951), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10853 ( .A1(n8890), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8445) );
  OAI211_X1 U10854 ( .C1(n8955), .C2(n8940), .A(n8446), .B(n8445), .ZN(n8447)
         );
  NAND2_X1 U10855 ( .A1(n12930), .A2(n13041), .ZN(n8964) );
  NAND2_X2 U10856 ( .A1(n8965), .A2(n8964), .ZN(n12922) );
  NAND2_X1 U10857 ( .A1(n8465), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10858 ( .A1(n10766), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10859 ( .A1(n8488), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10860 ( .A1(n8454), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8448) );
  INV_X1 U10861 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U10862 ( .A1(n9776), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10863 ( .A1(n8463), .A2(n8452), .ZN(n8453) );
  MUX2_X1 U10864 ( .A(SI_0_), .B(n8453), .S(n10090), .Z(n13473) );
  MUX2_X1 U10865 ( .A(n13472), .B(n13473), .S(n9868), .Z(n15678) );
  INV_X1 U10866 ( .A(n15678), .ZN(n12170) );
  NAND2_X1 U10867 ( .A1(n8465), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10868 ( .A1(n8488), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10869 ( .A1(n10766), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10870 ( .A1(n8454), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8455) );
  INV_X1 U10871 ( .A(n15674), .ZN(n15431) );
  NAND2_X1 U10872 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8460) );
  INV_X1 U10873 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8459) );
  INV_X1 U10874 ( .A(n8461), .ZN(n8462) );
  XNOR2_X1 U10875 ( .A(n8464), .B(n8463), .ZN(n9527) );
  NAND2_X1 U10876 ( .A1(n15651), .A2(n12180), .ZN(n10179) );
  NAND2_X1 U10877 ( .A1(n10179), .A2(n12179), .ZN(n15635) );
  NAND2_X1 U10878 ( .A1(n8465), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10879 ( .A1(n10766), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10880 ( .A1(n8488), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8466) );
  INV_X1 U10881 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8471) );
  XNOR2_X2 U10882 ( .A(n8472), .B(n8471), .ZN(n9886) );
  INV_X1 U10883 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10884 ( .A1(n8465), .A2(n8475), .ZN(n8479) );
  NAND2_X1 U10885 ( .A1(n10766), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10886 ( .A1(n8488), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U10887 ( .A1(n8454), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8476) );
  OR2_X1 U10888 ( .A1(n12152), .A2(SI_3_), .ZN(n8486) );
  XNOR2_X1 U10889 ( .A(n8481), .B(n8480), .ZN(n9492) );
  OR2_X1 U10890 ( .A1(n8749), .A2(n9492), .ZN(n8485) );
  INV_X1 U10891 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10892 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6719), .ZN(n8482) );
  NAND2_X1 U10893 ( .A1(n8725), .A2(n10062), .ZN(n8484) );
  NAND2_X1 U10894 ( .A1(n15636), .A2(n10366), .ZN(n12190) );
  INV_X1 U10895 ( .A(n15636), .ZN(n10799) );
  NAND2_X1 U10896 ( .A1(n10799), .A2(n15630), .ZN(n12191) );
  NAND2_X1 U10897 ( .A1(n15629), .A2(n15628), .ZN(n8487) );
  NAND2_X1 U10898 ( .A1(n8487), .A2(n12190), .ZN(n10784) );
  NAND2_X1 U10899 ( .A1(n8951), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8494) );
  BUF_X2 U10900 ( .A(n8488), .Z(n8890) );
  NAND2_X1 U10901 ( .A1(n8890), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8493) );
  INV_X1 U10902 ( .A(n8489), .ZN(n8503) );
  NAND2_X1 U10903 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8490) );
  NAND2_X1 U10904 ( .A1(n8503), .A2(n8490), .ZN(n10524) );
  NAND2_X1 U10905 ( .A1(n8465), .A2(n10524), .ZN(n8492) );
  NAND2_X1 U10906 ( .A1(n10766), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8491) );
  OR2_X1 U10907 ( .A1(n12152), .A2(SI_4_), .ZN(n8500) );
  XNOR2_X1 U10908 ( .A(n8496), .B(n8495), .ZN(n9495) );
  OR2_X1 U10909 ( .A1(n8749), .A2(n9495), .ZN(n8499) );
  OR2_X1 U10910 ( .A1(n8512), .A2(n8619), .ZN(n8497) );
  XNOR2_X1 U10911 ( .A(n8497), .B(n8511), .ZN(n15437) );
  NAND2_X1 U10912 ( .A1(n8725), .A2(n15437), .ZN(n8498) );
  NAND2_X1 U10913 ( .A1(n15623), .A2(n10525), .ZN(n12194) );
  INV_X1 U10914 ( .A(n15623), .ZN(n10372) );
  INV_X1 U10915 ( .A(n10525), .ZN(n15703) );
  NAND2_X1 U10916 ( .A1(n10372), .A2(n15703), .ZN(n12195) );
  NAND2_X1 U10917 ( .A1(n12194), .A2(n12195), .ZN(n10783) );
  INV_X1 U10918 ( .A(n10783), .ZN(n12328) );
  NAND2_X1 U10919 ( .A1(n10784), .A2(n12328), .ZN(n8501) );
  NAND2_X1 U10920 ( .A1(n8501), .A2(n12194), .ZN(n15606) );
  NAND2_X1 U10921 ( .A1(n10766), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10922 ( .A1(n8951), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8507) );
  INV_X1 U10923 ( .A(n8502), .ZN(n8521) );
  NAND2_X1 U10924 ( .A1(n8503), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U10925 ( .A1(n8521), .A2(n8504), .ZN(n15618) );
  NAND2_X1 U10926 ( .A1(n8465), .A2(n15618), .ZN(n8506) );
  NAND2_X1 U10927 ( .A1(n8890), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8505) );
  NAND4_X1 U10928 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(n12199) );
  OR2_X1 U10929 ( .A1(n12152), .A2(SI_5_), .ZN(n8518) );
  XNOR2_X1 U10930 ( .A(n8510), .B(n8509), .ZN(n9498) );
  OR2_X1 U10931 ( .A1(n8749), .A2(n9498), .ZN(n8517) );
  NAND2_X1 U10932 ( .A1(n8512), .A2(n8511), .ZN(n8514) );
  NAND2_X1 U10933 ( .A1(n8514), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8513) );
  MUX2_X1 U10934 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8513), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8515) );
  NAND2_X1 U10935 ( .A1(n8515), .A2(n8618), .ZN(n10646) );
  NAND2_X1 U10936 ( .A1(n8725), .A2(n10646), .ZN(n8516) );
  NAND2_X1 U10937 ( .A1(n15606), .A2(n15607), .ZN(n8519) );
  INV_X1 U10938 ( .A(n12199), .ZN(n10826) );
  NAND2_X1 U10939 ( .A1(n10826), .A2(n15617), .ZN(n12168) );
  NAND2_X1 U10940 ( .A1(n8519), .A2(n12168), .ZN(n11002) );
  NAND2_X1 U10941 ( .A1(n8951), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10942 ( .A1(n8890), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8525) );
  INV_X1 U10943 ( .A(n8520), .ZN(n8533) );
  NAND2_X1 U10944 ( .A1(n8521), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10945 ( .A1(n8533), .A2(n8522), .ZN(n10818) );
  NAND2_X1 U10946 ( .A1(n8465), .A2(n10818), .ZN(n8524) );
  NAND2_X1 U10947 ( .A1(n10766), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10948 ( .A1(n8618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8527) );
  OR2_X1 U10949 ( .A1(n12152), .A2(n9538), .ZN(n8531) );
  XNOR2_X1 U10950 ( .A(n9550), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8528) );
  XNOR2_X1 U10951 ( .A(n8529), .B(n8528), .ZN(n9539) );
  OR2_X1 U10952 ( .A1(n8749), .A2(n9539), .ZN(n8530) );
  OAI211_X1 U10953 ( .C1(n9868), .C2(n15459), .A(n8531), .B(n8530), .ZN(n10823) );
  NAND2_X1 U10954 ( .A1(n15611), .A2(n10823), .ZN(n12210) );
  INV_X1 U10955 ( .A(n10823), .ZN(n15712) );
  NAND2_X1 U10956 ( .A1(n11109), .A2(n15712), .ZN(n12205) );
  NAND2_X1 U10957 ( .A1(n11002), .A2(n12326), .ZN(n8532) );
  NAND2_X1 U10958 ( .A1(n8532), .A2(n12210), .ZN(n11043) );
  NAND2_X1 U10959 ( .A1(n8951), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10960 ( .A1(n8890), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10961 ( .A1(n8533), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10962 ( .A1(n8548), .A2(n8534), .ZN(n11049) );
  NAND2_X1 U10963 ( .A1(n8465), .A2(n11049), .ZN(n8536) );
  NAND2_X1 U10964 ( .A1(n10766), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8535) );
  OR2_X1 U10965 ( .A1(n12152), .A2(SI_7_), .ZN(n8546) );
  NAND2_X1 U10966 ( .A1(n8540), .A2(n8539), .ZN(n8541) );
  AND2_X1 U10967 ( .A1(n8542), .A2(n8541), .ZN(n9489) );
  OR2_X1 U10968 ( .A1(n8749), .A2(n9489), .ZN(n8545) );
  OR2_X1 U10969 ( .A1(n8555), .A2(n8619), .ZN(n8543) );
  XNOR2_X1 U10970 ( .A(n8543), .B(n8554), .ZN(n15470) );
  NAND2_X1 U10971 ( .A1(n8725), .A2(n15470), .ZN(n8544) );
  NAND2_X1 U10972 ( .A1(n11228), .A2(n11051), .ZN(n12212) );
  INV_X1 U10973 ( .A(n11051), .ZN(n15717) );
  NAND2_X1 U10974 ( .A1(n15597), .A2(n15717), .ZN(n12213) );
  NAND2_X1 U10975 ( .A1(n12212), .A2(n12213), .ZN(n12207) );
  INV_X1 U10976 ( .A(n12207), .ZN(n12327) );
  NAND2_X1 U10977 ( .A1(n11043), .A2(n12327), .ZN(n8547) );
  NAND2_X1 U10978 ( .A1(n8547), .A2(n12212), .ZN(n15602) );
  NAND2_X1 U10979 ( .A1(n10766), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10980 ( .A1(n8951), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10981 ( .A1(n8548), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10982 ( .A1(n8564), .A2(n8549), .ZN(n15600) );
  NAND2_X1 U10983 ( .A1(n8465), .A2(n15600), .ZN(n8551) );
  NAND2_X1 U10984 ( .A1(n8890), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8550) );
  NAND4_X1 U10985 ( .A1(n8553), .A2(n8552), .A3(n8551), .A4(n8550), .ZN(n12216) );
  NAND2_X1 U10986 ( .A1(n8555), .A2(n8554), .ZN(n8574) );
  NAND2_X1 U10987 ( .A1(n8574), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8556) );
  XNOR2_X1 U10988 ( .A(n8556), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10654) );
  INV_X1 U10989 ( .A(SI_8_), .ZN(n9521) );
  OR2_X1 U10990 ( .A1(n12152), .A2(n9521), .ZN(n8562) );
  OR2_X1 U10991 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NAND2_X1 U10992 ( .A1(n8560), .A2(n8559), .ZN(n9522) );
  OR2_X1 U10993 ( .A1(n8749), .A2(n9522), .ZN(n8561) );
  OAI211_X1 U10994 ( .C1(n9868), .C2(n15487), .A(n8562), .B(n8561), .ZN(n12218) );
  XNOR2_X1 U10995 ( .A(n12216), .B(n12218), .ZN(n15601) );
  INV_X1 U10996 ( .A(n12216), .ZN(n12217) );
  NAND2_X1 U10997 ( .A1(n12217), .A2(n12218), .ZN(n8563) );
  NAND2_X1 U10998 ( .A1(n8951), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10999 ( .A1(n8890), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U11000 ( .A1(n8564), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U11001 ( .A1(n8581), .A2(n8565), .ZN(n11437) );
  NAND2_X1 U11002 ( .A1(n8465), .A2(n11437), .ZN(n8567) );
  NAND2_X1 U11003 ( .A1(n10766), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8566) );
  OR2_X1 U11004 ( .A1(n8571), .A2(n8570), .ZN(n8572) );
  AND2_X1 U11005 ( .A1(n8573), .A2(n8572), .ZN(n9523) );
  OR2_X1 U11006 ( .A1(n8749), .A2(n9523), .ZN(n8580) );
  OR2_X1 U11007 ( .A1(n12152), .A2(SI_9_), .ZN(n8579) );
  NAND2_X1 U11008 ( .A1(n8576), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8575) );
  MUX2_X1 U11009 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8575), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8577) );
  NAND2_X1 U11010 ( .A1(n8577), .A2(n8606), .ZN(n15510) );
  NAND2_X1 U11011 ( .A1(n8725), .A2(n15510), .ZN(n8578) );
  INV_X1 U11012 ( .A(n11434), .ZN(n11252) );
  NOR2_X1 U11013 ( .A1(n15598), .A2(n11252), .ZN(n12223) );
  NAND2_X1 U11014 ( .A1(n15598), .A2(n11252), .ZN(n12225) );
  NAND2_X1 U11015 ( .A1(n10766), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U11016 ( .A1(n8951), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U11017 ( .A1(n8581), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U11018 ( .A1(n8596), .A2(n8582), .ZN(n11540) );
  NAND2_X1 U11019 ( .A1(n8465), .A2(n11540), .ZN(n8584) );
  NAND2_X1 U11020 ( .A1(n8890), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8583) );
  OR2_X1 U11021 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  NAND2_X1 U11022 ( .A1(n8590), .A2(n8589), .ZN(n9519) );
  NAND2_X1 U11023 ( .A1(n7160), .A2(n9519), .ZN(n8595) );
  OR2_X1 U11024 ( .A1(n12152), .A2(SI_10_), .ZN(n8594) );
  NAND2_X1 U11025 ( .A1(n8606), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8592) );
  INV_X1 U11026 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11027 ( .A1(n8725), .A2(n13091), .ZN(n8593) );
  INV_X1 U11028 ( .A(n11541), .ZN(n11447) );
  NAND2_X1 U11029 ( .A1(n11647), .A2(n11447), .ZN(n12230) );
  NAND2_X1 U11030 ( .A1(n11658), .A2(n11541), .ZN(n12229) );
  NAND2_X1 U11031 ( .A1(n8951), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U11032 ( .A1(n10766), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U11033 ( .A1(n8596), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11034 ( .A1(n8623), .A2(n8597), .ZN(n11655) );
  NAND2_X1 U11035 ( .A1(n8465), .A2(n11655), .ZN(n8599) );
  NAND2_X1 U11036 ( .A1(n8890), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8598) );
  OR2_X1 U11037 ( .A1(n8603), .A2(n8602), .ZN(n8604) );
  NAND2_X1 U11038 ( .A1(n8605), .A2(n8604), .ZN(n9537) );
  NAND2_X1 U11039 ( .A1(n9537), .A2(n7160), .ZN(n8610) );
  OAI21_X1 U11040 ( .B1(n8606), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8608) );
  INV_X1 U11041 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U11042 ( .A(n8608), .B(n8607), .ZN(n15528) );
  AOI22_X1 U11043 ( .A1(n8947), .A2(n9536), .B1(n8725), .B2(n15528), .ZN(n8609) );
  NAND2_X1 U11044 ( .A1(n8610), .A2(n8609), .ZN(n11650) );
  INV_X1 U11045 ( .A(n11650), .ZN(n11660) );
  NAND2_X1 U11046 ( .A1(n11696), .A2(n11660), .ZN(n12232) );
  NAND2_X1 U11047 ( .A1(n11688), .A2(n11650), .ZN(n12236) );
  NAND2_X1 U11048 ( .A1(n11558), .A2(n12335), .ZN(n8611) );
  NAND2_X1 U11049 ( .A1(n8611), .A2(n12232), .ZN(n11528) );
  OR2_X1 U11050 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U11051 ( .A1(n8615), .A2(n8614), .ZN(n9540) );
  OR2_X1 U11052 ( .A1(n9540), .A2(n8749), .ZN(n8622) );
  INV_X1 U11053 ( .A(n8616), .ZN(n8617) );
  NOR2_X1 U11054 ( .A1(n8618), .A2(n8617), .ZN(n8634) );
  OR2_X1 U11055 ( .A1(n8634), .A2(n8619), .ZN(n8620) );
  XNOR2_X1 U11056 ( .A(n8620), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U11057 ( .A1(n8947), .A2(SI_12_), .B1(n8725), .B2(n13096), .ZN(
        n8621) );
  NAND2_X1 U11058 ( .A1(n8622), .A2(n8621), .ZN(n11694) );
  NAND2_X1 U11059 ( .A1(n8951), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11060 ( .A1(n10766), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11061 ( .A1(n8623), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11062 ( .A1(n8639), .A2(n8624), .ZN(n11695) );
  NAND2_X1 U11063 ( .A1(n8465), .A2(n11695), .ZN(n8626) );
  NAND2_X1 U11064 ( .A1(n8890), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8625) );
  OR2_X1 U11065 ( .A1(n11694), .A2(n12994), .ZN(n12238) );
  NAND2_X1 U11066 ( .A1(n11694), .A2(n12994), .ZN(n12240) );
  NAND2_X1 U11067 ( .A1(n12238), .A2(n12240), .ZN(n12337) );
  NAND2_X1 U11068 ( .A1(n8630), .A2(n10154), .ZN(n8631) );
  NAND2_X1 U11069 ( .A1(n8632), .A2(n8631), .ZN(n9563) );
  NAND2_X1 U11070 ( .A1(n9563), .A2(n7160), .ZN(n8638) );
  INV_X1 U11071 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U11072 ( .A1(n8634), .A2(n8633), .ZN(n8649) );
  NAND2_X1 U11073 ( .A1(n8649), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8636) );
  INV_X1 U11074 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8635) );
  XNOR2_X1 U11075 ( .A(n8636), .B(n8635), .ZN(n15564) );
  AOI22_X1 U11076 ( .A1(n8947), .A2(n9564), .B1(n8725), .B2(n15564), .ZN(n8637) );
  NAND2_X1 U11077 ( .A1(n8638), .A2(n8637), .ZN(n12995) );
  NAND2_X1 U11078 ( .A1(n8951), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U11079 ( .A1(n8639), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U11080 ( .A1(n8654), .A2(n8640), .ZN(n12998) );
  NAND2_X1 U11081 ( .A1(n8465), .A2(n12998), .ZN(n8643) );
  NAND2_X1 U11082 ( .A1(n8890), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11083 ( .A1(n10766), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8641) );
  NOR2_X1 U11084 ( .A1(n12995), .A2(n12893), .ZN(n12249) );
  NAND2_X1 U11085 ( .A1(n12995), .A2(n12893), .ZN(n11620) );
  OR2_X1 U11086 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  NAND2_X1 U11087 ( .A1(n8648), .A2(n8647), .ZN(n9606) );
  NAND2_X1 U11088 ( .A1(n9606), .A2(n7160), .ZN(n8653) );
  INV_X1 U11089 ( .A(SI_14_), .ZN(n9607) );
  NAND2_X1 U11090 ( .A1(n8662), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8651) );
  INV_X1 U11091 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8650) );
  XNOR2_X1 U11092 ( .A(n8651), .B(n8650), .ZN(n15583) );
  AOI22_X1 U11093 ( .A1(n8947), .A2(n9607), .B1(n8725), .B2(n15583), .ZN(n8652) );
  NAND2_X1 U11094 ( .A1(n10766), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U11095 ( .A1(n8951), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11096 ( .A1(n8654), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U11097 ( .A1(n8666), .A2(n8655), .ZN(n12896) );
  NAND2_X1 U11098 ( .A1(n8465), .A2(n12896), .ZN(n8657) );
  NAND2_X1 U11099 ( .A1(n8890), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8656) );
  NAND4_X1 U11100 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n12992) );
  NAND2_X1 U11101 ( .A1(n13448), .A2(n12992), .ZN(n12244) );
  XNOR2_X1 U11102 ( .A(n8661), .B(n8660), .ZN(n9637) );
  NAND2_X1 U11103 ( .A1(n9637), .A2(n7160), .ZN(n8665) );
  OAI21_X1 U11104 ( .B1(n8662), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8663) );
  XNOR2_X1 U11105 ( .A(n8663), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U11106 ( .A1(n8947), .A2(SI_15_), .B1(n8725), .B2(n13101), .ZN(
        n8664) );
  NAND2_X1 U11107 ( .A1(n8665), .A2(n8664), .ZN(n13029) );
  NAND2_X1 U11108 ( .A1(n8951), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11109 ( .A1(n10766), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11110 ( .A1(n8666), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11111 ( .A1(n8680), .A2(n8667), .ZN(n13318) );
  NAND2_X1 U11112 ( .A1(n8465), .A2(n13318), .ZN(n8669) );
  NAND2_X1 U11113 ( .A1(n8890), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8668) );
  NAND4_X1 U11114 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n13042) );
  OR2_X1 U11115 ( .A1(n13029), .A2(n13302), .ZN(n12257) );
  NAND2_X1 U11116 ( .A1(n13029), .A2(n13302), .ZN(n12243) );
  OR2_X1 U11117 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U11118 ( .A1(n8675), .A2(n8674), .ZN(n9710) );
  OR2_X1 U11119 ( .A1(n9710), .A2(n8749), .ZN(n8679) );
  NAND2_X1 U11120 ( .A1(n8676), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8677) );
  XNOR2_X1 U11121 ( .A(n8677), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U11122 ( .A1(n8947), .A2(SI_16_), .B1(n8725), .B2(n13103), .ZN(
        n8678) );
  NAND2_X1 U11123 ( .A1(n8679), .A2(n8678), .ZN(n12949) );
  NAND2_X1 U11124 ( .A1(n8951), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U11125 ( .A1(n8890), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U11126 ( .A1(n8680), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11127 ( .A1(n8697), .A2(n8681), .ZN(n13306) );
  NAND2_X1 U11128 ( .A1(n8465), .A2(n13306), .ZN(n8683) );
  NAND2_X1 U11129 ( .A1(n10766), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8682) );
  OR2_X1 U11130 ( .A1(n12949), .A2(n13315), .ZN(n12258) );
  NAND2_X1 U11131 ( .A1(n12949), .A2(n13315), .ZN(n12259) );
  NAND2_X1 U11132 ( .A1(n12258), .A2(n12259), .ZN(n13298) );
  INV_X1 U11133 ( .A(n13298), .ZN(n13304) );
  NAND2_X1 U11134 ( .A1(n13305), .A2(n13304), .ZN(n13303) );
  NAND2_X1 U11135 ( .A1(n13303), .A2(n12259), .ZN(n13292) );
  OR2_X1 U11136 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  NAND2_X1 U11137 ( .A1(n8689), .A2(n8688), .ZN(n9839) );
  OR2_X1 U11138 ( .A1(n9839), .A2(n8749), .ZN(n8696) );
  NAND2_X1 U11139 ( .A1(n8690), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8692) );
  MUX2_X1 U11140 ( .A(n8692), .B(P3_IR_REG_31__SCAN_IN), .S(n8691), .Z(n8694)
         );
  INV_X1 U11141 ( .A(n8693), .ZN(n8707) );
  NAND2_X1 U11142 ( .A1(n8694), .A2(n8707), .ZN(n14862) );
  AOI22_X1 U11143 ( .A1(n8947), .A2(SI_17_), .B1(n8725), .B2(n13054), .ZN(
        n8695) );
  NAND2_X1 U11144 ( .A1(n8696), .A2(n8695), .ZN(n13373) );
  NAND2_X1 U11145 ( .A1(n8951), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11146 ( .A1(n10766), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U11147 ( .A1(n8697), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11148 ( .A1(n8711), .A2(n8698), .ZN(n13293) );
  NAND2_X1 U11149 ( .A1(n8465), .A2(n13293), .ZN(n8700) );
  NAND2_X1 U11150 ( .A1(n8890), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8699) );
  OR2_X1 U11151 ( .A1(n13373), .A2(n13301), .ZN(n12265) );
  NAND2_X1 U11152 ( .A1(n13373), .A2(n13301), .ZN(n13275) );
  NAND2_X1 U11153 ( .A1(n12265), .A2(n13275), .ZN(n8868) );
  NAND2_X1 U11154 ( .A1(n13292), .A2(n13291), .ZN(n13290) );
  OR2_X1 U11155 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  NAND2_X1 U11156 ( .A1(n8706), .A2(n8705), .ZN(n10081) );
  OR2_X1 U11157 ( .A1(n10081), .A2(n8749), .ZN(n8710) );
  NAND2_X1 U11158 ( .A1(n8707), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8708) );
  XNOR2_X1 U11159 ( .A(n8708), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U11160 ( .A1(n8947), .A2(SI_18_), .B1(n8725), .B2(n14869), .ZN(
        n8709) );
  NAND2_X1 U11161 ( .A1(n8711), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11162 ( .A1(n8728), .A2(n8712), .ZN(n13279) );
  NAND2_X1 U11163 ( .A1(n13279), .A2(n8465), .ZN(n8716) );
  NAND2_X1 U11164 ( .A1(n10766), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11165 ( .A1(n8951), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11166 ( .A1(n8890), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11167 ( .A1(n13278), .A2(n13256), .ZN(n12268) );
  INV_X1 U11168 ( .A(n13276), .ZN(n8865) );
  INV_X1 U11169 ( .A(n13275), .ZN(n12267) );
  NOR2_X1 U11170 ( .A1(n8865), .A2(n12267), .ZN(n8717) );
  OR2_X1 U11171 ( .A1(n8719), .A2(n8718), .ZN(n8720) );
  NAND2_X1 U11172 ( .A1(n8721), .A2(n8720), .ZN(n10155) );
  OR2_X1 U11173 ( .A1(n10155), .A2(n8749), .ZN(n8727) );
  INV_X1 U11174 ( .A(n8829), .ZN(n8723) );
  NAND2_X1 U11175 ( .A1(n8723), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8724) );
  AOI22_X1 U11176 ( .A1(n8947), .A2(SI_19_), .B1(n13058), .B2(n8725), .ZN(
        n8726) );
  NAND2_X1 U11177 ( .A1(n8727), .A2(n8726), .ZN(n12909) );
  NAND2_X1 U11178 ( .A1(n8728), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U11179 ( .A1(n8739), .A2(n8729), .ZN(n13263) );
  NAND2_X1 U11180 ( .A1(n13263), .A2(n8465), .ZN(n8732) );
  AOI22_X1 U11181 ( .A1(n8951), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n8890), .B2(
        P3_REG0_REG_19__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11182 ( .A1(n10766), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8730) );
  OR2_X1 U11183 ( .A1(n12909), .A2(n13274), .ZN(n12275) );
  NAND2_X1 U11184 ( .A1(n12909), .A2(n13274), .ZN(n12276) );
  NAND2_X1 U11185 ( .A1(n8734), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11186 ( .A1(n8736), .A2(n8735), .ZN(n10346) );
  OR2_X1 U11187 ( .A1(n10346), .A2(n8749), .ZN(n8738) );
  OR2_X1 U11188 ( .A1(n12152), .A2(n10345), .ZN(n8737) );
  NAND2_X1 U11189 ( .A1(n8739), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11190 ( .A1(n8752), .A2(n8740), .ZN(n13245) );
  NAND2_X1 U11191 ( .A1(n13245), .A2(n8465), .ZN(n8743) );
  AOI22_X1 U11192 ( .A1(n10766), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n8951), 
        .B2(P3_REG2_REG_20__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11193 ( .A1(n8890), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8741) );
  XNOR2_X1 U11194 ( .A(n13247), .B(n13257), .ZN(n13241) );
  OR2_X1 U11195 ( .A1(n13247), .A2(n13257), .ZN(n12165) );
  OR2_X1 U11196 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  NAND2_X1 U11197 ( .A1(n8748), .A2(n8747), .ZN(n10416) );
  OR2_X1 U11198 ( .A1(n10416), .A2(n8749), .ZN(n8751) );
  INV_X1 U11199 ( .A(SI_21_), .ZN(n10415) );
  OR2_X1 U11200 ( .A1(n12152), .A2(n10415), .ZN(n8750) );
  NAND2_X1 U11201 ( .A1(n8752), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11202 ( .A1(n8761), .A2(n8753), .ZN(n13233) );
  NAND2_X1 U11203 ( .A1(n13233), .A2(n8465), .ZN(n8756) );
  AOI22_X1 U11204 ( .A1(n10766), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8951), 
        .B2(P3_REG2_REG_21__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11205 ( .A1(n8890), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11206 ( .A1(n12933), .A2(n13238), .ZN(n12282) );
  XNOR2_X1 U11207 ( .A(n8758), .B(n8757), .ZN(n10547) );
  NAND2_X1 U11208 ( .A1(n10547), .A2(n7160), .ZN(n8760) );
  OR2_X1 U11209 ( .A1(n12152), .A2(n7129), .ZN(n8759) );
  NAND2_X1 U11210 ( .A1(n8761), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11211 ( .A1(n8772), .A2(n8762), .ZN(n13221) );
  NAND2_X1 U11212 ( .A1(n13221), .A2(n8465), .ZN(n8767) );
  INV_X1 U11213 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U11214 ( .A1(n8890), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11215 ( .A1(n8951), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8763) );
  OAI211_X1 U11216 ( .C1(n8955), .C2(n13351), .A(n8764), .B(n8763), .ZN(n8765)
         );
  INV_X1 U11217 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U11218 ( .A1(n13220), .A2(n13199), .ZN(n12286) );
  XNOR2_X1 U11219 ( .A(n8769), .B(n8768), .ZN(n10815) );
  NAND2_X1 U11220 ( .A1(n10815), .A2(n7160), .ZN(n8771) );
  INV_X1 U11221 ( .A(SI_23_), .ZN(n10817) );
  OR2_X1 U11222 ( .A1(n12152), .A2(n10817), .ZN(n8770) );
  NAND2_X1 U11223 ( .A1(n8772), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11224 ( .A1(n8783), .A2(n8773), .ZN(n13208) );
  NAND2_X1 U11225 ( .A1(n13208), .A2(n8465), .ZN(n8778) );
  INV_X1 U11226 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U11227 ( .A1(n8890), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11228 ( .A1(n8951), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8774) );
  OAI211_X1 U11229 ( .C1(n8955), .C2(n13347), .A(n8775), .B(n8774), .ZN(n8776)
         );
  INV_X1 U11230 ( .A(n8776), .ZN(n8777) );
  NAND2_X1 U11231 ( .A1(n13209), .A2(n13217), .ZN(n8779) );
  XNOR2_X1 U11232 ( .A(n8780), .B(n11791), .ZN(n11218) );
  NAND2_X1 U11233 ( .A1(n11218), .A2(n7160), .ZN(n8782) );
  INV_X1 U11234 ( .A(SI_24_), .ZN(n11219) );
  OR2_X1 U11235 ( .A1(n12152), .A2(n11219), .ZN(n8781) );
  NAND2_X1 U11236 ( .A1(n8783), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11237 ( .A1(n8795), .A2(n8784), .ZN(n13191) );
  NAND2_X1 U11238 ( .A1(n13191), .A2(n8465), .ZN(n8789) );
  INV_X1 U11239 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U11240 ( .A1(n8951), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11241 ( .A1(n8890), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8785) );
  OAI211_X1 U11242 ( .C1(n8955), .C2(n13341), .A(n8786), .B(n8785), .ZN(n8787)
         );
  INV_X1 U11243 ( .A(n8787), .ZN(n8788) );
  INV_X1 U11244 ( .A(n13184), .ZN(n8790) );
  NAND2_X1 U11245 ( .A1(n12976), .A2(n13200), .ZN(n12293) );
  NAND2_X1 U11246 ( .A1(n13180), .A2(n12293), .ZN(n13174) );
  XNOR2_X1 U11247 ( .A(n14151), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8791) );
  XNOR2_X1 U11248 ( .A(n8792), .B(n8791), .ZN(n11378) );
  NAND2_X1 U11249 ( .A1(n11378), .A2(n7160), .ZN(n8794) );
  OR2_X1 U11250 ( .A1(n12152), .A2(n11379), .ZN(n8793) );
  NAND2_X1 U11251 ( .A1(n8795), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11252 ( .A1(n8807), .A2(n8796), .ZN(n13175) );
  NAND2_X1 U11253 ( .A1(n13175), .A2(n8465), .ZN(n8802) );
  INV_X1 U11254 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11255 ( .A1(n8890), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11256 ( .A1(n8951), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U11257 ( .C1(n8955), .C2(n8799), .A(n8798), .B(n8797), .ZN(n8800)
         );
  INV_X1 U11258 ( .A(n8800), .ZN(n8801) );
  NAND2_X1 U11259 ( .A1(n13335), .A2(n13157), .ZN(n12163) );
  NAND2_X1 U11260 ( .A1(n12162), .A2(n12163), .ZN(n8880) );
  INV_X1 U11261 ( .A(n12163), .ZN(n8803) );
  XNOR2_X1 U11262 ( .A(n14145), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8804) );
  INV_X1 U11263 ( .A(SI_26_), .ZN(n11483) );
  OR2_X1 U11264 ( .A1(n12152), .A2(n11483), .ZN(n8806) );
  NAND2_X1 U11265 ( .A1(n8807), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11266 ( .A1(n8818), .A2(n8808), .ZN(n13162) );
  NAND2_X1 U11267 ( .A1(n13162), .A2(n8465), .ZN(n8813) );
  INV_X1 U11268 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13333) );
  NAND2_X1 U11269 ( .A1(n8951), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11270 ( .A1(n8890), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8809) );
  OAI211_X1 U11271 ( .C1(n13333), .C2(n8955), .A(n8810), .B(n8809), .ZN(n8811)
         );
  INV_X1 U11272 ( .A(n8811), .ZN(n8812) );
  NAND2_X1 U11273 ( .A1(n13025), .A2(n13169), .ZN(n12299) );
  XNOR2_X1 U11274 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8814) );
  XNOR2_X1 U11275 ( .A(n8815), .B(n8814), .ZN(n11517) );
  NAND2_X1 U11276 ( .A1(n11517), .A2(n7160), .ZN(n8817) );
  NAND2_X1 U11277 ( .A1(n8947), .A2(SI_27_), .ZN(n8816) );
  NAND2_X1 U11278 ( .A1(n8818), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11279 ( .A1(n8820), .A2(n8819), .ZN(n13149) );
  NAND2_X1 U11280 ( .A1(n13149), .A2(n8465), .ZN(n8825) );
  INV_X1 U11281 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13329) );
  NAND2_X1 U11282 ( .A1(n8890), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11283 ( .A1(n8951), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U11284 ( .C1(n8955), .C2(n13329), .A(n8822), .B(n8821), .ZN(n8823)
         );
  INV_X1 U11285 ( .A(n8823), .ZN(n8824) );
  INV_X1 U11286 ( .A(n13141), .ZN(n8826) );
  NAND2_X1 U11287 ( .A1(n13148), .A2(n13158), .ZN(n8963) );
  NAND2_X1 U11288 ( .A1(n13137), .A2(n8963), .ZN(n8827) );
  XOR2_X1 U11289 ( .A(n12922), .B(n8827), .Z(n13133) );
  NAND2_X1 U11290 ( .A1(n8899), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8830) );
  INV_X1 U11291 ( .A(n8831), .ZN(n8832) );
  NAND2_X1 U11292 ( .A1(n8832), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11293 ( .A1(n12359), .A2(n10344), .ZN(n8837) );
  AOI21_X1 U11294 ( .B1(n8837), .B2(n13058), .A(n12171), .ZN(n8840) );
  NAND2_X1 U11295 ( .A1(n12176), .A2(n10344), .ZN(n8838) );
  NAND2_X1 U11296 ( .A1(n8843), .A2(n8838), .ZN(n8934) );
  INV_X1 U11297 ( .A(n8934), .ZN(n8839) );
  OR2_X1 U11298 ( .A1(n8840), .A2(n8839), .ZN(n10162) );
  NAND2_X1 U11299 ( .A1(n15672), .A2(n10194), .ZN(n8842) );
  INV_X1 U11300 ( .A(n10344), .ZN(n8886) );
  AND2_X1 U11301 ( .A1(n8886), .A2(n13089), .ZN(n8841) );
  NAND2_X1 U11302 ( .A1(n12359), .A2(n8841), .ZN(n8933) );
  AND2_X1 U11303 ( .A1(n10344), .A2(n13058), .ZN(n12323) );
  NAND2_X1 U11304 ( .A1(n8843), .A2(n12323), .ZN(n15719) );
  INV_X1 U11305 ( .A(n13335), .ZN(n8881) );
  NAND2_X1 U11306 ( .A1(n15652), .A2(n15678), .ZN(n15657) );
  NAND2_X1 U11307 ( .A1(n10181), .A2(n15657), .ZN(n15656) );
  NAND2_X1 U11308 ( .A1(n15674), .A2(n15650), .ZN(n15639) );
  NAND2_X1 U11309 ( .A1(n15656), .A2(n15639), .ZN(n8845) );
  NAND2_X1 U11310 ( .A1(n15624), .A2(n15646), .ZN(n8846) );
  NAND2_X1 U11311 ( .A1(n10799), .A2(n10366), .ZN(n8848) );
  NAND2_X1 U11312 ( .A1(n15626), .A2(n8848), .ZN(n10797) );
  NOR2_X1 U11313 ( .A1(n7631), .A2(n7630), .ZN(n15610) );
  INV_X1 U11314 ( .A(n15617), .ZN(n12198) );
  NAND2_X1 U11315 ( .A1(n10826), .A2(n12198), .ZN(n8849) );
  NAND2_X1 U11316 ( .A1(n11109), .A2(n10823), .ZN(n8850) );
  NAND2_X1 U11317 ( .A1(n11044), .A2(n12207), .ZN(n8852) );
  NAND2_X1 U11318 ( .A1(n15597), .A2(n11051), .ZN(n8851) );
  AND2_X1 U11319 ( .A1(n12216), .A2(n12218), .ZN(n8853) );
  XNOR2_X1 U11320 ( .A(n15598), .B(n11434), .ZN(n12332) );
  NAND2_X1 U11321 ( .A1(n12229), .A2(n12230), .ZN(n12226) );
  NAND2_X1 U11322 ( .A1(n11444), .A2(n12226), .ZN(n11443) );
  NAND2_X1 U11323 ( .A1(n11647), .A2(n11541), .ZN(n8854) );
  NAND2_X1 U11324 ( .A1(n11443), .A2(n8854), .ZN(n11559) );
  NAND2_X1 U11325 ( .A1(n11696), .A2(n11650), .ZN(n8855) );
  NAND2_X1 U11326 ( .A1(n11559), .A2(n8855), .ZN(n8857) );
  NAND2_X1 U11327 ( .A1(n11660), .A2(n11688), .ZN(n8856) );
  NAND2_X1 U11328 ( .A1(n8857), .A2(n8856), .ZN(n11521) );
  NAND2_X1 U11329 ( .A1(n11521), .A2(n12337), .ZN(n8859) );
  INV_X1 U11330 ( .A(n12994), .ZN(n13043) );
  NAND2_X1 U11331 ( .A1(n11694), .A2(n13043), .ZN(n8858) );
  NOR2_X1 U11332 ( .A1(n12995), .A2(n12849), .ZN(n8861) );
  NAND2_X1 U11333 ( .A1(n12995), .A2(n12849), .ZN(n8860) );
  INV_X1 U11334 ( .A(n12992), .ZN(n13314) );
  OR2_X1 U11335 ( .A1(n13029), .A2(n13042), .ZN(n8862) );
  NAND2_X1 U11336 ( .A1(n13311), .A2(n8862), .ZN(n8864) );
  NAND2_X1 U11337 ( .A1(n13029), .A2(n13042), .ZN(n8863) );
  NAND2_X1 U11338 ( .A1(n8864), .A2(n8863), .ZN(n13299) );
  NAND2_X1 U11339 ( .A1(n12949), .A2(n13287), .ZN(n13284) );
  NAND2_X1 U11340 ( .A1(n13373), .A2(n12954), .ZN(n8867) );
  AND2_X1 U11341 ( .A1(n13284), .A2(n8867), .ZN(n13267) );
  AND2_X1 U11342 ( .A1(n13267), .A2(n8865), .ZN(n8866) );
  NAND2_X1 U11343 ( .A1(n13285), .A2(n8866), .ZN(n13271) );
  INV_X1 U11344 ( .A(n13256), .ZN(n13288) );
  OR2_X1 U11345 ( .A1(n13278), .A2(n13288), .ZN(n8870) );
  INV_X1 U11346 ( .A(n8867), .ZN(n8869) );
  OR2_X1 U11347 ( .A1(n8869), .A2(n8868), .ZN(n13268) );
  OR2_X1 U11348 ( .A1(n13276), .A2(n13268), .ZN(n13270) );
  AND2_X1 U11349 ( .A1(n8870), .A2(n13270), .ZN(n13253) );
  AND2_X1 U11350 ( .A1(n13253), .A2(n13261), .ZN(n8871) );
  NAND2_X1 U11351 ( .A1(n13271), .A2(n8871), .ZN(n13259) );
  INV_X1 U11352 ( .A(n13274), .ZN(n12982) );
  NAND2_X1 U11353 ( .A1(n12909), .A2(n12982), .ZN(n8872) );
  NAND2_X1 U11354 ( .A1(n13259), .A2(n8872), .ZN(n13237) );
  AND2_X1 U11355 ( .A1(n13247), .A2(n13228), .ZN(n8873) );
  NAND2_X1 U11356 ( .A1(n12281), .A2(n12282), .ZN(n13231) );
  OR2_X1 U11357 ( .A1(n12933), .A2(n13002), .ZN(n8874) );
  NAND2_X1 U11358 ( .A1(n13226), .A2(n8874), .ZN(n13215) );
  NAND2_X1 U11359 ( .A1(n13220), .A2(n13229), .ZN(n8875) );
  OR2_X1 U11360 ( .A1(n13220), .A2(n13229), .ZN(n8876) );
  INV_X1 U11361 ( .A(n13204), .ZN(n8877) );
  INV_X1 U11362 ( .A(n13209), .ZN(n13343) );
  NAND2_X1 U11363 ( .A1(n13185), .A2(n13184), .ZN(n13183) );
  INV_X1 U11364 ( .A(n13200), .ZN(n8878) );
  NAND2_X1 U11365 ( .A1(n12976), .A2(n8878), .ZN(n8879) );
  NAND2_X1 U11366 ( .A1(n13183), .A2(n8879), .ZN(n13167) );
  NAND2_X1 U11367 ( .A1(n13167), .A2(n8880), .ZN(n13171) );
  NAND2_X1 U11368 ( .A1(n13407), .A2(n13169), .ZN(n8882) );
  NAND2_X1 U11369 ( .A1(n12359), .A2(n13058), .ZN(n8971) );
  NAND2_X1 U11370 ( .A1(n12171), .A2(n8886), .ZN(n12357) );
  NAND3_X1 U11371 ( .A1(n8942), .A2(n8887), .A3(n15671), .ZN(n8898) );
  INV_X1 U11372 ( .A(n13469), .ZN(n9869) );
  INV_X1 U11373 ( .A(n6678), .ZN(n8888) );
  NAND2_X1 U11374 ( .A1(n9869), .A2(n8888), .ZN(n9880) );
  NAND2_X2 U11375 ( .A1(n12359), .A2(n12171), .ZN(n12292) );
  INV_X1 U11376 ( .A(n13117), .ZN(n8889) );
  NAND2_X1 U11377 ( .A1(n8889), .A2(n8465), .ZN(n10771) );
  INV_X1 U11378 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U11379 ( .A1(n8951), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11380 ( .A1(n8890), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8891) );
  OAI211_X1 U11381 ( .C1(n8955), .C2(n8984), .A(n8892), .B(n8891), .ZN(n8893)
         );
  INV_X1 U11382 ( .A(n8893), .ZN(n8894) );
  NAND2_X1 U11383 ( .A1(n9880), .A2(n9868), .ZN(n8895) );
  NOR2_X1 U11384 ( .A1(n12928), .A2(n15673), .ZN(n8896) );
  INV_X1 U11385 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11386 ( .A1(n8902), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8903) );
  INV_X1 U11387 ( .A(n8904), .ZN(n8905) );
  NAND2_X1 U11388 ( .A1(n8905), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8906) );
  MUX2_X1 U11389 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8906), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8907) );
  NAND2_X1 U11390 ( .A1(n8907), .A2(n8902), .ZN(n11381) );
  NAND2_X1 U11391 ( .A1(n6756), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8909) );
  XNOR2_X1 U11392 ( .A(n8909), .B(n8908), .ZN(n11221) );
  NOR2_X1 U11393 ( .A1(n11381), .A2(n11221), .ZN(n8910) );
  XNOR2_X1 U11394 ( .A(n11221), .B(P3_B_REG_SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11395 ( .A1(n8911), .A2(n11381), .ZN(n8912) );
  NOR2_X1 U11396 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8916) );
  NOR4_X1 U11397 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8915) );
  NOR4_X1 U11398 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8914) );
  NOR4_X1 U11399 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8913) );
  NAND4_X1 U11400 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n8922)
         );
  NOR4_X1 U11401 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8920) );
  NOR4_X1 U11402 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8919) );
  NOR4_X1 U11403 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8918) );
  NOR4_X1 U11404 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8917) );
  NAND4_X1 U11405 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n8921)
         );
  NOR2_X1 U11406 ( .A1(n8922), .A2(n8921), .ZN(n8923) );
  NOR2_X1 U11407 ( .A1(n9547), .A2(n8923), .ZN(n8969) );
  NOR2_X1 U11408 ( .A1(n10794), .A2(n8969), .ZN(n8932) );
  INV_X1 U11409 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11410 ( .A1(n8928), .A2(n9511), .ZN(n8926) );
  INV_X1 U11411 ( .A(n8924), .ZN(n11484) );
  NAND2_X1 U11412 ( .A1(n11484), .A2(n11381), .ZN(n8925) );
  INV_X1 U11413 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8927) );
  NAND2_X1 U11414 ( .A1(n8928), .A2(n8927), .ZN(n8930) );
  NAND2_X1 U11415 ( .A1(n11484), .A2(n11221), .ZN(n8929) );
  XNOR2_X1 U11416 ( .A(n10788), .B(n8968), .ZN(n8931) );
  OR2_X1 U11417 ( .A1(n12292), .A2(n10194), .ZN(n10164) );
  NAND2_X1 U11418 ( .A1(n12292), .A2(n8933), .ZN(n10787) );
  NAND2_X1 U11419 ( .A1(n10164), .A2(n10787), .ZN(n10785) );
  NAND2_X1 U11420 ( .A1(n10785), .A2(n10788), .ZN(n8938) );
  INV_X1 U11421 ( .A(n10194), .ZN(n12322) );
  NAND3_X1 U11422 ( .A1(n8971), .A2(n8934), .A3(n12322), .ZN(n8935) );
  NAND2_X1 U11423 ( .A1(n8935), .A2(n12292), .ZN(n8936) );
  INV_X1 U11424 ( .A(n10788), .ZN(n10786) );
  NAND2_X1 U11425 ( .A1(n8936), .A2(n10786), .ZN(n8937) );
  MUX2_X1 U11426 ( .A(n8940), .B(n13397), .S(n15764), .Z(n8941) );
  NAND2_X1 U11427 ( .A1(n8941), .A2(n6795), .ZN(P3_U3487) );
  OAI21_X1 U11428 ( .B1(n13041), .B2(n13400), .A(n8942), .ZN(n8950) );
  INV_X1 U11429 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U11430 ( .A1(n8944), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U11431 ( .A1(n8946), .A2(n8945), .ZN(n12143) );
  XNOR2_X1 U11432 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12141) );
  XNOR2_X1 U11433 ( .A(n12143), .B(n12141), .ZN(n13462) );
  NAND2_X1 U11434 ( .A1(n13462), .A2(n7160), .ZN(n8949) );
  NAND2_X1 U11435 ( .A1(n8947), .A2(SI_29_), .ZN(n8948) );
  NAND2_X1 U11436 ( .A1(n8949), .A2(n8948), .ZN(n8977) );
  OR2_X1 U11437 ( .A1(n8977), .A2(n12928), .ZN(n12311) );
  NAND2_X1 U11438 ( .A1(n8977), .A2(n12928), .ZN(n12310) );
  XNOR2_X1 U11439 ( .A(n8950), .B(n12313), .ZN(n8962) );
  NOR2_X1 U11440 ( .A1(n13041), .A2(n15637), .ZN(n8960) );
  INV_X1 U11441 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11442 ( .A1(n8890), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U11443 ( .A1(n8951), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8952) );
  OAI211_X1 U11444 ( .C1(n8955), .C2(n8954), .A(n8953), .B(n8952), .ZN(n8956)
         );
  INV_X1 U11445 ( .A(n8956), .ZN(n8957) );
  AND2_X1 U11446 ( .A1(n10771), .A2(n8957), .ZN(n12154) );
  INV_X1 U11447 ( .A(P3_B_REG_SCAN_IN), .ZN(n9200) );
  NOR2_X1 U11448 ( .A1(n13469), .A2(n9200), .ZN(n8958) );
  OR2_X1 U11449 ( .A1(n15673), .A2(n8958), .ZN(n13114) );
  AND2_X1 U11450 ( .A1(n8964), .A2(n8963), .ZN(n12307) );
  INV_X1 U11451 ( .A(n8965), .ZN(n12306) );
  XOR2_X1 U11452 ( .A(n12313), .B(n12159), .Z(n13126) );
  NOR2_X1 U11453 ( .A1(n13121), .A2(n8966), .ZN(n8983) );
  NOR2_X1 U11454 ( .A1(n10788), .A2(n8969), .ZN(n8967) );
  NAND2_X1 U11455 ( .A1(n8967), .A2(n8968), .ZN(n10196) );
  INV_X1 U11456 ( .A(n10162), .ZN(n8972) );
  INV_X1 U11457 ( .A(n8969), .ZN(n8970) );
  NAND3_X1 U11458 ( .A1(n10172), .A2(n8970), .A3(n10788), .ZN(n10191) );
  OR2_X1 U11459 ( .A1(n8971), .A2(n12353), .ZN(n10186) );
  OAI22_X1 U11460 ( .A1(n10196), .A2(n8972), .B1(n10191), .B2(n10186), .ZN(
        n8973) );
  INV_X1 U11461 ( .A(n10794), .ZN(n10195) );
  NAND2_X1 U11462 ( .A1(n8973), .A2(n10195), .ZN(n8976) );
  OR2_X1 U11463 ( .A1(n12292), .A2(n12322), .ZN(n8974) );
  NOR2_X1 U11464 ( .A1(n10794), .A2(n8974), .ZN(n10168) );
  INV_X1 U11465 ( .A(n10191), .ZN(n10185) );
  NAND2_X1 U11466 ( .A1(n10168), .A2(n10185), .ZN(n8975) );
  OR2_X1 U11467 ( .A1(n8983), .A2(n15742), .ZN(n8982) );
  INV_X1 U11468 ( .A(n8977), .ZN(n13124) );
  INV_X1 U11469 ( .A(n13449), .ZN(n8980) );
  INV_X1 U11470 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8978) );
  NOR2_X1 U11471 ( .A1(n15740), .A2(n8978), .ZN(n8979) );
  AOI21_X1 U11472 ( .B1(n8977), .B2(n8980), .A(n8979), .ZN(n8981) );
  NAND2_X1 U11473 ( .A1(n8982), .A2(n8981), .ZN(P3_U3456) );
  OR2_X1 U11474 ( .A1(n8983), .A2(n15761), .ZN(n8988) );
  INV_X1 U11475 ( .A(n13390), .ZN(n8986) );
  NOR2_X1 U11476 ( .A1(n15764), .A2(n8984), .ZN(n8985) );
  NAND2_X1 U11477 ( .A1(n8988), .A2(n8987), .ZN(P3_U3488) );
  INV_X1 U11478 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9014) );
  XOR2_X1 U11479 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n9070) );
  INV_X1 U11480 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9012) );
  XOR2_X1 U11481 ( .A(n9012), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n9067) );
  INV_X1 U11482 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9830) );
  INV_X1 U11483 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n8989) );
  XOR2_X1 U11484 ( .A(n8989), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n9017) );
  INV_X1 U11485 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9704) );
  XNOR2_X1 U11486 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n15520), .ZN(n9059) );
  XNOR2_X1 U11487 ( .A(n15499), .B(n9632), .ZN(n9021) );
  XOR2_X1 U11488 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n9341), .Z(n9030) );
  NAND2_X1 U11489 ( .A1(n9030), .A2(n9029), .ZN(n8992) );
  NAND2_X1 U11490 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8993), .ZN(n8994) );
  NAND2_X1 U11491 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8995), .ZN(n8997) );
  NAND2_X1 U11492 ( .A1(n9023), .A2(n9024), .ZN(n8996) );
  NAND2_X1 U11493 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8998), .ZN(n9000) );
  INV_X1 U11494 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U11495 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15466), .ZN(n9001) );
  INV_X1 U11496 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15481) );
  NAND2_X1 U11497 ( .A1(n9002), .A2(n15481), .ZN(n9004) );
  XNOR2_X1 U11498 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9002), .ZN(n9051) );
  NAND2_X1 U11499 ( .A1(n9051), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11500 ( .A1(n9021), .A2(n9022), .ZN(n9005) );
  NAND2_X1 U11501 ( .A1(n9007), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9009) );
  XOR2_X1 U11502 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n9007), .Z(n9019) );
  INV_X1 U11503 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11504 ( .A1(n9019), .A2(n9020), .ZN(n9008) );
  NAND2_X1 U11505 ( .A1(n9009), .A2(n9008), .ZN(n9018) );
  NAND2_X1 U11506 ( .A1(n9017), .A2(n9018), .ZN(n9010) );
  NOR2_X1 U11507 ( .A1(n9070), .A2(n9071), .ZN(n9013) );
  AOI21_X1 U11508 ( .B1(n9014), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9013), .ZN(
        n9015) );
  INV_X1 U11509 ( .A(n9015), .ZN(n9074) );
  INV_X1 U11510 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9016) );
  XOR2_X1 U11511 ( .A(n9016), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n9075) );
  XOR2_X1 U11512 ( .A(n9074), .B(n9075), .Z(n9073) );
  INV_X1 U11513 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15230) );
  INV_X1 U11514 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15229) );
  XOR2_X1 U11515 ( .A(n9018), .B(n9017), .Z(n9065) );
  INV_X1 U11516 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9063) );
  XOR2_X1 U11517 ( .A(n9020), .B(n9019), .Z(n14788) );
  XOR2_X1 U11518 ( .A(n9022), .B(n9021), .Z(n9055) );
  XNOR2_X1 U11519 ( .A(n9024), .B(n9023), .ZN(n9038) );
  INV_X1 U11520 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9037) );
  XNOR2_X1 U11521 ( .A(n9025), .B(n9026), .ZN(n9027) );
  NAND2_X1 U11522 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9027), .ZN(n9028) );
  AOI21_X1 U11523 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n9231), .A(n9026), .ZN(
        n15769) );
  INV_X1 U11524 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15768) );
  NOR2_X1 U11525 ( .A1(n15769), .A2(n15768), .ZN(n15777) );
  XNOR2_X1 U11526 ( .A(n9030), .B(n9029), .ZN(n9032) );
  NAND2_X1 U11527 ( .A1(n9031), .A2(n9032), .ZN(n9034) );
  NAND2_X1 U11528 ( .A1(n14780), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11529 ( .A1(n9034), .A2(n9033), .ZN(n15773) );
  XNOR2_X1 U11530 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9035), .ZN(n15774) );
  NAND2_X1 U11531 ( .A1(n15773), .A2(n15774), .ZN(n9036) );
  NOR2_X1 U11532 ( .A1(n15773), .A2(n15774), .ZN(n15772) );
  AOI21_X1 U11533 ( .B1(n9037), .B2(n9036), .A(n15772), .ZN(n15766) );
  NAND2_X1 U11534 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9038), .ZN(n9039) );
  NOR2_X1 U11535 ( .A1(n9043), .A2(n9042), .ZN(n9045) );
  NAND2_X1 U11536 ( .A1(n9046), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9050) );
  XNOR2_X1 U11537 ( .A(n9047), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n9048) );
  XOR2_X1 U11538 ( .A(n9049), .B(n9048), .Z(n14781) );
  XOR2_X1 U11539 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9051), .Z(n15771) );
  NAND2_X1 U11540 ( .A1(n15770), .A2(n15771), .ZN(n9054) );
  NAND2_X1 U11541 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9052), .ZN(n9053) );
  NOR2_X1 U11542 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14783), .ZN(n9056) );
  XNOR2_X1 U11543 ( .A(n9059), .B(n9058), .ZN(n9061) );
  NAND2_X1 U11544 ( .A1(n9060), .A2(n9061), .ZN(n9062) );
  NOR2_X1 U11545 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n15000), .ZN(n9066) );
  XOR2_X1 U11546 ( .A(n9068), .B(n9067), .Z(n15005) );
  NAND2_X1 U11547 ( .A1(n15004), .A2(n15005), .ZN(n9069) );
  NOR2_X1 U11548 ( .A1(n15004), .A2(n15005), .ZN(n15003) );
  XOR2_X1 U11549 ( .A(n9071), .B(n9070), .Z(n15009) );
  NAND2_X1 U11550 ( .A1(n15008), .A2(n15009), .ZN(n9072) );
  INV_X1 U11551 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U11552 ( .A1(n9075), .A2(n9074), .ZN(n9076) );
  INV_X1 U11553 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9077) );
  XNOR2_X1 U11554 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n9077), .ZN(n9081) );
  XNOR2_X1 U11555 ( .A(n9082), .B(n9081), .ZN(n9079) );
  NOR2_X1 U11556 ( .A1(n9078), .A2(n9079), .ZN(n15015) );
  INV_X1 U11557 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n9080) );
  XOR2_X1 U11558 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9080), .Z(n9084) );
  INV_X1 U11559 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15028) );
  XOR2_X1 U11560 ( .A(n9084), .B(n9088), .Z(n9086) );
  NAND2_X1 U11561 ( .A1(n9085), .A2(n9086), .ZN(n9087) );
  INV_X1 U11562 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14861) );
  NAND2_X1 U11563 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n9088), .ZN(n9090) );
  NOR2_X1 U11564 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n9088), .ZN(n9089) );
  XOR2_X1 U11565 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9091), .Z(n9092) );
  NOR2_X1 U11566 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9091), .ZN(n9094) );
  INV_X1 U11567 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15043) );
  XNOR2_X1 U11568 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n15043), .ZN(n9096) );
  XNOR2_X1 U11569 ( .A(n9097), .B(n9096), .ZN(n9095) );
  NOR2_X1 U11570 ( .A1(n9097), .A2(n9096), .ZN(n9098) );
  AOI21_X1 U11571 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15043), .A(n9098), .ZN(
        n9101) );
  XNOR2_X1 U11572 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9099) );
  XOR2_X1 U11573 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(n9099), .Z(n9100) );
  INV_X1 U11574 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n10414) );
  XNOR2_X1 U11575 ( .A(n10414), .B(keyinput_f71), .ZN(n9108) );
  AOI22_X1 U11576 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f119), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n9102) );
  OAI221_X1 U11577 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f119), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n9102), .ZN(n9107) );
  AOI22_X1 U11578 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_f104), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n9103) );
  OAI221_X1 U11579 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_f104), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n9103), .ZN(n9106) );
  AOI22_X1 U11580 ( .A1(keyinput_f72), .A2(P3_DATAO_REG_24__SCAN_IN), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n9104) );
  OAI221_X1 U11581 ( .B1(keyinput_f72), .B2(P3_DATAO_REG_24__SCAN_IN), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n9104), .ZN(n9105) );
  NOR4_X1 U11582 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n9136)
         );
  AOI22_X1 U11583 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(keyinput_f61), .ZN(n9109) );
  OAI221_X1 U11584 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P3_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n9109), .ZN(n9116) );
  AOI22_X1 U11585 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f118), .B1(SI_10_), .B2(keyinput_f22), .ZN(n9110) );
  OAI221_X1 U11586 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f118), .C1(
        SI_10_), .C2(keyinput_f22), .A(n9110), .ZN(n9115) );
  AOI22_X1 U11587 ( .A1(keyinput_f76), .A2(P3_DATAO_REG_20__SCAN_IN), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_f125), .ZN(n9111) );
  OAI221_X1 U11588 ( .B1(keyinput_f76), .B2(P3_DATAO_REG_20__SCAN_IN), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_f125), .A(n9111), .ZN(n9114) );
  AOI22_X1 U11589 ( .A1(keyinput_f69), .A2(P3_DATAO_REG_27__SCAN_IN), .B1(
        SI_29_), .B2(keyinput_f3), .ZN(n9112) );
  OAI221_X1 U11590 ( .B1(keyinput_f69), .B2(P3_DATAO_REG_27__SCAN_IN), .C1(
        SI_29_), .C2(keyinput_f3), .A(n9112), .ZN(n9113) );
  NOR4_X1 U11591 ( .A1(n9116), .A2(n9115), .A3(n9114), .A4(n9113), .ZN(n9135)
         );
  AOI22_X1 U11592 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput_f98), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n9117) );
  OAI221_X1 U11593 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_f98), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n9117), .ZN(n9124) );
  AOI22_X1 U11594 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9118) );
  OAI221_X1 U11595 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9118), .ZN(n9123) );
  AOI22_X1 U11596 ( .A1(keyinput_f84), .A2(P3_DATAO_REG_12__SCAN_IN), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_f122), .ZN(n9119) );
  OAI221_X1 U11597 ( .B1(keyinput_f84), .B2(P3_DATAO_REG_12__SCAN_IN), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_f122), .A(n9119), .ZN(n9122) );
  AOI22_X1 U11598 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(SI_12_), 
        .B2(keyinput_f20), .ZN(n9120) );
  OAI221_X1 U11599 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(SI_12_), .C2(keyinput_f20), .A(n9120), .ZN(n9121) );
  NOR4_X1 U11600 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n9134)
         );
  AOI22_X1 U11601 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f108), .B1(SI_6_), 
        .B2(keyinput_f26), .ZN(n9125) );
  OAI221_X1 U11602 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .C1(SI_6_), 
        .C2(keyinput_f26), .A(n9125), .ZN(n9132) );
  AOI22_X1 U11603 ( .A1(SI_8_), .A2(keyinput_f24), .B1(SI_19_), .B2(
        keyinput_f13), .ZN(n9126) );
  OAI221_X1 U11604 ( .B1(SI_8_), .B2(keyinput_f24), .C1(SI_19_), .C2(
        keyinput_f13), .A(n9126), .ZN(n9131) );
  AOI22_X1 U11605 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n9127) );
  OAI221_X1 U11606 ( .B1(SI_25_), .B2(keyinput_f7), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n9127), .ZN(n9130) );
  AOI22_X1 U11607 ( .A1(SI_13_), .A2(keyinput_f19), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n9128) );
  OAI221_X1 U11608 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n9128), .ZN(n9129) );
  NOR4_X1 U11609 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9133)
         );
  NAND4_X1 U11610 ( .A1(n9136), .A2(n9135), .A3(n9134), .A4(n9133), .ZN(n9257)
         );
  AOI22_X1 U11611 ( .A1(P3_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n9137) );
  OAI221_X1 U11612 ( .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        SI_23_), .C2(keyinput_f9), .A(n9137), .ZN(n9144) );
  AOI22_X1 U11613 ( .A1(SI_1_), .A2(keyinput_f31), .B1(SI_3_), .B2(
        keyinput_f29), .ZN(n9138) );
  OAI221_X1 U11614 ( .B1(SI_1_), .B2(keyinput_f31), .C1(SI_3_), .C2(
        keyinput_f29), .A(n9138), .ZN(n9143) );
  AOI22_X1 U11615 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f124), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n9139) );
  OAI221_X1 U11616 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f124), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n9139), .ZN(n9142) );
  AOI22_X1 U11617 ( .A1(keyinput_f87), .A2(P3_DATAO_REG_9__SCAN_IN), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_f116), .ZN(n9140) );
  OAI221_X1 U11618 ( .B1(keyinput_f87), .B2(P3_DATAO_REG_9__SCAN_IN), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_f116), .A(n9140), .ZN(n9141) );
  NOR4_X1 U11619 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n9172)
         );
  AOI22_X1 U11620 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f110), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n9145) );
  OAI221_X1 U11621 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f110), .C1(SI_2_), 
        .C2(keyinput_f30), .A(n9145), .ZN(n9152) );
  AOI22_X1 U11622 ( .A1(SI_15_), .A2(keyinput_f17), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n9146) );
  OAI221_X1 U11623 ( .B1(SI_15_), .B2(keyinput_f17), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n9146), .ZN(n9151) );
  AOI22_X1 U11624 ( .A1(keyinput_f65), .A2(P3_DATAO_REG_31__SCAN_IN), .B1(
        SI_20_), .B2(keyinput_f12), .ZN(n9147) );
  OAI221_X1 U11625 ( .B1(keyinput_f65), .B2(P3_DATAO_REG_31__SCAN_IN), .C1(
        SI_20_), .C2(keyinput_f12), .A(n9147), .ZN(n9150) );
  AOI22_X1 U11626 ( .A1(keyinput_f85), .A2(P3_DATAO_REG_11__SCAN_IN), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f126), .ZN(n9148) );
  OAI221_X1 U11627 ( .B1(keyinput_f85), .B2(P3_DATAO_REG_11__SCAN_IN), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f126), .A(n9148), .ZN(n9149) );
  NOR4_X1 U11628 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(n9171)
         );
  AOI22_X1 U11629 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_f123), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n9153) );
  OAI221_X1 U11630 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_f123), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n9153), .ZN(n9160) );
  AOI22_X1 U11631 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f115), .B1(SI_26_), 
        .B2(keyinput_f6), .ZN(n9154) );
  OAI221_X1 U11632 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f115), .C1(SI_26_), .C2(keyinput_f6), .A(n9154), .ZN(n9159) );
  AOI22_X1 U11633 ( .A1(keyinput_f86), .A2(P3_DATAO_REG_10__SCAN_IN), .B1(
        SI_9_), .B2(keyinput_f23), .ZN(n9155) );
  OAI221_X1 U11634 ( .B1(keyinput_f86), .B2(P3_DATAO_REG_10__SCAN_IN), .C1(
        SI_9_), .C2(keyinput_f23), .A(n9155), .ZN(n9158) );
  AOI22_X1 U11635 ( .A1(keyinput_f66), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(
        keyinput_f90), .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n9156) );
  OAI221_X1 U11636 ( .B1(keyinput_f66), .B2(P3_DATAO_REG_30__SCAN_IN), .C1(
        keyinput_f90), .C2(P3_DATAO_REG_6__SCAN_IN), .A(n9156), .ZN(n9157) );
  NOR4_X1 U11637 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n9170)
         );
  AOI22_X1 U11638 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        SI_14_), .B2(keyinput_f18), .ZN(n9161) );
  OAI221_X1 U11639 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        SI_14_), .C2(keyinput_f18), .A(n9161), .ZN(n9168) );
  AOI22_X1 U11640 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput_f83), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_f121), .ZN(n9162) );
  OAI221_X1 U11641 ( .B1(P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_f121), .A(n9162), .ZN(n9167) );
  AOI22_X1 U11642 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_f99), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n9163) );
  OAI221_X1 U11643 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_f99), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n9163), .ZN(n9166) );
  AOI22_X1 U11644 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_f101), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f112), .ZN(n9164) );
  OAI221_X1 U11645 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_f101), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f112), .A(n9164), .ZN(n9165) );
  NOR4_X1 U11646 ( .A1(n9168), .A2(n9167), .A3(n9166), .A4(n9165), .ZN(n9169)
         );
  NAND4_X1 U11647 ( .A1(n9172), .A2(n9171), .A3(n9170), .A4(n9169), .ZN(n9256)
         );
  AOI22_X1 U11648 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_f117), .ZN(n9173) );
  OAI221_X1 U11649 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_f117), .A(n9173), .ZN(n9180) );
  AOI22_X1 U11650 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_4_), .B2(
        keyinput_f28), .ZN(n9174) );
  OAI221_X1 U11651 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_4_), .C2(
        keyinput_f28), .A(n9174), .ZN(n9179) );
  AOI22_X1 U11652 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput_f96), .B1(
        keyinput_f81), .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n9175) );
  OAI221_X1 U11653 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_f96), .C1(
        keyinput_f81), .C2(P3_DATAO_REG_15__SCAN_IN), .A(n9175), .ZN(n9178) );
  AOI22_X1 U11654 ( .A1(keyinput_f68), .A2(P3_DATAO_REG_28__SCAN_IN), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n9176) );
  OAI221_X1 U11655 ( .B1(keyinput_f68), .B2(P3_DATAO_REG_28__SCAN_IN), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n9176), .ZN(n9177) );
  NOR4_X1 U11656 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), .ZN(n9211)
         );
  AOI22_X1 U11657 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f127), .B1(SI_27_), .B2(keyinput_f5), .ZN(n9181) );
  OAI221_X1 U11658 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f127), .C1(
        SI_27_), .C2(keyinput_f5), .A(n9181), .ZN(n9188) );
  AOI22_X1 U11659 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n9182) );
  OAI221_X1 U11660 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_17_), .C2(
        keyinput_f15), .A(n9182), .ZN(n9187) );
  AOI22_X1 U11661 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n9183) );
  OAI221_X1 U11662 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n9183), .ZN(n9186) );
  INV_X1 U11663 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U11664 ( .A1(n9967), .A2(keyinput_f93), .B1(n15466), .B2(
        keyinput_f103), .ZN(n9184) );
  OAI221_X1 U11665 ( .B1(n9967), .B2(keyinput_f93), .C1(n15466), .C2(
        keyinput_f103), .A(n9184), .ZN(n9185) );
  NOR4_X1 U11666 ( .A1(n9188), .A2(n9187), .A3(n9186), .A4(n9185), .ZN(n9210)
         );
  INV_X1 U11667 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11668 ( .A1(n9977), .A2(keyinput_f78), .B1(n13033), .B2(
        keyinput_f63), .ZN(n9189) );
  OAI221_X1 U11669 ( .B1(n9977), .B2(keyinput_f78), .C1(n13033), .C2(
        keyinput_f63), .A(n9189), .ZN(n9197) );
  INV_X1 U11670 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U11671 ( .A1(n10343), .A2(keyinput_f73), .B1(n11693), .B2(
        keyinput_f46), .ZN(n9190) );
  OAI221_X1 U11672 ( .B1(n10343), .B2(keyinput_f73), .C1(n11693), .C2(
        keyinput_f46), .A(n9190), .ZN(n9196) );
  INV_X1 U11673 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U11674 ( .A1(n9711), .A2(keyinput_f16), .B1(n10644), .B2(
        keyinput_f39), .ZN(n9191) );
  OAI221_X1 U11675 ( .B1(n9711), .B2(keyinput_f16), .C1(n10644), .C2(
        keyinput_f39), .A(n9191), .ZN(n9195) );
  XNOR2_X1 U11676 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f113), .ZN(n9193) );
  XNOR2_X1 U11677 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_f54), .ZN(n9192)
         );
  NAND2_X1 U11678 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  NOR4_X1 U11679 ( .A1(n9197), .A2(n9196), .A3(n9195), .A4(n9194), .ZN(n9209)
         );
  INV_X1 U11680 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n9328) );
  AOI22_X1 U11681 ( .A1(n11219), .A2(keyinput_f8), .B1(keyinput_f67), .B2(
        n9328), .ZN(n9198) );
  OAI221_X1 U11682 ( .B1(n11219), .B2(keyinput_f8), .C1(n9328), .C2(
        keyinput_f67), .A(n9198), .ZN(n9203) );
  AOI22_X1 U11683 ( .A1(n9200), .A2(keyinput_f64), .B1(keyinput_f120), .B2(
        n10149), .ZN(n9199) );
  OAI221_X1 U11684 ( .B1(n9200), .B2(keyinput_f64), .C1(n10149), .C2(
        keyinput_f120), .A(n9199), .ZN(n9202) );
  XNOR2_X1 U11685 ( .A(n7302), .B(keyinput_f107), .ZN(n9201) );
  OR3_X1 U11686 ( .A1(n9203), .A2(n9202), .A3(n9201), .ZN(n9207) );
  AOI22_X1 U11687 ( .A1(n9536), .A2(keyinput_f21), .B1(keyinput_f100), .B2(
        n9325), .ZN(n9204) );
  OAI221_X1 U11688 ( .B1(n9536), .B2(keyinput_f21), .C1(n9325), .C2(
        keyinput_f100), .A(n9204), .ZN(n9206) );
  INV_X1 U11689 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14779) );
  XNOR2_X1 U11690 ( .A(n14779), .B(keyinput_f33), .ZN(n9205) );
  NOR3_X1 U11691 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(n9208) );
  NAND4_X1 U11692 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n9255)
         );
  INV_X1 U11693 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9393) );
  INV_X1 U11694 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U11695 ( .A1(n9393), .A2(keyinput_f62), .B1(keyinput_f70), .B2(
        n10574), .ZN(n9212) );
  OAI221_X1 U11696 ( .B1(n9393), .B2(keyinput_f62), .C1(n10574), .C2(
        keyinput_f70), .A(n9212), .ZN(n9220) );
  INV_X1 U11697 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U11698 ( .A1(n13470), .A2(keyinput_f4), .B1(n13012), .B2(
        keyinput_f60), .ZN(n9213) );
  OAI221_X1 U11699 ( .B1(n13470), .B2(keyinput_f4), .C1(n13012), .C2(
        keyinput_f60), .A(n9213), .ZN(n9219) );
  XNOR2_X1 U11700 ( .A(SI_7_), .B(keyinput_f25), .ZN(n9217) );
  XNOR2_X1 U11701 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n9216)
         );
  XNOR2_X1 U11702 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_f44), .ZN(n9215)
         );
  XNOR2_X1 U11703 ( .A(SI_22_), .B(keyinput_f10), .ZN(n9214) );
  NAND4_X1 U11704 ( .A1(n9217), .A2(n9216), .A3(n9215), .A4(n9214), .ZN(n9218)
         );
  NOR3_X1 U11705 ( .A1(n9220), .A2(n9219), .A3(n9218), .ZN(n9253) );
  INV_X1 U11706 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11707 ( .A1(n9971), .A2(keyinput_f79), .B1(n15499), .B2(
        keyinput_f105), .ZN(n9221) );
  OAI221_X1 U11708 ( .B1(n9971), .B2(keyinput_f79), .C1(n15499), .C2(
        keyinput_f105), .A(n9221), .ZN(n9229) );
  INV_X1 U11709 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10158) );
  INV_X1 U11710 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U11711 ( .A1(n10158), .A2(keyinput_f74), .B1(keyinput_f92), .B2(
        n9973), .ZN(n9222) );
  OAI221_X1 U11712 ( .B1(n10158), .B2(keyinput_f74), .C1(n9973), .C2(
        keyinput_f92), .A(n9222), .ZN(n9228) );
  INV_X1 U11713 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11714 ( .A1(n10069), .A2(keyinput_f49), .B1(keyinput_f88), .B2(
        n9991), .ZN(n9223) );
  OAI221_X1 U11715 ( .B1(n10069), .B2(keyinput_f49), .C1(n9991), .C2(
        keyinput_f88), .A(n9223), .ZN(n9227) );
  INV_X1 U11716 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9388) );
  XOR2_X1 U11717 ( .A(n9388), .B(keyinput_f45), .Z(n9225) );
  XNOR2_X1 U11718 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f114), .ZN(n9224) );
  NAND2_X1 U11719 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NOR4_X1 U11720 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(n9252)
         );
  INV_X1 U11721 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U11722 ( .A1(n9987), .A2(keyinput_f77), .B1(n9231), .B2(
        keyinput_f97), .ZN(n9230) );
  OAI221_X1 U11723 ( .B1(n9987), .B2(keyinput_f77), .C1(n9231), .C2(
        keyinput_f97), .A(n9230), .ZN(n9240) );
  AOI22_X1 U11724 ( .A1(n15520), .A2(keyinput_f106), .B1(keyinput_f102), .B2(
        n9264), .ZN(n9232) );
  OAI221_X1 U11725 ( .B1(n15520), .B2(keyinput_f106), .C1(n9264), .C2(
        keyinput_f102), .A(n9232), .ZN(n9239) );
  INV_X1 U11726 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U11727 ( .A1(n12953), .A2(keyinput_f48), .B1(n9234), .B2(
        keyinput_f50), .ZN(n9233) );
  OAI221_X1 U11728 ( .B1(n12953), .B2(keyinput_f48), .C1(n9234), .C2(
        keyinput_f50), .A(n9233), .ZN(n9238) );
  INV_X1 U11729 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U11730 ( .A1(n9236), .A2(keyinput_f36), .B1(keyinput_f75), .B2(
        n10084), .ZN(n9235) );
  OAI221_X1 U11731 ( .B1(n9236), .B2(keyinput_f36), .C1(n10084), .C2(
        keyinput_f75), .A(n9235), .ZN(n9237) );
  NOR4_X1 U11732 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n9251)
         );
  INV_X1 U11733 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11734 ( .A1(n10082), .A2(keyinput_f14), .B1(keyinput_f82), .B2(
        n9981), .ZN(n9241) );
  OAI221_X1 U11735 ( .B1(n10082), .B2(keyinput_f14), .C1(n9981), .C2(
        keyinput_f82), .A(n9241), .ZN(n9244) );
  XNOR2_X1 U11736 ( .A(n9432), .B(keyinput_f109), .ZN(n9243) );
  INV_X1 U11737 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10006) );
  XNOR2_X1 U11738 ( .A(n10006), .B(keyinput_f94), .ZN(n9242) );
  OR3_X1 U11739 ( .A1(n9244), .A2(n9243), .A3(n9242), .ZN(n9249) );
  INV_X1 U11740 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n9989) );
  INV_X1 U11741 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11742 ( .A1(n9989), .A2(keyinput_f95), .B1(keyinput_f91), .B2(
        n9979), .ZN(n9245) );
  OAI221_X1 U11743 ( .B1(n9989), .B2(keyinput_f95), .C1(n9979), .C2(
        keyinput_f91), .A(n9245), .ZN(n9248) );
  INV_X1 U11744 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U11745 ( .A1(n10415), .A2(keyinput_f11), .B1(n12991), .B2(
        keyinput_f56), .ZN(n9246) );
  OAI221_X1 U11746 ( .B1(n10415), .B2(keyinput_f11), .C1(n12991), .C2(
        keyinput_f56), .A(n9246), .ZN(n9247) );
  NOR3_X1 U11747 ( .A1(n9249), .A2(n9248), .A3(n9247), .ZN(n9250) );
  NAND4_X1 U11748 ( .A1(n9253), .A2(n9252), .A3(n9251), .A4(n9250), .ZN(n9254)
         );
  OR4_X1 U11749 ( .A1(n9257), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n9260)
         );
  AOI21_X1 U11750 ( .B1(keyinput_f32), .B2(n9260), .A(keyinput_g32), .ZN(n9262) );
  INV_X1 U11751 ( .A(keyinput_f32), .ZN(n9259) );
  INV_X1 U11752 ( .A(keyinput_g32), .ZN(n9258) );
  AOI21_X1 U11753 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9261) );
  MUX2_X1 U11754 ( .A(n9262), .B(n9261), .S(SI_0_), .Z(n9263) );
  INV_X1 U11755 ( .A(n9263), .ZN(n9427) );
  XNOR2_X1 U11756 ( .A(n9264), .B(keyinput_g102), .ZN(n9271) );
  AOI22_X1 U11757 ( .A1(P3_DATAO_REG_19__SCAN_IN), .A2(keyinput_g77), .B1(
        SI_9_), .B2(keyinput_g23), .ZN(n9265) );
  OAI221_X1 U11758 ( .B1(P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .C1(
        SI_9_), .C2(keyinput_g23), .A(n9265), .ZN(n9270) );
  AOI22_X1 U11759 ( .A1(SI_13_), .A2(keyinput_g19), .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n9266) );
  OAI221_X1 U11760 ( .B1(SI_13_), .B2(keyinput_g19), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n9266), .ZN(n9269) );
  AOI22_X1 U11761 ( .A1(P3_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_g97), .ZN(n9267) );
  OAI221_X1 U11762 ( .B1(P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        P3_ADDR_REG_0__SCAN_IN), .C2(keyinput_g97), .A(n9267), .ZN(n9268) );
  NOR4_X1 U11763 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9299)
         );
  AOI22_X1 U11764 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_6_), 
        .B2(keyinput_g26), .ZN(n9272) );
  OAI221_X1 U11765 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(SI_6_), .C2(keyinput_g26), .A(n9272), .ZN(n9279) );
  AOI22_X1 U11766 ( .A1(P3_DATAO_REG_3__SCAN_IN), .A2(keyinput_g93), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9273) );
  OAI221_X1 U11767 ( .B1(P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_g93), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9273), .ZN(n9278) );
  AOI22_X1 U11768 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_g113), .B1(SI_18_), 
        .B2(keyinput_g14), .ZN(n9274) );
  OAI221_X1 U11769 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_g113), .C1(SI_18_), .C2(keyinput_g14), .A(n9274), .ZN(n9277) );
  AOI22_X1 U11770 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_g117), .B1(SI_14_), .B2(keyinput_g18), .ZN(n9275) );
  OAI221_X1 U11771 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_g117), .C1(
        SI_14_), .C2(keyinput_g18), .A(n9275), .ZN(n9276) );
  NOR4_X1 U11772 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(n9298)
         );
  AOI22_X1 U11773 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9280) );
  OAI221_X1 U11774 ( .B1(SI_8_), .B2(keyinput_g24), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9280), .ZN(n9287) );
  AOI22_X1 U11775 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n9281) );
  OAI221_X1 U11776 ( .B1(P3_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n9281), .ZN(n9286) );
  AOI22_X1 U11777 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_g104), .B1(
        SI_10_), .B2(keyinput_g22), .ZN(n9282) );
  OAI221_X1 U11778 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_10_), .C2(keyinput_g22), .A(n9282), .ZN(n9285) );
  AOI22_X1 U11779 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        SI_1_), .B2(keyinput_g31), .ZN(n9283) );
  OAI221_X1 U11780 ( .B1(P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        SI_1_), .C2(keyinput_g31), .A(n9283), .ZN(n9284) );
  NOR4_X1 U11781 ( .A1(n9287), .A2(n9286), .A3(n9285), .A4(n9284), .ZN(n9297)
         );
  AOI22_X1 U11782 ( .A1(SI_28_), .A2(keyinput_g4), .B1(P3_B_REG_SCAN_IN), .B2(
        keyinput_g64), .ZN(n9288) );
  OAI221_X1 U11783 ( .B1(SI_28_), .B2(keyinput_g4), .C1(P3_B_REG_SCAN_IN), 
        .C2(keyinput_g64), .A(n9288), .ZN(n9295) );
  AOI22_X1 U11784 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput_g98), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n9289) );
  OAI221_X1 U11785 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_g98), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n9289), .ZN(n9294) );
  AOI22_X1 U11786 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .ZN(n9290) );
  OAI221_X1 U11787 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        P3_WR_REG_SCAN_IN), .C2(keyinput_g0), .A(n9290), .ZN(n9293) );
  AOI22_X1 U11788 ( .A1(P3_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        SI_29_), .B2(keyinput_g3), .ZN(n9291) );
  OAI221_X1 U11789 ( .B1(P3_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        SI_29_), .C2(keyinput_g3), .A(n9291), .ZN(n9292) );
  NOR4_X1 U11790 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n9296)
         );
  NAND4_X1 U11791 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), .ZN(n9425)
         );
  AOI22_X1 U11792 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n9300) );
  OAI221_X1 U11793 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_4_), .C2(keyinput_g28), .A(n9300), .ZN(n9307) );
  AOI22_X1 U11794 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9301) );
  OAI221_X1 U11795 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n9301), .ZN(n9306) );
  AOI22_X1 U11796 ( .A1(P3_DATAO_REG_18__SCAN_IN), .A2(keyinput_g78), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_g101), .ZN(n9302) );
  OAI221_X1 U11797 ( .B1(P3_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_g101), .A(n9302), .ZN(n9305) );
  AOI22_X1 U11798 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g123), .B1(SI_15_), .B2(keyinput_g17), .ZN(n9303) );
  OAI221_X1 U11799 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g123), .C1(
        SI_15_), .C2(keyinput_g17), .A(n9303), .ZN(n9304) );
  NOR4_X1 U11800 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n9339)
         );
  AOI22_X1 U11801 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g124), .B1(SI_3_), 
        .B2(keyinput_g29), .ZN(n9308) );
  OAI221_X1 U11802 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g124), .C1(SI_3_), .C2(keyinput_g29), .A(n9308), .ZN(n9315) );
  AOI22_X1 U11803 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g110), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .ZN(n9309) );
  OAI221_X1 U11804 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g110), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n9309), .ZN(n9314) );
  AOI22_X1 U11805 ( .A1(P3_DATAO_REG_25__SCAN_IN), .A2(keyinput_g71), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n9310) );
  OAI221_X1 U11806 ( .B1(P3_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n9310), .ZN(n9313) );
  AOI22_X1 U11807 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g122), .B1(SI_17_), .B2(keyinput_g15), .ZN(n9311) );
  OAI221_X1 U11808 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g122), .C1(
        SI_17_), .C2(keyinput_g15), .A(n9311), .ZN(n9312) );
  NOR4_X1 U11809 ( .A1(n9315), .A2(n9314), .A3(n9313), .A4(n9312), .ZN(n9338)
         );
  AOI22_X1 U11810 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P3_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .ZN(n9316) );
  OAI221_X1 U11811 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        P3_DATAO_REG_24__SCAN_IN), .C2(keyinput_g72), .A(n9316), .ZN(n9323) );
  AOI22_X1 U11812 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_g125), .B1(SI_27_), .B2(keyinput_g5), .ZN(n9317) );
  OAI221_X1 U11813 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_g125), .C1(
        SI_27_), .C2(keyinput_g5), .A(n9317), .ZN(n9322) );
  AOI22_X1 U11814 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g112), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_g126), .ZN(n9318) );
  OAI221_X1 U11815 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g112), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_g126), .A(n9318), .ZN(n9321) );
  AOI22_X1 U11816 ( .A1(SI_16_), .A2(keyinput_g16), .B1(SI_12_), .B2(
        keyinput_g20), .ZN(n9319) );
  OAI221_X1 U11817 ( .B1(SI_16_), .B2(keyinput_g16), .C1(SI_12_), .C2(
        keyinput_g20), .A(n9319), .ZN(n9320) );
  NOR4_X1 U11818 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(n9337)
         );
  AOI22_X1 U11819 ( .A1(n9431), .A2(keyinput_g121), .B1(keyinput_g100), .B2(
        n9325), .ZN(n9324) );
  OAI221_X1 U11820 ( .B1(n9431), .B2(keyinput_g121), .C1(n9325), .C2(
        keyinput_g100), .A(n9324), .ZN(n9335) );
  AOI22_X1 U11821 ( .A1(n9328), .A2(keyinput_g67), .B1(n9327), .B2(
        keyinput_g35), .ZN(n9326) );
  OAI221_X1 U11822 ( .B1(n9328), .B2(keyinput_g67), .C1(n9327), .C2(
        keyinput_g35), .A(n9326), .ZN(n9334) );
  XOR2_X1 U11823 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_g43), .Z(n9331) );
  XNOR2_X1 U11824 ( .A(SI_5_), .B(keyinput_g27), .ZN(n9330) );
  XNOR2_X1 U11825 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g114), .ZN(n9329) );
  NAND3_X1 U11826 ( .A1(n9331), .A2(n9330), .A3(n9329), .ZN(n9333) );
  XNOR2_X1 U11827 ( .A(n9991), .B(keyinput_g88), .ZN(n9332) );
  NOR4_X1 U11828 ( .A1(n9335), .A2(n9334), .A3(n9333), .A4(n9332), .ZN(n9336)
         );
  NAND4_X1 U11829 ( .A1(n9339), .A2(n9338), .A3(n9337), .A4(n9336), .ZN(n9424)
         );
  AOI22_X1 U11830 ( .A1(n13012), .A2(keyinput_g60), .B1(keyinput_g99), .B2(
        n9341), .ZN(n9340) );
  OAI221_X1 U11831 ( .B1(n13012), .B2(keyinput_g60), .C1(n9341), .C2(
        keyinput_g99), .A(n9340), .ZN(n9349) );
  INV_X1 U11832 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10004) );
  INV_X1 U11833 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11834 ( .A1(n10004), .A2(keyinput_g96), .B1(n9963), .B2(
        keyinput_g89), .ZN(n9342) );
  OAI221_X1 U11835 ( .B1(n10004), .B2(keyinput_g96), .C1(n9963), .C2(
        keyinput_g89), .A(n9342), .ZN(n9348) );
  INV_X1 U11836 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U11837 ( .A1(n9975), .A2(keyinput_g80), .B1(n8424), .B2(
        keyinput_g53), .ZN(n9343) );
  OAI221_X1 U11838 ( .B1(n9975), .B2(keyinput_g80), .C1(n8424), .C2(
        keyinput_g53), .A(n9343), .ZN(n9347) );
  INV_X1 U11839 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9345) );
  AOI22_X1 U11840 ( .A1(n9345), .A2(keyinput_g38), .B1(P3_U3151), .B2(
        keyinput_g34), .ZN(n9344) );
  OAI221_X1 U11841 ( .B1(n9345), .B2(keyinput_g38), .C1(P3_U3151), .C2(
        keyinput_g34), .A(n9344), .ZN(n9346) );
  NOR4_X1 U11842 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), .ZN(n9381)
         );
  AOI22_X1 U11843 ( .A1(n10084), .A2(keyinput_g75), .B1(n9973), .B2(
        keyinput_g92), .ZN(n9350) );
  OAI221_X1 U11844 ( .B1(n10084), .B2(keyinput_g75), .C1(n9973), .C2(
        keyinput_g92), .A(n9350), .ZN(n9358) );
  INV_X1 U11845 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U11846 ( .A1(n15466), .A2(keyinput_g103), .B1(keyinput_g69), .B2(
        n10765), .ZN(n9351) );
  OAI221_X1 U11847 ( .B1(n15466), .B2(keyinput_g103), .C1(n10765), .C2(
        keyinput_g69), .A(n9351), .ZN(n9357) );
  AOI22_X1 U11848 ( .A1(n7129), .A2(keyinput_g10), .B1(keyinput_g118), .B2(
        n9822), .ZN(n9352) );
  OAI221_X1 U11849 ( .B1(n7129), .B2(keyinput_g10), .C1(n9822), .C2(
        keyinput_g118), .A(n9352), .ZN(n9355) );
  XNOR2_X1 U11850 ( .A(n9989), .B(keyinput_g95), .ZN(n9354) );
  XNOR2_X1 U11851 ( .A(n9602), .B(keyinput_g115), .ZN(n9353) );
  OR3_X1 U11852 ( .A1(n9355), .A2(n9354), .A3(n9353), .ZN(n9356) );
  NOR3_X1 U11853 ( .A1(n9358), .A2(n9357), .A3(n9356), .ZN(n9380) );
  AOI22_X1 U11854 ( .A1(n10343), .A2(keyinput_g73), .B1(n8475), .B2(
        keyinput_g40), .ZN(n9359) );
  OAI221_X1 U11855 ( .B1(n10343), .B2(keyinput_g73), .C1(n8475), .C2(
        keyinput_g40), .A(n9359), .ZN(n9367) );
  AOI22_X1 U11856 ( .A1(n11693), .A2(keyinput_g46), .B1(keyinput_g21), .B2(
        n9536), .ZN(n9360) );
  OAI221_X1 U11857 ( .B1(n11693), .B2(keyinput_g46), .C1(n9536), .C2(
        keyinput_g21), .A(n9360), .ZN(n9366) );
  INV_X1 U11858 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n9965) );
  XNOR2_X1 U11859 ( .A(n9965), .B(keyinput_g90), .ZN(n9365) );
  XNOR2_X1 U11860 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g127), .ZN(n9363)
         );
  XNOR2_X1 U11861 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n9362)
         );
  XNOR2_X1 U11862 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g108), .ZN(n9361) );
  NAND3_X1 U11863 ( .A1(n9363), .A2(n9362), .A3(n9361), .ZN(n9364) );
  NOR4_X1 U11864 ( .A1(n9367), .A2(n9366), .A3(n9365), .A4(n9364), .ZN(n9379)
         );
  INV_X1 U11865 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11866 ( .A1(n11379), .A2(keyinput_g7), .B1(keyinput_g86), .B2(
        n9969), .ZN(n9368) );
  OAI221_X1 U11867 ( .B1(n11379), .B2(keyinput_g7), .C1(n9969), .C2(
        keyinput_g86), .A(n9368), .ZN(n9377) );
  INV_X1 U11868 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9370) );
  AOI22_X1 U11869 ( .A1(n15520), .A2(keyinput_g106), .B1(n9370), .B2(
        keyinput_g55), .ZN(n9369) );
  OAI221_X1 U11870 ( .B1(n15520), .B2(keyinput_g106), .C1(n9370), .C2(
        keyinput_g55), .A(n9369), .ZN(n9376) );
  XNOR2_X1 U11871 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g109), .ZN(n9374) );
  XNOR2_X1 U11872 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_g116), .ZN(n9373) );
  XNOR2_X1 U11873 ( .A(SI_7_), .B(keyinput_g25), .ZN(n9372) );
  XNOR2_X1 U11874 ( .A(SI_31_), .B(keyinput_g1), .ZN(n9371) );
  NAND4_X1 U11875 ( .A1(n9374), .A2(n9373), .A3(n9372), .A4(n9371), .ZN(n9375)
         );
  NOR3_X1 U11876 ( .A1(n9377), .A2(n9376), .A3(n9375), .ZN(n9378) );
  NAND4_X1 U11877 ( .A1(n9381), .A2(n9380), .A3(n9379), .A4(n9378), .ZN(n9423)
         );
  INV_X1 U11878 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U11879 ( .A1(n11483), .A2(keyinput_g6), .B1(keyinput_g65), .B2(
        n10773), .ZN(n9382) );
  OAI221_X1 U11880 ( .B1(n11483), .B2(keyinput_g6), .C1(n10773), .C2(
        keyinput_g65), .A(n9382), .ZN(n9391) );
  AOI22_X1 U11881 ( .A1(n11219), .A2(keyinput_g8), .B1(keyinput_g9), .B2(
        n10817), .ZN(n9383) );
  OAI221_X1 U11882 ( .B1(n11219), .B2(keyinput_g8), .C1(n10817), .C2(
        keyinput_g9), .A(n9383), .ZN(n9386) );
  XNOR2_X1 U11883 ( .A(n9979), .B(keyinput_g91), .ZN(n9385) );
  XOR2_X1 U11884 ( .A(SI_2_), .B(keyinput_g30), .Z(n9384) );
  OR3_X1 U11885 ( .A1(n9386), .A2(n9385), .A3(n9384), .ZN(n9390) );
  AOI22_X1 U11886 ( .A1(n10345), .A2(keyinput_g12), .B1(n9388), .B2(
        keyinput_g45), .ZN(n9387) );
  OAI221_X1 U11887 ( .B1(n10345), .B2(keyinput_g12), .C1(n9388), .C2(
        keyinput_g45), .A(n9387), .ZN(n9389) );
  NOR3_X1 U11888 ( .A1(n9391), .A2(n9390), .A3(n9389), .ZN(n9421) );
  AOI22_X1 U11889 ( .A1(n10146), .A2(keyinput_g119), .B1(n9393), .B2(
        keyinput_g62), .ZN(n9392) );
  OAI221_X1 U11890 ( .B1(n10146), .B2(keyinput_g119), .C1(n9393), .C2(
        keyinput_g62), .A(n9392), .ZN(n9400) );
  AOI22_X1 U11891 ( .A1(n14779), .A2(keyinput_g33), .B1(n15499), .B2(
        keyinput_g105), .ZN(n9394) );
  OAI221_X1 U11892 ( .B1(n14779), .B2(keyinput_g33), .C1(n15499), .C2(
        keyinput_g105), .A(n9394), .ZN(n9399) );
  INV_X1 U11893 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U11894 ( .A1(n10006), .A2(keyinput_g94), .B1(n9985), .B2(
        keyinput_g85), .ZN(n9395) );
  OAI221_X1 U11895 ( .B1(n10006), .B2(keyinput_g94), .C1(n9985), .C2(
        keyinput_g85), .A(n9395), .ZN(n9398) );
  AOI22_X1 U11896 ( .A1(n8433), .A2(keyinput_g51), .B1(keyinput_g74), .B2(
        n10158), .ZN(n9396) );
  OAI221_X1 U11897 ( .B1(n8433), .B2(keyinput_g51), .C1(n10158), .C2(
        keyinput_g74), .A(n9396), .ZN(n9397) );
  NOR4_X1 U11898 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n9420)
         );
  INV_X1 U11899 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11900 ( .A1(n9983), .A2(keyinput_g83), .B1(n10156), .B2(
        keyinput_g13), .ZN(n9401) );
  OAI221_X1 U11901 ( .B1(n9983), .B2(keyinput_g83), .C1(n10156), .C2(
        keyinput_g13), .A(n9401), .ZN(n9408) );
  INV_X1 U11902 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n10832) );
  INV_X1 U11903 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U11904 ( .A1(n10832), .A2(keyinput_g66), .B1(n11654), .B2(
        keyinput_g58), .ZN(n9402) );
  OAI221_X1 U11905 ( .B1(n10832), .B2(keyinput_g66), .C1(n11654), .C2(
        keyinput_g58), .A(n9402), .ZN(n9407) );
  AOI22_X1 U11906 ( .A1(n12953), .A2(keyinput_g48), .B1(keyinput_g49), .B2(
        n10069), .ZN(n9403) );
  OAI221_X1 U11907 ( .B1(n12953), .B2(keyinput_g48), .C1(n10069), .C2(
        keyinput_g49), .A(n9403), .ZN(n9406) );
  AOI22_X1 U11908 ( .A1(n10415), .A2(keyinput_g11), .B1(keyinput_g120), .B2(
        n10149), .ZN(n9404) );
  OAI221_X1 U11909 ( .B1(n10415), .B2(keyinput_g11), .C1(n10149), .C2(
        keyinput_g120), .A(n9404), .ZN(n9405) );
  NOR4_X1 U11910 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n9405), .ZN(n9419)
         );
  AOI22_X1 U11911 ( .A1(n10574), .A2(keyinput_g70), .B1(n12991), .B2(
        keyinput_g56), .ZN(n9409) );
  OAI221_X1 U11912 ( .B1(n10574), .B2(keyinput_g70), .C1(n12991), .C2(
        keyinput_g56), .A(n9409), .ZN(n9417) );
  INV_X1 U11913 ( .A(SI_30_), .ZN(n13460) );
  AOI22_X1 U11914 ( .A1(n13460), .A2(keyinput_g2), .B1(n12943), .B2(
        keyinput_g47), .ZN(n9410) );
  OAI221_X1 U11915 ( .B1(n13460), .B2(keyinput_g2), .C1(n12943), .C2(
        keyinput_g47), .A(n9410), .ZN(n9416) );
  XNOR2_X1 U11916 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_g41), .ZN(n9414)
         );
  XNOR2_X1 U11917 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g111), .ZN(n9413) );
  XNOR2_X1 U11918 ( .A(n14775), .B(keyinput_g107), .ZN(n9412) );
  XNOR2_X1 U11919 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .ZN(n9411)
         );
  NAND4_X1 U11920 ( .A1(n9414), .A2(n9413), .A3(n9412), .A4(n9411), .ZN(n9415)
         );
  NOR3_X1 U11921 ( .A1(n9417), .A2(n9416), .A3(n9415), .ZN(n9418) );
  NAND4_X1 U11922 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(n9422)
         );
  NOR4_X1 U11923 ( .A1(n9425), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(n9426)
         );
  NOR2_X1 U11924 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  INV_X1 U11925 ( .A(n9742), .ZN(n11425) );
  NOR2_X1 U11926 ( .A1(n9475), .A2(n11425), .ZN(n9744) );
  INV_X1 U11927 ( .A(n9429), .ZN(n10161) );
  INV_X1 U11928 ( .A(n9574), .ZN(n9435) );
  INV_X1 U11929 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9439) );
  NOR2_X1 U11930 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9575) );
  NOR2_X1 U11931 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9442) );
  OAI21_X1 U11932 ( .B1(n10551), .B2(n9447), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9443) );
  MUX2_X1 U11933 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9443), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9449) );
  NAND2_X1 U11934 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  NAND2_X1 U11935 ( .A1(n9451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9453) );
  XNOR2_X1 U11936 ( .A(n9453), .B(n9452), .ZN(n9812) );
  INV_X1 U11937 ( .A(n9571), .ZN(n9454) );
  INV_X2 U11938 ( .A(n9715), .ZN(n13509) );
  NAND2_X1 U11939 ( .A1(n13509), .A2(n6854), .ZN(n9457) );
  XNOR2_X1 U11940 ( .A(n10539), .B(n9457), .ZN(n13575) );
  INV_X2 U11941 ( .A(n13493), .ZN(n13525) );
  NAND2_X1 U11942 ( .A1(n13525), .A2(n15291), .ZN(n13576) );
  NAND2_X1 U11943 ( .A1(n13572), .A2(n13509), .ZN(n9455) );
  AND2_X1 U11944 ( .A1(n13576), .A2(n9455), .ZN(n9456) );
  INV_X1 U11945 ( .A(n10539), .ZN(n9458) );
  NAND2_X1 U11946 ( .A1(n9458), .A2(n9457), .ZN(n9459) );
  NAND2_X1 U11947 ( .A1(n13574), .A2(n9459), .ZN(n9460) );
  XNOR2_X1 U11948 ( .A(n13493), .B(n15282), .ZN(n9461) );
  NAND2_X1 U11949 ( .A1(n13509), .A2(n13703), .ZN(n9462) );
  XNOR2_X1 U11950 ( .A(n9461), .B(n9462), .ZN(n10540) );
  NAND2_X1 U11951 ( .A1(n9460), .A2(n10540), .ZN(n10546) );
  INV_X1 U11952 ( .A(n9461), .ZN(n9463) );
  NAND2_X1 U11953 ( .A1(n9463), .A2(n9462), .ZN(n9464) );
  NAND2_X1 U11954 ( .A1(n10546), .A2(n9464), .ZN(n9474) );
  XNOR2_X1 U11955 ( .A(n13505), .B(n12387), .ZN(n10453) );
  AND2_X1 U11956 ( .A1(n13509), .A2(n13702), .ZN(n9465) );
  NAND2_X1 U11957 ( .A1(n10453), .A2(n9465), .ZN(n10447) );
  INV_X1 U11958 ( .A(n10453), .ZN(n9467) );
  INV_X1 U11959 ( .A(n9465), .ZN(n9466) );
  NAND2_X1 U11960 ( .A1(n9467), .A2(n9466), .ZN(n9468) );
  NAND2_X1 U11961 ( .A1(n10447), .A2(n9468), .ZN(n9473) );
  INV_X1 U11962 ( .A(n9469), .ZN(n9470) );
  INV_X1 U11963 ( .A(n9741), .ZN(n9471) );
  NAND3_X1 U11964 ( .A1(n15343), .A2(n9471), .A3(n15403), .ZN(n9472) );
  OR2_X2 U11965 ( .A1(n9484), .A2(n9472), .ZN(n13653) );
  INV_X1 U11966 ( .A(n10449), .ZN(n10450) );
  AOI211_X1 U11967 ( .C1(n9474), .C2(n9473), .A(n13653), .B(n10450), .ZN(n9487) );
  NAND2_X1 U11968 ( .A1(n9484), .A2(n9479), .ZN(n9477) );
  AND3_X1 U11969 ( .A1(n9475), .A2(n9742), .A3(n12667), .ZN(n9476) );
  NAND2_X1 U11970 ( .A1(n9477), .A2(n9476), .ZN(n10443) );
  NAND2_X1 U11971 ( .A1(n10443), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13674) );
  MUX2_X1 U11972 ( .A(n13649), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n9486) );
  NOR2_X1 U11973 ( .A1(n15292), .A2(n11216), .ZN(n10568) );
  NAND2_X1 U11974 ( .A1(n15343), .A2(n10568), .ZN(n9478) );
  INV_X1 U11975 ( .A(n9479), .ZN(n9480) );
  INV_X1 U11976 ( .A(n13668), .ZN(n13662) );
  AOI22_X1 U11977 ( .A1(n13991), .A2(n13703), .B1(n13988), .B2(n13701), .ZN(
        n10869) );
  NAND2_X1 U11978 ( .A1(n15343), .A2(n9482), .ZN(n9483) );
  OAI22_X1 U11979 ( .A1(n13662), .A2(n15363), .B1(n10869), .B2(n13646), .ZN(
        n9485) );
  OR3_X1 U11980 ( .A1(n9487), .A2(n9486), .A3(n9485), .ZN(P2_U3190) );
  NOR2_X1 U11981 ( .A1(n10090), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12136) );
  INV_X2 U11982 ( .A(n12136), .ZN(n14150) );
  INV_X1 U11983 ( .A(n10112), .ZN(n9516) );
  AND2_X1 U11984 ( .A1(n10090), .A2(P2_U3088), .ZN(n14138) );
  INV_X2 U11985 ( .A(n14138), .ZN(n14152) );
  OAI222_X1 U11986 ( .A1(P2_U3088), .A2(n15152), .B1(n14150), .B2(n9516), .C1(
        n9488), .C2(n14152), .ZN(P2_U3325) );
  NAND2_X1 U11987 ( .A1(n11804), .A2(P3_U3151), .ZN(n13471) );
  INV_X1 U11988 ( .A(SI_7_), .ZN(n9491) );
  AND2_X1 U11989 ( .A1(n10090), .A2(P3_U3151), .ZN(n13455) );
  INV_X2 U11990 ( .A(n13455), .ZN(n13468) );
  INV_X1 U11991 ( .A(n9489), .ZN(n9490) );
  OAI222_X1 U11992 ( .A1(P3_U3151), .A2(n15470), .B1(n13471), .B2(n9491), .C1(
        n13468), .C2(n9490), .ZN(P3_U3288) );
  INV_X1 U11993 ( .A(SI_3_), .ZN(n9494) );
  INV_X1 U11994 ( .A(n9492), .ZN(n9493) );
  OAI222_X1 U11995 ( .A1(P3_U3151), .A2(n10062), .B1(n13471), .B2(n9494), .C1(
        n13468), .C2(n9493), .ZN(P3_U3292) );
  INV_X1 U11996 ( .A(SI_4_), .ZN(n9497) );
  INV_X1 U11997 ( .A(n9495), .ZN(n9496) );
  OAI222_X1 U11998 ( .A1(P3_U3151), .A2(n15437), .B1(n13471), .B2(n9497), .C1(
        n13468), .C2(n9496), .ZN(P3_U3291) );
  INV_X1 U11999 ( .A(SI_5_), .ZN(n9500) );
  INV_X1 U12000 ( .A(n9498), .ZN(n9499) );
  OAI222_X1 U12001 ( .A1(P3_U3151), .A2(n10646), .B1(n13471), .B2(n9500), .C1(
        n13468), .C2(n9499), .ZN(P3_U3290) );
  OAI222_X1 U12002 ( .A1(P2_U3088), .A2(n13711), .B1(n14150), .B2(n10091), 
        .C1(n9501), .C2(n14152), .ZN(P2_U3326) );
  INV_X1 U12003 ( .A(n10263), .ZN(n9507) );
  INV_X1 U12004 ( .A(n9853), .ZN(n15165) );
  OAI222_X1 U12005 ( .A1(n14152), .A2(n9502), .B1(n14150), .B2(n9507), .C1(
        P2_U3088), .C2(n15165), .ZN(P2_U3324) );
  NAND2_X1 U12006 ( .A1(n11804), .A2(P1_U3086), .ZN(n14771) );
  INV_X1 U12007 ( .A(n14771), .ZN(n11440) );
  INV_X1 U12008 ( .A(n11440), .ZN(n14764) );
  AND2_X1 U12009 ( .A1(n10090), .A2(P1_U3086), .ZN(n14758) );
  INV_X2 U12010 ( .A(n14758), .ZN(n14768) );
  NAND2_X1 U12011 ( .A1(n9503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9504) );
  MUX2_X1 U12012 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9504), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9505) );
  INV_X1 U12013 ( .A(n14324), .ZN(n9506) );
  OAI222_X1 U12014 ( .A1(n14764), .A2(n9508), .B1(n14768), .B2(n9507), .C1(
        P1_U3086), .C2(n9506), .ZN(P1_U3352) );
  INV_X1 U12015 ( .A(n9509), .ZN(n9548) );
  NAND2_X1 U12016 ( .A1(n9548), .A2(n10788), .ZN(n9510) );
  OAI21_X1 U12017 ( .B1(n9548), .B2(n9511), .A(n9510), .ZN(P3_U3377) );
  NAND2_X1 U12018 ( .A1(n10172), .A2(n9548), .ZN(n9512) );
  OAI21_X1 U12019 ( .B1(n9548), .B2(n8927), .A(n9512), .ZN(P3_U3376) );
  OR2_X1 U12020 ( .A1(n9513), .A2(n10407), .ZN(n9514) );
  XNOR2_X1 U12021 ( .A(n9514), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10113) );
  INV_X1 U12022 ( .A(n10113), .ZN(n9611) );
  OAI222_X1 U12023 ( .A1(P1_U3086), .A2(n9611), .B1(n14768), .B2(n9516), .C1(
        n9515), .C2(n14764), .ZN(P1_U3353) );
  INV_X1 U12024 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U12025 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14775), .ZN(n9517) );
  INV_X1 U12026 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10093) );
  OAI222_X1 U12027 ( .A1(P1_U3086), .A2(n10094), .B1(n14768), .B2(n10091), 
        .C1(n10093), .C2(n14764), .ZN(P1_U3354) );
  CLKBUF_X1 U12028 ( .A(n13471), .Z(n11518) );
  INV_X1 U12029 ( .A(SI_10_), .ZN(n9520) );
  OAI222_X1 U12030 ( .A1(P3_U3151), .A2(n13091), .B1(n11518), .B2(n9520), .C1(
        n13468), .C2(n9519), .ZN(P3_U3285) );
  OAI222_X1 U12031 ( .A1(n13468), .A2(n9522), .B1(n11518), .B2(n9521), .C1(
        P3_U3151), .C2(n15487), .ZN(P3_U3287) );
  INV_X1 U12032 ( .A(SI_9_), .ZN(n9525) );
  INV_X1 U12033 ( .A(n9523), .ZN(n9524) );
  OAI222_X1 U12034 ( .A1(P3_U3151), .A2(n15510), .B1(n11518), .B2(n9525), .C1(
        n13468), .C2(n9524), .ZN(P3_U3286) );
  OAI222_X1 U12035 ( .A1(n13468), .A2(n9527), .B1(n11518), .B2(n9526), .C1(
        P3_U3151), .C2(n6680), .ZN(P3_U3294) );
  INV_X1 U12036 ( .A(n10420), .ZN(n9534) );
  NAND2_X1 U12037 ( .A1(n9529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9528) );
  MUX2_X1 U12038 ( .A(n9528), .B(P1_IR_REG_31__SCAN_IN), .S(n9530), .Z(n9532)
         );
  INV_X1 U12039 ( .A(n9529), .ZN(n9531) );
  NAND2_X1 U12040 ( .A1(n9531), .A2(n9530), .ZN(n9551) );
  NAND2_X1 U12041 ( .A1(n9532), .A2(n9551), .ZN(n9626) );
  OAI222_X1 U12042 ( .A1(n14764), .A2(n9533), .B1(n14768), .B2(n9534), .C1(
        P1_U3086), .C2(n9626), .ZN(P1_U3351) );
  INV_X1 U12043 ( .A(n9854), .ZN(n10050) );
  OAI222_X1 U12044 ( .A1(n14152), .A2(n9535), .B1(n14150), .B2(n9534), .C1(
        P2_U3088), .C2(n10050), .ZN(P2_U3323) );
  OAI222_X1 U12045 ( .A1(n15528), .A2(P3_U3151), .B1(n13468), .B2(n9537), .C1(
        n11518), .C2(n9536), .ZN(P3_U3284) );
  OAI222_X1 U12046 ( .A1(P3_U3151), .A2(n15459), .B1(n13468), .B2(n9539), .C1(
        n9538), .C2(n11518), .ZN(P3_U3289) );
  OAI222_X1 U12047 ( .A1(n11518), .A2(n9541), .B1(n13468), .B2(n9540), .C1(
        n15546), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12048 ( .A(n10580), .ZN(n9545) );
  NAND2_X1 U12049 ( .A1(n9551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9542) );
  XNOR2_X1 U12050 ( .A(n9542), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10581) );
  INV_X1 U12051 ( .A(n10581), .ZN(n9543) );
  OAI222_X1 U12052 ( .A1(n14764), .A2(n9544), .B1(n14768), .B2(n9545), .C1(
        P1_U3086), .C2(n9543), .ZN(P1_U3350) );
  INV_X1 U12053 ( .A(n9855), .ZN(n15182) );
  OAI222_X1 U12054 ( .A1(n14152), .A2(n9546), .B1(n14150), .B2(n9545), .C1(
        P2_U3088), .C2(n15182), .ZN(P2_U3322) );
  AND2_X1 U12055 ( .A1(n9549), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12056 ( .A1(n9549), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12057 ( .A1(n9549), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12058 ( .A1(n9549), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12059 ( .A1(n9549), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12060 ( .A1(n9549), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12061 ( .A1(n9549), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12062 ( .A1(n9549), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12063 ( .A1(n9549), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12064 ( .A1(n9549), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12065 ( .A1(n9549), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12066 ( .A1(n9549), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12067 ( .A1(n9549), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12068 ( .A1(n9549), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12069 ( .A1(n9549), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12070 ( .A1(n9549), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12071 ( .A1(n9549), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12072 ( .A1(n9549), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12073 ( .A1(n9549), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12074 ( .A1(n9549), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12075 ( .A1(n9549), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12076 ( .A1(n9549), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12077 ( .A1(n9549), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12078 ( .A1(n9549), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12079 ( .A1(n9549), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12080 ( .A1(n9549), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12081 ( .A1(n9549), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12082 ( .A1(n9549), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12083 ( .A1(n9549), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12084 ( .A1(n9549), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  INV_X1 U12085 ( .A(n9922), .ZN(n9863) );
  INV_X1 U12086 ( .A(n10712), .ZN(n9557) );
  OAI222_X1 U12087 ( .A1(P2_U3088), .A2(n9863), .B1(n14150), .B2(n9557), .C1(
        n9550), .C2(n14152), .ZN(P2_U3321) );
  INV_X1 U12088 ( .A(n9551), .ZN(n9553) );
  INV_X1 U12089 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U12090 ( .A1(n9553), .A2(n9552), .ZN(n9555) );
  NAND2_X1 U12091 ( .A1(n9555), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9554) );
  MUX2_X1 U12092 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9554), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9556) );
  AND2_X1 U12093 ( .A1(n9556), .A2(n9596), .ZN(n10713) );
  INV_X1 U12094 ( .A(n10713), .ZN(n9683) );
  OAI222_X1 U12095 ( .A1(n14764), .A2(n9558), .B1(n14768), .B2(n9557), .C1(
        n9683), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12096 ( .A(n10904), .ZN(n9561) );
  INV_X1 U12097 ( .A(n9924), .ZN(n15197) );
  OAI222_X1 U12098 ( .A1(n14152), .A2(n9559), .B1(n14150), .B2(n9561), .C1(
        P2_U3088), .C2(n15197), .ZN(P2_U3320) );
  NAND2_X1 U12099 ( .A1(n9596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9560) );
  XNOR2_X1 U12100 ( .A(n9560), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10905) );
  INV_X1 U12101 ( .A(n10905), .ZN(n9659) );
  OAI222_X1 U12102 ( .A1(n14764), .A2(n9562), .B1(n14768), .B2(n9561), .C1(
        P1_U3086), .C2(n9659), .ZN(P1_U3348) );
  OAI222_X1 U12103 ( .A1(P3_U3151), .A2(n15564), .B1(n11518), .B2(n9564), .C1(
        n13468), .C2(n9563), .ZN(P3_U3282) );
  INV_X1 U12104 ( .A(n9568), .ZN(n11644) );
  NAND3_X1 U12105 ( .A1(n11644), .A2(n12838), .A3(P1_B_REG_SCAN_IN), .ZN(n9566) );
  INV_X1 U12106 ( .A(P1_B_REG_SCAN_IN), .ZN(n14399) );
  AOI21_X1 U12107 ( .B1(n9568), .B2(n14399), .A(n14769), .ZN(n9565) );
  NAND2_X1 U12108 ( .A1(n9566), .A2(n9565), .ZN(n9768) );
  NAND2_X1 U12109 ( .A1(n14161), .A2(n9768), .ZN(n15075) );
  INV_X1 U12110 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9570) );
  INV_X1 U12111 ( .A(n9754), .ZN(n9569) );
  AOI22_X1 U12112 ( .A1(n15075), .A2(n9570), .B1(n9569), .B2(n9571), .ZN(
        P1_U3445) );
  INV_X1 U12113 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U12114 ( .A1(n12838), .A2(n14769), .ZN(n9756) );
  INV_X1 U12115 ( .A(n9756), .ZN(n9572) );
  AOI22_X1 U12116 ( .A1(n15075), .A2(n9573), .B1(n9572), .B2(n9571), .ZN(
        P1_U3446) );
  INV_X1 U12117 ( .A(n9812), .ZN(n9579) );
  NAND2_X1 U12118 ( .A1(n9579), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12132) );
  NAND2_X1 U12119 ( .A1(n9803), .A2(n12132), .ZN(n9589) );
  NAND2_X1 U12120 ( .A1(n14773), .A2(n12092), .ZN(n11915) );
  OR2_X1 U12121 ( .A1(n11915), .A2(n9579), .ZN(n9586) );
  NAND2_X1 U12122 ( .A1(n9586), .A2(n10092), .ZN(n9587) );
  AND2_X1 U12123 ( .A1(n9589), .A2(n9587), .ZN(n14343) );
  INV_X1 U12124 ( .A(n9587), .ZN(n9588) );
  NAND2_X1 U12125 ( .A1(n9589), .A2(n9588), .ZN(n9629) );
  INV_X1 U12126 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9797) );
  INV_X1 U12127 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U12128 ( .A1(n6679), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9592) );
  OR2_X1 U12129 ( .A1(n6688), .A2(n9592), .ZN(n9945) );
  AOI21_X1 U12130 ( .B1(n6679), .B2(n9797), .A(n9945), .ZN(n9593) );
  XNOR2_X1 U12131 ( .A(n9593), .B(n7302), .ZN(n9594) );
  AOI22_X1 U12132 ( .A1(n9631), .A2(n9594), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9595) );
  OAI21_X1 U12133 ( .B1(n15042), .B2(n7100), .A(n9595), .ZN(P1_U3243) );
  INV_X1 U12134 ( .A(n10909), .ZN(n9599) );
  NAND2_X1 U12135 ( .A1(n9597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9603) );
  XNOR2_X1 U12136 ( .A(n9603), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10910) );
  INV_X1 U12137 ( .A(n10910), .ZN(n9663) );
  OAI222_X1 U12138 ( .A1(n14764), .A2(n9598), .B1(n14768), .B2(n9599), .C1(
        P1_U3086), .C2(n9663), .ZN(P1_U3347) );
  INV_X1 U12139 ( .A(n9925), .ZN(n10037) );
  OAI222_X1 U12140 ( .A1(n14152), .A2(n9600), .B1(n14150), .B2(n9599), .C1(
        P2_U3088), .C2(n10037), .ZN(P2_U3319) );
  INV_X1 U12141 ( .A(n10353), .ZN(n9941) );
  OAI222_X1 U12142 ( .A1(P2_U3088), .A2(n9941), .B1(n14150), .B2(n10919), .C1(
        n9601), .C2(n14152), .ZN(P2_U3318) );
  NAND2_X1 U12143 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  XNOR2_X1 U12144 ( .A(n9821), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10920) );
  INV_X1 U12145 ( .A(n10920), .ZN(n9664) );
  OAI222_X1 U12146 ( .A1(n14764), .A2(n9605), .B1(n14768), .B2(n10919), .C1(
        n9664), .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U12147 ( .A1(P3_U3151), .A2(n15583), .B1(n11518), .B2(n9607), .C1(
        n13468), .C2(n9606), .ZN(P3_U3281) );
  CLKBUF_X2 U12148 ( .A(P1_U4016), .Z(n14319) );
  NOR2_X1 U12149 ( .A1(n14343), .A2(n14319), .ZN(P1_U3085) );
  INV_X1 U12150 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11122) );
  MUX2_X1 U12151 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11122), .S(n10113), .Z(
        n9610) );
  INV_X1 U12152 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11127) );
  MUX2_X1 U12153 ( .A(n11127), .B(P1_REG2_REG_1__SCAN_IN), .S(n10094), .Z(
        n9608) );
  AND2_X1 U12154 ( .A1(n14775), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U12155 ( .A1(n9608), .A2(n9684), .ZN(n9949) );
  OR2_X1 U12156 ( .A1(n10094), .A2(n11127), .ZN(n9948) );
  NAND2_X1 U12157 ( .A1(n9949), .A2(n9948), .ZN(n9609) );
  NAND2_X1 U12158 ( .A1(n9610), .A2(n9609), .ZN(n9952) );
  INV_X1 U12159 ( .A(n9952), .ZN(n14330) );
  NOR2_X1 U12160 ( .A1(n9611), .A2(n11122), .ZN(n14329) );
  INV_X1 U12161 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U12162 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10122), .S(n14324), .Z(
        n14331) );
  OAI21_X1 U12163 ( .B1(n14330), .B2(n14329), .A(n14331), .ZN(n14338) );
  NAND2_X1 U12164 ( .A1(n14324), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14337) );
  INV_X1 U12165 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10478) );
  MUX2_X1 U12166 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10478), .S(n9626), .Z(
        n14336) );
  AOI21_X1 U12167 ( .B1(n14338), .B2(n14337), .A(n14336), .ZN(n14340) );
  NOR2_X1 U12168 ( .A1(n9626), .A2(n10478), .ZN(n9732) );
  INV_X1 U12169 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11147) );
  MUX2_X1 U12170 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11147), .S(n10581), .Z(
        n9731) );
  OAI21_X1 U12171 ( .B1(n14340), .B2(n9732), .A(n9731), .ZN(n9730) );
  NAND2_X1 U12172 ( .A1(n10581), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9676) );
  INV_X1 U12173 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9612) );
  MUX2_X1 U12174 ( .A(n9612), .B(P1_REG2_REG_6__SCAN_IN), .S(n10713), .Z(n9675) );
  AOI21_X1 U12175 ( .B1(n9730), .B2(n9676), .A(n9675), .ZN(n9678) );
  NOR2_X1 U12176 ( .A1(n9683), .A2(n9612), .ZN(n9652) );
  INV_X1 U12177 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9613) );
  MUX2_X1 U12178 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9613), .S(n10905), .Z(n9614) );
  OAI21_X1 U12179 ( .B1(n9678), .B2(n9652), .A(n9614), .ZN(n9655) );
  NAND2_X1 U12180 ( .A1(n10905), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9618) );
  INV_X1 U12181 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9615) );
  MUX2_X1 U12182 ( .A(n9615), .B(P1_REG2_REG_8__SCAN_IN), .S(n10910), .Z(n9617) );
  AOI21_X1 U12183 ( .B1(n9655), .B2(n9618), .A(n9617), .ZN(n9700) );
  NOR2_X1 U12184 ( .A1(n6688), .A2(n6679), .ZN(n9616) );
  NAND3_X1 U12185 ( .A1(n9655), .A2(n9618), .A3(n9617), .ZN(n9619) );
  NAND2_X1 U12186 ( .A1(n14389), .A2(n9619), .ZN(n9636) );
  INV_X1 U12187 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15144) );
  MUX2_X1 U12188 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n15144), .S(n10910), .Z(
        n9628) );
  INV_X1 U12189 ( .A(n9626), .ZN(n14344) );
  INV_X1 U12190 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10121) );
  MUX2_X1 U12191 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10121), .S(n14324), .Z(
        n9625) );
  INV_X1 U12192 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10107) );
  MUX2_X1 U12193 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10107), .S(n10113), .Z(
        n9623) );
  INV_X1 U12194 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9806) );
  MUX2_X1 U12195 ( .A(n9806), .B(P1_REG1_REG_1__SCAN_IN), .S(n10094), .Z(n9621) );
  AND2_X1 U12196 ( .A1(n14775), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U12197 ( .A1(n9621), .A2(n9620), .ZN(n9954) );
  OR2_X1 U12198 ( .A1(n10094), .A2(n9806), .ZN(n9953) );
  NAND2_X1 U12199 ( .A1(n9954), .A2(n9953), .ZN(n9622) );
  NAND2_X1 U12200 ( .A1(n10113), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U12201 ( .A1(n14326), .A2(n14325), .ZN(n9624) );
  NAND2_X1 U12202 ( .A1(n9625), .A2(n9624), .ZN(n14347) );
  NAND2_X1 U12203 ( .A1(n14324), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14346) );
  INV_X1 U12204 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15136) );
  MUX2_X1 U12205 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15136), .S(n9626), .Z(
        n14348) );
  AOI21_X1 U12206 ( .B1(n14347), .B2(n14346), .A(n14348), .ZN(n14345) );
  INV_X1 U12207 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15138) );
  MUX2_X1 U12208 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15138), .S(n10581), .Z(
        n9726) );
  NAND2_X1 U12209 ( .A1(n9725), .A2(n9726), .ZN(n9724) );
  OAI21_X1 U12210 ( .B1(n10581), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9724), .ZN(
        n9674) );
  INV_X1 U12211 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15140) );
  MUX2_X1 U12212 ( .A(n15140), .B(P1_REG1_REG_6__SCAN_IN), .S(n10713), .Z(
        n9673) );
  NOR2_X1 U12213 ( .A1(n9674), .A2(n9673), .ZN(n9672) );
  INV_X1 U12214 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15142) );
  MUX2_X1 U12215 ( .A(n15142), .B(P1_REG1_REG_7__SCAN_IN), .S(n10905), .Z(
        n9647) );
  NOR2_X1 U12216 ( .A1(n9648), .A2(n9647), .ZN(n9646) );
  AOI21_X1 U12217 ( .B1(n10905), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9646), .ZN(
        n9627) );
  NAND2_X1 U12218 ( .A1(n9627), .A2(n9628), .ZN(n9695) );
  OAI21_X1 U12219 ( .B1(n9628), .B2(n9627), .A(n9695), .ZN(n9630) );
  INV_X1 U12220 ( .A(n6679), .ZN(n12128) );
  NAND2_X1 U12221 ( .A1(n9630), .A2(n14383), .ZN(n9635) );
  AND2_X1 U12222 ( .A1(n9631), .A2(n6688), .ZN(n14387) );
  NAND2_X1 U12223 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11321) );
  OAI21_X1 U12224 ( .B1(n15042), .B2(n9632), .A(n11321), .ZN(n9633) );
  AOI21_X1 U12225 ( .B1(n10910), .B2(n14387), .A(n9633), .ZN(n9634) );
  OAI211_X1 U12226 ( .C1(n9700), .C2(n9636), .A(n9635), .B(n9634), .ZN(
        P1_U3251) );
  INV_X1 U12227 ( .A(n13101), .ZN(n14822) );
  INV_X1 U12228 ( .A(n9637), .ZN(n9639) );
  OAI222_X1 U12229 ( .A1(n14822), .A2(P3_U3151), .B1(n13468), .B2(n9639), .C1(
        n9638), .C2(n11518), .ZN(P3_U3280) );
  INV_X1 U12230 ( .A(n10933), .ZN(n9644) );
  INV_X1 U12231 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12232 ( .A1(n9821), .A2(n9640), .ZN(n9641) );
  NAND2_X1 U12233 ( .A1(n9641), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9642) );
  XNOR2_X1 U12234 ( .A(n9642), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10934) );
  INV_X1 U12235 ( .A(n10934), .ZN(n9827) );
  OAI222_X1 U12236 ( .A1(n14764), .A2(n9643), .B1(n14768), .B2(n9644), .C1(
        P1_U3086), .C2(n9827), .ZN(P1_U3345) );
  INV_X1 U12237 ( .A(n10380), .ZN(n10361) );
  OAI222_X1 U12238 ( .A1(n14152), .A2(n9645), .B1(n14150), .B2(n9644), .C1(
        P2_U3088), .C2(n10361), .ZN(P2_U3317) );
  NAND2_X1 U12239 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11066) );
  AOI211_X1 U12240 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n15036), .ZN(n9649)
         );
  INV_X1 U12241 ( .A(n9649), .ZN(n9650) );
  NAND2_X1 U12242 ( .A1(n11066), .A2(n9650), .ZN(n9651) );
  AOI21_X1 U12243 ( .B1(n14343), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9651), .ZN(
        n9658) );
  INV_X1 U12244 ( .A(n9652), .ZN(n9654) );
  MUX2_X1 U12245 ( .A(n9613), .B(P1_REG2_REG_7__SCAN_IN), .S(n10905), .Z(n9653) );
  NAND2_X1 U12246 ( .A1(n9654), .A2(n9653), .ZN(n9656) );
  OAI211_X1 U12247 ( .C1(n9678), .C2(n9656), .A(n14389), .B(n9655), .ZN(n9657)
         );
  OAI211_X1 U12248 ( .C1(n15038), .C2(n9659), .A(n9658), .B(n9657), .ZN(
        P1_U3250) );
  INV_X1 U12249 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15146) );
  NAND2_X1 U12250 ( .A1(n9663), .A2(n15144), .ZN(n9693) );
  MUX2_X1 U12251 ( .A(n15146), .B(P1_REG1_REG_9__SCAN_IN), .S(n10920), .Z(
        n9694) );
  AOI21_X1 U12252 ( .B1(n15146), .B2(n9664), .A(n9697), .ZN(n9662) );
  INV_X1 U12253 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9660) );
  MUX2_X1 U12254 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9660), .S(n10934), .Z(
        n9661) );
  NAND2_X1 U12255 ( .A1(n9662), .A2(n9661), .ZN(n9826) );
  OAI211_X1 U12256 ( .C1(n9662), .C2(n9661), .A(n9826), .B(n14383), .ZN(n9671)
         );
  NAND2_X1 U12257 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11577)
         );
  INV_X1 U12258 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9665) );
  NOR2_X1 U12259 ( .A1(n9663), .A2(n9615), .ZN(n9699) );
  MUX2_X1 U12260 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9665), .S(n10920), .Z(n9698) );
  OAI21_X1 U12261 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9706) );
  OAI21_X1 U12262 ( .B1(n9665), .B2(n9664), .A(n9706), .ZN(n9667) );
  INV_X1 U12263 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10937) );
  MUX2_X1 U12264 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10937), .S(n10934), .Z(
        n9666) );
  NAND2_X1 U12265 ( .A1(n9667), .A2(n9666), .ZN(n9833) );
  OAI211_X1 U12266 ( .C1(n9667), .C2(n9666), .A(n14389), .B(n9833), .ZN(n9668)
         );
  NAND2_X1 U12267 ( .A1(n11577), .A2(n9668), .ZN(n9669) );
  AOI21_X1 U12268 ( .B1(n14343), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9669), .ZN(
        n9670) );
  OAI211_X1 U12269 ( .C1(n15038), .C2(n9827), .A(n9671), .B(n9670), .ZN(
        P1_U3253) );
  AOI211_X1 U12270 ( .C1(n9674), .C2(n9673), .A(n9672), .B(n15036), .ZN(n9680)
         );
  AND3_X1 U12271 ( .A1(n9730), .A2(n9676), .A3(n9675), .ZN(n9677) );
  NOR3_X1 U12272 ( .A1(n15034), .A2(n9678), .A3(n9677), .ZN(n9679) );
  NOR2_X1 U12273 ( .A1(n9680), .A2(n9679), .ZN(n9682) );
  AND2_X1 U12274 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10730) );
  AOI21_X1 U12275 ( .B1(n14343), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10730), .ZN(
        n9681) );
  OAI211_X1 U12276 ( .C1(n9683), .C2(n15038), .A(n9682), .B(n9681), .ZN(
        P1_U3249) );
  INV_X1 U12277 ( .A(n9684), .ZN(n9944) );
  MUX2_X1 U12278 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n11127), .S(n10094), .Z(
        n9686) );
  INV_X1 U12279 ( .A(n9949), .ZN(n9685) );
  AOI211_X1 U12280 ( .C1(n9944), .C2(n9686), .A(n9685), .B(n15034), .ZN(n9690)
         );
  MUX2_X1 U12281 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9806), .S(n10094), .Z(n9687) );
  OAI21_X1 U12282 ( .B1(n9797), .B2(n7302), .A(n9687), .ZN(n9688) );
  AND3_X1 U12283 ( .A1(n14383), .A2(n9954), .A3(n9688), .ZN(n9689) );
  NOR2_X1 U12284 ( .A1(n9690), .A2(n9689), .ZN(n9692) );
  AOI22_X1 U12285 ( .A1(n14343), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9691) );
  OAI211_X1 U12286 ( .C1(n10094), .C2(n15038), .A(n9692), .B(n9691), .ZN(
        P1_U3244) );
  AND3_X1 U12287 ( .A1(n9695), .A2(n9694), .A3(n9693), .ZN(n9696) );
  OAI21_X1 U12288 ( .B1(n9697), .B2(n9696), .A(n14383), .ZN(n9709) );
  NOR3_X1 U12289 ( .A1(n9700), .A2(n9699), .A3(n9698), .ZN(n9701) );
  NOR2_X1 U12290 ( .A1(n9701), .A2(n15034), .ZN(n9707) );
  NAND2_X1 U12291 ( .A1(n14387), .A2(n10920), .ZN(n9703) );
  NAND2_X1 U12292 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9702) );
  OAI211_X1 U12293 ( .C1(n9704), .C2(n15042), .A(n9703), .B(n9702), .ZN(n9705)
         );
  AOI21_X1 U12294 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9708) );
  NAND2_X1 U12295 ( .A1(n9709), .A2(n9708), .ZN(P1_U3252) );
  INV_X1 U12296 ( .A(n13103), .ZN(n14840) );
  OAI222_X1 U12297 ( .A1(P3_U3151), .A2(n14840), .B1(n11518), .B2(n9711), .C1(
        n13468), .C2(n9710), .ZN(P3_U3279) );
  XNOR2_X1 U12298 ( .A(n9712), .B(n9713), .ZN(n15286) );
  NAND2_X1 U12299 ( .A1(n10670), .A2(n15282), .ZN(n9714) );
  NAND2_X1 U12300 ( .A1(n9715), .A2(n9714), .ZN(n9716) );
  NOR2_X1 U12301 ( .A1(n9716), .A2(n10863), .ZN(n15284) );
  INV_X1 U12302 ( .A(n15284), .ZN(n9717) );
  OAI21_X1 U12303 ( .B1(n10538), .B2(n15403), .A(n9717), .ZN(n9722) );
  XNOR2_X1 U12304 ( .A(n12611), .B(n9718), .ZN(n9720) );
  AOI22_X1 U12305 ( .A1(n13991), .A2(n6854), .B1(n13988), .B2(n13702), .ZN(
        n10537) );
  INV_X1 U12306 ( .A(n10537), .ZN(n9719) );
  AOI21_X1 U12307 ( .B1(n9720), .B2(n15293), .A(n9719), .ZN(n15290) );
  INV_X1 U12308 ( .A(n15290), .ZN(n9721) );
  AOI211_X1 U12309 ( .C1(n15286), .C2(n15390), .A(n9722), .B(n9721), .ZN(
        n15357) );
  NAND2_X1 U12310 ( .A1(n15424), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9723) );
  OAI21_X1 U12311 ( .B1(n15357), .B2(n15424), .A(n9723), .ZN(P2_U3501) );
  OAI21_X1 U12312 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9737) );
  NAND2_X1 U12313 ( .A1(n14387), .A2(n10581), .ZN(n9728) );
  NAND2_X1 U12314 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9727) );
  OAI211_X1 U12315 ( .C1(n9729), .C2(n15042), .A(n9728), .B(n9727), .ZN(n9736)
         );
  INV_X1 U12316 ( .A(n9730), .ZN(n9734) );
  NOR3_X1 U12317 ( .A1(n14340), .A2(n9732), .A3(n9731), .ZN(n9733) );
  NOR3_X1 U12318 ( .A1(n15034), .A2(n9734), .A3(n9733), .ZN(n9735) );
  AOI211_X1 U12319 ( .C1(n14383), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9738)
         );
  INV_X1 U12320 ( .A(n9738), .ZN(P1_U3248) );
  INV_X1 U12321 ( .A(n10948), .ZN(n9823) );
  INV_X1 U12322 ( .A(n11081), .ZN(n11073) );
  OAI222_X1 U12323 ( .A1(n14152), .A2(n9739), .B1(n14150), .B2(n9823), .C1(
        P2_U3088), .C2(n11073), .ZN(P2_U3316) );
  AOI21_X1 U12324 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9743) );
  OR2_X1 U12325 ( .A1(n9744), .A2(n9743), .ZN(n9751) );
  NOR2_X1 U12326 ( .A1(n8293), .A2(P2_U3088), .ZN(n14137) );
  NAND2_X1 U12327 ( .A1(n9745), .A2(n14141), .ZN(n15214) );
  INV_X1 U12328 ( .A(n14141), .ZN(n12668) );
  INV_X1 U12329 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U12330 ( .A1(n15274), .A2(n9746), .ZN(n9747) );
  AND2_X1 U12331 ( .A1(n9751), .A2(n8293), .ZN(n15151) );
  OAI211_X1 U12332 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15214), .A(n9747), .B(
        n15265), .ZN(n9748) );
  INV_X1 U12333 ( .A(n9748), .ZN(n9750) );
  AOI22_X1 U12334 ( .A1(n15270), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15274), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9749) );
  MUX2_X1 U12335 ( .A(n9750), .B(n9749), .S(n13713), .Z(n9753) );
  NOR2_X2 U12336 ( .A1(n9751), .A2(P2_U3088), .ZN(n15266) );
  AOI22_X1 U12337 ( .A1(n15266), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9752) );
  NAND2_X1 U12338 ( .A1(n9753), .A2(n9752), .ZN(P2_U3214) );
  OR2_X1 U12339 ( .A1(n9768), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U12340 ( .A1(n9757), .A2(n9756), .ZN(n10214) );
  INV_X1 U12341 ( .A(n10214), .ZN(n9769) );
  NOR4_X1 U12342 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9766) );
  NOR4_X1 U12343 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9765) );
  OR4_X1 U12344 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9763) );
  NOR4_X1 U12345 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9761) );
  NOR4_X1 U12346 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9760) );
  NOR4_X1 U12347 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9759) );
  NOR4_X1 U12348 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9758) );
  NAND4_X1 U12349 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(n9762)
         );
  NOR4_X1 U12350 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9763), .A4(n9762), .ZN(n9764) );
  AND3_X1 U12351 ( .A1(n9766), .A2(n9765), .A3(n9764), .ZN(n9767) );
  NAND3_X1 U12352 ( .A1(n10470), .A2(n9769), .A3(n9804), .ZN(n9801) );
  NAND2_X1 U12353 ( .A1(n9770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U12354 ( .A1(n9772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U12355 ( .A1(n15055), .A2(n14390), .ZN(n10460) );
  NAND2_X1 U12356 ( .A1(n9801), .A2(n10460), .ZN(n14162) );
  NAND2_X1 U12357 ( .A1(n12089), .A2(n11166), .ZN(n9802) );
  INV_X1 U12358 ( .A(n9802), .ZN(n9774) );
  NOR2_X1 U12359 ( .A1(n9803), .A2(n15126), .ZN(n9775) );
  NAND2_X1 U12360 ( .A1(n10090), .A2(SI_0_), .ZN(n9777) );
  XNOR2_X1 U12361 ( .A(n9777), .B(n9776), .ZN(n14774) );
  MUX2_X1 U12362 ( .A(n7302), .B(n14774), .S(n10092), .Z(n10238) );
  AND2_X4 U12363 ( .A1(n9792), .A2(n11016), .ZN(n12804) );
  XNOR2_X2 U12364 ( .A(n9779), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U12365 ( .A1(n6674), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9790) );
  NAND2_X4 U12366 ( .A1(n9784), .A2(n9786), .ZN(n11900) );
  INV_X1 U12367 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9783) );
  INV_X2 U12368 ( .A(n9784), .ZN(n14762) );
  INV_X1 U12369 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9785) );
  OR2_X1 U12370 ( .A1(n10120), .A2(n9785), .ZN(n9788) );
  NAND2_X4 U12371 ( .A1(n14762), .A2(n9786), .ZN(n11902) );
  INV_X1 U12372 ( .A(n9813), .ZN(n9791) );
  INV_X1 U12373 ( .A(n10238), .ZN(n10250) );
  NAND2_X1 U12374 ( .A1(n14320), .A2(n11309), .ZN(n9796) );
  NAND2_X1 U12375 ( .A1(n12804), .A2(n10250), .ZN(n9795) );
  OAI211_X1 U12376 ( .C1(n9797), .C2(n9813), .A(n9796), .B(n9795), .ZN(n10085)
         );
  AND2_X1 U12377 ( .A1(n9799), .A2(n10085), .ZN(n10089) );
  INV_X1 U12378 ( .A(n10089), .ZN(n9798) );
  OAI21_X1 U12379 ( .B1(n9799), .B2(n10085), .A(n9798), .ZN(n9943) );
  NAND3_X1 U12380 ( .A1(n14161), .A2(n11915), .A3(n15126), .ZN(n9800) );
  INV_X1 U12381 ( .A(n11915), .ZN(n10119) );
  AND2_X1 U12382 ( .A1(n10119), .A2(n9802), .ZN(n9814) );
  NOR2_X1 U12383 ( .A1(n9803), .A2(n9814), .ZN(n12129) );
  NAND2_X1 U12384 ( .A1(n12129), .A2(n9804), .ZN(n10216) );
  OR2_X1 U12385 ( .A1(n10216), .A2(n10214), .ZN(n10471) );
  NOR2_X2 U12386 ( .A1(n10471), .A2(n10254), .ZN(n14953) );
  NAND2_X1 U12387 ( .A1(n6675), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9810) );
  INV_X1 U12388 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11128) );
  OR2_X1 U12389 ( .A1(n11900), .A2(n11128), .ZN(n9809) );
  INV_X1 U12390 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9805) );
  OR2_X1 U12391 ( .A1(n10120), .A2(n9805), .ZN(n9808) );
  OR2_X1 U12392 ( .A1(n11902), .A2(n9806), .ZN(n9807) );
  INV_X1 U12393 ( .A(n14318), .ZN(n9811) );
  INV_X1 U12394 ( .A(n6688), .ZN(n10118) );
  NOR2_X1 U12395 ( .A1(n9811), .A2(n14401), .ZN(n15063) );
  AOI22_X1 U12396 ( .A1(n9943), .A2(n14951), .B1(n14953), .B2(n15063), .ZN(
        n9818) );
  NAND2_X1 U12397 ( .A1(n9813), .A2(n9812), .ZN(n9815) );
  NOR2_X1 U12398 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  NAND2_X1 U12399 ( .A1(n14162), .A2(n9816), .ZN(n10292) );
  OR2_X1 U12400 ( .A1(n10292), .A2(P1_U3086), .ZN(n10211) );
  NAND2_X1 U12401 ( .A1(n10211), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9817) );
  OAI211_X1 U12402 ( .C1(n14300), .C2(n10238), .A(n9818), .B(n9817), .ZN(
        P1_U3232) );
  OR2_X1 U12403 ( .A1(n9819), .A2(n10407), .ZN(n9820) );
  NAND2_X1 U12404 ( .A1(n9821), .A2(n9820), .ZN(n10078) );
  XNOR2_X1 U12405 ( .A(n9822), .B(n10078), .ZN(n10949) );
  INV_X1 U12406 ( .A(n10949), .ZN(n9824) );
  OAI222_X1 U12407 ( .A1(n9825), .A2(n14764), .B1(P1_U3086), .B2(n9824), .C1(
        n14768), .C2(n9823), .ZN(P1_U3344) );
  INV_X1 U12408 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10956) );
  MUX2_X1 U12409 ( .A(n10956), .B(P1_REG1_REG_11__SCAN_IN), .S(n10949), .Z(
        n9829) );
  OAI21_X1 U12410 ( .B1(n9660), .B2(n9827), .A(n9826), .ZN(n9828) );
  AOI21_X1 U12411 ( .B1(n9829), .B2(n9828), .A(n10140), .ZN(n9838) );
  NAND2_X1 U12412 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14955)
         );
  OAI21_X1 U12413 ( .B1(n15042), .B2(n9830), .A(n14955), .ZN(n9836) );
  NAND2_X1 U12414 ( .A1(n10934), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9832) );
  INV_X1 U12415 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10990) );
  MUX2_X1 U12416 ( .A(n10990), .B(P1_REG2_REG_11__SCAN_IN), .S(n10949), .Z(
        n9831) );
  AOI21_X1 U12417 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n10131) );
  AND3_X1 U12418 ( .A1(n9833), .A2(n9832), .A3(n9831), .ZN(n9834) );
  NOR3_X1 U12419 ( .A1(n10131), .A2(n9834), .A3(n15034), .ZN(n9835) );
  AOI211_X1 U12420 ( .C1(n14387), .C2(n10949), .A(n9836), .B(n9835), .ZN(n9837) );
  OAI21_X1 U12421 ( .B1(n9838), .B2(n15036), .A(n9837), .ZN(P1_U3254) );
  OAI222_X1 U12422 ( .A1(P3_U3151), .A2(n14862), .B1(n11518), .B2(n9840), .C1(
        n13468), .C2(n9839), .ZN(P3_U3278) );
  NAND2_X1 U12423 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10607) );
  INV_X1 U12424 ( .A(n10607), .ZN(n9849) );
  INV_X1 U12425 ( .A(n13711), .ZN(n13710) );
  XNOR2_X1 U12426 ( .A(n13711), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n13706) );
  INV_X1 U12427 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9841) );
  MUX2_X1 U12428 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9841), .S(n15152), .Z(
        n15158) );
  AOI21_X1 U12429 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n9852), .A(n15157), .ZN(
        n15170) );
  INV_X1 U12430 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9842) );
  MUX2_X1 U12431 ( .A(n9842), .B(P2_REG2_REG_3__SCAN_IN), .S(n9853), .Z(n15169) );
  NOR2_X1 U12432 ( .A1(n15170), .A2(n15169), .ZN(n15168) );
  INV_X1 U12433 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10744) );
  MUX2_X1 U12434 ( .A(n10744), .B(P2_REG2_REG_4__SCAN_IN), .S(n9854), .Z(
        n10039) );
  NOR2_X1 U12435 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  INV_X1 U12436 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9843) );
  MUX2_X1 U12437 ( .A(n9843), .B(P2_REG2_REG_5__SCAN_IN), .S(n9855), .Z(n15184) );
  NAND2_X1 U12438 ( .A1(n9855), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9846) );
  INV_X1 U12439 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9844) );
  MUX2_X1 U12440 ( .A(n9844), .B(P2_REG2_REG_6__SCAN_IN), .S(n9922), .Z(n9845)
         );
  AOI21_X1 U12441 ( .B1(n15187), .B2(n9846), .A(n9845), .ZN(n9918) );
  AND3_X1 U12442 ( .A1(n15187), .A2(n9846), .A3(n9845), .ZN(n9847) );
  NOR3_X1 U12443 ( .A1(n9918), .A2(n9847), .A3(n15221), .ZN(n9848) );
  AOI211_X1 U12444 ( .C1(n15266), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n9849), .B(
        n9848), .ZN(n9862) );
  NAND2_X1 U12445 ( .A1(n13710), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9851) );
  INV_X1 U12446 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15412) );
  NAND2_X1 U12447 ( .A1(n13711), .A2(n15412), .ZN(n9850) );
  NAND4_X1 U12448 ( .A1(n9851), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .A4(n9850), .ZN(n13715) );
  NAND2_X1 U12449 ( .A1(n13715), .A2(n9851), .ZN(n15154) );
  XNOR2_X1 U12450 ( .A(n15152), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U12451 ( .A1(n15154), .A2(n15155), .B1(n9852), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n15173) );
  INV_X1 U12452 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15414) );
  MUX2_X1 U12453 ( .A(n15414), .B(P2_REG1_REG_3__SCAN_IN), .S(n9853), .Z(
        n15172) );
  OR2_X1 U12454 ( .A1(n15173), .A2(n15172), .ZN(n15175) );
  NAND2_X1 U12455 ( .A1(n9853), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10044) );
  INV_X1 U12456 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15416) );
  MUX2_X1 U12457 ( .A(n15416), .B(P2_REG1_REG_4__SCAN_IN), .S(n9854), .Z(
        n10043) );
  AOI21_X1 U12458 ( .B1(n15175), .B2(n10044), .A(n10043), .ZN(n10046) );
  AOI21_X1 U12459 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n9854), .A(n10046), .ZN(
        n15189) );
  INV_X1 U12460 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15418) );
  MUX2_X1 U12461 ( .A(n15418), .B(P2_REG1_REG_5__SCAN_IN), .S(n9855), .Z(
        n15188) );
  OR2_X1 U12462 ( .A1(n15189), .A2(n15188), .ZN(n15191) );
  NAND2_X1 U12463 ( .A1(n9855), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9858) );
  INV_X1 U12464 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9856) );
  MUX2_X1 U12465 ( .A(n9856), .B(P2_REG1_REG_6__SCAN_IN), .S(n9922), .Z(n9857)
         );
  AOI21_X1 U12466 ( .B1(n15191), .B2(n9858), .A(n9857), .ZN(n9921) );
  INV_X1 U12467 ( .A(n9921), .ZN(n9860) );
  NAND3_X1 U12468 ( .A1(n15191), .A2(n9858), .A3(n9857), .ZN(n9859) );
  NAND3_X1 U12469 ( .A1(n15270), .A2(n9860), .A3(n9859), .ZN(n9861) );
  OAI211_X1 U12470 ( .C1(n15265), .C2(n9863), .A(n9862), .B(n9861), .ZN(
        P2_U3220) );
  MUX2_X1 U12471 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n6678), .Z(n10056) );
  XNOR2_X1 U12472 ( .A(n10056), .B(n10062), .ZN(n10057) );
  MUX2_X1 U12473 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6678), .Z(n9864) );
  XNOR2_X1 U12474 ( .A(n9864), .B(n6680), .ZN(n10008) );
  INV_X1 U12475 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15683) );
  INV_X1 U12476 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n15743) );
  MUX2_X1 U12477 ( .A(n15683), .B(n15743), .S(n6678), .Z(n9992) );
  NAND2_X1 U12478 ( .A1(n9992), .A2(n13472), .ZN(n10007) );
  OAI22_X1 U12479 ( .A1(n10008), .A2(n10007), .B1(n9864), .B2(n6680), .ZN(
        n9900) );
  MUX2_X1 U12480 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n6678), .Z(n9865) );
  XOR2_X1 U12481 ( .A(n9886), .B(n9865), .Z(n9901) );
  INV_X1 U12482 ( .A(n9886), .ZN(n9915) );
  INV_X1 U12483 ( .A(n9865), .ZN(n9866) );
  AOI22_X1 U12484 ( .A1(n9900), .A2(n9901), .B1(n9915), .B2(n9866), .ZN(n10058) );
  XOR2_X1 U12485 ( .A(n10057), .B(n10058), .Z(n9899) );
  NOR2_X2 U12486 ( .A1(n13044), .A2(n9869), .ZN(n15588) );
  NAND2_X1 U12487 ( .A1(n12320), .A2(n10160), .ZN(n9867) );
  AND2_X1 U12488 ( .A1(n9868), .A2(n9867), .ZN(n9877) );
  OR2_X1 U12489 ( .A1(n10160), .A2(P3_U3151), .ZN(n12362) );
  NAND2_X1 U12490 ( .A1(n10794), .A2(n12362), .ZN(n9878) );
  INV_X1 U12491 ( .A(n9882), .ZN(n9870) );
  MUX2_X1 U12492 ( .A(n9870), .B(n13044), .S(n9869), .Z(n15584) );
  INV_X1 U12493 ( .A(n15584), .ZN(n14870) );
  INV_X1 U12494 ( .A(n10062), .ZN(n9897) );
  NAND2_X1 U12495 ( .A1(n9882), .A2(n6678), .ZN(n15488) );
  INV_X1 U12496 ( .A(n13472), .ZN(n9871) );
  NAND2_X1 U12497 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9871), .ZN(n9996) );
  INV_X1 U12498 ( .A(n9996), .ZN(n9872) );
  OAI21_X1 U12499 ( .B1(n6680), .B2(n9872), .A(n7623), .ZN(n10013) );
  INV_X1 U12500 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U12501 ( .A1(n10015), .A2(n7623), .ZN(n9903) );
  INV_X1 U12502 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U12503 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n9873), .S(n9886), .Z(n9904)
         );
  NAND2_X1 U12504 ( .A1(n9886), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12505 ( .A1(n9902), .A2(n9874), .ZN(n10063) );
  NAND2_X1 U12506 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n9875), .ZN(n10064) );
  OAI21_X1 U12507 ( .B1(n9875), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10064), .ZN(
        n9876) );
  NAND2_X1 U12508 ( .A1(n15586), .A2(n9876), .ZN(n9895) );
  INV_X1 U12509 ( .A(n9877), .ZN(n9879) );
  NOR2_X1 U12510 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8475), .ZN(n10371) );
  AOI21_X1 U12511 ( .B1(n15581), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10371), .ZN(
        n9894) );
  INV_X1 U12512 ( .A(n9880), .ZN(n9881) );
  NOR2_X1 U12513 ( .A1(n13472), .A2(n15683), .ZN(n9995) );
  NAND2_X1 U12514 ( .A1(n8461), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9883) );
  INV_X1 U12515 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U12516 ( .A1(n9908), .A2(n9909), .ZN(n9907) );
  NAND2_X1 U12517 ( .A1(n9886), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9887) );
  INV_X1 U12518 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9889) );
  AOI21_X1 U12519 ( .B1(n9890), .B2(n9889), .A(n10052), .ZN(n9891) );
  INV_X1 U12520 ( .A(n9891), .ZN(n9892) );
  NAND2_X1 U12521 ( .A1(n14879), .A2(n9892), .ZN(n9893) );
  NAND3_X1 U12522 ( .A1(n9895), .A2(n9894), .A3(n9893), .ZN(n9896) );
  AOI21_X1 U12523 ( .B1(n14870), .B2(n9897), .A(n9896), .ZN(n9898) );
  OAI21_X1 U12524 ( .B1(n9899), .B2(n15549), .A(n9898), .ZN(P3_U3185) );
  XOR2_X1 U12525 ( .A(n9901), .B(n9900), .Z(n9917) );
  OAI21_X1 U12526 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9905) );
  NAND2_X1 U12527 ( .A1(n15586), .A2(n9905), .ZN(n9913) );
  INV_X1 U12528 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10309) );
  NOR2_X1 U12529 ( .A1(n10309), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9906) );
  AOI21_X1 U12530 ( .B1(n15581), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n9906), .ZN(
        n9912) );
  OAI21_X1 U12531 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(n9910) );
  NAND2_X1 U12532 ( .A1(n14879), .A2(n9910), .ZN(n9911) );
  NAND3_X1 U12533 ( .A1(n9913), .A2(n9912), .A3(n9911), .ZN(n9914) );
  AOI21_X1 U12534 ( .B1(n14870), .B2(n9915), .A(n9914), .ZN(n9916) );
  OAI21_X1 U12535 ( .B1(n9917), .B2(n15549), .A(n9916), .ZN(P3_U3184) );
  INV_X1 U12536 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9919) );
  MUX2_X1 U12537 ( .A(n9919), .B(P2_REG2_REG_7__SCAN_IN), .S(n9924), .Z(n15204) );
  NOR2_X1 U12538 ( .A1(n15205), .A2(n15204), .ZN(n15203) );
  AOI21_X1 U12539 ( .B1(n9924), .B2(P2_REG2_REG_7__SCAN_IN), .A(n15203), .ZN(
        n10027) );
  INV_X1 U12540 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9920) );
  MUX2_X1 U12541 ( .A(n9920), .B(P2_REG2_REG_8__SCAN_IN), .S(n9925), .Z(n10026) );
  NOR2_X1 U12542 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  INV_X1 U12543 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9934) );
  NOR3_X1 U12544 ( .A1(n9936), .A2(n9934), .A3(n15221), .ZN(n9927) );
  AOI21_X1 U12545 ( .B1(n9922), .B2(P2_REG1_REG_6__SCAN_IN), .A(n9921), .ZN(
        n15201) );
  INV_X1 U12546 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U12547 ( .A(n9923), .B(P2_REG1_REG_7__SCAN_IN), .S(n9924), .Z(n15200) );
  NOR2_X1 U12548 ( .A1(n15201), .A2(n15200), .ZN(n15199) );
  AOI21_X1 U12549 ( .B1(n9924), .B2(P2_REG1_REG_7__SCAN_IN), .A(n15199), .ZN(
        n10031) );
  INV_X1 U12550 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15420) );
  MUX2_X1 U12551 ( .A(n15420), .B(P2_REG1_REG_8__SCAN_IN), .S(n9925), .Z(
        n10030) );
  NOR2_X1 U12552 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  AOI21_X1 U12553 ( .B1(n9925), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10029), .ZN(
        n9931) );
  INV_X1 U12554 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9928) );
  NOR3_X1 U12555 ( .A1(n9931), .A2(n9928), .A3(n15214), .ZN(n9926) );
  NOR3_X1 U12556 ( .A1(n9927), .A2(n15268), .A3(n9926), .ZN(n9942) );
  NAND2_X1 U12557 ( .A1(n9941), .A2(n9928), .ZN(n9930) );
  MUX2_X1 U12558 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9928), .S(n10353), .Z(n9929) );
  NAND2_X1 U12559 ( .A1(n9931), .A2(n9929), .ZN(n10347) );
  OAI21_X1 U12560 ( .B1(n9931), .B2(n9930), .A(n10347), .ZN(n9933) );
  INV_X1 U12561 ( .A(n15266), .ZN(n15231) );
  INV_X1 U12562 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14784) );
  NAND2_X1 U12563 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10880) );
  OAI21_X1 U12564 ( .B1(n15231), .B2(n14784), .A(n10880), .ZN(n9932) );
  AOI21_X1 U12565 ( .B1(n9933), .B2(n15270), .A(n9932), .ZN(n9940) );
  NOR3_X1 U12566 ( .A1(n9936), .A2(n10353), .A3(P2_REG2_REG_9__SCAN_IN), .ZN(
        n9938) );
  MUX2_X1 U12567 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9934), .S(n10353), .Z(n9935) );
  NAND2_X1 U12568 ( .A1(n9936), .A2(n9935), .ZN(n10352) );
  INV_X1 U12569 ( .A(n10352), .ZN(n9937) );
  OAI21_X1 U12570 ( .B1(n9938), .B2(n9937), .A(n15274), .ZN(n9939) );
  OAI211_X1 U12571 ( .C1(n9942), .C2(n9941), .A(n9940), .B(n9939), .ZN(
        P2_U3223) );
  MUX2_X1 U12572 ( .A(n9944), .B(n9943), .S(n6679), .Z(n9947) );
  NAND2_X1 U12573 ( .A1(n9945), .A2(n7302), .ZN(n9946) );
  OAI211_X1 U12574 ( .C1(n9947), .C2(n6688), .A(n14319), .B(n9946), .ZN(n14354) );
  AOI22_X1 U12575 ( .A1(n14343), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9960) );
  MUX2_X1 U12576 ( .A(n11122), .B(P1_REG2_REG_2__SCAN_IN), .S(n10113), .Z(
        n9950) );
  NAND3_X1 U12577 ( .A1(n9950), .A2(n9949), .A3(n9948), .ZN(n9951) );
  NAND3_X1 U12578 ( .A1(n14389), .A2(n9952), .A3(n9951), .ZN(n9959) );
  MUX2_X1 U12579 ( .A(n10107), .B(P1_REG1_REG_2__SCAN_IN), .S(n10113), .Z(
        n9955) );
  NAND3_X1 U12580 ( .A1(n9955), .A2(n9954), .A3(n9953), .ZN(n9956) );
  NAND3_X1 U12581 ( .A1(n14383), .A2(n14326), .A3(n9956), .ZN(n9958) );
  NAND2_X1 U12582 ( .A1(n14387), .A2(n10113), .ZN(n9957) );
  AND4_X1 U12583 ( .A1(n9960), .A2(n9959), .A3(n9958), .A4(n9957), .ZN(n9961)
         );
  NAND2_X1 U12584 ( .A1(n14354), .A2(n9961), .ZN(P1_U3245) );
  NAND2_X1 U12585 ( .A1(n15597), .A2(P3_U3897), .ZN(n9962) );
  OAI21_X1 U12586 ( .B1(P3_U3897), .B2(n9963), .A(n9962), .ZN(P3_U3498) );
  NAND2_X1 U12587 ( .A1(n11109), .A2(P3_U3897), .ZN(n9964) );
  OAI21_X1 U12588 ( .B1(P3_U3897), .B2(n9965), .A(n9964), .ZN(P3_U3497) );
  NAND2_X1 U12589 ( .A1(n10799), .A2(P3_U3897), .ZN(n9966) );
  OAI21_X1 U12590 ( .B1(P3_U3897), .B2(n9967), .A(n9966), .ZN(P3_U3494) );
  NAND2_X1 U12591 ( .A1(n11647), .A2(P3_U3897), .ZN(n9968) );
  OAI21_X1 U12592 ( .B1(P3_U3897), .B2(n9969), .A(n9968), .ZN(P3_U3501) );
  NAND2_X1 U12593 ( .A1(n12954), .A2(P3_U3897), .ZN(n9970) );
  OAI21_X1 U12594 ( .B1(P3_U3897), .B2(n9971), .A(n9970), .ZN(P3_U3508) );
  NAND2_X1 U12595 ( .A1(n10372), .A2(P3_U3897), .ZN(n9972) );
  OAI21_X1 U12596 ( .B1(P3_U3897), .B2(n9973), .A(n9972), .ZN(P3_U3495) );
  NAND2_X1 U12597 ( .A1(n13287), .A2(P3_U3897), .ZN(n9974) );
  OAI21_X1 U12598 ( .B1(P3_U3897), .B2(n9975), .A(n9974), .ZN(P3_U3507) );
  NAND2_X1 U12599 ( .A1(n13288), .A2(P3_U3897), .ZN(n9976) );
  OAI21_X1 U12600 ( .B1(P3_U3897), .B2(n9977), .A(n9976), .ZN(P3_U3509) );
  NAND2_X1 U12601 ( .A1(n12199), .A2(P3_U3897), .ZN(n9978) );
  OAI21_X1 U12602 ( .B1(P3_U3897), .B2(n9979), .A(n9978), .ZN(P3_U3496) );
  NAND2_X1 U12603 ( .A1(n12992), .A2(P3_U3897), .ZN(n9980) );
  OAI21_X1 U12604 ( .B1(P3_U3897), .B2(n9981), .A(n9980), .ZN(P3_U3505) );
  NAND2_X1 U12605 ( .A1(n12893), .A2(P3_U3897), .ZN(n9982) );
  OAI21_X1 U12606 ( .B1(P3_U3897), .B2(n9983), .A(n9982), .ZN(P3_U3504) );
  NAND2_X1 U12607 ( .A1(n11688), .A2(P3_U3897), .ZN(n9984) );
  OAI21_X1 U12608 ( .B1(P3_U3897), .B2(n9985), .A(n9984), .ZN(P3_U3502) );
  NAND2_X1 U12609 ( .A1(n12982), .A2(P3_U3897), .ZN(n9986) );
  OAI21_X1 U12610 ( .B1(P3_U3897), .B2(n9987), .A(n9986), .ZN(P3_U3510) );
  NAND2_X1 U12611 ( .A1(n15431), .A2(P3_U3897), .ZN(n9988) );
  OAI21_X1 U12612 ( .B1(P3_U3897), .B2(n9989), .A(n9988), .ZN(P3_U3492) );
  NAND2_X1 U12613 ( .A1(n12216), .A2(P3_U3897), .ZN(n9990) );
  OAI21_X1 U12614 ( .B1(P3_U3897), .B2(n9991), .A(n9990), .ZN(P3_U3499) );
  NOR3_X1 U12615 ( .A1(n15586), .A2(n14879), .A3(n15588), .ZN(n10002) );
  INV_X1 U12616 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15675) );
  INV_X1 U12617 ( .A(n9992), .ZN(n9993) );
  NAND3_X1 U12618 ( .A1(n15588), .A2(n9993), .A3(n9871), .ZN(n9994) );
  OAI21_X1 U12619 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15675), .A(n9994), .ZN(
        n9999) );
  INV_X1 U12620 ( .A(n9995), .ZN(n9997) );
  OAI22_X1 U12621 ( .A1(n15594), .A2(n9997), .B1(n9996), .B2(n15488), .ZN(
        n9998) );
  AOI211_X1 U12622 ( .C1(n15581), .C2(P3_ADDR_REG_0__SCAN_IN), .A(n9999), .B(
        n9998), .ZN(n10001) );
  NAND2_X1 U12623 ( .A1(n14870), .A2(n13472), .ZN(n10000) );
  OAI211_X1 U12624 ( .C1(n10002), .C2(n10007), .A(n10001), .B(n10000), .ZN(
        P3_U3182) );
  NAND2_X1 U12625 ( .A1(n15652), .A2(P3_U3897), .ZN(n10003) );
  OAI21_X1 U12626 ( .B1(P3_U3897), .B2(n10004), .A(n10003), .ZN(P3_U3491) );
  NAND2_X1 U12627 ( .A1(n15655), .A2(P3_U3897), .ZN(n10005) );
  OAI21_X1 U12628 ( .B1(P3_U3897), .B2(n10006), .A(n10005), .ZN(P3_U3493) );
  XOR2_X1 U12629 ( .A(n10008), .B(n10007), .Z(n10024) );
  NAND2_X1 U12630 ( .A1(n10009), .A2(n15668), .ZN(n10010) );
  NAND2_X1 U12631 ( .A1(n10011), .A2(n10010), .ZN(n10022) );
  NAND2_X1 U12632 ( .A1(n10013), .A2(n10012), .ZN(n10014) );
  AND2_X1 U12633 ( .A1(n10015), .A2(n10014), .ZN(n10018) );
  NAND2_X1 U12634 ( .A1(n15581), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U12635 ( .A1(P3_U3151), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n10016) );
  OAI211_X1 U12636 ( .C1(n15488), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10021) );
  NOR2_X1 U12637 ( .A1(n15584), .A2(n6680), .ZN(n10020) );
  AOI211_X1 U12638 ( .C1(n14879), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10023) );
  OAI21_X1 U12639 ( .B1(n15549), .B2(n10024), .A(n10023), .ZN(P3_U3183) );
  AOI211_X1 U12640 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n15221), .ZN(
        n10028) );
  INV_X1 U12641 ( .A(n10028), .ZN(n10034) );
  AOI211_X1 U12642 ( .C1(n10031), .C2(n10030), .A(n10029), .B(n15214), .ZN(
        n10032) );
  INV_X1 U12643 ( .A(n10032), .ZN(n10033) );
  NAND2_X1 U12644 ( .A1(n10034), .A2(n10033), .ZN(n10035) );
  AND2_X1 U12645 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10692) );
  AOI211_X1 U12646 ( .C1(n15266), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10035), .B(
        n10692), .ZN(n10036) );
  OAI21_X1 U12647 ( .B1(n10037), .B2(n15265), .A(n10036), .ZN(P2_U3222) );
  NAND2_X1 U12648 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10451) );
  AOI211_X1 U12649 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n15221), .ZN(
        n10041) );
  INV_X1 U12650 ( .A(n10041), .ZN(n10042) );
  NAND2_X1 U12651 ( .A1(n10451), .A2(n10042), .ZN(n10048) );
  AND3_X1 U12652 ( .A1(n15175), .A2(n10044), .A3(n10043), .ZN(n10045) );
  NOR3_X1 U12653 ( .A1(n15214), .A2(n10046), .A3(n10045), .ZN(n10047) );
  AOI211_X1 U12654 ( .C1(n15266), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10048), .B(
        n10047), .ZN(n10049) );
  OAI21_X1 U12655 ( .B1(n10050), .B2(n15265), .A(n10049), .ZN(P2_U3218) );
  INV_X1 U12656 ( .A(n10051), .ZN(n10053) );
  INV_X1 U12657 ( .A(n15437), .ZN(n10067) );
  INV_X1 U12658 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U12659 ( .A1(n10067), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n10054), 
        .B2(n15437), .ZN(n15439) );
  INV_X1 U12660 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15620) );
  AOI21_X1 U12661 ( .B1(n10055), .B2(n15620), .A(n10619), .ZN(n10076) );
  OAI22_X1 U12662 ( .A1(n10058), .A2(n10057), .B1(n10056), .B2(n10062), .ZN(
        n15436) );
  MUX2_X1 U12663 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n6678), .Z(n10059) );
  XNOR2_X1 U12664 ( .A(n10059), .B(n10067), .ZN(n15435) );
  INV_X1 U12665 ( .A(n10059), .ZN(n10060) );
  AOI22_X1 U12666 ( .A1(n15436), .A2(n15435), .B1(n10067), .B2(n10060), .ZN(
        n10649) );
  MUX2_X1 U12667 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n6678), .Z(n10647) );
  XNOR2_X1 U12668 ( .A(n10647), .B(n10646), .ZN(n10648) );
  XNOR2_X1 U12669 ( .A(n10649), .B(n10648), .ZN(n10061) );
  NAND2_X1 U12670 ( .A1(n10061), .A2(n15588), .ZN(n10075) );
  INV_X1 U12671 ( .A(n10646), .ZN(n10618) );
  INV_X1 U12672 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U12673 ( .A1(n10067), .A2(n15749), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n15437), .ZN(n15442) );
  NAND2_X1 U12674 ( .A1(n10063), .A2(n10062), .ZN(n10065) );
  NAND2_X1 U12675 ( .A1(n10065), .A2(n10064), .ZN(n15441) );
  NAND2_X1 U12676 ( .A1(n15442), .A2(n15441), .ZN(n10066) );
  XNOR2_X1 U12677 ( .A(n10618), .B(n10631), .ZN(n10068) );
  NAND2_X1 U12678 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n10068), .ZN(n10632) );
  OAI21_X1 U12679 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n10068), .A(n10632), .ZN(
        n10073) );
  INV_X1 U12680 ( .A(n15581), .ZN(n15519) );
  NOR2_X1 U12681 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10069), .ZN(n10705) );
  INV_X1 U12682 ( .A(n10705), .ZN(n10070) );
  OAI21_X1 U12683 ( .B1(n15519), .B2(n9264), .A(n10070), .ZN(n10072) );
  NOR2_X1 U12684 ( .A1(n15584), .A2(n10646), .ZN(n10071) );
  AOI211_X1 U12685 ( .C1(n15586), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10074) );
  OAI211_X1 U12686 ( .C1(n10076), .C2(n15594), .A(n10075), .B(n10074), .ZN(
        P3_U3187) );
  INV_X1 U12687 ( .A(n15226), .ZN(n11084) );
  INV_X1 U12688 ( .A(n11270), .ZN(n10079) );
  OAI222_X1 U12689 ( .A1(P2_U3088), .A2(n11084), .B1(n14150), .B2(n10079), 
        .C1(n10077), .C2(n14152), .ZN(P2_U3315) );
  OAI21_X1 U12690 ( .B1(n10078), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10147) );
  XNOR2_X1 U12691 ( .A(n10147), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11271) );
  INV_X1 U12692 ( .A(n11271), .ZN(n10137) );
  OAI222_X1 U12693 ( .A1(n14764), .A2(n10080), .B1(n14768), .B2(n10079), .C1(
        n10137), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12694 ( .A(n14869), .ZN(n13090) );
  OAI222_X1 U12695 ( .A1(P3_U3151), .A2(n13090), .B1(n11518), .B2(n10082), 
        .C1(n13468), .C2(n10081), .ZN(P3_U3277) );
  NAND2_X1 U12696 ( .A1(n13002), .A2(P3_U3897), .ZN(n10083) );
  OAI21_X1 U12697 ( .B1(P3_U3897), .B2(n10084), .A(n10083), .ZN(P3_U3512) );
  INV_X1 U12698 ( .A(n10085), .ZN(n10087) );
  OR2_X1 U12699 ( .A1(n10092), .A2(n10094), .ZN(n10095) );
  NAND2_X1 U12700 ( .A1(n12804), .A2(n10244), .ZN(n10099) );
  NAND2_X1 U12701 ( .A1(n14318), .A2(n11309), .ZN(n10098) );
  NOR2_X1 U12702 ( .A1(n6686), .A2(n11129), .ZN(n10101) );
  AOI21_X1 U12703 ( .B1(n12817), .B2(n14318), .A(n10101), .ZN(n10102) );
  NAND2_X1 U12704 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  OAI21_X1 U12705 ( .B1(n10103), .B2(n10102), .A(n10104), .ZN(n10206) );
  NOR2_X2 U12706 ( .A1(n10207), .A2(n10206), .ZN(n10205) );
  INV_X1 U12707 ( .A(n10104), .ZN(n10105) );
  NAND2_X1 U12708 ( .A1(n6674), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10111) );
  INV_X1 U12709 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11118) );
  OR2_X1 U12710 ( .A1(n11900), .A2(n11118), .ZN(n10110) );
  INV_X1 U12711 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10106) );
  OR2_X1 U12712 ( .A1(n10120), .A2(n10106), .ZN(n10109) );
  NAND2_X1 U12713 ( .A1(n10112), .A2(n6685), .ZN(n10114) );
  AOI22_X1 U12714 ( .A1(n11309), .A2(n14317), .B1(n12804), .B2(n11934), .ZN(
        n10115) );
  XNOR2_X1 U12715 ( .A(n10115), .B(n12824), .ZN(n10288) );
  AOI22_X1 U12716 ( .A1(n12817), .A2(n14317), .B1(n11309), .B2(n11934), .ZN(
        n10287) );
  XNOR2_X1 U12717 ( .A(n10288), .B(n10287), .ZN(n10116) );
  AOI21_X1 U12718 ( .B1(n10117), .B2(n10116), .A(n6812), .ZN(n10129) );
  INV_X1 U12719 ( .A(n14953), .ZN(n14294) );
  NAND2_X1 U12720 ( .A1(n11884), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10126) );
  OR2_X1 U12721 ( .A1(n11900), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10125) );
  OR2_X1 U12722 ( .A1(n11902), .A2(n10121), .ZN(n10124) );
  OR2_X1 U12723 ( .A1(n10273), .A2(n10122), .ZN(n10123) );
  AOI22_X1 U12724 ( .A1(n14563), .A2(n14318), .B1(n14316), .B2(n14565), .ZN(
        n10229) );
  OAI22_X1 U12725 ( .A1(n14300), .A2(n7180), .B1(n14294), .B2(n10229), .ZN(
        n10127) );
  AOI21_X1 U12726 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10211), .A(n10127), .ZN(
        n10128) );
  OAI21_X1 U12727 ( .B1(n10129), .B2(n14277), .A(n10128), .ZN(P1_U3237) );
  INV_X1 U12728 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10130) );
  MUX2_X1 U12729 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10130), .S(n11271), .Z(
        n10133) );
  AOI21_X1 U12730 ( .B1(n10949), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10131), 
        .ZN(n10132) );
  NAND2_X1 U12731 ( .A1(n10132), .A2(n10133), .ZN(n10314) );
  OAI21_X1 U12732 ( .B1(n10133), .B2(n10132), .A(n10314), .ZN(n10144) );
  INV_X1 U12733 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10134) );
  NOR2_X1 U12734 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10134), .ZN(n10135) );
  AOI21_X1 U12735 ( .B1(n14343), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10135), 
        .ZN(n10136) );
  OAI21_X1 U12736 ( .B1(n15038), .B2(n10137), .A(n10136), .ZN(n10143) );
  NOR2_X1 U12737 ( .A1(n10949), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10138) );
  INV_X1 U12738 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14812) );
  MUX2_X1 U12739 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n14812), .S(n11271), .Z(
        n10139) );
  OAI21_X1 U12740 ( .B1(n10140), .B2(n10138), .A(n10139), .ZN(n10310) );
  OR3_X1 U12741 ( .A1(n10140), .A2(n10139), .A3(n10138), .ZN(n10141) );
  AOI21_X1 U12742 ( .B1(n10310), .B2(n10141), .A(n15036), .ZN(n10142) );
  AOI211_X1 U12743 ( .C1(n14389), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10145) );
  INV_X1 U12744 ( .A(n10145), .ZN(P1_U3255) );
  INV_X1 U12745 ( .A(n11277), .ZN(n10153) );
  NAND2_X1 U12746 ( .A1(n10147), .A2(n10146), .ZN(n10148) );
  NAND2_X1 U12747 ( .A1(n10148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10150) );
  NAND2_X1 U12748 ( .A1(n10150), .A2(n10149), .ZN(n10338) );
  OR2_X1 U12749 ( .A1(n10150), .A2(n10149), .ZN(n10151) );
  INV_X1 U12750 ( .A(n11278), .ZN(n11178) );
  OAI222_X1 U12751 ( .A1(n14771), .A2(n10152), .B1(n14768), .B2(n10153), .C1(
        n11178), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12752 ( .A(n15234), .ZN(n11086) );
  OAI222_X1 U12753 ( .A1(n14152), .A2(n10154), .B1(n14150), .B2(n10153), .C1(
        n11086), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI222_X1 U12754 ( .A1(n13471), .A2(n10156), .B1(P3_U3151), .B2(n13089), 
        .C1(n13468), .C2(n10155), .ZN(P3_U3276) );
  NAND2_X1 U12755 ( .A1(n13229), .A2(P3_U3897), .ZN(n10157) );
  OAI21_X1 U12756 ( .B1(P3_U3897), .B2(n10158), .A(n10157), .ZN(P3_U3513) );
  INV_X1 U12757 ( .A(n10186), .ZN(n10159) );
  NAND2_X1 U12758 ( .A1(n10196), .A2(n10159), .ZN(n10166) );
  AND2_X1 U12759 ( .A1(n10161), .A2(n10160), .ZN(n10165) );
  NAND2_X1 U12760 ( .A1(n10191), .A2(n10162), .ZN(n10163) );
  NAND4_X1 U12761 ( .A1(n10166), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10167) );
  NAND2_X1 U12762 ( .A1(n10167), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10170) );
  NAND2_X1 U12763 ( .A1(n10168), .A2(n10196), .ZN(n10169) );
  NOR2_X1 U12764 ( .A1(n13037), .A2(P3_U3151), .ZN(n15434) );
  INV_X1 U12765 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10204) );
  INV_X1 U12766 ( .A(n12353), .ZN(n10171) );
  NAND2_X1 U12767 ( .A1(n10172), .A2(n10171), .ZN(n10174) );
  AOI21_X1 U12768 ( .B1(n12171), .B2(n10344), .A(n10194), .ZN(n10173) );
  MUX2_X1 U12769 ( .A(n12179), .B(n15639), .S(n12848), .Z(n10300) );
  NAND2_X1 U12770 ( .A1(n10175), .A2(n12848), .ZN(n10176) );
  OR2_X1 U12771 ( .A1(n15674), .A2(n10176), .ZN(n10177) );
  NAND2_X1 U12772 ( .A1(n15657), .A2(n12848), .ZN(n10178) );
  NAND2_X1 U12773 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  INV_X1 U12774 ( .A(n15651), .ZN(n10182) );
  INV_X4 U12775 ( .A(n12848), .ZN(n12921) );
  NAND3_X1 U12776 ( .A1(n10182), .A2(n15658), .A3(n12921), .ZN(n10183) );
  OAI211_X1 U12777 ( .C1(n10184), .C2(n15657), .A(n10301), .B(n10183), .ZN(
        n10190) );
  NAND2_X1 U12778 ( .A1(n10185), .A2(n15672), .ZN(n10188) );
  OR2_X1 U12779 ( .A1(n10196), .A2(n10186), .ZN(n10187) );
  NAND2_X1 U12780 ( .A1(n10188), .A2(n10187), .ZN(n10189) );
  NAND2_X1 U12781 ( .A1(n10190), .A2(n15432), .ZN(n10203) );
  INV_X1 U12782 ( .A(n12323), .ZN(n15663) );
  NAND2_X1 U12783 ( .A1(n10191), .A2(n15663), .ZN(n10193) );
  NOR2_X1 U12784 ( .A1(n10794), .A2(n15718), .ZN(n10192) );
  NAND2_X1 U12785 ( .A1(n10195), .A2(n10194), .ZN(n10197) );
  OR2_X1 U12786 ( .A1(n10197), .A2(n15637), .ZN(n12358) );
  NOR2_X2 U12787 ( .A1(n12358), .A2(n10196), .ZN(n13020) );
  INV_X1 U12788 ( .A(n15652), .ZN(n10200) );
  INV_X1 U12789 ( .A(n10196), .ZN(n10199) );
  INV_X1 U12790 ( .A(n10197), .ZN(n10198) );
  NAND3_X1 U12791 ( .A1(n10199), .A2(n15654), .A3(n10198), .ZN(n13023) );
  OAI22_X1 U12792 ( .A1(n13035), .A2(n10200), .B1(n15624), .B2(n13023), .ZN(
        n10201) );
  AOI21_X1 U12793 ( .B1(n15429), .B2(n10175), .A(n10201), .ZN(n10202) );
  OAI211_X1 U12794 ( .C1(n15434), .C2(n10204), .A(n10203), .B(n10202), .ZN(
        P3_U3162) );
  AOI21_X1 U12795 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10213) );
  INV_X1 U12796 ( .A(n14563), .ZN(n14460) );
  NOR2_X1 U12797 ( .A1(n14294), .A2(n14460), .ZN(n14265) );
  NAND2_X1 U12798 ( .A1(n14953), .A2(n14565), .ZN(n14262) );
  INV_X1 U12799 ( .A(n14262), .ZN(n10208) );
  AOI22_X1 U12800 ( .A1(n14265), .A2(n14320), .B1(n10208), .B2(n14317), .ZN(
        n10209) );
  OAI21_X1 U12801 ( .B1(n11129), .B2(n14300), .A(n10209), .ZN(n10210) );
  AOI21_X1 U12802 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10211), .A(n10210), .ZN(
        n10212) );
  OAI21_X1 U12803 ( .B1(n10213), .B2(n14277), .A(n10212), .ZN(P1_U3222) );
  NAND2_X1 U12804 ( .A1(n10214), .A2(n10460), .ZN(n10215) );
  OR2_X1 U12805 ( .A1(n10216), .A2(n10215), .ZN(n10255) );
  INV_X2 U12806 ( .A(n15135), .ZN(n15113) );
  NAND2_X1 U12807 ( .A1(n11928), .A2(n14773), .ZN(n10217) );
  NAND2_X1 U12808 ( .A1(n12824), .A2(n10217), .ZN(n10474) );
  OR2_X1 U12809 ( .A1(n10474), .A2(n14390), .ZN(n11018) );
  OR2_X1 U12810 ( .A1(n11911), .A2(n11166), .ZN(n15064) );
  OR2_X1 U12811 ( .A1(n15064), .A2(n14773), .ZN(n15119) );
  OR2_X1 U12812 ( .A1(n14318), .A2(n10244), .ZN(n10218) );
  NAND2_X1 U12813 ( .A1(n10234), .A2(n10218), .ZN(n10222) );
  NAND2_X1 U12814 ( .A1(n7180), .A2(n14317), .ZN(n10220) );
  AND2_X2 U12815 ( .A1(n10220), .A2(n11937), .ZN(n11857) );
  INV_X1 U12816 ( .A(n11857), .ZN(n10221) );
  INV_X1 U12817 ( .A(n10223), .ZN(n11125) );
  NAND2_X1 U12818 ( .A1(n11129), .A2(n10238), .ZN(n10237) );
  INV_X1 U12819 ( .A(n10270), .ZN(n10224) );
  AOI211_X1 U12820 ( .C1(n11934), .C2(n10237), .A(n14630), .B(n10224), .ZN(
        n11120) );
  AOI21_X1 U12821 ( .B1(n15116), .B2(n11934), .A(n11120), .ZN(n10232) );
  INV_X1 U12822 ( .A(n11925), .ZN(n10225) );
  NAND2_X1 U12823 ( .A1(n11929), .A2(n10225), .ZN(n11927) );
  NAND2_X1 U12824 ( .A1(n14318), .A2(n11129), .ZN(n11930) );
  AND2_X2 U12825 ( .A1(n11927), .A2(n11930), .ZN(n10226) );
  OAI21_X1 U12826 ( .B1(n11857), .B2(n10226), .A(n10272), .ZN(n10231) );
  NAND2_X1 U12827 ( .A1(n14773), .A2(n14390), .ZN(n10228) );
  OR2_X1 U12828 ( .A1(n12089), .A2(n11912), .ZN(n10227) );
  INV_X1 U12829 ( .A(n10229), .ZN(n10230) );
  AOI21_X1 U12830 ( .B1(n10231), .B2(n14792), .A(n10230), .ZN(n11121) );
  OAI211_X1 U12831 ( .C1(n14732), .C2(n11125), .A(n10232), .B(n11121), .ZN(
        n10260) );
  NAND2_X1 U12832 ( .A1(n10260), .A2(n15113), .ZN(n10233) );
  OAI21_X1 U12833 ( .B1(n15113), .B2(n10106), .A(n10233), .ZN(P1_U3465) );
  INV_X1 U12834 ( .A(n10248), .ZN(n10236) );
  INV_X1 U12835 ( .A(n10234), .ZN(n10235) );
  AOI21_X1 U12836 ( .B1(n10236), .B2(n11856), .A(n10235), .ZN(n11134) );
  OAI21_X1 U12837 ( .B1(n11856), .B2(n15128), .A(n14460), .ZN(n10242) );
  NOR2_X1 U12838 ( .A1(n10219), .A2(n14401), .ZN(n10241) );
  OAI21_X1 U12839 ( .B1(n11129), .B2(n10238), .A(n10237), .ZN(n10243) );
  XOR2_X1 U12840 ( .A(n14318), .B(n10243), .Z(n10239) );
  NOR3_X1 U12841 ( .A1(n10239), .A2(n15128), .A3(n14320), .ZN(n10240) );
  NOR2_X1 U12842 ( .A1(n10243), .A2(n14630), .ZN(n11131) );
  AOI21_X1 U12843 ( .B1(n15116), .B2(n10244), .A(n11131), .ZN(n10245) );
  OAI211_X1 U12844 ( .C1(n14732), .C2(n11134), .A(n11126), .B(n10245), .ZN(
        n10258) );
  NAND2_X1 U12845 ( .A1(n10258), .A2(n15113), .ZN(n10246) );
  OAI21_X1 U12846 ( .B1(n15113), .B2(n9805), .A(n10246), .ZN(P1_U3462) );
  NOR2_X1 U12847 ( .A1(n15134), .A2(n14792), .ZN(n10252) );
  INV_X1 U12848 ( .A(n15063), .ZN(n10251) );
  INV_X1 U12849 ( .A(n10476), .ZN(n10249) );
  NAND2_X1 U12850 ( .A1(n10250), .A2(n10249), .ZN(n15062) );
  OAI211_X1 U12851 ( .C1(n10252), .C2(n15066), .A(n10251), .B(n15062), .ZN(
        n10256) );
  NAND2_X1 U12852 ( .A1(n10256), .A2(n15113), .ZN(n10253) );
  OAI21_X1 U12853 ( .B1(n15113), .B2(n9785), .A(n10253), .ZN(P1_U3459) );
  NAND2_X1 U12854 ( .A1(n10256), .A2(n15150), .ZN(n10257) );
  OAI21_X1 U12855 ( .B1(n15150), .B2(n9797), .A(n10257), .ZN(P1_U3528) );
  NAND2_X1 U12856 ( .A1(n10258), .A2(n15150), .ZN(n10259) );
  OAI21_X1 U12857 ( .B1(n15150), .B2(n9806), .A(n10259), .ZN(P1_U3529) );
  NAND2_X1 U12858 ( .A1(n10260), .A2(n15150), .ZN(n10261) );
  OAI21_X1 U12859 ( .B1(n15150), .B2(n10107), .A(n10261), .ZN(P1_U3530) );
  INV_X1 U12860 ( .A(n15119), .ZN(n15097) );
  OR2_X1 U12861 ( .A1(n14317), .A2(n11934), .ZN(n10262) );
  NAND2_X1 U12862 ( .A1(n10263), .A2(n11892), .ZN(n10265) );
  AOI22_X1 U12863 ( .A1(n6671), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11852), 
        .B2(n14324), .ZN(n10264) );
  NAND2_X1 U12864 ( .A1(n10267), .A2(n10266), .ZN(n10473) );
  OR2_X1 U12865 ( .A1(n10267), .A2(n10266), .ZN(n10268) );
  NAND2_X1 U12866 ( .A1(n10473), .A2(n10268), .ZN(n11706) );
  INV_X1 U12867 ( .A(n11941), .ZN(n11707) );
  NAND2_X1 U12868 ( .A1(n11941), .A2(n10270), .ZN(n10269) );
  NAND2_X1 U12869 ( .A1(n10269), .A2(n15055), .ZN(n10271) );
  NOR2_X2 U12870 ( .A1(n11941), .A2(n10270), .ZN(n10479) );
  OR2_X1 U12871 ( .A1(n10271), .A2(n10479), .ZN(n11711) );
  OAI21_X1 U12872 ( .B1(n11707), .B2(n15126), .A(n11711), .ZN(n10282) );
  NAND2_X1 U12873 ( .A1(n10272), .A2(n11937), .ZN(n10463) );
  XNOR2_X1 U12874 ( .A(n10463), .B(n10266), .ZN(n10281) );
  INV_X1 U12875 ( .A(n11018), .ZN(n15123) );
  NAND2_X1 U12876 ( .A1(n11706), .A2(n15123), .ZN(n10280) );
  NAND2_X1 U12877 ( .A1(n11884), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10277) );
  OR2_X1 U12878 ( .A1(n11902), .A2(n15136), .ZN(n10276) );
  OR2_X1 U12879 ( .A1(n10273), .A2(n10478), .ZN(n10275) );
  XNOR2_X1 U12880 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10462) );
  OR2_X1 U12881 ( .A1(n11900), .A2(n10462), .ZN(n10274) );
  OR2_X1 U12882 ( .A1(n11946), .A2(n14401), .ZN(n10279) );
  NAND2_X1 U12883 ( .A1(n14317), .A2(n14563), .ZN(n10278) );
  AND2_X1 U12884 ( .A1(n10279), .A2(n10278), .ZN(n10293) );
  OAI211_X1 U12885 ( .C1(n15128), .C2(n10281), .A(n10280), .B(n10293), .ZN(
        n11704) );
  AOI211_X1 U12886 ( .C1(n15097), .C2(n11706), .A(n10282), .B(n11704), .ZN(
        n10284) );
  OR2_X1 U12887 ( .A1(n10284), .A2(n15148), .ZN(n10283) );
  OAI21_X1 U12888 ( .B1(n15150), .B2(n10121), .A(n10283), .ZN(P1_U3531) );
  INV_X1 U12889 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10286) );
  OR2_X1 U12890 ( .A1(n10284), .A2(n15135), .ZN(n10285) );
  OAI21_X1 U12891 ( .B1(n15113), .B2(n10286), .A(n10285), .ZN(P1_U3468) );
  AOI22_X1 U12892 ( .A1(n11941), .A2(n12804), .B1(n11309), .B2(n14316), .ZN(
        n10289) );
  XNOR2_X1 U12893 ( .A(n10289), .B(n12824), .ZN(n10418) );
  XOR2_X1 U12894 ( .A(n10419), .B(n10418), .Z(n10290) );
  OAI211_X1 U12895 ( .C1(n10291), .C2(n10290), .A(n10417), .B(n14951), .ZN(
        n10299) );
  INV_X1 U12896 ( .A(n14958), .ZN(n14296) );
  INV_X1 U12897 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10297) );
  INV_X1 U12898 ( .A(n10293), .ZN(n10294) );
  NAND2_X1 U12899 ( .A1(n14953), .A2(n10294), .ZN(n10295) );
  NAND2_X1 U12900 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14321) );
  NAND2_X1 U12901 ( .A1(n10295), .A2(n14321), .ZN(n10296) );
  AOI21_X1 U12902 ( .B1(n14296), .B2(n10297), .A(n10296), .ZN(n10298) );
  OAI211_X1 U12903 ( .C1(n11707), .C2(n14300), .A(n10299), .B(n10298), .ZN(
        P1_U3218) );
  XNOR2_X1 U12904 ( .A(n10306), .B(n12848), .ZN(n10362) );
  XNOR2_X1 U12905 ( .A(n10362), .B(n15624), .ZN(n10303) );
  NAND2_X1 U12906 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  NAND2_X1 U12907 ( .A1(n10302), .A2(n10303), .ZN(n10365) );
  OAI21_X1 U12908 ( .B1(n10303), .B2(n10302), .A(n10365), .ZN(n10304) );
  NAND2_X1 U12909 ( .A1(n10304), .A2(n15432), .ZN(n10308) );
  OAI22_X1 U12910 ( .A1(n13035), .A2(n15674), .B1(n15636), .B2(n13023), .ZN(
        n10305) );
  AOI21_X1 U12911 ( .B1(n10306), .B2(n15429), .A(n10305), .ZN(n10307) );
  OAI211_X1 U12912 ( .C1(n15434), .C2(n10309), .A(n10308), .B(n10307), .ZN(
        P3_U3177) );
  OAI21_X1 U12913 ( .B1(n11271), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10310), 
        .ZN(n10312) );
  INV_X1 U12914 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14984) );
  MUX2_X1 U12915 ( .A(n14984), .B(P1_REG1_REG_13__SCAN_IN), .S(n11278), .Z(
        n10311) );
  NOR2_X1 U12916 ( .A1(n10312), .A2(n10311), .ZN(n11169) );
  AOI211_X1 U12917 ( .C1(n10312), .C2(n10311), .A(n15036), .B(n11169), .ZN(
        n10313) );
  INV_X1 U12918 ( .A(n10313), .ZN(n10321) );
  NAND2_X1 U12919 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14248)
         );
  INV_X1 U12920 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11177) );
  MUX2_X1 U12921 ( .A(n11177), .B(P1_REG2_REG_13__SCAN_IN), .S(n11278), .Z(
        n10316) );
  OAI21_X1 U12922 ( .B1(n11271), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10314), 
        .ZN(n10315) );
  NOR2_X1 U12923 ( .A1(n10315), .A2(n10316), .ZN(n14368) );
  AOI211_X1 U12924 ( .C1(n10316), .C2(n10315), .A(n14368), .B(n15034), .ZN(
        n10317) );
  INV_X1 U12925 ( .A(n10317), .ZN(n10318) );
  NAND2_X1 U12926 ( .A1(n14248), .A2(n10318), .ZN(n10319) );
  AOI21_X1 U12927 ( .B1(n14343), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10319), 
        .ZN(n10320) );
  OAI211_X1 U12928 ( .C1(n15038), .C2(n11178), .A(n10321), .B(n10320), .ZN(
        P1_U3256) );
  XNOR2_X1 U12929 ( .A(n10322), .B(n12618), .ZN(n10781) );
  INV_X1 U12930 ( .A(n10855), .ZN(n10324) );
  INV_X1 U12931 ( .A(n10395), .ZN(n10323) );
  AOI211_X1 U12932 ( .C1(n12411), .C2(n10324), .A(n13922), .B(n10323), .ZN(
        n10774) );
  XNOR2_X1 U12933 ( .A(n10325), .B(n10326), .ZN(n10329) );
  NAND2_X1 U12934 ( .A1(n13988), .A2(n13698), .ZN(n10328) );
  NAND2_X1 U12935 ( .A1(n13991), .A2(n13700), .ZN(n10327) );
  AND2_X1 U12936 ( .A1(n10328), .A2(n10327), .ZN(n10609) );
  OAI21_X1 U12937 ( .B1(n10329), .B2(n13950), .A(n10609), .ZN(n10778) );
  AOI211_X1 U12938 ( .C1(n15390), .C2(n10781), .A(n10774), .B(n10778), .ZN(
        n10335) );
  AOI22_X1 U12939 ( .A1(n14059), .A2(n12411), .B1(n15424), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10330) );
  OAI21_X1 U12940 ( .B1(n10335), .B2(n15424), .A(n10330), .ZN(P2_U3505) );
  INV_X1 U12941 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10331) );
  OAI22_X1 U12942 ( .A1(n10332), .A2(n14132), .B1(n15409), .B2(n10331), .ZN(
        n10333) );
  INV_X1 U12943 ( .A(n10333), .ZN(n10334) );
  OAI21_X1 U12944 ( .B1(n10335), .B2(n15407), .A(n10334), .ZN(P2_U3448) );
  NAND2_X1 U12945 ( .A1(n13044), .A2(P3_DATAO_REG_24__SCAN_IN), .ZN(n10336) );
  OAI21_X1 U12946 ( .B1(n13200), .B2(n13044), .A(n10336), .ZN(P3_U3515) );
  INV_X1 U12947 ( .A(n11384), .ZN(n10340) );
  INV_X1 U12948 ( .A(n13723), .ZN(n13733) );
  OAI222_X1 U12949 ( .A1(n14152), .A2(n10337), .B1(n14150), .B2(n10340), .C1(
        n13733), .C2(P2_U3088), .ZN(P2_U3313) );
  NAND2_X1 U12950 ( .A1(n10338), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10339) );
  INV_X1 U12951 ( .A(n14361), .ZN(n11180) );
  OAI222_X1 U12952 ( .A1(n14771), .A2(n10341), .B1(n14768), .B2(n10340), .C1(
        n11180), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12953 ( .A(n13217), .ZN(n13186) );
  NAND2_X1 U12954 ( .A1(n13186), .A2(P3_U3897), .ZN(n10342) );
  OAI21_X1 U12955 ( .B1(P3_U3897), .B2(n10343), .A(n10342), .ZN(P3_U3514) );
  OAI222_X1 U12956 ( .A1(n13468), .A2(n10346), .B1(n11518), .B2(n10345), .C1(
        P3_U3151), .C2(n10344), .ZN(P3_U3275) );
  OAI21_X1 U12957 ( .B1(n10353), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10347), .ZN(
        n10349) );
  INV_X1 U12958 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15422) );
  MUX2_X1 U12959 ( .A(n15422), .B(P2_REG1_REG_10__SCAN_IN), .S(n10380), .Z(
        n10348) );
  AOI21_X1 U12960 ( .B1(n10349), .B2(n10348), .A(n15214), .ZN(n10350) );
  NAND2_X1 U12961 ( .A1(n10350), .A2(n10377), .ZN(n10360) );
  NAND2_X1 U12962 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11327)
         );
  INV_X1 U12963 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10351) );
  MUX2_X1 U12964 ( .A(n10351), .B(P2_REG2_REG_10__SCAN_IN), .S(n10380), .Z(
        n10355) );
  OAI21_X1 U12965 ( .B1(n10353), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10352), .ZN(
        n10354) );
  NOR2_X1 U12966 ( .A1(n10354), .A2(n10355), .ZN(n10379) );
  AOI211_X1 U12967 ( .C1(n10355), .C2(n10354), .A(n10379), .B(n15221), .ZN(
        n10356) );
  INV_X1 U12968 ( .A(n10356), .ZN(n10357) );
  NAND2_X1 U12969 ( .A1(n11327), .A2(n10357), .ZN(n10358) );
  AOI21_X1 U12970 ( .B1(n15266), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10358), 
        .ZN(n10359) );
  OAI211_X1 U12971 ( .C1(n15265), .C2(n10361), .A(n10360), .B(n10359), .ZN(
        P2_U3224) );
  INV_X1 U12972 ( .A(n10362), .ZN(n10363) );
  NAND2_X1 U12973 ( .A1(n10363), .A2(n15624), .ZN(n10364) );
  XNOR2_X1 U12974 ( .A(n10366), .B(n12921), .ZN(n10526) );
  AOI21_X1 U12975 ( .B1(n10368), .B2(n10367), .A(n13027), .ZN(n10369) );
  NAND2_X1 U12976 ( .A1(n10369), .A2(n10529), .ZN(n10374) );
  OAI22_X1 U12977 ( .A1(n13035), .A2(n15624), .B1(n15630), .B2(n13040), .ZN(
        n10370) );
  AOI211_X1 U12978 ( .C1(n15430), .C2(n10372), .A(n10371), .B(n10370), .ZN(
        n10373) );
  OAI211_X1 U12979 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11233), .A(n10374), .B(
        n10373), .ZN(P3_U3158) );
  NAND2_X1 U12980 ( .A1(n10380), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10376) );
  INV_X1 U12981 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15425) );
  MUX2_X1 U12982 ( .A(n15425), .B(P2_REG1_REG_11__SCAN_IN), .S(n11081), .Z(
        n10375) );
  AOI21_X1 U12983 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n11080) );
  NAND3_X1 U12984 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n10378) );
  NAND2_X1 U12985 ( .A1(n10378), .A2(n15270), .ZN(n10388) );
  INV_X1 U12986 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11072) );
  MUX2_X1 U12987 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11072), .S(n11081), .Z(
        n10381) );
  NAND2_X1 U12988 ( .A1(n10382), .A2(n10381), .ZN(n15220) );
  OAI21_X1 U12989 ( .B1(n10382), .B2(n10381), .A(n15220), .ZN(n10383) );
  NAND2_X1 U12990 ( .A1(n10383), .A2(n15274), .ZN(n10387) );
  NAND2_X1 U12991 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11209)
         );
  INV_X1 U12992 ( .A(n11209), .ZN(n10385) );
  NOR2_X1 U12993 ( .A1(n15265), .A2(n11073), .ZN(n10384) );
  AOI211_X1 U12994 ( .C1(n15266), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10385), 
        .B(n10384), .ZN(n10386) );
  OAI211_X1 U12995 ( .C1(n11080), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        P2_U3225) );
  INV_X1 U12996 ( .A(n11454), .ZN(n10392) );
  OR2_X1 U12997 ( .A1(n10389), .A2(n10407), .ZN(n10390) );
  XNOR2_X1 U12998 ( .A(n10390), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11455) );
  INV_X1 U12999 ( .A(n11455), .ZN(n15024) );
  OAI222_X1 U13000 ( .A1(n14771), .A2(n10391), .B1(n14768), .B2(n10392), .C1(
        n15024), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13001 ( .A(n15244), .ZN(n13735) );
  OAI222_X1 U13002 ( .A1(n14152), .A2(n10393), .B1(n14150), .B2(n10392), .C1(
        n13735), .C2(P2_U3088), .ZN(P2_U3312) );
  XOR2_X1 U13003 ( .A(n10394), .B(n12620), .Z(n10813) );
  NAND2_X1 U13004 ( .A1(n10395), .A2(n12424), .ZN(n10396) );
  NAND2_X1 U13005 ( .A1(n10396), .A2(n11160), .ZN(n10397) );
  NOR2_X1 U13006 ( .A1(n10758), .A2(n10397), .ZN(n10806) );
  XNOR2_X1 U13007 ( .A(n10398), .B(n12620), .ZN(n10399) );
  AOI22_X1 U13008 ( .A1(n13991), .A2(n13699), .B1(n13988), .B2(n13697), .ZN(
        n10519) );
  OAI21_X1 U13009 ( .B1(n10399), .B2(n13950), .A(n10519), .ZN(n10810) );
  AOI211_X1 U13010 ( .C1(n15390), .C2(n10813), .A(n10806), .B(n10810), .ZN(
        n10404) );
  AOI22_X1 U13011 ( .A1(n14059), .A2(n12424), .B1(n15424), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10400) );
  OAI21_X1 U13012 ( .B1(n10404), .B2(n15424), .A(n10400), .ZN(P2_U3506) );
  INV_X1 U13013 ( .A(n12424), .ZN(n10523) );
  INV_X1 U13014 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10401) );
  OAI22_X1 U13015 ( .A1(n10523), .A2(n14132), .B1(n15409), .B2(n10401), .ZN(
        n10402) );
  INV_X1 U13016 ( .A(n10402), .ZN(n10403) );
  OAI21_X1 U13017 ( .B1(n10404), .B2(n15407), .A(n10403), .ZN(P2_U3451) );
  INV_X1 U13018 ( .A(n11596), .ZN(n10412) );
  NOR2_X1 U13019 ( .A1(n10405), .A2(n10407), .ZN(n10406) );
  MUX2_X1 U13020 ( .A(n10407), .B(n10406), .S(P1_IR_REG_16__SCAN_IN), .Z(
        n10409) );
  INV_X1 U13021 ( .A(n10551), .ZN(n10408) );
  OAI222_X1 U13022 ( .A1(n14771), .A2(n10410), .B1(n14768), .B2(n10412), .C1(
        n11372), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U13023 ( .A1(P2_U3088), .A2(n15264), .B1(n14150), .B2(n10412), 
        .C1(n10411), .C2(n14152), .ZN(P2_U3311) );
  INV_X1 U13024 ( .A(n13157), .ZN(n13187) );
  NAND2_X1 U13025 ( .A1(n13187), .A2(P3_U3897), .ZN(n10413) );
  OAI21_X1 U13026 ( .B1(P3_U3897), .B2(n10414), .A(n10413), .ZN(P3_U3516) );
  OAI222_X1 U13027 ( .A1(n13468), .A2(n10416), .B1(n11518), .B2(n10415), .C1(
        P3_U3151), .C2(n12176), .ZN(P3_U3274) );
  NAND2_X1 U13028 ( .A1(n10420), .A2(n11892), .ZN(n10422) );
  AOI22_X1 U13029 ( .A1(n11853), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11852), 
        .B2(n14344), .ZN(n10421) );
  OR2_X1 U13030 ( .A1(n11947), .A2(n6686), .ZN(n10424) );
  INV_X1 U13031 ( .A(n11946), .ZN(n14315) );
  NAND2_X1 U13032 ( .A1(n14315), .A2(n12817), .ZN(n10423) );
  NAND2_X1 U13033 ( .A1(n10424), .A2(n10423), .ZN(n10575) );
  OAI22_X1 U13034 ( .A1(n11947), .A2(n12823), .B1(n11946), .B2(n6686), .ZN(
        n10427) );
  XNOR2_X1 U13035 ( .A(n10427), .B(n12824), .ZN(n10578) );
  XNOR2_X1 U13036 ( .A(n10579), .B(n10578), .ZN(n10439) );
  INV_X1 U13037 ( .A(n11947), .ZN(n15077) );
  NAND2_X1 U13038 ( .A1(n14316), .A2(n14563), .ZN(n10435) );
  AOI21_X1 U13039 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10428) );
  NOR2_X1 U13040 ( .A1(n10428), .A2(n10594), .ZN(n10593) );
  NAND2_X1 U13041 ( .A1(n11889), .A2(n10593), .ZN(n10433) );
  OR2_X1 U13042 ( .A1(n11902), .A2(n15138), .ZN(n10432) );
  OR2_X1 U13043 ( .A1(n10273), .A2(n11147), .ZN(n10431) );
  INV_X1 U13044 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10429) );
  OR2_X1 U13045 ( .A1(n6689), .A2(n10429), .ZN(n10430) );
  NAND4_X1 U13046 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n14314) );
  NAND2_X1 U13047 ( .A1(n14314), .A2(n14565), .ZN(n10434) );
  NAND2_X1 U13048 ( .A1(n10435), .A2(n10434), .ZN(n15076) );
  AND2_X1 U13049 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14342) );
  AOI21_X1 U13050 ( .B1(n14953), .B2(n15076), .A(n14342), .ZN(n10436) );
  OAI21_X1 U13051 ( .B1(n14958), .B2(n10462), .A(n10436), .ZN(n10437) );
  AOI21_X1 U13052 ( .B1(n14950), .B2(n15077), .A(n10437), .ZN(n10438) );
  OAI21_X1 U13053 ( .B1(n10439), .B2(n14277), .A(n10438), .ZN(P1_U3230) );
  NAND2_X1 U13054 ( .A1(n13676), .A2(n13922), .ZN(n13663) );
  INV_X1 U13055 ( .A(n13663), .ZN(n13641) );
  NAND2_X1 U13056 ( .A1(n13641), .A2(n13705), .ZN(n10442) );
  AOI21_X1 U13057 ( .B1(n13705), .B2(n13922), .A(n13653), .ZN(n10440) );
  NOR2_X1 U13058 ( .A1(n10440), .A2(n13668), .ZN(n10441) );
  MUX2_X1 U13059 ( .A(n10442), .B(n10441), .S(n12367), .Z(n10445) );
  INV_X1 U13060 ( .A(n13988), .ZN(n15294) );
  NOR2_X1 U13061 ( .A1(n13646), .A2(n15294), .ZN(n13549) );
  OR2_X1 U13062 ( .A1(n10443), .A2(P2_U3088), .ZN(n13578) );
  AOI22_X1 U13063 ( .A1(n13549), .A2(n6854), .B1(n13578), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10444) );
  NAND2_X1 U13064 ( .A1(n10445), .A2(n10444), .ZN(P2_U3204) );
  XNOR2_X1 U13065 ( .A(n13505), .B(n12401), .ZN(n10491) );
  INV_X1 U13066 ( .A(n10446), .ZN(n11160) );
  NAND2_X1 U13067 ( .A1(n13922), .A2(n13701), .ZN(n10484) );
  XNOR2_X1 U13068 ( .A(n10491), .B(n10484), .ZN(n10448) );
  INV_X1 U13069 ( .A(n10448), .ZN(n10454) );
  INV_X1 U13070 ( .A(n10487), .ZN(n10493) );
  AOI21_X1 U13071 ( .B1(n10450), .B2(n10454), .A(n10493), .ZN(n10459) );
  INV_X1 U13072 ( .A(n12401), .ZN(n15368) );
  NAND2_X1 U13073 ( .A1(n13549), .A2(n13700), .ZN(n10452) );
  OAI211_X1 U13074 ( .C1(n15368), .C2(n13662), .A(n10452), .B(n10451), .ZN(
        n10457) );
  NAND3_X1 U13075 ( .A1(n13641), .A2(n10454), .A3(n10453), .ZN(n10455) );
  INV_X1 U13076 ( .A(n13659), .ZN(n13630) );
  AOI21_X1 U13077 ( .B1(n10455), .B2(n13630), .A(n12390), .ZN(n10456) );
  AOI211_X1 U13078 ( .C1(n13649), .C2(n10742), .A(n10457), .B(n10456), .ZN(
        n10458) );
  OAI21_X1 U13079 ( .B1(n10459), .B2(n13653), .A(n10458), .ZN(P2_U3202) );
  INV_X1 U13080 ( .A(n10460), .ZN(n10461) );
  INV_X1 U13081 ( .A(n14633), .ZN(n15070) );
  INV_X1 U13082 ( .A(n10462), .ZN(n10469) );
  NAND2_X1 U13083 ( .A1(n10463), .A2(n11936), .ZN(n10465) );
  INV_X1 U13084 ( .A(n14316), .ZN(n11940) );
  NAND2_X1 U13085 ( .A1(n11941), .A2(n11940), .ZN(n10464) );
  XNOR2_X1 U13086 ( .A(n15077), .B(n11946), .ZN(n11859) );
  INV_X1 U13087 ( .A(n11859), .ZN(n10466) );
  XNOR2_X1 U13088 ( .A(n10962), .B(n10466), .ZN(n10467) );
  NAND2_X1 U13089 ( .A1(n10467), .A2(n14792), .ZN(n15080) );
  INV_X1 U13090 ( .A(n15080), .ZN(n10468) );
  AOI211_X1 U13091 ( .C1(n15070), .C2(n10469), .A(n15076), .B(n10468), .ZN(
        n10483) );
  OR2_X1 U13092 ( .A1(n11941), .A2(n14316), .ZN(n10472) );
  XNOR2_X1 U13093 ( .A(n10898), .B(n11859), .ZN(n15082) );
  INV_X1 U13094 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U13095 ( .A1(n14636), .A2(n10475), .ZN(n15067) );
  NOR2_X1 U13096 ( .A1(n10476), .A2(n12089), .ZN(n10477) );
  OAI22_X1 U13097 ( .A1(n14614), .A2(n11947), .B1(n10478), .B2(n14636), .ZN(
        n10481) );
  NAND2_X1 U13098 ( .A1(n11947), .A2(n10479), .ZN(n11137) );
  OAI211_X1 U13099 ( .C1(n11947), .C2(n10479), .A(n15055), .B(n11137), .ZN(
        n15078) );
  NOR2_X1 U13100 ( .A1(n14654), .A2(n15078), .ZN(n10480) );
  AOI211_X1 U13101 ( .C1(n15082), .C2(n14656), .A(n10481), .B(n10480), .ZN(
        n10482) );
  OAI21_X1 U13102 ( .B1(n10483), .B2(n15074), .A(n10482), .ZN(P1_U3289) );
  INV_X1 U13103 ( .A(n10491), .ZN(n10485) );
  NAND2_X1 U13104 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  XNOR2_X1 U13105 ( .A(n15377), .B(n13493), .ZN(n10498) );
  NAND2_X1 U13106 ( .A1(n13922), .A2(n13700), .ZN(n10499) );
  XNOR2_X1 U13107 ( .A(n10498), .B(n10499), .ZN(n10492) );
  INV_X1 U13108 ( .A(n15377), .ZN(n10858) );
  INV_X1 U13109 ( .A(n13646), .ZN(n13671) );
  NAND2_X1 U13110 ( .A1(n13988), .A2(n13699), .ZN(n10489) );
  NAND2_X1 U13111 ( .A1(n13991), .A2(n13701), .ZN(n10488) );
  NAND2_X1 U13112 ( .A1(n10489), .A2(n10488), .ZN(n10850) );
  NAND2_X1 U13113 ( .A1(n13671), .A2(n10850), .ZN(n10490) );
  NAND2_X1 U13114 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15181) );
  OAI211_X1 U13115 ( .C1(n13662), .C2(n10858), .A(n10490), .B(n15181), .ZN(
        n10496) );
  AOI22_X1 U13116 ( .A1(n13641), .A2(n13701), .B1(n13676), .B2(n10491), .ZN(
        n10494) );
  NOR3_X1 U13117 ( .A1(n10494), .A2(n10493), .A3(n10492), .ZN(n10495) );
  AOI211_X1 U13118 ( .C1(n13649), .C2(n10856), .A(n10496), .B(n10495), .ZN(
        n10497) );
  OAI21_X1 U13119 ( .B1(n10502), .B2(n13653), .A(n10497), .ZN(P2_U3199) );
  INV_X1 U13120 ( .A(n10498), .ZN(n10500) );
  NAND2_X1 U13121 ( .A1(n10500), .A2(n10499), .ZN(n10501) );
  XNOR2_X1 U13122 ( .A(n12411), .B(n13505), .ZN(n10503) );
  AND2_X1 U13123 ( .A1(n13509), .A2(n13699), .ZN(n10504) );
  NAND2_X1 U13124 ( .A1(n10503), .A2(n10504), .ZN(n10514) );
  INV_X1 U13125 ( .A(n10503), .ZN(n10513) );
  INV_X1 U13126 ( .A(n10504), .ZN(n10505) );
  NAND2_X1 U13127 ( .A1(n10513), .A2(n10505), .ZN(n10506) );
  NAND2_X1 U13128 ( .A1(n10514), .A2(n10506), .ZN(n10613) );
  INV_X1 U13129 ( .A(n10613), .ZN(n10507) );
  XNOR2_X1 U13130 ( .A(n12424), .B(n13505), .ZN(n10686) );
  AND2_X1 U13131 ( .A1(n13509), .A2(n13698), .ZN(n10508) );
  NAND2_X1 U13132 ( .A1(n10686), .A2(n10508), .ZN(n10684) );
  INV_X1 U13133 ( .A(n10686), .ZN(n10510) );
  INV_X1 U13134 ( .A(n10508), .ZN(n10509) );
  NAND2_X1 U13135 ( .A1(n10510), .A2(n10509), .ZN(n10511) );
  AND2_X1 U13136 ( .A1(n10684), .A2(n10511), .ZN(n10515) );
  INV_X1 U13137 ( .A(n10515), .ZN(n10512) );
  AOI21_X1 U13138 ( .B1(n10610), .B2(n10512), .A(n13653), .ZN(n10518) );
  NOR3_X1 U13139 ( .A1(n13663), .A2(n12413), .A3(n10513), .ZN(n10517) );
  NAND2_X1 U13140 ( .A1(n10516), .A2(n10515), .ZN(n10688) );
  OAI21_X1 U13141 ( .B1(n10518), .B2(n10517), .A(n10688), .ZN(n10522) );
  NAND2_X1 U13142 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15196) );
  OAI21_X1 U13143 ( .B1(n13646), .B2(n10519), .A(n15196), .ZN(n10520) );
  AOI21_X1 U13144 ( .B1(n13649), .B2(n10807), .A(n10520), .ZN(n10521) );
  OAI211_X1 U13145 ( .C1(n10523), .C2(n13662), .A(n10522), .B(n10521), .ZN(
        P2_U3185) );
  INV_X1 U13146 ( .A(n10524), .ZN(n10796) );
  XNOR2_X1 U13147 ( .A(n10525), .B(n12848), .ZN(n10700) );
  XNOR2_X1 U13148 ( .A(n10700), .B(n15623), .ZN(n10531) );
  INV_X1 U13149 ( .A(n10526), .ZN(n10527) );
  NAND2_X1 U13150 ( .A1(n10799), .A2(n10527), .ZN(n10528) );
  OAI21_X1 U13151 ( .B1(n10531), .B2(n10530), .A(n10703), .ZN(n10532) );
  NAND2_X1 U13152 ( .A1(n10532), .A2(n15432), .ZN(n10536) );
  NAND2_X1 U13153 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15448) );
  INV_X1 U13154 ( .A(n15448), .ZN(n10534) );
  OAI22_X1 U13155 ( .A1(n13035), .A2(n15636), .B1(n15703), .B2(n13040), .ZN(
        n10533) );
  AOI211_X1 U13156 ( .C1(n15430), .C2(n12199), .A(n10534), .B(n10533), .ZN(
        n10535) );
  OAI211_X1 U13157 ( .C1(n10796), .C2(n11233), .A(n10536), .B(n10535), .ZN(
        P3_U3170) );
  OAI22_X1 U13158 ( .A1(n13662), .A2(n10538), .B1(n10537), .B2(n13646), .ZN(
        n10544) );
  AOI22_X1 U13159 ( .A1(n13641), .A2(n6854), .B1(n13676), .B2(n10539), .ZN(
        n10542) );
  INV_X1 U13160 ( .A(n13574), .ZN(n10541) );
  NOR3_X1 U13161 ( .A1(n10542), .A2(n10541), .A3(n10540), .ZN(n10543) );
  AOI211_X1 U13162 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n13578), .A(n10544), .B(
        n10543), .ZN(n10545) );
  OAI21_X1 U13163 ( .B1(n10546), .B2(n13653), .A(n10545), .ZN(P2_U3209) );
  INV_X1 U13164 ( .A(n10547), .ZN(n10549) );
  OAI22_X1 U13165 ( .A1(n12359), .A2(P3_U3151), .B1(SI_22_), .B2(n13471), .ZN(
        n10548) );
  AOI21_X1 U13166 ( .B1(n10549), .B2(n13455), .A(n10548), .ZN(P3_U3273) );
  INV_X1 U13167 ( .A(n11851), .ZN(n10553) );
  OAI222_X1 U13168 ( .A1(P2_U3088), .A2(n13739), .B1(n14150), .B2(n10553), 
        .C1(n10550), .C2(n14152), .ZN(P2_U3310) );
  NAND2_X1 U13169 ( .A1(n10551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10552) );
  XNOR2_X1 U13170 ( .A(n10552), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14376) );
  INV_X1 U13171 ( .A(n14376), .ZN(n14373) );
  OAI222_X1 U13172 ( .A1(n14764), .A2(n10554), .B1(n14768), .B2(n10553), .C1(
        n14373), .C2(P1_U3086), .ZN(P1_U3338) );
  XNOR2_X1 U13173 ( .A(n10555), .B(n12622), .ZN(n10889) );
  NAND3_X1 U13174 ( .A1(n10556), .A2(n15343), .A3(n12667), .ZN(n10557) );
  OR2_X1 U13175 ( .A1(n10558), .A2(n10557), .ZN(n10559) );
  NAND2_X1 U13176 ( .A1(n12646), .A2(n12666), .ZN(n10669) );
  INV_X1 U13177 ( .A(n10669), .ZN(n10560) );
  NAND2_X1 U13178 ( .A1(n15303), .A2(n10560), .ZN(n15300) );
  OAI21_X1 U13179 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(n10565) );
  OAI22_X1 U13180 ( .A1(n12430), .A2(n13953), .B1(n15294), .B2(n12454), .ZN(
        n10564) );
  AOI21_X1 U13181 ( .B1(n10565), .B2(n15293), .A(n10564), .ZN(n10566) );
  NAND2_X1 U13182 ( .A1(n10890), .A2(n15303), .ZN(n10572) );
  INV_X1 U13183 ( .A(n10839), .ZN(n10567) );
  AOI211_X1 U13184 ( .C1(n12441), .C2(n10757), .A(n10446), .B(n10567), .ZN(
        n10891) );
  NAND2_X1 U13185 ( .A1(n15303), .A2(n10568), .ZN(n13998) );
  AOI22_X1 U13186 ( .A1(n15305), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10879), 
        .B2(n15283), .ZN(n10569) );
  OAI21_X1 U13187 ( .B1(n7193), .B2(n13998), .A(n10569), .ZN(n10570) );
  AOI21_X1 U13188 ( .B1(n10891), .B2(n15285), .A(n10570), .ZN(n10571) );
  OAI211_X1 U13189 ( .C1(n10889), .C2(n15300), .A(n10572), .B(n10571), .ZN(
        P2_U3256) );
  NAND2_X1 U13190 ( .A1(n13143), .A2(P3_U3897), .ZN(n10573) );
  OAI21_X1 U13191 ( .B1(P3_U3897), .B2(n10574), .A(n10573), .ZN(P3_U3517) );
  NAND2_X1 U13192 ( .A1(n10580), .A2(n11892), .ZN(n10583) );
  AOI22_X1 U13193 ( .A1(n11853), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11852), 
        .B2(n10581), .ZN(n10582) );
  NAND2_X1 U13194 ( .A1(n10583), .A2(n10582), .ZN(n15084) );
  NAND2_X1 U13195 ( .A1(n15084), .A2(n12804), .ZN(n10585) );
  NAND2_X1 U13196 ( .A1(n10585), .A2(n10584), .ZN(n10586) );
  XNOR2_X1 U13197 ( .A(n10586), .B(n12824), .ZN(n10590) );
  NAND2_X1 U13198 ( .A1(n15084), .A2(n7074), .ZN(n10588) );
  NAND2_X1 U13199 ( .A1(n12817), .A2(n14314), .ZN(n10587) );
  NAND2_X1 U13200 ( .A1(n10588), .A2(n10587), .ZN(n10589) );
  NOR2_X1 U13201 ( .A1(n10590), .A2(n10589), .ZN(n10710) );
  NAND2_X1 U13202 ( .A1(n10590), .A2(n10589), .ZN(n10709) );
  INV_X1 U13203 ( .A(n10709), .ZN(n10591) );
  NOR2_X1 U13204 ( .A1(n10710), .A2(n10591), .ZN(n10592) );
  XNOR2_X1 U13205 ( .A(n10711), .B(n10592), .ZN(n10605) );
  INV_X1 U13206 ( .A(n10593), .ZN(n11140) );
  OR2_X1 U13207 ( .A1(n11946), .A2(n14460), .ZN(n10601) );
  NAND2_X1 U13208 ( .A1(n11807), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10599) );
  OR2_X1 U13209 ( .A1(n10273), .A2(n9612), .ZN(n10598) );
  NAND2_X1 U13210 ( .A1(n10594), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10721) );
  OAI21_X1 U13211 ( .B1(n10594), .B2(P1_REG3_REG_6__SCAN_IN), .A(n10721), .ZN(
        n15050) );
  OR2_X1 U13212 ( .A1(n11900), .A2(n15050), .ZN(n10597) );
  INV_X1 U13213 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10595) );
  OR2_X1 U13214 ( .A1(n6689), .A2(n10595), .ZN(n10596) );
  NAND4_X1 U13215 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n14313) );
  NAND2_X1 U13216 ( .A1(n14313), .A2(n14565), .ZN(n10600) );
  NAND2_X1 U13217 ( .A1(n10601), .A2(n10600), .ZN(n11145) );
  AOI22_X1 U13218 ( .A1(n14953), .A2(n11145), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10603) );
  NAND2_X1 U13219 ( .A1(n14950), .A2(n15084), .ZN(n10602) );
  OAI211_X1 U13220 ( .C1(n14958), .C2(n11140), .A(n10603), .B(n10602), .ZN(
        n10604) );
  AOI21_X1 U13221 ( .B1(n10605), .B2(n14951), .A(n10604), .ZN(n10606) );
  INV_X1 U13222 ( .A(n10606), .ZN(P1_U3227) );
  NAND2_X1 U13223 ( .A1(n13668), .A2(n12411), .ZN(n10608) );
  OAI211_X1 U13224 ( .C1(n10609), .C2(n13646), .A(n10608), .B(n10607), .ZN(
        n10615) );
  INV_X1 U13225 ( .A(n10610), .ZN(n10611) );
  AOI211_X1 U13226 ( .C1(n10613), .C2(n10612), .A(n13653), .B(n10611), .ZN(
        n10614) );
  AOI211_X1 U13227 ( .C1(n13649), .C2(n10775), .A(n10615), .B(n10614), .ZN(
        n10616) );
  INV_X1 U13228 ( .A(n10616), .ZN(P2_U3211) );
  INV_X1 U13229 ( .A(n15470), .ZN(n10636) );
  NOR2_X1 U13230 ( .A1(n10618), .A2(n10617), .ZN(n10620) );
  AOI22_X1 U13231 ( .A1(n10652), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n7301), .B2(
        n15459), .ZN(n15454) );
  NOR2_X1 U13232 ( .A1(n10636), .A2(n10621), .ZN(n10622) );
  INV_X1 U13233 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15474) );
  INV_X1 U13234 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13235 ( .A1(n10654), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n10623), 
        .B2(n15487), .ZN(n15491) );
  INV_X1 U13236 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15505) );
  NOR2_X1 U13237 ( .A1(n10625), .A2(n10626), .ZN(n10627) );
  NAND2_X1 U13238 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n13091), .ZN(n10628) );
  OAI21_X1 U13239 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13091), .A(n10628), 
        .ZN(n10629) );
  AOI21_X1 U13240 ( .B1(n10630), .B2(n10629), .A(n13046), .ZN(n10668) );
  INV_X1 U13241 ( .A(n13091), .ZN(n10659) );
  INV_X1 U13242 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U13243 ( .A1(n10659), .A2(n15762), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n13091), .ZN(n10643) );
  INV_X1 U13244 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U13245 ( .A1(n10654), .A2(n15757), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15487), .ZN(n15486) );
  INV_X1 U13246 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15753) );
  AOI22_X1 U13247 ( .A1(n10652), .A2(n15753), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15459), .ZN(n15458) );
  NAND2_X1 U13248 ( .A1(n10646), .A2(n10631), .ZN(n10633) );
  NAND2_X1 U13249 ( .A1(n10633), .A2(n10632), .ZN(n15457) );
  NAND2_X1 U13250 ( .A1(n15458), .A2(n15457), .ZN(n10634) );
  NAND2_X1 U13251 ( .A1(n15470), .A2(n10635), .ZN(n10638) );
  NAND2_X1 U13252 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15469), .ZN(n10637) );
  NAND2_X1 U13253 ( .A1(n10638), .A2(n10637), .ZN(n15485) );
  NAND2_X1 U13254 ( .A1(n15486), .A2(n15485), .ZN(n10639) );
  NAND2_X1 U13255 ( .A1(n15510), .A2(n10640), .ZN(n10641) );
  NAND2_X1 U13256 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15509), .ZN(n15508) );
  NAND2_X1 U13257 ( .A1(n10641), .A2(n15508), .ZN(n10642) );
  NAND2_X1 U13258 ( .A1(n10643), .A2(n10642), .ZN(n13092) );
  OAI21_X1 U13259 ( .B1(n10643), .B2(n10642), .A(n13092), .ZN(n10666) );
  NOR2_X1 U13260 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10644), .ZN(n11539) );
  AOI21_X1 U13261 ( .B1(n15581), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11539), 
        .ZN(n10664) );
  INV_X1 U13262 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15759) );
  MUX2_X1 U13263 ( .A(n15505), .B(n15759), .S(n6678), .Z(n10657) );
  INV_X1 U13264 ( .A(n10657), .ZN(n10645) );
  NAND2_X1 U13265 ( .A1(n10645), .A2(n15510), .ZN(n15500) );
  MUX2_X1 U13266 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n6678), .Z(n10655) );
  OR2_X1 U13267 ( .A1(n10655), .A2(n15487), .ZN(n10656) );
  OAI22_X1 U13268 ( .A1(n10649), .A2(n10648), .B1(n10647), .B2(n10646), .ZN(
        n15452) );
  MUX2_X1 U13269 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6678), .Z(n10650) );
  XNOR2_X1 U13270 ( .A(n10650), .B(n10652), .ZN(n15451) );
  INV_X1 U13271 ( .A(n10650), .ZN(n10651) );
  AOI22_X1 U13272 ( .A1(n15452), .A2(n15451), .B1(n10652), .B2(n10651), .ZN(
        n15468) );
  MUX2_X1 U13273 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6678), .Z(n10653) );
  XNOR2_X1 U13274 ( .A(n10653), .B(n15470), .ZN(n15467) );
  OAI22_X1 U13275 ( .A1(n15468), .A2(n15467), .B1(n10653), .B2(n15470), .ZN(
        n15484) );
  XNOR2_X1 U13276 ( .A(n10655), .B(n10654), .ZN(n15483) );
  NAND2_X1 U13277 ( .A1(n15484), .A2(n15483), .ZN(n15482) );
  NAND2_X1 U13278 ( .A1(n10656), .A2(n15482), .ZN(n15503) );
  NAND2_X1 U13279 ( .A1(n15500), .A2(n15503), .ZN(n10658) );
  NAND2_X1 U13280 ( .A1(n10657), .A2(n10625), .ZN(n15501) );
  NAND2_X1 U13281 ( .A1(n10658), .A2(n15501), .ZN(n10661) );
  MUX2_X1 U13282 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n6678), .Z(n13060) );
  XNOR2_X1 U13283 ( .A(n13060), .B(n10659), .ZN(n10660) );
  NAND2_X1 U13284 ( .A1(n10661), .A2(n10660), .ZN(n13062) );
  OAI21_X1 U13285 ( .B1(n10661), .B2(n10660), .A(n13062), .ZN(n10662) );
  NAND2_X1 U13286 ( .A1(n10662), .A2(n15588), .ZN(n10663) );
  OAI211_X1 U13287 ( .C1(n15584), .C2(n13091), .A(n10664), .B(n10663), .ZN(
        n10665) );
  AOI21_X1 U13288 ( .B1(n10666), .B2(n15586), .A(n10665), .ZN(n10667) );
  OAI21_X1 U13289 ( .B1(n10668), .B2(n15594), .A(n10667), .ZN(P3_U3192) );
  XNOR2_X1 U13290 ( .A(n12612), .B(n13572), .ZN(n15354) );
  INV_X1 U13291 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10681) );
  INV_X1 U13292 ( .A(n10670), .ZN(n10671) );
  AOI211_X1 U13293 ( .C1(n12367), .C2(n12363), .A(n13922), .B(n10671), .ZN(
        n15350) );
  AOI22_X1 U13294 ( .A1(n15281), .A2(n12363), .B1(n15285), .B2(n15350), .ZN(
        n10680) );
  OAI21_X1 U13295 ( .B1(n10673), .B2(n12612), .A(n10672), .ZN(n10674) );
  NAND2_X1 U13296 ( .A1(n10674), .A2(n15293), .ZN(n10678) );
  NAND2_X1 U13297 ( .A1(n13988), .A2(n13703), .ZN(n10676) );
  NAND2_X1 U13298 ( .A1(n13991), .A2(n13705), .ZN(n10675) );
  NAND2_X1 U13299 ( .A1(n10676), .A2(n10675), .ZN(n13573) );
  INV_X1 U13300 ( .A(n13573), .ZN(n10677) );
  NAND2_X1 U13301 ( .A1(n10678), .A2(n10677), .ZN(n15349) );
  AOI22_X1 U13302 ( .A1(n15303), .A2(n15349), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15283), .ZN(n10679) );
  OAI211_X1 U13303 ( .C1(n10681), .C2(n15303), .A(n10680), .B(n10679), .ZN(
        n10682) );
  AOI21_X1 U13304 ( .B1(n15354), .B2(n15287), .A(n10682), .ZN(n10683) );
  INV_X1 U13305 ( .A(n10683), .ZN(P2_U3264) );
  XNOR2_X1 U13306 ( .A(n12428), .B(n13505), .ZN(n10882) );
  NAND2_X1 U13307 ( .A1(n13922), .A2(n13697), .ZN(n10874) );
  XNOR2_X1 U13308 ( .A(n10882), .B(n10874), .ZN(n10689) );
  AND2_X1 U13309 ( .A1(n10689), .A2(n10684), .ZN(n10685) );
  NAND3_X1 U13310 ( .A1(n13641), .A2(n13698), .A3(n10686), .ZN(n10687) );
  OAI21_X1 U13311 ( .B1(n10688), .B2(n13653), .A(n10687), .ZN(n10691) );
  INV_X1 U13312 ( .A(n10689), .ZN(n10690) );
  NAND2_X1 U13313 ( .A1(n10691), .A2(n10690), .ZN(n10697) );
  AOI21_X1 U13314 ( .B1(n13549), .B2(n13695), .A(n10692), .ZN(n10696) );
  AOI22_X1 U13315 ( .A1(n10693), .A2(n13649), .B1(n13659), .B2(n13698), .ZN(
        n10695) );
  NAND2_X1 U13316 ( .A1(n13668), .A2(n12428), .ZN(n10694) );
  AND4_X1 U13317 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10698) );
  OAI21_X1 U13318 ( .B1(n10877), .B2(n13653), .A(n10698), .ZN(P2_U3193) );
  NAND2_X1 U13319 ( .A1(n13044), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10699) );
  OAI21_X1 U13320 ( .B1(n12928), .B2(n13044), .A(n10699), .ZN(P3_U3520) );
  XNOR2_X1 U13321 ( .A(n15617), .B(n12921), .ZN(n10819) );
  XNOR2_X1 U13322 ( .A(n10819), .B(n12199), .ZN(n10821) );
  INV_X1 U13323 ( .A(n10700), .ZN(n10701) );
  NAND2_X1 U13324 ( .A1(n10701), .A2(n15623), .ZN(n10702) );
  XOR2_X1 U13325 ( .A(n10822), .B(n10821), .Z(n10708) );
  OAI22_X1 U13326 ( .A1(n13035), .A2(n15623), .B1(n12198), .B2(n13040), .ZN(
        n10704) );
  AOI211_X1 U13327 ( .C1(n15430), .C2(n11109), .A(n10705), .B(n10704), .ZN(
        n10707) );
  NAND2_X1 U13328 ( .A1(n13037), .A2(n15618), .ZN(n10706) );
  OAI211_X1 U13329 ( .C1(n10708), .C2(n13027), .A(n10707), .B(n10706), .ZN(
        P3_U3167) );
  NAND2_X1 U13330 ( .A1(n10712), .A2(n11892), .ZN(n10715) );
  AOI22_X1 U13331 ( .A1(n11853), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11852), 
        .B2(n10713), .ZN(n10714) );
  NAND2_X1 U13332 ( .A1(n10715), .A2(n10714), .ZN(n15053) );
  INV_X1 U13333 ( .A(n14313), .ZN(n10970) );
  NOR2_X1 U13334 ( .A1(n10970), .A2(n12826), .ZN(n10716) );
  AOI21_X1 U13335 ( .B1(n15053), .B2(n7074), .A(n10716), .ZN(n11054) );
  AOI22_X1 U13336 ( .A1(n15053), .A2(n12804), .B1(n11309), .B2(n14313), .ZN(
        n10717) );
  XNOR2_X1 U13337 ( .A(n10717), .B(n12824), .ZN(n11055) );
  XOR2_X1 U13338 ( .A(n11054), .B(n11055), .Z(n10718) );
  OAI211_X1 U13339 ( .C1(n10719), .C2(n10718), .A(n11059), .B(n14951), .ZN(
        n10734) );
  NAND2_X1 U13340 ( .A1(n14314), .A2(n14563), .ZN(n10729) );
  NAND2_X1 U13341 ( .A1(n6675), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10727) );
  OR2_X1 U13342 ( .A1(n11902), .A2(n15142), .ZN(n10726) );
  AND2_X1 U13343 ( .A1(n10721), .A2(n10720), .ZN(n10722) );
  OR2_X1 U13344 ( .A1(n10722), .A2(n10913), .ZN(n11096) );
  OR2_X1 U13345 ( .A1(n11900), .A2(n11096), .ZN(n10725) );
  INV_X1 U13346 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10723) );
  OR2_X1 U13347 ( .A1(n6689), .A2(n10723), .ZN(n10724) );
  NAND4_X1 U13348 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n14312) );
  NAND2_X1 U13349 ( .A1(n14312), .A2(n14565), .ZN(n10728) );
  NAND2_X1 U13350 ( .A1(n10729), .A2(n10728), .ZN(n15049) );
  AOI21_X1 U13351 ( .B1(n14953), .B2(n15049), .A(n10730), .ZN(n10731) );
  OAI21_X1 U13352 ( .B1(n14958), .B2(n15050), .A(n10731), .ZN(n10732) );
  AOI21_X1 U13353 ( .B1(n14950), .B2(n15053), .A(n10732), .ZN(n10733) );
  NAND2_X1 U13354 ( .A1(n10734), .A2(n10733), .ZN(P1_U3239) );
  XNOR2_X1 U13355 ( .A(n10735), .B(n10737), .ZN(n15372) );
  XNOR2_X1 U13356 ( .A(n10737), .B(n10736), .ZN(n10739) );
  AOI22_X1 U13357 ( .A1(n13991), .A2(n13702), .B1(n13988), .B2(n13700), .ZN(
        n10738) );
  OAI21_X1 U13358 ( .B1(n10739), .B2(n13950), .A(n10738), .ZN(n10740) );
  AOI21_X1 U13359 ( .B1(n15376), .B2(n15372), .A(n10740), .ZN(n15369) );
  INV_X1 U13360 ( .A(n15300), .ZN(n11040) );
  INV_X1 U13361 ( .A(n10741), .ZN(n10864) );
  OAI211_X1 U13362 ( .C1(n10864), .C2(n15368), .A(n11160), .B(n10852), .ZN(
        n15367) );
  INV_X1 U13363 ( .A(n10742), .ZN(n10743) );
  OAI22_X1 U13364 ( .A1(n15303), .A2(n10744), .B1(n10743), .B2(n15298), .ZN(
        n10745) );
  AOI21_X1 U13365 ( .B1(n15281), .B2(n12401), .A(n10745), .ZN(n10746) );
  OAI21_X1 U13366 ( .B1(n13907), .B2(n15367), .A(n10746), .ZN(n10747) );
  AOI21_X1 U13367 ( .B1(n11040), .B2(n15372), .A(n10747), .ZN(n10748) );
  OAI21_X1 U13368 ( .B1(n15305), .B2(n15369), .A(n10748), .ZN(P2_U3261) );
  XOR2_X1 U13369 ( .A(n12621), .B(n10749), .Z(n15388) );
  INV_X1 U13370 ( .A(n15388), .ZN(n10763) );
  INV_X1 U13371 ( .A(n10750), .ZN(n10751) );
  AOI21_X1 U13372 ( .B1(n12621), .B2(n10752), .A(n10751), .ZN(n10755) );
  NAND2_X1 U13373 ( .A1(n15388), .A2(n15376), .ZN(n10754) );
  AOI22_X1 U13374 ( .A1(n13991), .A2(n13698), .B1(n13988), .B2(n13695), .ZN(
        n10753) );
  OAI211_X1 U13375 ( .C1(n10755), .C2(n13950), .A(n10754), .B(n10753), .ZN(
        n15386) );
  NAND2_X1 U13376 ( .A1(n15386), .A2(n15303), .ZN(n10762) );
  OAI22_X1 U13377 ( .A1(n15303), .A2(n9920), .B1(n10756), .B2(n15298), .ZN(
        n10760) );
  OAI211_X1 U13378 ( .C1(n15385), .C2(n10758), .A(n11160), .B(n10757), .ZN(
        n15384) );
  NOR2_X1 U13379 ( .A1(n13907), .A2(n15384), .ZN(n10759) );
  AOI211_X1 U13380 ( .C1(n15281), .C2(n12428), .A(n10760), .B(n10759), .ZN(
        n10761) );
  OAI211_X1 U13381 ( .C1(n10763), .C2(n15300), .A(n10762), .B(n10761), .ZN(
        P2_U3257) );
  NAND2_X1 U13382 ( .A1(n12925), .A2(P3_U3897), .ZN(n10764) );
  OAI21_X1 U13383 ( .B1(P3_U3897), .B2(n10765), .A(n10764), .ZN(P3_U3518) );
  NAND2_X1 U13384 ( .A1(n8890), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U13385 ( .A1(n10766), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10768) );
  NAND2_X1 U13386 ( .A1(n8951), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10767) );
  AND3_X1 U13387 ( .A1(n10769), .A2(n10768), .A3(n10767), .ZN(n10770) );
  NAND2_X1 U13388 ( .A1(n10771), .A2(n10770), .ZN(n13116) );
  NAND2_X1 U13389 ( .A1(n13116), .A2(P3_U3897), .ZN(n10772) );
  OAI21_X1 U13390 ( .B1(P3_U3897), .B2(n10773), .A(n10772), .ZN(P3_U3522) );
  INV_X1 U13391 ( .A(n10774), .ZN(n10777) );
  AOI22_X1 U13392 ( .A1(n15281), .A2(n12411), .B1(n15283), .B2(n10775), .ZN(
        n10776) );
  OAI21_X1 U13393 ( .B1(n10777), .B2(n13907), .A(n10776), .ZN(n10780) );
  MUX2_X1 U13394 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10778), .S(n15303), .Z(
        n10779) );
  AOI211_X1 U13395 ( .C1(n15287), .C2(n10781), .A(n10780), .B(n10779), .ZN(
        n10782) );
  INV_X1 U13396 ( .A(n10782), .ZN(P2_U3259) );
  XNOR2_X1 U13397 ( .A(n10784), .B(n10783), .ZN(n15704) );
  INV_X1 U13398 ( .A(n15704), .ZN(n10804) );
  NAND2_X1 U13399 ( .A1(n10786), .A2(n10785), .ZN(n10790) );
  NAND2_X1 U13400 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  AND2_X1 U13401 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  AND2_X1 U13402 ( .A1(n12171), .A2(n12323), .ZN(n15616) );
  NAND2_X1 U13403 ( .A1(n15682), .A2(n15616), .ZN(n11453) );
  INV_X1 U13404 ( .A(n11453), .ZN(n15666) );
  OAI22_X1 U13405 ( .A1(n13320), .A2(n15703), .B1(n10796), .B2(n15676), .ZN(
        n10803) );
  XNOR2_X1 U13406 ( .A(n10797), .B(n12328), .ZN(n10798) );
  NAND2_X1 U13407 ( .A1(n10798), .A2(n15671), .ZN(n10801) );
  AOI22_X1 U13408 ( .A1(n10799), .A2(n15653), .B1(n15654), .B2(n12199), .ZN(
        n10800) );
  OAI211_X1 U13409 ( .C1(n15704), .C2(n15662), .A(n10801), .B(n10800), .ZN(
        n15706) );
  MUX2_X1 U13410 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15706), .S(n15682), .Z(
        n10802) );
  AOI211_X1 U13411 ( .C1(n10804), .C2(n15666), .A(n10803), .B(n10802), .ZN(
        n10805) );
  INV_X1 U13412 ( .A(n10805), .ZN(P3_U3229) );
  INV_X1 U13413 ( .A(n10806), .ZN(n10809) );
  AOI22_X1 U13414 ( .A1(n15281), .A2(n12424), .B1(n10807), .B2(n15283), .ZN(
        n10808) );
  OAI21_X1 U13415 ( .B1(n13907), .B2(n10809), .A(n10808), .ZN(n10812) );
  MUX2_X1 U13416 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10810), .S(n15303), .Z(
        n10811) );
  AOI211_X1 U13417 ( .C1(n15287), .C2(n10813), .A(n10812), .B(n10811), .ZN(
        n10814) );
  INV_X1 U13418 ( .A(n10814), .ZN(P2_U3258) );
  NAND2_X1 U13419 ( .A1(n10815), .A2(n13455), .ZN(n10816) );
  OAI211_X1 U13420 ( .C1(n10817), .C2(n13471), .A(n10816), .B(n12362), .ZN(
        P3_U3272) );
  INV_X1 U13421 ( .A(n10818), .ZN(n11004) );
  AND2_X1 U13422 ( .A1(n10819), .A2(n10826), .ZN(n10820) );
  XNOR2_X1 U13423 ( .A(n10823), .B(n12848), .ZN(n11108) );
  XNOR2_X1 U13424 ( .A(n15611), .B(n11108), .ZN(n10824) );
  NAND2_X1 U13425 ( .A1(n10825), .A2(n10824), .ZN(n11111) );
  OAI211_X1 U13426 ( .C1(n10825), .C2(n10824), .A(n11111), .B(n15432), .ZN(
        n10830) );
  NAND2_X1 U13427 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15464) );
  INV_X1 U13428 ( .A(n15464), .ZN(n10828) );
  OAI22_X1 U13429 ( .A1(n13035), .A2(n10826), .B1(n15712), .B2(n13040), .ZN(
        n10827) );
  AOI211_X1 U13430 ( .C1(n15430), .C2(n15597), .A(n10828), .B(n10827), .ZN(
        n10829) );
  OAI211_X1 U13431 ( .C1(n11004), .C2(n11233), .A(n10830), .B(n10829), .ZN(
        P3_U3179) );
  INV_X1 U13432 ( .A(n12154), .ZN(n12147) );
  NAND2_X1 U13433 ( .A1(n12147), .A2(P3_U3897), .ZN(n10831) );
  OAI21_X1 U13434 ( .B1(P3_U3897), .B2(n10832), .A(n10831), .ZN(P3_U3521) );
  XNOR2_X1 U13435 ( .A(n10833), .B(n12624), .ZN(n15391) );
  INV_X1 U13436 ( .A(n15391), .ZN(n10847) );
  OAI21_X1 U13437 ( .B1(n12624), .B2(n10835), .A(n10834), .ZN(n10836) );
  NAND2_X1 U13438 ( .A1(n10836), .A2(n15293), .ZN(n10838) );
  AOI22_X1 U13439 ( .A1(n13991), .A2(n13695), .B1(n13988), .B2(n13693), .ZN(
        n10837) );
  NAND2_X1 U13440 ( .A1(n10838), .A2(n10837), .ZN(n15397) );
  INV_X1 U13441 ( .A(n15393), .ZN(n10844) );
  NAND2_X1 U13442 ( .A1(n15393), .A2(n10839), .ZN(n10840) );
  NAND2_X1 U13443 ( .A1(n10840), .A2(n11160), .ZN(n10841) );
  NOR2_X1 U13444 ( .A1(n11036), .A2(n10841), .ZN(n15395) );
  NAND2_X1 U13445 ( .A1(n15395), .A2(n15285), .ZN(n10843) );
  AOI22_X1 U13446 ( .A1(n15305), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11326), 
        .B2(n15283), .ZN(n10842) );
  OAI211_X1 U13447 ( .C1(n10844), .C2(n13998), .A(n10843), .B(n10842), .ZN(
        n10845) );
  AOI21_X1 U13448 ( .B1(n15397), .B2(n15303), .A(n10845), .ZN(n10846) );
  OAI21_X1 U13449 ( .B1(n14004), .B2(n10847), .A(n10846), .ZN(P2_U3255) );
  XNOR2_X1 U13450 ( .A(n10848), .B(n12616), .ZN(n15374) );
  XNOR2_X1 U13451 ( .A(n10849), .B(n12616), .ZN(n10851) );
  AOI21_X1 U13452 ( .B1(n10851), .B2(n15293), .A(n10850), .ZN(n15381) );
  MUX2_X1 U13453 ( .A(n9843), .B(n15381), .S(n15303), .Z(n10861) );
  NAND2_X1 U13454 ( .A1(n10852), .A2(n15377), .ZN(n10853) );
  NAND2_X1 U13455 ( .A1(n10853), .A2(n11160), .ZN(n10854) );
  NOR2_X1 U13456 ( .A1(n10855), .A2(n10854), .ZN(n15379) );
  INV_X1 U13457 ( .A(n10856), .ZN(n10857) );
  OAI22_X1 U13458 ( .A1(n13998), .A2(n10858), .B1(n15298), .B2(n10857), .ZN(
        n10859) );
  AOI21_X1 U13459 ( .B1(n15285), .B2(n15379), .A(n10859), .ZN(n10860) );
  OAI211_X1 U13460 ( .C1(n14004), .C2(n15374), .A(n10861), .B(n10860), .ZN(
        P2_U3260) );
  XNOR2_X1 U13461 ( .A(n10867), .B(n10862), .ZN(n15358) );
  INV_X1 U13462 ( .A(n10863), .ZN(n10865) );
  AOI211_X1 U13463 ( .C1(n12387), .C2(n10865), .A(n13922), .B(n10864), .ZN(
        n15360) );
  OAI22_X1 U13464 ( .A1(n13998), .A2(n15363), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15298), .ZN(n10866) );
  AOI21_X1 U13465 ( .B1(n15285), .B2(n15360), .A(n10866), .ZN(n10873) );
  XNOR2_X1 U13466 ( .A(n10868), .B(n10867), .ZN(n10871) );
  INV_X1 U13467 ( .A(n10869), .ZN(n10870) );
  AOI21_X1 U13468 ( .B1(n10871), .B2(n15293), .A(n10870), .ZN(n15362) );
  MUX2_X1 U13469 ( .A(n9842), .B(n15362), .S(n15303), .Z(n10872) );
  OAI211_X1 U13470 ( .C1(n14004), .C2(n15358), .A(n10873), .B(n10872), .ZN(
        P2_U3262) );
  INV_X1 U13471 ( .A(n10882), .ZN(n10875) );
  NAND2_X1 U13472 ( .A1(n10875), .A2(n10874), .ZN(n10876) );
  NAND2_X1 U13473 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  XNOR2_X1 U13474 ( .A(n12441), .B(n13505), .ZN(n11192) );
  NAND2_X1 U13475 ( .A1(n13922), .A2(n13695), .ZN(n11193) );
  XNOR2_X1 U13476 ( .A(n11192), .B(n11193), .ZN(n10883) );
  INV_X1 U13477 ( .A(n13549), .ZN(n13657) );
  AOI22_X1 U13478 ( .A1(n10879), .A2(n13649), .B1(n13659), .B2(n13697), .ZN(
        n10881) );
  OAI211_X1 U13479 ( .C1(n12454), .C2(n13657), .A(n10881), .B(n10880), .ZN(
        n10887) );
  INV_X1 U13480 ( .A(n10877), .ZN(n10885) );
  AOI22_X1 U13481 ( .A1(n13641), .A2(n13697), .B1(n13676), .B2(n10882), .ZN(
        n10884) );
  NOR3_X1 U13482 ( .A1(n10885), .A2(n10884), .A3(n10883), .ZN(n10886) );
  AOI211_X1 U13483 ( .C1(n12441), .C2(n13668), .A(n10887), .B(n10886), .ZN(
        n10888) );
  OAI21_X1 U13484 ( .B1(n11196), .B2(n13653), .A(n10888), .ZN(P2_U3203) );
  INV_X1 U13485 ( .A(n10889), .ZN(n10892) );
  AOI211_X1 U13486 ( .C1(n10892), .C2(n15399), .A(n10891), .B(n10890), .ZN(
        n10897) );
  AOI22_X1 U13487 ( .A1(n14059), .A2(n12441), .B1(n15424), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10893) );
  OAI21_X1 U13488 ( .B1(n10897), .B2(n15424), .A(n10893), .ZN(P2_U3508) );
  INV_X1 U13489 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10894) );
  NOR2_X1 U13490 ( .A1(n15409), .A2(n10894), .ZN(n10895) );
  AOI21_X1 U13491 ( .B1(n8335), .B2(n12441), .A(n10895), .ZN(n10896) );
  OAI21_X1 U13492 ( .B1(n10897), .B2(n15407), .A(n10896), .ZN(P2_U3457) );
  NAND2_X1 U13493 ( .A1(n10898), .A2(n11946), .ZN(n10899) );
  XNOR2_X1 U13494 ( .A(n15084), .B(n14314), .ZN(n11861) );
  INV_X1 U13495 ( .A(n11861), .ZN(n11135) );
  OR2_X1 U13496 ( .A1(n15084), .A2(n14314), .ZN(n10900) );
  NAND2_X1 U13497 ( .A1(n10901), .A2(n10900), .ZN(n15044) );
  XNOR2_X1 U13498 ( .A(n15053), .B(n14313), .ZN(n11860) );
  INV_X1 U13499 ( .A(n11860), .ZN(n15045) );
  NAND2_X1 U13500 ( .A1(n15044), .A2(n15045), .ZN(n10903) );
  OR2_X1 U13501 ( .A1(n15053), .A2(n14313), .ZN(n10902) );
  NAND2_X1 U13502 ( .A1(n10903), .A2(n10902), .ZN(n11094) );
  NAND2_X1 U13503 ( .A1(n10904), .A2(n11892), .ZN(n10907) );
  AOI22_X1 U13504 ( .A1(n11853), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11852), 
        .B2(n10905), .ZN(n10906) );
  XNOR2_X1 U13505 ( .A(n11963), .B(n14312), .ZN(n11863) );
  INV_X1 U13506 ( .A(n11863), .ZN(n11099) );
  OR2_X1 U13507 ( .A1(n11963), .A2(n14312), .ZN(n10908) );
  NAND2_X1 U13508 ( .A1(n10909), .A2(n11892), .ZN(n10912) );
  AOI22_X1 U13509 ( .A1(n11853), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11852), 
        .B2(n10910), .ZN(n10911) );
  NAND2_X1 U13510 ( .A1(n11884), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10918) );
  OR2_X1 U13511 ( .A1(n10273), .A2(n9615), .ZN(n10917) );
  OR2_X1 U13512 ( .A1(n11902), .A2(n15144), .ZN(n10916) );
  NAND2_X1 U13513 ( .A1(n10913), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10924) );
  OR2_X1 U13514 ( .A1(n10913), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U13515 ( .A1(n10924), .A2(n10914), .ZN(n11322) );
  OR2_X1 U13516 ( .A1(n11900), .A2(n11322), .ZN(n10915) );
  NAND4_X1 U13517 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n14311) );
  INV_X1 U13518 ( .A(n14311), .ZN(n10974) );
  XNOR2_X1 U13519 ( .A(n15107), .B(n10974), .ZN(n11865) );
  OR2_X1 U13520 ( .A1(n10919), .A2(n11817), .ZN(n10922) );
  AOI22_X1 U13521 ( .A1(n11853), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10920), 
        .B2(n11852), .ZN(n10921) );
  NAND2_X1 U13522 ( .A1(n6675), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10930) );
  OR2_X1 U13523 ( .A1(n11902), .A2(n15146), .ZN(n10929) );
  INV_X1 U13524 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13525 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  NAND2_X1 U13526 ( .A1(n10939), .A2(n10925), .ZN(n11497) );
  OR2_X1 U13527 ( .A1(n11900), .A2(n11497), .ZN(n10928) );
  INV_X1 U13528 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10926) );
  OR2_X1 U13529 ( .A1(n6689), .A2(n10926), .ZN(n10927) );
  NAND4_X1 U13530 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n14310) );
  XNOR2_X1 U13531 ( .A(n15115), .B(n11492), .ZN(n11867) );
  NAND2_X1 U13532 ( .A1(n11015), .A2(n11867), .ZN(n10932) );
  OR2_X1 U13533 ( .A1(n15115), .A2(n14310), .ZN(n10931) );
  NAND2_X1 U13534 ( .A1(n10933), .A2(n11892), .ZN(n10936) );
  AOI22_X1 U13535 ( .A1(n10934), .A2(n11852), .B1(n11853), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U13536 ( .A1(n11807), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10945) );
  OR2_X1 U13537 ( .A1(n10273), .A2(n10937), .ZN(n10944) );
  NAND2_X1 U13538 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  NAND2_X1 U13539 ( .A1(n10953), .A2(n10940), .ZN(n11576) );
  OR2_X1 U13540 ( .A1(n11900), .A2(n11576), .ZN(n10943) );
  INV_X1 U13541 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10941) );
  OR2_X1 U13542 ( .A1(n6689), .A2(n10941), .ZN(n10942) );
  NAND4_X1 U13543 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n14309) );
  INV_X1 U13544 ( .A(n14309), .ZN(n11573) );
  OR2_X1 U13545 ( .A1(n11984), .A2(n11573), .ZN(n10976) );
  NAND2_X1 U13546 ( .A1(n11984), .A2(n11573), .ZN(n10946) );
  NAND2_X1 U13547 ( .A1(n10976), .A2(n10946), .ZN(n11866) );
  OR2_X1 U13548 ( .A1(n11984), .A2(n14309), .ZN(n10947) );
  NAND2_X1 U13549 ( .A1(n10948), .A2(n11892), .ZN(n10951) );
  AOI22_X1 U13550 ( .A1(n10949), .A2(n11852), .B1(n11853), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U13551 ( .A1(n6674), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10960) );
  AND2_X1 U13552 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  OR2_X1 U13553 ( .A1(n10954), .A2(n10978), .ZN(n14957) );
  OR2_X1 U13554 ( .A1(n11900), .A2(n14957), .ZN(n10959) );
  INV_X1 U13555 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10955) );
  OR2_X1 U13556 ( .A1(n6689), .A2(n10955), .ZN(n10958) );
  OR2_X1 U13557 ( .A1(n11902), .A2(n10956), .ZN(n10957) );
  NAND4_X1 U13558 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n14308) );
  XNOR2_X1 U13559 ( .A(n14986), .B(n14308), .ZN(n11869) );
  INV_X1 U13560 ( .A(n11869), .ZN(n11268) );
  XNOR2_X1 U13561 ( .A(n11269), .B(n11268), .ZN(n14985) );
  INV_X1 U13562 ( .A(n14985), .ZN(n10995) );
  NAND2_X1 U13563 ( .A1(n11947), .A2(n14315), .ZN(n10961) );
  NAND2_X1 U13564 ( .A1(n10962), .A2(n10961), .ZN(n10964) );
  OR2_X1 U13565 ( .A1(n11947), .A2(n14315), .ZN(n10963) );
  INV_X1 U13566 ( .A(n14314), .ZN(n10966) );
  OR2_X1 U13567 ( .A1(n15084), .A2(n10966), .ZN(n10965) );
  NAND2_X1 U13568 ( .A1(n11144), .A2(n10965), .ZN(n10968) );
  NAND2_X1 U13569 ( .A1(n15084), .A2(n10966), .ZN(n10967) );
  AND2_X1 U13570 ( .A1(n15053), .A2(n10970), .ZN(n10969) );
  OR2_X1 U13571 ( .A1(n15053), .A2(n10970), .ZN(n10971) );
  INV_X1 U13572 ( .A(n14312), .ZN(n11260) );
  NOR2_X1 U13573 ( .A1(n11963), .A2(n11260), .ZN(n10973) );
  NAND2_X1 U13574 ( .A1(n11963), .A2(n11260), .ZN(n10972) );
  NAND2_X1 U13575 ( .A1(n15115), .A2(n11492), .ZN(n10975) );
  INV_X1 U13576 ( .A(n11866), .ZN(n11357) );
  OAI211_X1 U13577 ( .C1(n10977), .C2(n11869), .A(n11290), .B(n14792), .ZN(
        n10988) );
  NAND2_X1 U13578 ( .A1(n14309), .A2(n14563), .ZN(n10986) );
  NAND2_X1 U13579 ( .A1(n6675), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10984) );
  OR2_X1 U13580 ( .A1(n11902), .A2(n14812), .ZN(n10983) );
  NAND2_X1 U13581 ( .A1(n10978), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11282) );
  OR2_X1 U13582 ( .A1(n10978), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10979) );
  NAND2_X1 U13583 ( .A1(n11282), .A2(n10979), .ZN(n14799) );
  OR2_X1 U13584 ( .A1(n11900), .A2(n14799), .ZN(n10982) );
  INV_X1 U13585 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10980) );
  OR2_X1 U13586 ( .A1(n6689), .A2(n10980), .ZN(n10981) );
  NAND4_X1 U13587 ( .A1(n10984), .A2(n10983), .A3(n10982), .A4(n10981), .ZN(
        n14307) );
  NAND2_X1 U13588 ( .A1(n14307), .A2(n14565), .ZN(n10985) );
  NAND2_X1 U13589 ( .A1(n10986), .A2(n10985), .ZN(n14954) );
  INV_X1 U13590 ( .A(n14954), .ZN(n10987) );
  NAND2_X1 U13591 ( .A1(n10988), .A2(n10987), .ZN(n14991) );
  INV_X1 U13592 ( .A(n11984), .ZN(n15127) );
  INV_X1 U13593 ( .A(n15115), .ZN(n11485) );
  INV_X1 U13594 ( .A(n15053), .ZN(n15092) );
  AOI21_X1 U13595 ( .B1(n11352), .B2(n14986), .A(n14630), .ZN(n10989) );
  NAND2_X1 U13596 ( .A1(n10989), .A2(n14802), .ZN(n14987) );
  OAI22_X1 U13597 ( .A1(n14636), .A2(n10990), .B1(n14957), .B2(n14633), .ZN(
        n10991) );
  AOI21_X1 U13598 ( .B1(n14986), .B2(n15052), .A(n10991), .ZN(n10992) );
  OAI21_X1 U13599 ( .B1(n14987), .B2(n14654), .A(n10992), .ZN(n10993) );
  AOI21_X1 U13600 ( .B1(n14991), .B2(n14636), .A(n10993), .ZN(n10994) );
  OAI21_X1 U13601 ( .B1(n15067), .B2(n10995), .A(n10994), .ZN(P1_U3282) );
  NAND2_X1 U13602 ( .A1(n10996), .A2(n12326), .ZN(n10997) );
  NAND3_X1 U13603 ( .A1(n10998), .A2(n15671), .A3(n10997), .ZN(n11000) );
  AOI22_X1 U13604 ( .A1(n15597), .A2(n15654), .B1(n15653), .B2(n12199), .ZN(
        n10999) );
  NAND2_X1 U13605 ( .A1(n11000), .A2(n10999), .ZN(n15713) );
  MUX2_X1 U13606 ( .A(n15713), .B(P3_REG2_REG_6__SCAN_IN), .S(n15649), .Z(
        n11001) );
  INV_X1 U13607 ( .A(n11001), .ZN(n11007) );
  XNOR2_X1 U13608 ( .A(n11002), .B(n12326), .ZN(n15715) );
  INV_X1 U13609 ( .A(n15662), .ZN(n15645) );
  NAND2_X1 U13610 ( .A1(n15682), .A2(n15645), .ZN(n11003) );
  OAI22_X1 U13611 ( .A1(n13320), .A2(n15712), .B1(n11004), .B2(n15676), .ZN(
        n11005) );
  AOI21_X1 U13612 ( .B1(n15715), .B2(n15631), .A(n11005), .ZN(n11006) );
  NAND2_X1 U13613 ( .A1(n11007), .A2(n11006), .ZN(P3_U3227) );
  INV_X1 U13614 ( .A(n11008), .ZN(n11011) );
  INV_X1 U13615 ( .A(n11867), .ZN(n11010) );
  OAI21_X1 U13616 ( .B1(n11011), .B2(n11010), .A(n11009), .ZN(n11014) );
  NAND2_X1 U13617 ( .A1(n14311), .A2(n14563), .ZN(n11013) );
  NAND2_X1 U13618 ( .A1(n14309), .A2(n14565), .ZN(n11012) );
  NAND2_X1 U13619 ( .A1(n11013), .A2(n11012), .ZN(n11495) );
  AOI21_X1 U13620 ( .B1(n11014), .B2(n14792), .A(n11495), .ZN(n15118) );
  XOR2_X1 U13621 ( .A(n11015), .B(n11867), .Z(n15120) );
  INV_X1 U13622 ( .A(n15120), .ZN(n15122) );
  OR2_X1 U13623 ( .A1(n11016), .A2(n11166), .ZN(n11916) );
  INV_X1 U13624 ( .A(n11916), .ZN(n11017) );
  NAND2_X1 U13625 ( .A1(n14636), .A2(n11017), .ZN(n11705) );
  OAI21_X1 U13626 ( .B1(n15074), .B2(n11018), .A(n11705), .ZN(n14641) );
  NAND2_X1 U13627 ( .A1(n15122), .A2(n14641), .ZN(n11023) );
  OAI21_X1 U13628 ( .B1(n11485), .B2(n11258), .A(n15055), .ZN(n11019) );
  NOR2_X1 U13629 ( .A1(n11019), .A2(n11350), .ZN(n15114) );
  NOR2_X1 U13630 ( .A1(n11485), .A2(n14614), .ZN(n11021) );
  OAI22_X1 U13631 ( .A1(n14636), .A2(n9665), .B1(n11497), .B2(n14633), .ZN(
        n11020) );
  AOI211_X1 U13632 ( .C1(n15114), .C2(n15058), .A(n11021), .B(n11020), .ZN(
        n11022) );
  OAI211_X1 U13633 ( .C1(n15074), .C2(n15118), .A(n11023), .B(n11022), .ZN(
        P1_U3284) );
  INV_X1 U13634 ( .A(n13750), .ZN(n13744) );
  INV_X1 U13635 ( .A(n11840), .ZN(n11027) );
  OAI222_X1 U13636 ( .A1(P2_U3088), .A2(n13744), .B1(n14150), .B2(n11027), 
        .C1(n11024), .C2(n14152), .ZN(P2_U3309) );
  NAND2_X1 U13637 ( .A1(n11025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11026) );
  XNOR2_X1 U13638 ( .A(n11026), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14380) );
  INV_X1 U13639 ( .A(n14380), .ZN(n15037) );
  OAI222_X1 U13640 ( .A1(n14764), .A2(n11028), .B1(n14768), .B2(n11027), .C1(
        n15037), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI21_X1 U13641 ( .B1(n11030), .B2(n12625), .A(n11029), .ZN(n11031) );
  NAND2_X1 U13642 ( .A1(n11031), .A2(n15293), .ZN(n11035) );
  XNOR2_X1 U13643 ( .A(n11032), .B(n12625), .ZN(n15400) );
  NAND2_X1 U13644 ( .A1(n15400), .A2(n15376), .ZN(n11034) );
  AOI22_X1 U13645 ( .A1(n13991), .A2(n13694), .B1(n13988), .B2(n13692), .ZN(
        n11033) );
  NAND3_X1 U13646 ( .A1(n11035), .A2(n11034), .A3(n11033), .ZN(n15406) );
  INV_X1 U13647 ( .A(n15406), .ZN(n11042) );
  OAI211_X1 U13648 ( .C1(n15404), .C2(n11036), .A(n11160), .B(n11158), .ZN(
        n15401) );
  AOI22_X1 U13649 ( .A1(n15305), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11207), 
        .B2(n15283), .ZN(n11038) );
  NAND2_X1 U13650 ( .A1(n12459), .A2(n15281), .ZN(n11037) );
  OAI211_X1 U13651 ( .C1(n15401), .C2(n13907), .A(n11038), .B(n11037), .ZN(
        n11039) );
  AOI21_X1 U13652 ( .B1(n15400), .B2(n11040), .A(n11039), .ZN(n11041) );
  OAI21_X1 U13653 ( .B1(n11042), .B2(n15305), .A(n11041), .ZN(P2_U3254) );
  XNOR2_X1 U13654 ( .A(n11043), .B(n12327), .ZN(n11046) );
  INV_X1 U13655 ( .A(n11046), .ZN(n15720) );
  XNOR2_X1 U13656 ( .A(n11044), .B(n12207), .ZN(n11048) );
  OAI22_X1 U13657 ( .A1(n12217), .A2(n15673), .B1(n15611), .B2(n15637), .ZN(
        n11045) );
  AOI21_X1 U13658 ( .B1(n11046), .B2(n15645), .A(n11045), .ZN(n11047) );
  OAI21_X1 U13659 ( .B1(n11048), .B2(n15641), .A(n11047), .ZN(n15722) );
  NAND2_X1 U13660 ( .A1(n15722), .A2(n15682), .ZN(n11053) );
  INV_X1 U13661 ( .A(n13320), .ZN(n13246) );
  INV_X1 U13662 ( .A(n11049), .ZN(n11117) );
  OAI22_X1 U13663 ( .A1(n15682), .A2(n15474), .B1(n11117), .B2(n15676), .ZN(
        n11050) );
  AOI21_X1 U13664 ( .B1(n13246), .B2(n11051), .A(n11050), .ZN(n11052) );
  OAI211_X1 U13665 ( .C1(n15720), .C2(n11453), .A(n11053), .B(n11052), .ZN(
        P3_U3226) );
  INV_X1 U13666 ( .A(n11054), .ZN(n11057) );
  INV_X1 U13667 ( .A(n11055), .ZN(n11056) );
  NAND2_X1 U13668 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  NOR2_X1 U13669 ( .A1(n11260), .A2(n12826), .ZN(n11060) );
  AOI21_X1 U13670 ( .B1(n11963), .B2(n7074), .A(n11060), .ZN(n11312) );
  AOI22_X1 U13671 ( .A1(n11963), .A2(n12804), .B1(n11309), .B2(n14312), .ZN(
        n11061) );
  XNOR2_X1 U13672 ( .A(n11061), .B(n12824), .ZN(n11311) );
  XOR2_X1 U13673 ( .A(n11312), .B(n11311), .Z(n11062) );
  OAI211_X1 U13674 ( .C1(n11063), .C2(n11062), .A(n11316), .B(n14951), .ZN(
        n11070) );
  NAND2_X1 U13675 ( .A1(n14313), .A2(n14563), .ZN(n11065) );
  NAND2_X1 U13676 ( .A1(n14311), .A2(n14565), .ZN(n11064) );
  NAND2_X1 U13677 ( .A1(n11065), .A2(n11064), .ZN(n11102) );
  INV_X1 U13678 ( .A(n11066), .ZN(n11068) );
  NOR2_X1 U13679 ( .A1(n14958), .A2(n11096), .ZN(n11067) );
  AOI211_X1 U13680 ( .C1(n14953), .C2(n11102), .A(n11068), .B(n11067), .ZN(
        n11069) );
  OAI211_X1 U13681 ( .C1(n7176), .C2(n14300), .A(n11070), .B(n11069), .ZN(
        P1_U3213) );
  INV_X1 U13682 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11077) );
  NOR2_X1 U13683 ( .A1(n11086), .A2(n11077), .ZN(n11071) );
  AOI21_X1 U13684 ( .B1(n11077), .B2(n11086), .A(n11071), .ZN(n15239) );
  INV_X1 U13685 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U13686 ( .A1(n11073), .A2(n11072), .ZN(n15218) );
  OR2_X1 U13687 ( .A1(n15226), .A2(n11076), .ZN(n11075) );
  NAND2_X1 U13688 ( .A1(n15226), .A2(n11076), .ZN(n11074) );
  AND2_X1 U13689 ( .A1(n11075), .A2(n11074), .ZN(n15219) );
  AOI21_X1 U13690 ( .B1(n15220), .B2(n15218), .A(n15219), .ZN(n15217) );
  AOI21_X1 U13691 ( .B1(n11076), .B2(n11084), .A(n15217), .ZN(n15240) );
  OAI21_X1 U13692 ( .B1(n11077), .B2(n11086), .A(n15238), .ZN(n13722) );
  OAI211_X1 U13693 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n11078), .A(n15274), 
        .B(n13724), .ZN(n11093) );
  NAND2_X1 U13694 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11585)
         );
  NOR2_X1 U13695 ( .A1(n13723), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11079) );
  AOI21_X1 U13696 ( .B1(n13723), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11079), 
        .ZN(n11089) );
  INV_X1 U13697 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11087) );
  INV_X1 U13698 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15211) );
  AOI21_X1 U13699 ( .B1(n11081), .B2(P2_REG1_REG_11__SCAN_IN), .A(n11080), 
        .ZN(n15210) );
  OR2_X1 U13700 ( .A1(n11084), .A2(n15211), .ZN(n11082) );
  OAI211_X1 U13701 ( .C1(P2_REG1_REG_12__SCAN_IN), .C2(n15226), .A(n15210), 
        .B(n11082), .ZN(n15216) );
  INV_X1 U13702 ( .A(n15216), .ZN(n11083) );
  AOI21_X1 U13703 ( .B1(n15211), .B2(n11084), .A(n11083), .ZN(n15237) );
  NOR2_X1 U13704 ( .A1(n15234), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11085) );
  AOI21_X1 U13705 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n15234), .A(n11085), 
        .ZN(n15236) );
  NAND2_X1 U13706 ( .A1(n15237), .A2(n15236), .ZN(n15235) );
  OAI21_X1 U13707 ( .B1(n11087), .B2(n11086), .A(n15235), .ZN(n11088) );
  NAND2_X1 U13708 ( .A1(n11089), .A2(n11088), .ZN(n13732) );
  OAI211_X1 U13709 ( .C1(n11089), .C2(n11088), .A(n13732), .B(n15270), .ZN(
        n11090) );
  NAND2_X1 U13710 ( .A1(n11585), .A2(n11090), .ZN(n11091) );
  AOI21_X1 U13711 ( .B1(n15266), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n11091), 
        .ZN(n11092) );
  OAI211_X1 U13712 ( .C1(n15265), .C2(n13733), .A(n11093), .B(n11092), .ZN(
        P2_U3228) );
  XNOR2_X1 U13713 ( .A(n11094), .B(n11099), .ZN(n15098) );
  NAND2_X1 U13714 ( .A1(n15054), .A2(n11963), .ZN(n11095) );
  NAND3_X1 U13715 ( .A1(n11259), .A2(n15055), .A3(n11095), .ZN(n15099) );
  INV_X1 U13716 ( .A(n11096), .ZN(n11097) );
  AOI22_X1 U13717 ( .A1(n11963), .A2(n15052), .B1(n11097), .B2(n15070), .ZN(
        n11098) );
  OAI21_X1 U13718 ( .B1(n15099), .B2(n14654), .A(n11098), .ZN(n11106) );
  XNOR2_X1 U13719 ( .A(n11100), .B(n11099), .ZN(n11101) );
  NAND2_X1 U13720 ( .A1(n11101), .A2(n14792), .ZN(n11104) );
  INV_X1 U13721 ( .A(n11102), .ZN(n11103) );
  NAND2_X1 U13722 ( .A1(n11104), .A2(n11103), .ZN(n15101) );
  MUX2_X1 U13723 ( .A(n15101), .B(P1_REG2_REG_7__SCAN_IN), .S(n15074), .Z(
        n11105) );
  AOI211_X1 U13724 ( .C1(n15098), .C2(n14641), .A(n11106), .B(n11105), .ZN(
        n11107) );
  INV_X1 U13725 ( .A(n11107), .ZN(P1_U3286) );
  NAND2_X1 U13726 ( .A1(n11109), .A2(n11108), .ZN(n11110) );
  XNOR2_X1 U13727 ( .A(n12207), .B(n12848), .ZN(n11222) );
  OAI211_X1 U13728 ( .C1(n11112), .C2(n11222), .A(n11225), .B(n15432), .ZN(
        n11116) );
  NAND2_X1 U13729 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n15479) );
  INV_X1 U13730 ( .A(n15479), .ZN(n11114) );
  OAI22_X1 U13731 ( .A1(n13035), .A2(n15611), .B1(n15717), .B2(n13040), .ZN(
        n11113) );
  AOI211_X1 U13732 ( .C1(n15430), .C2(n12216), .A(n11114), .B(n11113), .ZN(
        n11115) );
  OAI211_X1 U13733 ( .C1(n11117), .C2(n11233), .A(n11116), .B(n11115), .ZN(
        P3_U3153) );
  INV_X1 U13734 ( .A(n14641), .ZN(n14544) );
  OAI22_X1 U13735 ( .A1(n14614), .A2(n7180), .B1(n14633), .B2(n11118), .ZN(
        n11119) );
  AOI21_X1 U13736 ( .B1(n15058), .B2(n11120), .A(n11119), .ZN(n11124) );
  MUX2_X1 U13737 ( .A(n11122), .B(n11121), .S(n14636), .Z(n11123) );
  OAI211_X1 U13738 ( .C1(n14544), .C2(n11125), .A(n11124), .B(n11123), .ZN(
        P1_U3291) );
  MUX2_X1 U13739 ( .A(n11127), .B(n11126), .S(n14636), .Z(n11133) );
  OAI22_X1 U13740 ( .A1(n14614), .A2(n11129), .B1(n14633), .B2(n11128), .ZN(
        n11130) );
  AOI21_X1 U13741 ( .B1(n15058), .B2(n11131), .A(n11130), .ZN(n11132) );
  OAI211_X1 U13742 ( .C1(n14544), .C2(n11134), .A(n11133), .B(n11132), .ZN(
        P1_U3292) );
  XNOR2_X1 U13743 ( .A(n11136), .B(n11135), .ZN(n15090) );
  INV_X1 U13744 ( .A(n15090), .ZN(n11150) );
  NAND2_X1 U13745 ( .A1(n15084), .A2(n11137), .ZN(n11138) );
  NAND3_X1 U13746 ( .A1(n11139), .A2(n15055), .A3(n11138), .ZN(n15086) );
  INV_X1 U13747 ( .A(n15086), .ZN(n11143) );
  INV_X1 U13748 ( .A(n15084), .ZN(n11141) );
  OAI22_X1 U13749 ( .A1(n14614), .A2(n11141), .B1(n14633), .B2(n11140), .ZN(
        n11142) );
  AOI21_X1 U13750 ( .B1(n15058), .B2(n11143), .A(n11142), .ZN(n11149) );
  XNOR2_X1 U13751 ( .A(n11144), .B(n11861), .ZN(n11146) );
  AOI21_X1 U13752 ( .B1(n11146), .B2(n14792), .A(n11145), .ZN(n15087) );
  MUX2_X1 U13753 ( .A(n11147), .B(n15087), .S(n14636), .Z(n11148) );
  OAI211_X1 U13754 ( .C1(n11150), .C2(n14544), .A(n11149), .B(n11148), .ZN(
        P1_U3288) );
  XNOR2_X1 U13755 ( .A(n14912), .B(n11151), .ZN(n12628) );
  INV_X1 U13756 ( .A(n12628), .ZN(n11152) );
  XNOR2_X1 U13757 ( .A(n11153), .B(n11152), .ZN(n11154) );
  NAND2_X1 U13758 ( .A1(n11154), .A2(n15293), .ZN(n11156) );
  AOI22_X1 U13759 ( .A1(n13991), .A2(n13693), .B1(n13988), .B2(n13691), .ZN(
        n11155) );
  AND2_X1 U13760 ( .A1(n11156), .A2(n11155), .ZN(n14918) );
  XNOR2_X1 U13761 ( .A(n11157), .B(n12628), .ZN(n14916) );
  NAND2_X1 U13762 ( .A1(n11158), .A2(n14912), .ZN(n11159) );
  NAND3_X1 U13763 ( .A1(n11241), .A2(n11160), .A3(n11159), .ZN(n14914) );
  AOI22_X1 U13764 ( .A1(n15305), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11339), 
        .B2(n15283), .ZN(n11162) );
  NAND2_X1 U13765 ( .A1(n14912), .A2(n15281), .ZN(n11161) );
  OAI211_X1 U13766 ( .C1(n14914), .C2(n13907), .A(n11162), .B(n11161), .ZN(
        n11163) );
  AOI21_X1 U13767 ( .B1(n14916), .B2(n15287), .A(n11163), .ZN(n11164) );
  OAI21_X1 U13768 ( .B1(n14918), .B2(n15305), .A(n11164), .ZN(P2_U3253) );
  INV_X1 U13769 ( .A(n11831), .ZN(n11167) );
  OAI222_X1 U13770 ( .A1(n14152), .A2(n11165), .B1(n14150), .B2(n11167), .C1(
        P2_U3088), .C2(n13759), .ZN(P2_U3308) );
  OAI222_X1 U13771 ( .A1(n14764), .A2(n11168), .B1(n14768), .B2(n11167), .C1(
        n11166), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U13772 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14943)
         );
  INV_X1 U13773 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14978) );
  MUX2_X1 U13774 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14978), .S(n14361), .Z(
        n14357) );
  NAND2_X1 U13775 ( .A1(n14356), .A2(n14357), .ZN(n14355) );
  OAI21_X1 U13776 ( .B1(n14361), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14355), 
        .ZN(n11170) );
  XNOR2_X1 U13777 ( .A(n11170), .B(n15024), .ZN(n15019) );
  NOR2_X1 U13778 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15019), .ZN(n15018) );
  INV_X1 U13779 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U13780 ( .A1(n11372), .A2(n11172), .ZN(n11171) );
  OAI21_X1 U13781 ( .B1(n11372), .B2(n11172), .A(n11171), .ZN(n11173) );
  INV_X1 U13782 ( .A(n11173), .ZN(n11174) );
  OAI211_X1 U13783 ( .C1(n11175), .C2(n11174), .A(n11364), .B(n14383), .ZN(
        n11176) );
  AND2_X1 U13784 ( .A1(n14943), .A2(n11176), .ZN(n11190) );
  INV_X1 U13785 ( .A(n11372), .ZN(n11597) );
  INV_X1 U13786 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14362) );
  NOR2_X1 U13787 ( .A1(n11178), .A2(n11177), .ZN(n14363) );
  MUX2_X1 U13788 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14362), .S(n14361), .Z(
        n11179) );
  OAI21_X1 U13789 ( .B1(n14368), .B2(n14363), .A(n11179), .ZN(n14366) );
  OAI21_X1 U13790 ( .B1(n14362), .B2(n11180), .A(n14366), .ZN(n11181) );
  NOR2_X1 U13791 ( .A1(n11181), .A2(n11455), .ZN(n11183) );
  AOI21_X1 U13792 ( .B1(n11455), .B2(n11181), .A(n11183), .ZN(n11182) );
  INV_X1 U13793 ( .A(n11182), .ZN(n15021) );
  NOR2_X1 U13794 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15021), .ZN(n15020) );
  NOR2_X1 U13795 ( .A1(n11183), .A2(n15020), .ZN(n11186) );
  OAI21_X1 U13796 ( .B1(n11597), .B2(P1_REG2_REG_16__SCAN_IN), .A(n11186), 
        .ZN(n11184) );
  AOI21_X1 U13797 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n11597), .A(n11184), 
        .ZN(n11370) );
  NOR2_X1 U13798 ( .A1(n11372), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11185) );
  AOI211_X1 U13799 ( .C1(n11372), .C2(P1_REG2_REG_16__SCAN_IN), .A(n11186), 
        .B(n11185), .ZN(n11187) );
  NOR3_X1 U13800 ( .A1(n15034), .A2(n11370), .A3(n11187), .ZN(n11188) );
  AOI21_X1 U13801 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14343), .A(n11188), 
        .ZN(n11189) );
  OAI211_X1 U13802 ( .C1(n15038), .C2(n11372), .A(n11190), .B(n11189), .ZN(
        P1_U3259) );
  OAI222_X1 U13803 ( .A1(n14152), .A2(n11191), .B1(n14150), .B2(n11818), .C1(
        n12659), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13804 ( .A1(n14771), .A2(n11819), .B1(P1_U3086), .B2(n11912), 
        .C1(n14768), .C2(n11818), .ZN(P1_U3334) );
  INV_X1 U13805 ( .A(n11192), .ZN(n11194) );
  NAND2_X1 U13806 ( .A1(n11194), .A2(n11193), .ZN(n11195) );
  XNOR2_X1 U13807 ( .A(n15393), .B(n13493), .ZN(n11204) );
  AND2_X1 U13808 ( .A1(n13509), .A2(n13694), .ZN(n11197) );
  NAND2_X1 U13809 ( .A1(n11204), .A2(n11197), .ZN(n11202) );
  INV_X1 U13810 ( .A(n11204), .ZN(n11199) );
  INV_X1 U13811 ( .A(n11197), .ZN(n11198) );
  NAND2_X1 U13812 ( .A1(n11199), .A2(n11198), .ZN(n11200) );
  NAND2_X1 U13813 ( .A1(n11202), .A2(n11200), .ZN(n11333) );
  INV_X1 U13814 ( .A(n11333), .ZN(n11201) );
  XNOR2_X1 U13815 ( .A(n12459), .B(n13505), .ZN(n11342) );
  NAND2_X1 U13816 ( .A1(n13922), .A2(n13693), .ZN(n11337) );
  XNOR2_X1 U13817 ( .A(n11342), .B(n11337), .ZN(n11206) );
  AND2_X1 U13818 ( .A1(n11206), .A2(n11202), .ZN(n11203) );
  NAND3_X1 U13819 ( .A1(n11204), .A2(n13641), .A3(n13694), .ZN(n11205) );
  OAI21_X1 U13820 ( .B1(n11330), .B2(n13653), .A(n11205), .ZN(n11214) );
  INV_X1 U13821 ( .A(n11206), .ZN(n11213) );
  AOI22_X1 U13822 ( .A1(n11207), .A2(n13649), .B1(n13659), .B2(n13694), .ZN(
        n11211) );
  NAND2_X1 U13823 ( .A1(n12459), .A2(n13668), .ZN(n11210) );
  NAND2_X1 U13824 ( .A1(n13549), .A2(n13692), .ZN(n11208) );
  NAND4_X1 U13825 ( .A1(n11211), .A2(n11210), .A3(n11209), .A4(n11208), .ZN(
        n11212) );
  AOI21_X1 U13826 ( .B1(n11214), .B2(n11213), .A(n11212), .ZN(n11215) );
  OAI21_X1 U13827 ( .B1(n11341), .B2(n13653), .A(n11215), .ZN(P2_U3208) );
  INV_X1 U13828 ( .A(n11878), .ZN(n11217) );
  OAI222_X1 U13829 ( .A1(n14152), .A2(n6996), .B1(n14150), .B2(n11217), .C1(
        n11216), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI222_X1 U13830 ( .A1(n14764), .A2(n7478), .B1(P1_U3086), .B2(n12089), .C1(
        n14768), .C2(n11217), .ZN(P1_U3335) );
  INV_X1 U13831 ( .A(n11218), .ZN(n11220) );
  OAI222_X1 U13832 ( .A1(n11221), .A2(P3_U3151), .B1(n13468), .B2(n11220), 
        .C1(n11219), .C2(n11518), .ZN(P3_U3271) );
  INV_X1 U13833 ( .A(n15600), .ZN(n11234) );
  INV_X1 U13834 ( .A(n11222), .ZN(n11223) );
  NAND2_X1 U13835 ( .A1(n11223), .A2(n15597), .ZN(n11224) );
  XNOR2_X1 U13836 ( .A(n12218), .B(n12921), .ZN(n11427) );
  XNOR2_X1 U13837 ( .A(n11427), .B(n12216), .ZN(n11226) );
  OAI211_X1 U13838 ( .C1(n11227), .C2(n11226), .A(n11430), .B(n15432), .ZN(
        n11232) );
  NAND2_X1 U13839 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15497) );
  INV_X1 U13840 ( .A(n15497), .ZN(n11230) );
  INV_X1 U13841 ( .A(n12218), .ZN(n15603) );
  OAI22_X1 U13842 ( .A1(n13035), .A2(n11228), .B1(n15603), .B2(n13040), .ZN(
        n11229) );
  AOI211_X1 U13843 ( .C1(n15430), .C2(n15598), .A(n11230), .B(n11229), .ZN(
        n11231) );
  OAI211_X1 U13844 ( .C1(n11234), .C2(n11233), .A(n11232), .B(n11231), .ZN(
        P3_U3161) );
  NAND2_X1 U13845 ( .A1(n11236), .A2(n11235), .ZN(n12627) );
  XNOR2_X1 U13846 ( .A(n11237), .B(n12627), .ZN(n11238) );
  AOI22_X1 U13847 ( .A1(n13991), .A2(n13692), .B1(n13988), .B2(n13690), .ZN(
        n11512) );
  OAI21_X1 U13848 ( .B1(n11238), .B2(n13950), .A(n11512), .ZN(n11417) );
  INV_X1 U13849 ( .A(n11417), .ZN(n11246) );
  XOR2_X1 U13850 ( .A(n12627), .B(n11239), .Z(n11419) );
  INV_X1 U13851 ( .A(n11240), .ZN(n11411) );
  AOI211_X1 U13852 ( .C1(n12470), .C2(n11241), .A(n13922), .B(n11411), .ZN(
        n11418) );
  NAND2_X1 U13853 ( .A1(n11418), .A2(n15285), .ZN(n11243) );
  AOI22_X1 U13854 ( .A1(n15305), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11514), 
        .B2(n15283), .ZN(n11242) );
  OAI211_X1 U13855 ( .C1(n7204), .C2(n13998), .A(n11243), .B(n11242), .ZN(
        n11244) );
  AOI21_X1 U13856 ( .B1(n11419), .B2(n15287), .A(n11244), .ZN(n11245) );
  OAI21_X1 U13857 ( .B1(n11246), .B2(n15305), .A(n11245), .ZN(P2_U3252) );
  AOI21_X1 U13858 ( .B1(n11247), .B2(n12332), .A(n15641), .ZN(n11250) );
  OAI22_X1 U13859 ( .A1(n12217), .A2(n15637), .B1(n11658), .B2(n15673), .ZN(
        n11248) );
  AOI21_X1 U13860 ( .B1(n11250), .B2(n11249), .A(n11248), .ZN(n15729) );
  XNOR2_X1 U13861 ( .A(n11251), .B(n12332), .ZN(n15733) );
  NOR2_X1 U13862 ( .A1(n11252), .A2(n15718), .ZN(n15731) );
  AOI22_X1 U13863 ( .A1(n15731), .A2(n15679), .B1(n6668), .B2(n11437), .ZN(
        n11253) );
  OAI21_X1 U13864 ( .B1(n15505), .B2(n15682), .A(n11253), .ZN(n11254) );
  AOI21_X1 U13865 ( .B1(n15733), .B2(n15631), .A(n11254), .ZN(n11255) );
  OAI21_X1 U13866 ( .B1(n15729), .B2(n15649), .A(n11255), .ZN(P3_U3224) );
  XNOR2_X1 U13867 ( .A(n11256), .B(n11865), .ZN(n15109) );
  AND2_X1 U13868 ( .A1(n14636), .A2(n14792), .ZN(n14528) );
  INV_X1 U13869 ( .A(n14528), .ZN(n15068) );
  XNOR2_X1 U13870 ( .A(n11257), .B(n11865), .ZN(n15111) );
  NAND2_X1 U13871 ( .A1(n15111), .A2(n14656), .ZN(n11267) );
  AOI211_X1 U13872 ( .C1(n15107), .C2(n11259), .A(n14630), .B(n11258), .ZN(
        n15105) );
  INV_X1 U13873 ( .A(n15107), .ZN(n11264) );
  OAI22_X1 U13874 ( .A1(n11260), .A2(n14460), .B1(n11492), .B2(n14401), .ZN(
        n15106) );
  INV_X1 U13875 ( .A(n15106), .ZN(n11261) );
  OAI22_X1 U13876 ( .A1(n15074), .A2(n11261), .B1(n11322), .B2(n14633), .ZN(
        n11262) );
  AOI21_X1 U13877 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n15074), .A(n11262), .ZN(
        n11263) );
  OAI21_X1 U13878 ( .B1(n11264), .B2(n14614), .A(n11263), .ZN(n11265) );
  AOI21_X1 U13879 ( .B1(n15105), .B2(n15058), .A(n11265), .ZN(n11266) );
  OAI211_X1 U13880 ( .C1(n15109), .C2(n15068), .A(n11267), .B(n11266), .ZN(
        P1_U3285) );
  NAND2_X1 U13881 ( .A1(n11270), .A2(n11892), .ZN(n11273) );
  AOI22_X1 U13882 ( .A1(n11271), .A2(n11852), .B1(n11853), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11272) );
  OR2_X1 U13883 ( .A1(n14801), .A2(n12697), .ZN(n11291) );
  NAND2_X1 U13884 ( .A1(n14801), .A2(n12697), .ZN(n11274) );
  NAND2_X1 U13885 ( .A1(n11291), .A2(n11274), .ZN(n14791) );
  NAND2_X1 U13886 ( .A1(n14790), .A2(n14791), .ZN(n11276) );
  OR2_X1 U13887 ( .A1(n14801), .A2(n14307), .ZN(n11275) );
  NAND2_X1 U13888 ( .A1(n11276), .A2(n11275), .ZN(n11399) );
  NAND2_X1 U13889 ( .A1(n11277), .A2(n11892), .ZN(n11280) );
  AOI22_X1 U13890 ( .A1(n11278), .A2(n11852), .B1(n11853), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U13891 ( .A1(n11807), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11288) );
  OR2_X1 U13892 ( .A1(n10273), .A2(n11177), .ZN(n11287) );
  INV_X1 U13893 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U13894 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  NAND2_X1 U13895 ( .A1(n11294), .A2(n11283), .ZN(n14249) );
  OR2_X1 U13896 ( .A1(n11900), .A2(n14249), .ZN(n11286) );
  INV_X1 U13897 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11284) );
  OR2_X1 U13898 ( .A1(n6689), .A2(n11284), .ZN(n11285) );
  NAND4_X1 U13899 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n14306) );
  XNOR2_X1 U13900 ( .A(n14245), .B(n14306), .ZN(n11871) );
  INV_X1 U13901 ( .A(n11871), .ZN(n11398) );
  XNOR2_X1 U13902 ( .A(n11399), .B(n11398), .ZN(n14979) );
  INV_X1 U13903 ( .A(n14979), .ZN(n11308) );
  INV_X1 U13904 ( .A(n14308), .ZN(n12687) );
  OR2_X1 U13905 ( .A1(n14986), .A2(n12687), .ZN(n11289) );
  INV_X1 U13906 ( .A(n14791), .ZN(n14794) );
  OAI211_X1 U13907 ( .C1(n11292), .C2(n11871), .A(n11383), .B(n14792), .ZN(
        n11301) );
  AOI22_X1 U13908 ( .A1(n11807), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n11884), 
        .B2(P1_REG0_REG_14__SCAN_IN), .ZN(n11299) );
  INV_X1 U13909 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11293) );
  AND2_X1 U13910 ( .A1(n11294), .A2(n11293), .ZN(n11295) );
  OR2_X1 U13911 ( .A1(n11295), .A2(n11388), .ZN(n14934) );
  NAND2_X1 U13912 ( .A1(n6674), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11296) );
  OAI21_X1 U13913 ( .B1(n14934), .B2(n11900), .A(n11296), .ZN(n11297) );
  INV_X1 U13914 ( .A(n11297), .ZN(n11298) );
  OAI22_X1 U13915 ( .A1(n12713), .A2(n14401), .B1(n12697), .B2(n14460), .ZN(
        n14252) );
  INV_X1 U13916 ( .A(n14252), .ZN(n11300) );
  NAND2_X1 U13917 ( .A1(n11301), .A2(n11300), .ZN(n14983) );
  AOI21_X1 U13918 ( .B1(n14245), .B2(n6806), .A(n14630), .ZN(n11303) );
  NAND2_X1 U13919 ( .A1(n11303), .A2(n11394), .ZN(n14980) );
  OAI22_X1 U13920 ( .A1(n14636), .A2(n11177), .B1(n14249), .B2(n14633), .ZN(
        n11304) );
  AOI21_X1 U13921 ( .B1(n14245), .B2(n15052), .A(n11304), .ZN(n11305) );
  OAI21_X1 U13922 ( .B1(n14980), .B2(n14654), .A(n11305), .ZN(n11306) );
  AOI21_X1 U13923 ( .B1(n14983), .B2(n14636), .A(n11306), .ZN(n11307) );
  OAI21_X1 U13924 ( .B1(n15067), .B2(n11308), .A(n11307), .ZN(P1_U3280) );
  AOI22_X1 U13925 ( .A1(n15107), .A2(n12804), .B1(n11309), .B2(n14311), .ZN(
        n11310) );
  XNOR2_X1 U13926 ( .A(n11310), .B(n12824), .ZN(n11488) );
  AOI22_X1 U13927 ( .A1(n15107), .A2(n7074), .B1(n12817), .B2(n14311), .ZN(
        n11487) );
  XNOR2_X1 U13928 ( .A(n11488), .B(n11487), .ZN(n11319) );
  INV_X1 U13929 ( .A(n11311), .ZN(n11314) );
  INV_X1 U13930 ( .A(n11312), .ZN(n11313) );
  INV_X1 U13931 ( .A(n11489), .ZN(n11317) );
  AOI21_X1 U13932 ( .B1(n11319), .B2(n11318), .A(n11317), .ZN(n11325) );
  NAND2_X1 U13933 ( .A1(n14953), .A2(n15106), .ZN(n11320) );
  OAI211_X1 U13934 ( .C1(n14958), .C2(n11322), .A(n11321), .B(n11320), .ZN(
        n11323) );
  AOI21_X1 U13935 ( .B1(n15107), .B2(n14950), .A(n11323), .ZN(n11324) );
  OAI21_X1 U13936 ( .B1(n11325), .B2(n14277), .A(n11324), .ZN(P1_U3221) );
  AOI22_X1 U13937 ( .A1(n13649), .A2(n11326), .B1(n13549), .B2(n13693), .ZN(
        n11328) );
  OAI211_X1 U13938 ( .C1(n11329), .C2(n13630), .A(n11328), .B(n11327), .ZN(
        n11335) );
  INV_X1 U13939 ( .A(n11330), .ZN(n11331) );
  AOI211_X1 U13940 ( .C1(n11333), .C2(n11332), .A(n13653), .B(n11331), .ZN(
        n11334) );
  AOI211_X1 U13941 ( .C1(n15393), .C2(n13668), .A(n11335), .B(n11334), .ZN(
        n11336) );
  INV_X1 U13942 ( .A(n11336), .ZN(P2_U3189) );
  INV_X1 U13943 ( .A(n11342), .ZN(n11338) );
  XNOR2_X1 U13944 ( .A(n14912), .B(n13505), .ZN(n11505) );
  NAND2_X1 U13945 ( .A1(n13922), .A2(n13692), .ZN(n11506) );
  XNOR2_X1 U13946 ( .A(n11505), .B(n11506), .ZN(n11343) );
  AOI22_X1 U13947 ( .A1(n11339), .A2(n13649), .B1(n13659), .B2(n13693), .ZN(
        n11340) );
  NAND2_X1 U13948 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15227)
         );
  OAI211_X1 U13949 ( .C1(n12472), .C2(n13657), .A(n11340), .B(n15227), .ZN(
        n11347) );
  INV_X1 U13950 ( .A(n11341), .ZN(n11345) );
  AOI22_X1 U13951 ( .A1(n11342), .A2(n13676), .B1(n13641), .B2(n13693), .ZN(
        n11344) );
  NOR3_X1 U13952 ( .A1(n11345), .A2(n11344), .A3(n11343), .ZN(n11346) );
  AOI211_X1 U13953 ( .C1(n14912), .C2(n13668), .A(n11347), .B(n11346), .ZN(
        n11348) );
  OAI21_X1 U13954 ( .B1(n11508), .B2(n13653), .A(n11348), .ZN(P2_U3196) );
  XNOR2_X1 U13955 ( .A(n11349), .B(n11866), .ZN(n15133) );
  INV_X1 U13956 ( .A(n11350), .ZN(n11351) );
  AOI21_X1 U13957 ( .B1(n11351), .B2(n11984), .A(n14630), .ZN(n11353) );
  AOI22_X1 U13958 ( .A1(n11353), .A2(n11352), .B1(n14565), .B2(n14308), .ZN(
        n15125) );
  NAND2_X1 U13959 ( .A1(n14310), .A2(n14563), .ZN(n15124) );
  NOR2_X1 U13960 ( .A1(n15074), .A2(n15124), .ZN(n11355) );
  OAI22_X1 U13961 ( .A1(n14636), .A2(n10937), .B1(n11576), .B2(n14633), .ZN(
        n11354) );
  AOI211_X1 U13962 ( .C1(n11984), .C2(n15052), .A(n11355), .B(n11354), .ZN(
        n11356) );
  OAI21_X1 U13963 ( .B1(n15125), .B2(n14654), .A(n11356), .ZN(n11361) );
  NOR2_X1 U13964 ( .A1(n11358), .A2(n11357), .ZN(n15130) );
  INV_X1 U13965 ( .A(n11359), .ZN(n15129) );
  NOR3_X1 U13966 ( .A1(n15130), .A2(n15129), .A3(n15068), .ZN(n11360) );
  AOI211_X1 U13967 ( .C1(n14656), .C2(n15133), .A(n11361), .B(n11360), .ZN(
        n11362) );
  INV_X1 U13968 ( .A(n11362), .ZN(P1_U3283) );
  NAND2_X1 U13969 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14223)
         );
  NOR2_X1 U13970 ( .A1(n14376), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11363) );
  AOI21_X1 U13971 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14376), .A(n11363), 
        .ZN(n11366) );
  OAI21_X1 U13972 ( .B1(n11172), .B2(n11372), .A(n11364), .ZN(n11365) );
  NAND2_X1 U13973 ( .A1(n11365), .A2(n11366), .ZN(n14372) );
  OAI211_X1 U13974 ( .C1(n11366), .C2(n11365), .A(n14383), .B(n14372), .ZN(
        n11367) );
  NAND2_X1 U13975 ( .A1(n14223), .A2(n11367), .ZN(n11368) );
  AOI21_X1 U13976 ( .B1(n14343), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11368), 
        .ZN(n11377) );
  INV_X1 U13977 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U13978 ( .A1(n14376), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n11369), 
        .B2(n14373), .ZN(n11375) );
  INV_X1 U13979 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11373) );
  INV_X1 U13980 ( .A(n11370), .ZN(n11371) );
  OAI21_X1 U13981 ( .B1(n11373), .B2(n11372), .A(n11371), .ZN(n11374) );
  NAND2_X1 U13982 ( .A1(n11375), .A2(n11374), .ZN(n14377) );
  OAI211_X1 U13983 ( .C1(n11375), .C2(n11374), .A(n14389), .B(n14377), .ZN(
        n11376) );
  OAI211_X1 U13984 ( .C1(n15038), .C2(n14373), .A(n11377), .B(n11376), .ZN(
        P1_U3260) );
  INV_X1 U13985 ( .A(n11378), .ZN(n11380) );
  OAI222_X1 U13986 ( .A1(P3_U3151), .A2(n11381), .B1(n13468), .B2(n11380), 
        .C1(n11379), .C2(n11518), .ZN(P3_U3270) );
  INV_X1 U13987 ( .A(n14306), .ZN(n12707) );
  OR2_X1 U13988 ( .A1(n14245), .A2(n12707), .ZN(n11382) );
  NAND2_X1 U13989 ( .A1(n11384), .A2(n11892), .ZN(n11386) );
  AOI22_X1 U13990 ( .A1(n14361), .A2(n11852), .B1(n11853), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U13991 ( .A1(n14929), .A2(n12713), .ZN(n12001) );
  OAI211_X1 U13992 ( .C1(n11387), .C2(n12006), .A(n11463), .B(n14792), .ZN(
        n11393) );
  NOR2_X1 U13993 ( .A1(n11388), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11389) );
  OR2_X1 U13994 ( .A1(n11468), .A2(n11389), .ZN(n14292) );
  AOI22_X1 U13995 ( .A1(n11807), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n6674), 
        .B2(P1_REG2_REG_15__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U13996 ( .A1(n11884), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11390) );
  OAI211_X1 U13997 ( .C1(n14292), .C2(n11900), .A(n11391), .B(n11390), .ZN(
        n14304) );
  INV_X1 U13998 ( .A(n14304), .ZN(n12726) );
  OAI22_X1 U13999 ( .A1(n12726), .A2(n14401), .B1(n12707), .B2(n14460), .ZN(
        n14931) );
  INV_X1 U14000 ( .A(n14931), .ZN(n11392) );
  NAND2_X1 U14001 ( .A1(n11393), .A2(n11392), .ZN(n14977) );
  INV_X1 U14002 ( .A(n14977), .ZN(n11404) );
  OAI22_X1 U14003 ( .A1(n14636), .A2(n14362), .B1(n14934), .B2(n14633), .ZN(
        n11397) );
  INV_X1 U14004 ( .A(n14929), .ZN(n14975) );
  INV_X1 U14005 ( .A(n11394), .ZN(n11395) );
  OAI211_X1 U14006 ( .C1(n14975), .C2(n11395), .A(n15055), .B(n11466), .ZN(
        n14973) );
  NOR2_X1 U14007 ( .A1(n14973), .A2(n14654), .ZN(n11396) );
  AOI211_X1 U14008 ( .C1(n15052), .C2(n14929), .A(n11397), .B(n11396), .ZN(
        n11403) );
  OR2_X1 U14009 ( .A1(n14245), .A2(n14306), .ZN(n11400) );
  NAND2_X1 U14010 ( .A1(n11401), .A2(n12006), .ZN(n14971) );
  NAND3_X1 U14011 ( .A1(n14972), .A2(n14971), .A3(n14656), .ZN(n11402) );
  OAI211_X1 U14012 ( .C1(n15074), .C2(n11404), .A(n11403), .B(n11402), .ZN(
        P1_U3279) );
  XNOR2_X1 U14013 ( .A(n11405), .B(n11410), .ZN(n11406) );
  OAI222_X1 U14014 ( .A1(n11406), .A2(n13950), .B1(n15294), .B2(n13605), .C1(
        n13953), .C2(n12472), .ZN(n14908) );
  INV_X1 U14015 ( .A(n14908), .ZN(n11416) );
  INV_X1 U14016 ( .A(n11407), .ZN(n11408) );
  AOI21_X1 U14017 ( .B1(n11410), .B2(n11409), .A(n11408), .ZN(n14910) );
  OAI211_X1 U14018 ( .C1(n14907), .C2(n11411), .A(n11160), .B(n11640), .ZN(
        n14906) );
  AOI22_X1 U14019 ( .A1(n15305), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11584), 
        .B2(n15283), .ZN(n11413) );
  NAND2_X1 U14020 ( .A1(n12483), .A2(n15281), .ZN(n11412) );
  OAI211_X1 U14021 ( .C1(n14906), .C2(n13907), .A(n11413), .B(n11412), .ZN(
        n11414) );
  AOI21_X1 U14022 ( .B1(n14910), .B2(n15287), .A(n11414), .ZN(n11415) );
  OAI21_X1 U14023 ( .B1(n11416), .B2(n15305), .A(n11415), .ZN(P2_U3251) );
  AOI211_X1 U14024 ( .C1(n11419), .C2(n15390), .A(n11418), .B(n11417), .ZN(
        n11424) );
  AOI22_X1 U14025 ( .A1(n12470), .A2(n14059), .B1(n15424), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11420) );
  OAI21_X1 U14026 ( .B1(n11424), .B2(n15424), .A(n11420), .ZN(P2_U3512) );
  INV_X1 U14027 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11421) );
  NOR2_X1 U14028 ( .A1(n15409), .A2(n11421), .ZN(n11422) );
  AOI21_X1 U14029 ( .B1(n12470), .B2(n8335), .A(n11422), .ZN(n11423) );
  OAI21_X1 U14030 ( .B1(n11424), .B2(n15407), .A(n11423), .ZN(P2_U3469) );
  AND2_X1 U14031 ( .A1(n11425), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12661) );
  AOI21_X1 U14032 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14138), .A(n12661), 
        .ZN(n11426) );
  OAI21_X1 U14033 ( .B1(n11793), .B2(n14150), .A(n11426), .ZN(P2_U3304) );
  XNOR2_X1 U14034 ( .A(n11434), .B(n12848), .ZN(n11531) );
  XNOR2_X1 U14035 ( .A(n11531), .B(n15598), .ZN(n11433) );
  INV_X1 U14036 ( .A(n11427), .ZN(n11428) );
  NAND2_X1 U14037 ( .A1(n11428), .A2(n12216), .ZN(n11429) );
  INV_X1 U14038 ( .A(n11535), .ZN(n11431) );
  AOI21_X1 U14039 ( .B1(n11433), .B2(n11432), .A(n11431), .ZN(n11439) );
  AOI22_X1 U14040 ( .A1(n12216), .A2(n13020), .B1(n11434), .B2(n15429), .ZN(
        n11435) );
  NAND2_X1 U14041 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15517) );
  OAI211_X1 U14042 ( .C1(n11658), .C2(n13023), .A(n11435), .B(n15517), .ZN(
        n11436) );
  AOI21_X1 U14043 ( .B1(n11437), .B2(n13037), .A(n11436), .ZN(n11438) );
  OAI21_X1 U14044 ( .B1(n11439), .B2(n13027), .A(n11438), .ZN(P3_U3171) );
  NAND2_X1 U14045 ( .A1(n11440), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11441) );
  OAI211_X1 U14046 ( .C1(n11793), .C2(n14768), .A(n12132), .B(n11441), .ZN(
        P1_U3332) );
  INV_X1 U14047 ( .A(n12226), .ZN(n12334) );
  XNOR2_X1 U14048 ( .A(n11442), .B(n12334), .ZN(n15735) );
  OAI211_X1 U14049 ( .C1(n11444), .C2(n12226), .A(n11443), .B(n15671), .ZN(
        n11446) );
  AOI22_X1 U14050 ( .A1(n11688), .A2(n15654), .B1(n15653), .B2(n15598), .ZN(
        n11445) );
  OAI211_X1 U14051 ( .C1(n15662), .C2(n15735), .A(n11446), .B(n11445), .ZN(
        n15736) );
  NAND2_X1 U14052 ( .A1(n15736), .A2(n15682), .ZN(n11452) );
  NOR2_X1 U14053 ( .A1(n11447), .A2(n15718), .ZN(n15737) );
  INV_X1 U14054 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11449) );
  INV_X1 U14055 ( .A(n11540), .ZN(n11448) );
  OAI22_X1 U14056 ( .A1(n15682), .A2(n11449), .B1(n11448), .B2(n15676), .ZN(
        n11450) );
  AOI21_X1 U14057 ( .B1(n15679), .B2(n15737), .A(n11450), .ZN(n11451) );
  OAI211_X1 U14058 ( .C1(n15735), .C2(n11453), .A(n11452), .B(n11451), .ZN(
        P3_U3223) );
  NAND2_X1 U14059 ( .A1(n11454), .A2(n11892), .ZN(n11457) );
  AOI22_X1 U14060 ( .A1(n11853), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11852), 
        .B2(n11455), .ZN(n11456) );
  NAND2_X1 U14061 ( .A1(n12721), .A2(n12726), .ZN(n12014) );
  INV_X1 U14062 ( .A(n12713), .ZN(n14305) );
  NAND2_X1 U14063 ( .A1(n14929), .A2(n14305), .ZN(n11458) );
  NAND2_X1 U14064 ( .A1(n14972), .A2(n11458), .ZN(n11462) );
  INV_X1 U14065 ( .A(n11462), .ZN(n11460) );
  NAND2_X1 U14066 ( .A1(n11460), .A2(n11459), .ZN(n11612) );
  INV_X1 U14067 ( .A(n11612), .ZN(n11461) );
  AOI21_X1 U14068 ( .B1(n11876), .B2(n11462), .A(n11461), .ZN(n11552) );
  OAI21_X1 U14069 ( .B1(n11464), .B2(n11876), .A(n11595), .ZN(n11465) );
  INV_X1 U14070 ( .A(n11465), .ZN(n11550) );
  AOI21_X1 U14071 ( .B1(n12721), .B2(n11466), .A(n14630), .ZN(n11467) );
  OR2_X2 U14072 ( .A1(n11466), .A2(n12721), .ZN(n11613) );
  NAND2_X1 U14073 ( .A1(n11467), .A2(n11613), .ZN(n11548) );
  INV_X1 U14074 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U14075 ( .A1(n14305), .A2(n14563), .ZN(n11473) );
  OR2_X1 U14076 ( .A1(n11468), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U14077 ( .A1(n11601), .A2(n11469), .ZN(n14945) );
  AOI22_X1 U14078 ( .A1(n6675), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11884), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14079 ( .A1(n11807), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11470) );
  OAI211_X1 U14080 ( .C1(n14945), .C2(n11900), .A(n11471), .B(n11470), .ZN(
        n14431) );
  NAND2_X1 U14081 ( .A1(n14431), .A2(n14565), .ZN(n11472) );
  AND2_X1 U14082 ( .A1(n11473), .A2(n11472), .ZN(n14293) );
  OAI21_X1 U14083 ( .B1(n14292), .B2(n14633), .A(n14293), .ZN(n11474) );
  NAND2_X1 U14084 ( .A1(n11474), .A2(n14636), .ZN(n11475) );
  OAI21_X1 U14085 ( .B1(n14636), .B2(n11476), .A(n11475), .ZN(n11477) );
  AOI21_X1 U14086 ( .B1(n12721), .B2(n15052), .A(n11477), .ZN(n11478) );
  OAI21_X1 U14087 ( .B1(n11548), .B2(n14654), .A(n11478), .ZN(n11479) );
  AOI21_X1 U14088 ( .B1(n11550), .B2(n14528), .A(n11479), .ZN(n11480) );
  OAI21_X1 U14089 ( .B1(n11552), .B2(n15067), .A(n11480), .ZN(P1_U3278) );
  INV_X1 U14090 ( .A(n11481), .ZN(n11482) );
  OAI222_X1 U14091 ( .A1(P3_U3151), .A2(n11484), .B1(n11518), .B2(n11483), 
        .C1(n13468), .C2(n11482), .ZN(P3_U3269) );
  OAI22_X1 U14092 ( .A1(n11485), .A2(n12823), .B1(n11492), .B2(n6686), .ZN(
        n11486) );
  XOR2_X1 U14093 ( .A(n12824), .B(n11486), .Z(n11568) );
  INV_X1 U14094 ( .A(n11487), .ZN(n11491) );
  INV_X1 U14095 ( .A(n11488), .ZN(n11490) );
  NOR2_X1 U14096 ( .A1(n11492), .A2(n12826), .ZN(n11493) );
  AOI21_X1 U14097 ( .B1(n15115), .B2(n7074), .A(n11493), .ZN(n11566) );
  INV_X1 U14098 ( .A(n11566), .ZN(n11494) );
  XOR2_X1 U14099 ( .A(n11568), .B(n11569), .Z(n11500) );
  AOI22_X1 U14100 ( .A1(n14953), .A2(n11495), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11496) );
  OAI21_X1 U14101 ( .B1(n14958), .B2(n11497), .A(n11496), .ZN(n11498) );
  AOI21_X1 U14102 ( .B1(n15115), .B2(n14950), .A(n11498), .ZN(n11499) );
  OAI21_X1 U14103 ( .B1(n11500), .B2(n14277), .A(n11499), .ZN(P1_U3231) );
  XNOR2_X1 U14104 ( .A(n12470), .B(n13493), .ZN(n11501) );
  AND2_X1 U14105 ( .A1(n13509), .A2(n13691), .ZN(n11502) );
  NAND2_X1 U14106 ( .A1(n11501), .A2(n11502), .ZN(n11582) );
  INV_X1 U14107 ( .A(n11501), .ZN(n11587) );
  INV_X1 U14108 ( .A(n11502), .ZN(n11503) );
  NAND2_X1 U14109 ( .A1(n11587), .A2(n11503), .ZN(n11504) );
  NAND2_X1 U14110 ( .A1(n11582), .A2(n11504), .ZN(n11510) );
  INV_X1 U14111 ( .A(n11505), .ZN(n11507) );
  INV_X1 U14112 ( .A(n11583), .ZN(n11589) );
  AOI211_X1 U14113 ( .C1(n11510), .C2(n11509), .A(n13653), .B(n11589), .ZN(
        n11511) );
  INV_X1 U14114 ( .A(n11511), .ZN(n11516) );
  OAI22_X1 U14115 ( .A1(n13646), .A2(n11512), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15232), .ZN(n11513) );
  AOI21_X1 U14116 ( .B1(n13649), .B2(n11514), .A(n11513), .ZN(n11515) );
  OAI211_X1 U14117 ( .C1(n7204), .C2(n13662), .A(n11516), .B(n11515), .ZN(
        P2_U3206) );
  INV_X1 U14118 ( .A(n11517), .ZN(n11520) );
  OAI222_X1 U14119 ( .A1(P3_U3151), .A2(n13078), .B1(n13468), .B2(n11520), 
        .C1(n11519), .C2(n11518), .ZN(P3_U3268) );
  XNOR2_X1 U14120 ( .A(n11521), .B(n11527), .ZN(n11523) );
  OAI22_X1 U14121 ( .A1(n11696), .A2(n15637), .B1(n12849), .B2(n15673), .ZN(
        n11522) );
  AOI21_X1 U14122 ( .B1(n11523), .B2(n15671), .A(n11522), .ZN(n14894) );
  AND2_X1 U14123 ( .A1(n11694), .A2(n15677), .ZN(n14891) );
  INV_X1 U14124 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11525) );
  INV_X1 U14125 ( .A(n11695), .ZN(n11524) );
  OAI22_X1 U14126 ( .A1(n15682), .A2(n11525), .B1(n11524), .B2(n15676), .ZN(
        n11526) );
  AOI21_X1 U14127 ( .B1(n14891), .B2(n15679), .A(n11526), .ZN(n11530) );
  XNOR2_X1 U14128 ( .A(n11528), .B(n11527), .ZN(n14892) );
  NAND2_X1 U14129 ( .A1(n14892), .A2(n15631), .ZN(n11529) );
  OAI211_X1 U14130 ( .C1(n14894), .C2(n15649), .A(n11530), .B(n11529), .ZN(
        P3_U3221) );
  XNOR2_X1 U14131 ( .A(n11541), .B(n12921), .ZN(n11645) );
  XNOR2_X1 U14132 ( .A(n11645), .B(n11658), .ZN(n11538) );
  INV_X1 U14133 ( .A(n11531), .ZN(n11533) );
  INV_X1 U14134 ( .A(n15598), .ZN(n11532) );
  NAND2_X1 U14135 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  INV_X1 U14136 ( .A(n11649), .ZN(n11536) );
  AOI211_X1 U14137 ( .C1(n11538), .C2(n11537), .A(n13027), .B(n11536), .ZN(
        n11547) );
  AOI21_X1 U14138 ( .B1(n11688), .B2(n15430), .A(n11539), .ZN(n11545) );
  NAND2_X1 U14139 ( .A1(n13037), .A2(n11540), .ZN(n11544) );
  NAND2_X1 U14140 ( .A1(n11541), .A2(n15429), .ZN(n11543) );
  NAND2_X1 U14141 ( .A1(n13020), .A2(n15598), .ZN(n11542) );
  NAND4_X1 U14142 ( .A1(n11545), .A2(n11544), .A3(n11543), .A4(n11542), .ZN(
        n11546) );
  OR2_X1 U14143 ( .A1(n11547), .A2(n11546), .ZN(P3_U3157) );
  INV_X1 U14144 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11554) );
  INV_X1 U14145 ( .A(n12721), .ZN(n14301) );
  OAI211_X1 U14146 ( .C1(n14301), .C2(n15126), .A(n11548), .B(n14293), .ZN(
        n11549) );
  AOI21_X1 U14147 ( .B1(n11550), .B2(n14792), .A(n11549), .ZN(n11551) );
  OAI21_X1 U14148 ( .B1(n11552), .B2(n14732), .A(n11551), .ZN(n11555) );
  NAND2_X1 U14149 ( .A1(n11555), .A2(n15150), .ZN(n11553) );
  OAI21_X1 U14150 ( .B1(n15150), .B2(n11554), .A(n11553), .ZN(P1_U3543) );
  INV_X1 U14151 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U14152 ( .A1(n11555), .A2(n15113), .ZN(n11556) );
  OAI21_X1 U14153 ( .B1(n15113), .B2(n11557), .A(n11556), .ZN(P1_U3504) );
  INV_X1 U14154 ( .A(n15631), .ZN(n13250) );
  XNOR2_X1 U14155 ( .A(n11558), .B(n12335), .ZN(n14898) );
  INV_X1 U14156 ( .A(n14898), .ZN(n11565) );
  XOR2_X1 U14157 ( .A(n11559), .B(n12335), .Z(n11560) );
  OAI222_X1 U14158 ( .A1(n15673), .A2(n12994), .B1(n15637), .B2(n11658), .C1(
        n11560), .C2(n15641), .ZN(n14896) );
  NAND2_X1 U14159 ( .A1(n14896), .A2(n15682), .ZN(n11564) );
  NOR2_X1 U14160 ( .A1(n11650), .A2(n15718), .ZN(n14897) );
  INV_X1 U14161 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15523) );
  INV_X1 U14162 ( .A(n11655), .ZN(n11561) );
  OAI22_X1 U14163 ( .A1(n15682), .A2(n15523), .B1(n11561), .B2(n15676), .ZN(
        n11562) );
  AOI21_X1 U14164 ( .B1(n15679), .B2(n14897), .A(n11562), .ZN(n11563) );
  OAI211_X1 U14165 ( .C1(n13250), .C2(n11565), .A(n11564), .B(n11563), .ZN(
        P3_U3222) );
  NAND2_X1 U14166 ( .A1(n11984), .A2(n12804), .ZN(n11571) );
  NAND2_X1 U14167 ( .A1(n14309), .A2(n7074), .ZN(n11570) );
  NAND2_X1 U14168 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  XNOR2_X1 U14169 ( .A(n11572), .B(n12824), .ZN(n12689) );
  NOR2_X1 U14170 ( .A1(n11573), .A2(n12826), .ZN(n11574) );
  AOI21_X1 U14171 ( .B1(n11984), .B2(n7074), .A(n11574), .ZN(n12690) );
  XNOR2_X1 U14172 ( .A(n12689), .B(n12690), .ZN(n11575) );
  OAI211_X1 U14173 ( .C1(n6805), .C2(n11575), .A(n12692), .B(n14951), .ZN(
        n11581) );
  NOR2_X1 U14174 ( .A1(n14958), .A2(n11576), .ZN(n11579) );
  OAI21_X1 U14175 ( .B1(n14262), .B2(n12687), .A(n11577), .ZN(n11578) );
  AOI211_X1 U14176 ( .C1(n14265), .C2(n14310), .A(n11579), .B(n11578), .ZN(
        n11580) );
  OAI211_X1 U14177 ( .C1(n15127), .C2(n14300), .A(n11581), .B(n11580), .ZN(
        P1_U3217) );
  XNOR2_X1 U14178 ( .A(n12483), .B(n13505), .ZN(n11663) );
  NAND2_X1 U14179 ( .A1(n13922), .A2(n13690), .ZN(n11664) );
  XNOR2_X1 U14180 ( .A(n11663), .B(n11664), .ZN(n11590) );
  AOI22_X1 U14181 ( .A1(n11584), .A2(n13649), .B1(n13659), .B2(n13691), .ZN(
        n11586) );
  OAI211_X1 U14182 ( .C1(n13605), .C2(n13657), .A(n11586), .B(n11585), .ZN(
        n11593) );
  NOR3_X1 U14183 ( .A1(n11587), .A2(n12472), .A3(n13663), .ZN(n11588) );
  AOI21_X1 U14184 ( .B1(n11589), .B2(n13676), .A(n11588), .ZN(n11591) );
  NOR2_X1 U14185 ( .A1(n11591), .A2(n11590), .ZN(n11592) );
  AOI211_X1 U14186 ( .C1(n12483), .C2(n13668), .A(n11593), .B(n11592), .ZN(
        n11594) );
  OAI21_X1 U14187 ( .B1(n11667), .B2(n13653), .A(n11594), .ZN(P2_U3187) );
  INV_X1 U14188 ( .A(n14945), .ZN(n11610) );
  NAND2_X1 U14189 ( .A1(n11595), .A2(n12013), .ZN(n14430) );
  NAND2_X1 U14190 ( .A1(n11596), .A2(n11892), .ZN(n11599) );
  AOI22_X1 U14191 ( .A1(n11853), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11852), 
        .B2(n11597), .ZN(n11598) );
  XNOR2_X1 U14192 ( .A(n14940), .B(n14431), .ZN(n11874) );
  XNOR2_X1 U14193 ( .A(n14430), .B(n11874), .ZN(n11609) );
  INV_X1 U14194 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14195 ( .A1(n11601), .A2(n11600), .ZN(n11602) );
  AND2_X1 U14196 ( .A1(n11844), .A2(n11602), .ZN(n14647) );
  NAND2_X1 U14197 ( .A1(n14647), .A2(n11889), .ZN(n11607) );
  NAND2_X1 U14198 ( .A1(n11807), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U14199 ( .A1(n11884), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11603) );
  OAI211_X1 U14200 ( .C1(n10273), .C2(n11369), .A(n11604), .B(n11603), .ZN(
        n11605) );
  INV_X1 U14201 ( .A(n11605), .ZN(n11606) );
  NAND2_X1 U14202 ( .A1(n11607), .A2(n11606), .ZN(n14435) );
  INV_X1 U14203 ( .A(n14435), .ZN(n12737) );
  OAI22_X1 U14204 ( .A1(n12737), .A2(n14401), .B1(n12726), .B2(n14460), .ZN(
        n14942) );
  INV_X1 U14205 ( .A(n14942), .ZN(n11608) );
  OAI21_X1 U14206 ( .B1(n11609), .B2(n15128), .A(n11608), .ZN(n14968) );
  AOI21_X1 U14207 ( .B1(n11610), .B2(n15070), .A(n14968), .ZN(n11619) );
  OR2_X1 U14208 ( .A1(n12721), .A2(n14304), .ZN(n11611) );
  XNOR2_X1 U14209 ( .A(n14412), .B(n14429), .ZN(n14970) );
  INV_X1 U14210 ( .A(n14940), .ZN(n14967) );
  INV_X1 U14211 ( .A(n11613), .ZN(n11615) );
  NOR2_X2 U14212 ( .A1(n14940), .A2(n11613), .ZN(n14651) );
  INV_X1 U14213 ( .A(n14651), .ZN(n11614) );
  OAI211_X1 U14214 ( .C1(n14967), .C2(n11615), .A(n11614), .B(n15055), .ZN(
        n14966) );
  AOI22_X1 U14215 ( .A1(n14940), .A2(n15052), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n15074), .ZN(n11616) );
  OAI21_X1 U14216 ( .B1(n14966), .B2(n14654), .A(n11616), .ZN(n11617) );
  AOI21_X1 U14217 ( .B1(n14970), .B2(n14656), .A(n11617), .ZN(n11618) );
  OAI21_X1 U14218 ( .B1(n11619), .B2(n15074), .A(n11618), .ZN(P1_U3277) );
  INV_X1 U14219 ( .A(n11620), .ZN(n12248) );
  XNOR2_X1 U14220 ( .A(n11621), .B(n6705), .ZN(n11624) );
  NAND2_X1 U14221 ( .A1(n12992), .A2(n15654), .ZN(n11622) );
  OAI21_X1 U14222 ( .B1(n12994), .B2(n15637), .A(n11622), .ZN(n11623) );
  AOI21_X1 U14223 ( .B1(n11624), .B2(n15671), .A(n11623), .ZN(n14889) );
  NOR2_X1 U14224 ( .A1(n12995), .A2(n15718), .ZN(n14886) );
  INV_X1 U14225 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15559) );
  INV_X1 U14226 ( .A(n12998), .ZN(n11625) );
  OAI22_X1 U14227 ( .A1(n15682), .A2(n15559), .B1(n11625), .B2(n15676), .ZN(
        n11626) );
  AOI21_X1 U14228 ( .B1(n14886), .B2(n15679), .A(n11626), .ZN(n11629) );
  XNOR2_X1 U14229 ( .A(n11627), .B(n6705), .ZN(n14887) );
  NAND2_X1 U14230 ( .A1(n14887), .A2(n15631), .ZN(n11628) );
  OAI211_X1 U14231 ( .C1(n14889), .C2(n15649), .A(n11629), .B(n11628), .ZN(
        P3_U3220) );
  OAI222_X1 U14232 ( .A1(P2_U3088), .A2(n11631), .B1(n14150), .B2(n11790), 
        .C1(n11630), .C2(n14152), .ZN(P2_U3303) );
  INV_X1 U14233 ( .A(n11632), .ZN(n11633) );
  AOI21_X1 U14234 ( .B1(n11635), .B2(n11634), .A(n11633), .ZN(n14092) );
  XNOR2_X1 U14235 ( .A(n11636), .B(n11635), .ZN(n11637) );
  AOI222_X1 U14236 ( .A1(n11637), .A2(n15293), .B1(n13689), .B2(n13988), .C1(
        n13690), .C2(n13991), .ZN(n14091) );
  OAI21_X1 U14237 ( .B1(n11672), .B2(n15298), .A(n14091), .ZN(n11638) );
  NAND2_X1 U14238 ( .A1(n11638), .A2(n15303), .ZN(n11643) );
  INV_X1 U14239 ( .A(n13994), .ZN(n11639) );
  AOI211_X1 U14240 ( .C1(n14089), .C2(n11640), .A(n13922), .B(n11639), .ZN(
        n14088) );
  OAI22_X1 U14241 ( .A1(n7202), .A2(n13998), .B1(n7976), .B2(n15303), .ZN(
        n11641) );
  AOI21_X1 U14242 ( .B1(n14088), .B2(n15285), .A(n11641), .ZN(n11642) );
  OAI211_X1 U14243 ( .C1(n14092), .C2(n14004), .A(n11643), .B(n11642), .ZN(
        P2_U3250) );
  OAI222_X1 U14244 ( .A1(n14771), .A2(n11791), .B1(P1_U3086), .B2(n11644), 
        .C1(n14768), .C2(n11790), .ZN(P1_U3331) );
  INV_X1 U14245 ( .A(n11645), .ZN(n11646) );
  NAND2_X1 U14246 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  XNOR2_X1 U14247 ( .A(n11650), .B(n12921), .ZN(n11651) );
  NAND2_X1 U14248 ( .A1(n11652), .A2(n11651), .ZN(n11690) );
  NAND2_X1 U14249 ( .A1(n11689), .A2(n11690), .ZN(n11653) );
  XNOR2_X1 U14250 ( .A(n11653), .B(n11696), .ZN(n11662) );
  NOR2_X1 U14251 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11654), .ZN(n15526) );
  AOI21_X1 U14252 ( .B1(n13043), .B2(n15430), .A(n15526), .ZN(n11657) );
  NAND2_X1 U14253 ( .A1(n13037), .A2(n11655), .ZN(n11656) );
  OAI211_X1 U14254 ( .C1(n11658), .C2(n13035), .A(n11657), .B(n11656), .ZN(
        n11659) );
  AOI21_X1 U14255 ( .B1(n11660), .B2(n15429), .A(n11659), .ZN(n11661) );
  OAI21_X1 U14256 ( .B1(n11662), .B2(n13027), .A(n11661), .ZN(P3_U3176) );
  INV_X1 U14257 ( .A(n11663), .ZN(n11665) );
  NAND2_X1 U14258 ( .A1(n11665), .A2(n11664), .ZN(n11666) );
  XNOR2_X1 U14259 ( .A(n14089), .B(n13505), .ZN(n13474) );
  AOI22_X1 U14260 ( .A1(n11669), .A2(n13676), .B1(n13641), .B2(n13992), .ZN(
        n11677) );
  AND2_X1 U14261 ( .A1(n13509), .A2(n13992), .ZN(n11668) );
  INV_X1 U14262 ( .A(n13478), .ZN(n11676) );
  OAI22_X1 U14263 ( .A1(n13630), .A2(n11671), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11670), .ZN(n11674) );
  OAI22_X1 U14264 ( .A1(n13657), .A2(n13615), .B1(n13674), .B2(n11672), .ZN(
        n11673) );
  AOI211_X1 U14265 ( .C1(n14089), .C2(n13668), .A(n11674), .B(n11673), .ZN(
        n11675) );
  OAI21_X1 U14266 ( .B1(n11677), .B2(n11676), .A(n11675), .ZN(P2_U3213) );
  NAND2_X1 U14267 ( .A1(n11678), .A2(n12340), .ZN(n11679) );
  NAND3_X1 U14268 ( .A1(n11680), .A2(n15671), .A3(n11679), .ZN(n11682) );
  AOI22_X1 U14269 ( .A1(n12893), .A2(n15653), .B1(n15654), .B2(n13042), .ZN(
        n11681) );
  INV_X1 U14270 ( .A(n12340), .ZN(n11683) );
  XNOR2_X1 U14271 ( .A(n11684), .B(n11683), .ZN(n13385) );
  AOI22_X1 U14272 ( .A1(n15649), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n6668), 
        .B2(n12896), .ZN(n11685) );
  OAI21_X1 U14273 ( .B1(n13448), .B2(n13320), .A(n11685), .ZN(n11686) );
  AOI21_X1 U14274 ( .B1(n13385), .B2(n15631), .A(n11686), .ZN(n11687) );
  OAI21_X1 U14275 ( .B1(n13387), .B2(n15649), .A(n11687), .ZN(P3_U3219) );
  NAND2_X1 U14276 ( .A1(n11689), .A2(n11688), .ZN(n11691) );
  XNOR2_X1 U14277 ( .A(n11694), .B(n12921), .ZN(n12844) );
  XNOR2_X1 U14278 ( .A(n12844), .B(n12994), .ZN(n11692) );
  XNOR2_X1 U14279 ( .A(n12843), .B(n11692), .ZN(n11702) );
  NOR2_X1 U14280 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11693), .ZN(n15544) );
  AOI21_X1 U14281 ( .B1(n12893), .B2(n15430), .A(n15544), .ZN(n11700) );
  NAND2_X1 U14282 ( .A1(n11694), .A2(n15429), .ZN(n11699) );
  NAND2_X1 U14283 ( .A1(n13037), .A2(n11695), .ZN(n11698) );
  OR2_X1 U14284 ( .A1(n11696), .A2(n13035), .ZN(n11697) );
  NAND4_X1 U14285 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  AOI21_X1 U14286 ( .B1(n11702), .B2(n15432), .A(n11701), .ZN(n11703) );
  INV_X1 U14287 ( .A(n11703), .ZN(P3_U3164) );
  MUX2_X1 U14288 ( .A(n11704), .B(P1_REG2_REG_3__SCAN_IN), .S(n15074), .Z(
        n11713) );
  INV_X1 U14289 ( .A(n11705), .ZN(n15059) );
  NAND2_X1 U14290 ( .A1(n11706), .A2(n15059), .ZN(n11710) );
  OAI22_X1 U14291 ( .A1(n14614), .A2(n11707), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14633), .ZN(n11708) );
  INV_X1 U14292 ( .A(n11708), .ZN(n11709) );
  OAI211_X1 U14293 ( .C1(n14654), .C2(n11711), .A(n11710), .B(n11709), .ZN(
        n11712) );
  OR2_X1 U14294 ( .A1(n11713), .A2(n11712), .ZN(P1_U3290) );
  INV_X1 U14295 ( .A(n11761), .ZN(n14140) );
  OAI222_X1 U14296 ( .A1(n14771), .A2(n11762), .B1(n14768), .B2(n14140), .C1(
        n6688), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U14297 ( .A1(n14152), .A2(n11716), .B1(P2_U3088), .B2(n11715), 
        .C1(n14150), .C2(n11714), .ZN(P2_U3305) );
  INV_X1 U14298 ( .A(n11719), .ZN(n11720) );
  NAND2_X1 U14299 ( .A1(n11720), .A2(n13465), .ZN(n11721) );
  MUX2_X1 U14300 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11804), .Z(n11731) );
  XNOR2_X1 U14301 ( .A(n11731), .B(SI_30_), .ZN(n11733) );
  INV_X1 U14302 ( .A(n11733), .ZN(n11723) );
  INV_X1 U14303 ( .A(n12577), .ZN(n14763) );
  INV_X1 U14304 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12144) );
  INV_X1 U14305 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11725) );
  NOR2_X1 U14306 ( .A1(n11902), .A2(n11725), .ZN(n11730) );
  INV_X1 U14307 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n11726) );
  NOR2_X1 U14308 ( .A1(n10273), .A2(n11726), .ZN(n11729) );
  INV_X1 U14309 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11727) );
  NOR2_X1 U14310 ( .A1(n6689), .A2(n11727), .ZN(n11728) );
  INV_X1 U14311 ( .A(n11731), .ZN(n11732) );
  MUX2_X1 U14312 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11804), .Z(n11735) );
  XNOR2_X1 U14313 ( .A(n11735), .B(SI_31_), .ZN(n11736) );
  NAND2_X1 U14314 ( .A1(n14759), .A2(n11892), .ZN(n11739) );
  INV_X1 U14315 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14754) );
  OR2_X1 U14316 ( .A1(n11893), .A2(n14754), .ZN(n11738) );
  XOR2_X1 U14317 ( .A(n14402), .B(n14397), .Z(n12122) );
  INV_X1 U14318 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14319 ( .A1(n6674), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11741) );
  NAND2_X1 U14320 ( .A1(n11884), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11740) );
  OAI211_X1 U14321 ( .C1(n11902), .C2(n11742), .A(n11741), .B(n11740), .ZN(
        n14457) );
  INV_X1 U14322 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14761) );
  XOR2_X1 U14323 ( .A(n14457), .B(n14396), .Z(n11909) );
  INV_X1 U14324 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14765) );
  NOR2_X1 U14325 ( .A1(n6676), .A2(n14765), .ZN(n11743) );
  NAND2_X1 U14326 ( .A1(n11807), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11752) );
  INV_X1 U14327 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n11744) );
  OR2_X1 U14328 ( .A1(n10273), .A2(n11744), .ZN(n11751) );
  INV_X1 U14329 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11843) );
  INV_X1 U14330 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14261) );
  NAND2_X1 U14331 ( .A1(n11809), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U14332 ( .A1(n11784), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U14333 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n11899), .ZN(n11898) );
  INV_X1 U14334 ( .A(n11898), .ZN(n11745) );
  NAND2_X1 U14335 ( .A1(n11745), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11775) );
  INV_X1 U14336 ( .A(n11775), .ZN(n11746) );
  NAND2_X1 U14337 ( .A1(n11746), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11764) );
  INV_X1 U14338 ( .A(n11764), .ZN(n11747) );
  NAND2_X1 U14339 ( .A1(n11747), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14458) );
  OR2_X1 U14340 ( .A1(n11900), .A2(n14458), .ZN(n11750) );
  INV_X1 U14341 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n11748) );
  OR2_X1 U14342 ( .A1(n6689), .A2(n11748), .ZN(n11749) );
  XNOR2_X1 U14343 ( .A(n14666), .B(n14302), .ZN(n14450) );
  NAND2_X1 U14344 ( .A1(n12133), .A2(n11892), .ZN(n11754) );
  OR2_X1 U14345 ( .A1(n6676), .A2(n12134), .ZN(n11753) );
  AND2_X2 U14346 ( .A1(n11754), .A2(n11753), .ZN(n14495) );
  NAND2_X1 U14347 ( .A1(n11807), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11760) );
  INV_X1 U14348 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14497) );
  OR2_X1 U14349 ( .A1(n10273), .A2(n14497), .ZN(n11759) );
  INV_X1 U14350 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14156) );
  NAND2_X1 U14351 ( .A1(n11775), .A2(n14156), .ZN(n11755) );
  NAND2_X1 U14352 ( .A1(n11764), .A2(n11755), .ZN(n14496) );
  OR2_X1 U14353 ( .A1(n11900), .A2(n14496), .ZN(n11758) );
  INV_X1 U14354 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n11756) );
  OR2_X1 U14355 ( .A1(n6689), .A2(n11756), .ZN(n11757) );
  NOR2_X1 U14356 ( .A1(n14495), .A2(n14426), .ZN(n14447) );
  NAND2_X1 U14357 ( .A1(n11807), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11769) );
  INV_X1 U14358 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14476) );
  OR2_X1 U14359 ( .A1(n10273), .A2(n14476), .ZN(n11768) );
  INV_X1 U14360 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11763) );
  XNOR2_X1 U14361 ( .A(n11764), .B(n11763), .ZN(n14475) );
  OR2_X1 U14362 ( .A1(n11900), .A2(n14475), .ZN(n11767) );
  INV_X1 U14363 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n11765) );
  OR2_X1 U14364 ( .A1(n6689), .A2(n11765), .ZN(n11766) );
  NAND2_X1 U14365 ( .A1(n14674), .A2(n14461), .ZN(n14449) );
  NAND2_X1 U14366 ( .A1(n14144), .A2(n11892), .ZN(n11772) );
  OR2_X1 U14367 ( .A1(n6676), .A2(n14770), .ZN(n11771) );
  NAND2_X1 U14368 ( .A1(n6675), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11780) );
  INV_X1 U14369 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11773) );
  OR2_X1 U14370 ( .A1(n6689), .A2(n11773), .ZN(n11779) );
  INV_X1 U14371 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U14372 ( .A1(n11898), .A2(n14283), .ZN(n11774) );
  NAND2_X1 U14373 ( .A1(n11775), .A2(n11774), .ZN(n14505) );
  OR2_X1 U14374 ( .A1(n11900), .A2(n14505), .ZN(n11778) );
  INV_X1 U14375 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11776) );
  OR2_X1 U14376 ( .A1(n11902), .A2(n11776), .ZN(n11777) );
  NAND4_X1 U14377 ( .A1(n11780), .A2(n11779), .A3(n11778), .A4(n11777), .ZN(
        n14424) );
  INV_X1 U14378 ( .A(n14424), .ZN(n14205) );
  NAND2_X1 U14379 ( .A1(n14688), .A2(n14205), .ZN(n14446) );
  OR2_X1 U14380 ( .A1(n14688), .A2(n14205), .ZN(n11781) );
  NAND2_X1 U14381 ( .A1(n14446), .A2(n11781), .ZN(n14423) );
  NAND2_X1 U14382 ( .A1(n6675), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11789) );
  INV_X1 U14383 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11782) );
  OR2_X1 U14384 ( .A1(n11902), .A2(n11782), .ZN(n11788) );
  OAI21_X1 U14385 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11784), .A(n11783), 
        .ZN(n14537) );
  OR2_X1 U14386 ( .A1(n11900), .A2(n14537), .ZN(n11787) );
  INV_X1 U14387 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n11785) );
  OR2_X1 U14388 ( .A1(n6689), .A2(n11785), .ZN(n11786) );
  NAND4_X1 U14389 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n14303) );
  OR2_X1 U14390 ( .A1(n6676), .A2(n11791), .ZN(n11792) );
  INV_X1 U14391 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11794) );
  OR2_X1 U14392 ( .A1(n6676), .A2(n11794), .ZN(n11795) );
  NAND2_X2 U14393 ( .A1(n11796), .A2(n11795), .ZN(n14557) );
  NAND2_X1 U14394 ( .A1(n11807), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11803) );
  INV_X1 U14395 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n11797) );
  OR2_X1 U14396 ( .A1(n10273), .A2(n11797), .ZN(n11802) );
  OAI21_X1 U14397 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11809), .A(n11798), 
        .ZN(n14554) );
  OR2_X1 U14398 ( .A1(n11900), .A2(n14554), .ZN(n11801) );
  INV_X1 U14399 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11799) );
  OR2_X1 U14400 ( .A1(n6689), .A2(n11799), .ZN(n11800) );
  NAND4_X1 U14401 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n14566) );
  OR2_X1 U14402 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  XNOR2_X1 U14403 ( .A(n11806), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14772) );
  NAND2_X1 U14404 ( .A1(n11807), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11816) );
  INV_X1 U14405 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11808) );
  OR2_X1 U14406 ( .A1(n10273), .A2(n11808), .ZN(n11815) );
  INV_X1 U14407 ( .A(n11822), .ZN(n11811) );
  INV_X1 U14408 ( .A(n11809), .ZN(n11810) );
  OAI21_X1 U14409 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11811), .A(n11810), 
        .ZN(n14571) );
  OR2_X1 U14410 ( .A1(n11900), .A2(n14571), .ZN(n11814) );
  INV_X1 U14411 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11812) );
  OR2_X1 U14412 ( .A1(n6689), .A2(n11812), .ZN(n11813) );
  NAND4_X1 U14413 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n14420) );
  INV_X1 U14414 ( .A(n14420), .ZN(n14443) );
  XNOR2_X1 U14415 ( .A(n7346), .B(n14443), .ZN(n14575) );
  OR2_X1 U14416 ( .A1(n6676), .A2(n11819), .ZN(n11820) );
  OR2_X1 U14417 ( .A1(n11883), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11823) );
  AND2_X1 U14418 ( .A1(n11823), .A2(n11822), .ZN(n14589) );
  NAND2_X1 U14419 ( .A1(n14589), .A2(n11889), .ZN(n11829) );
  INV_X1 U14420 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11826) );
  NAND2_X1 U14421 ( .A1(n6674), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11825) );
  NAND2_X1 U14422 ( .A1(n11884), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11824) );
  OAI211_X1 U14423 ( .C1(n11826), .C2(n11902), .A(n11825), .B(n11824), .ZN(
        n11827) );
  INV_X1 U14424 ( .A(n11827), .ZN(n11828) );
  NAND2_X1 U14425 ( .A1(n11829), .A2(n11828), .ZN(n14564) );
  OR2_X1 U14426 ( .A1(n14590), .A2(n14564), .ZN(n14419) );
  NAND2_X1 U14427 ( .A1(n14590), .A2(n14564), .ZN(n11830) );
  AOI22_X1 U14428 ( .A1(n11853), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14390), 
        .B2(n11852), .ZN(n11832) );
  NOR2_X1 U14429 ( .A1(n11845), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11834) );
  OR2_X1 U14430 ( .A1(n11881), .A2(n11834), .ZN(n14611) );
  INV_X1 U14431 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U14432 ( .A1(n6674), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11836) );
  NAND2_X1 U14433 ( .A1(n11884), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11835) );
  OAI211_X1 U14434 ( .C1(n11837), .C2(n11902), .A(n11836), .B(n11835), .ZN(
        n11838) );
  INV_X1 U14435 ( .A(n11838), .ZN(n11839) );
  OAI21_X1 U14436 ( .B1(n14611), .B2(n11900), .A(n11839), .ZN(n14417) );
  INV_X1 U14437 ( .A(n14617), .ZN(n14609) );
  NAND2_X1 U14438 ( .A1(n11840), .A2(n11892), .ZN(n11842) );
  AOI22_X1 U14439 ( .A1(n11853), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11852), 
        .B2(n14380), .ZN(n11841) );
  AND2_X1 U14440 ( .A1(n11844), .A2(n11843), .ZN(n11846) );
  OR2_X1 U14441 ( .A1(n11846), .A2(n11845), .ZN(n14634) );
  INV_X1 U14442 ( .A(n14634), .ZN(n14273) );
  INV_X1 U14443 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14444 ( .A1(n11884), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11848) );
  INV_X1 U14445 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14635) );
  OR2_X1 U14446 ( .A1(n10273), .A2(n14635), .ZN(n11847) );
  OAI211_X1 U14447 ( .C1(n11849), .C2(n11902), .A(n11848), .B(n11847), .ZN(
        n11850) );
  AOI21_X1 U14448 ( .B1(n14273), .B2(n11889), .A(n11850), .ZN(n14416) );
  NAND2_X1 U14449 ( .A1(n11851), .A2(n11892), .ZN(n11855) );
  AOI22_X1 U14450 ( .A1(n11853), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11852), 
        .B2(n14376), .ZN(n11854) );
  NAND2_X1 U14451 ( .A1(n14652), .A2(n14435), .ZN(n14413) );
  NAND2_X1 U14452 ( .A1(n14415), .A2(n14413), .ZN(n14648) );
  INV_X1 U14453 ( .A(n12006), .ZN(n11873) );
  NAND4_X1 U14454 ( .A1(n11936), .A2(n11857), .A3(n11856), .A4(n15066), .ZN(
        n11858) );
  NOR2_X1 U14455 ( .A1(n11859), .A2(n11858), .ZN(n11862) );
  NAND4_X1 U14456 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11864) );
  OR4_X1 U14457 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11868) );
  NOR2_X1 U14458 ( .A1(n14791), .A2(n11868), .ZN(n11870) );
  NAND3_X1 U14459 ( .A1(n11871), .A2(n11870), .A3(n11869), .ZN(n11872) );
  NOR2_X1 U14460 ( .A1(n11873), .A2(n11872), .ZN(n11875) );
  NAND4_X1 U14461 ( .A1(n14648), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11877) );
  NOR4_X1 U14462 ( .A1(n14584), .A2(n14609), .A3(n14629), .A4(n11877), .ZN(
        n11890) );
  NAND2_X1 U14463 ( .A1(n11878), .A2(n11892), .ZN(n11880) );
  OR2_X1 U14464 ( .A1(n6676), .A2(n7478), .ZN(n11879) );
  NOR2_X1 U14465 ( .A1(n11881), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11882) );
  OR2_X1 U14466 ( .A1(n11883), .A2(n11882), .ZN(n14602) );
  INV_X1 U14467 ( .A(n14602), .ZN(n14240) );
  INV_X1 U14468 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11887) );
  NAND2_X1 U14469 ( .A1(n6675), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11886) );
  NAND2_X1 U14470 ( .A1(n11884), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11885) );
  OAI211_X1 U14471 ( .C1(n11902), .C2(n11887), .A(n11886), .B(n11885), .ZN(
        n11888) );
  AOI21_X1 U14472 ( .B1(n14240), .B2(n11889), .A(n11888), .ZN(n14441) );
  INV_X1 U14473 ( .A(n14441), .ZN(n14418) );
  XNOR2_X1 U14474 ( .A(n14440), .B(n14418), .ZN(n14599) );
  NAND4_X1 U14475 ( .A1(n14548), .A2(n14575), .A3(n11890), .A4(n14599), .ZN(
        n11891) );
  NOR3_X1 U14476 ( .A1(n14423), .A2(n14532), .A3(n11891), .ZN(n11907) );
  NAND2_X1 U14477 ( .A1(n12836), .A2(n11892), .ZN(n11895) );
  OR2_X1 U14478 ( .A1(n6676), .A2(n12839), .ZN(n11894) );
  NAND2_X1 U14479 ( .A1(n6674), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11906) );
  INV_X1 U14480 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11897) );
  OR2_X1 U14481 ( .A1(n6689), .A2(n11897), .ZN(n11905) );
  OAI21_X1 U14482 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11899), .A(n11898), 
        .ZN(n14521) );
  OR2_X1 U14483 ( .A1(n11900), .A2(n14521), .ZN(n11904) );
  INV_X1 U14484 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11901) );
  OR2_X1 U14485 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  NAND4_X1 U14486 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n14445) );
  XNOR2_X1 U14487 ( .A(n14694), .B(n14445), .ZN(n14422) );
  NAND4_X1 U14488 ( .A1(n14485), .A2(n14472), .A3(n11907), .A4(n14422), .ZN(
        n11908) );
  XOR2_X1 U14489 ( .A(n14390), .B(n11910), .Z(n12127) );
  NAND2_X1 U14490 ( .A1(n11912), .A2(n11911), .ZN(n11920) );
  INV_X1 U14491 ( .A(n11920), .ZN(n12126) );
  NAND2_X1 U14492 ( .A1(n14397), .A2(n11935), .ZN(n12116) );
  INV_X1 U14493 ( .A(n14402), .ZN(n12093) );
  INV_X1 U14494 ( .A(n14773), .ZN(n11913) );
  NAND2_X1 U14495 ( .A1(n11913), .A2(n12089), .ZN(n11914) );
  NAND2_X1 U14496 ( .A1(n11915), .A2(n11914), .ZN(n11917) );
  NAND2_X1 U14497 ( .A1(n11917), .A2(n11916), .ZN(n12121) );
  INV_X1 U14498 ( .A(n12121), .ZN(n11918) );
  NAND2_X1 U14499 ( .A1(n12093), .A2(n11918), .ZN(n11924) );
  NOR2_X1 U14500 ( .A1(n14397), .A2(n11935), .ZN(n12119) );
  XOR2_X1 U14501 ( .A(n12121), .B(n12119), .Z(n11919) );
  NAND4_X1 U14502 ( .A1(n11919), .A2(n14660), .A3(n14402), .A4(n11920), .ZN(
        n11923) );
  NAND2_X1 U14503 ( .A1(n12121), .A2(n11920), .ZN(n12118) );
  INV_X1 U14504 ( .A(n12118), .ZN(n11921) );
  NAND4_X1 U14505 ( .A1(n12116), .A2(n12093), .A3(n11921), .A4(n14397), .ZN(
        n11922) );
  OAI211_X1 U14506 ( .C1(n12116), .C2(n11924), .A(n11923), .B(n11922), .ZN(
        n12125) );
  MUX2_X1 U14507 ( .A(n14495), .B(n12830), .S(n12017), .Z(n12087) );
  INV_X1 U14508 ( .A(n12087), .ZN(n12088) );
  MUX2_X1 U14509 ( .A(n15053), .B(n14313), .S(n12097), .Z(n11962) );
  MUX2_X1 U14510 ( .A(n14314), .B(n15084), .S(n12097), .Z(n11957) );
  NAND2_X1 U14511 ( .A1(n11925), .A2(n11930), .ZN(n11926) );
  MUX2_X1 U14512 ( .A(n11927), .B(n11926), .S(n11935), .Z(n11933) );
  AND2_X1 U14513 ( .A1(n15066), .A2(n11928), .ZN(n11932) );
  MUX2_X1 U14514 ( .A(n11930), .B(n11929), .S(n11935), .Z(n11931) );
  OAI21_X1 U14515 ( .B1(n11937), .B2(n12017), .A(n11936), .ZN(n11938) );
  NAND2_X1 U14516 ( .A1(n11967), .A2(n14316), .ZN(n11943) );
  NAND2_X1 U14517 ( .A1(n12017), .A2(n11940), .ZN(n11942) );
  MUX2_X1 U14518 ( .A(n11943), .B(n11942), .S(n11941), .Z(n11944) );
  MUX2_X1 U14519 ( .A(n11947), .B(n11946), .S(n12017), .Z(n11949) );
  MUX2_X1 U14520 ( .A(n14315), .B(n15077), .S(n12017), .Z(n11948) );
  NAND2_X1 U14521 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  NAND2_X1 U14522 ( .A1(n11952), .A2(n11951), .ZN(n11956) );
  NAND2_X1 U14523 ( .A1(n11956), .A2(n11957), .ZN(n11954) );
  MUX2_X1 U14524 ( .A(n14314), .B(n15084), .S(n11967), .Z(n11953) );
  NAND2_X1 U14525 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  OAI21_X1 U14526 ( .B1(n11957), .B2(n11956), .A(n11955), .ZN(n11961) );
  NAND2_X1 U14527 ( .A1(n11961), .A2(n11962), .ZN(n11959) );
  MUX2_X1 U14528 ( .A(n15053), .B(n14313), .S(n11967), .Z(n11958) );
  NAND2_X1 U14529 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  OAI21_X1 U14530 ( .B1(n11962), .B2(n11961), .A(n11960), .ZN(n11966) );
  MUX2_X1 U14531 ( .A(n14312), .B(n11963), .S(n12097), .Z(n11965) );
  MUX2_X1 U14532 ( .A(n14312), .B(n11963), .S(n11967), .Z(n11964) );
  MUX2_X1 U14533 ( .A(n14311), .B(n15107), .S(n11967), .Z(n11971) );
  NAND2_X1 U14534 ( .A1(n11970), .A2(n11971), .ZN(n11969) );
  MUX2_X1 U14535 ( .A(n14311), .B(n15107), .S(n12097), .Z(n11968) );
  NAND2_X1 U14536 ( .A1(n11969), .A2(n11968), .ZN(n11975) );
  INV_X1 U14537 ( .A(n11971), .ZN(n11972) );
  NAND2_X1 U14538 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  MUX2_X1 U14539 ( .A(n15115), .B(n14310), .S(n11967), .Z(n11979) );
  NAND2_X1 U14540 ( .A1(n11978), .A2(n11979), .ZN(n11977) );
  MUX2_X1 U14541 ( .A(n15115), .B(n14310), .S(n12097), .Z(n11976) );
  NAND2_X1 U14542 ( .A1(n11977), .A2(n11976), .ZN(n11983) );
  INV_X1 U14543 ( .A(n11978), .ZN(n11981) );
  INV_X1 U14544 ( .A(n11979), .ZN(n11980) );
  NAND2_X1 U14545 ( .A1(n11981), .A2(n11980), .ZN(n11982) );
  MUX2_X1 U14546 ( .A(n14309), .B(n11984), .S(n11967), .Z(n11986) );
  MUX2_X1 U14547 ( .A(n14309), .B(n11984), .S(n12017), .Z(n11985) );
  INV_X1 U14548 ( .A(n11986), .ZN(n11987) );
  INV_X1 U14549 ( .A(n11967), .ZN(n12097) );
  MUX2_X1 U14550 ( .A(n14308), .B(n14986), .S(n12017), .Z(n11991) );
  NAND2_X1 U14551 ( .A1(n11990), .A2(n11991), .ZN(n11989) );
  MUX2_X1 U14552 ( .A(n14308), .B(n14986), .S(n11967), .Z(n11988) );
  NAND2_X1 U14553 ( .A1(n11989), .A2(n11988), .ZN(n11995) );
  INV_X1 U14554 ( .A(n11990), .ZN(n11993) );
  INV_X1 U14555 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14556 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  MUX2_X1 U14557 ( .A(n14307), .B(n14801), .S(n11967), .Z(n12000) );
  MUX2_X1 U14558 ( .A(n14306), .B(n14245), .S(n12097), .Z(n12004) );
  NAND2_X1 U14559 ( .A1(n12097), .A2(n14306), .ZN(n11997) );
  NAND2_X1 U14560 ( .A1(n14245), .A2(n11967), .ZN(n11996) );
  NAND3_X1 U14561 ( .A1(n12004), .A2(n11997), .A3(n11996), .ZN(n11998) );
  MUX2_X1 U14562 ( .A(n12697), .B(n7185), .S(n12097), .Z(n11999) );
  NAND2_X1 U14563 ( .A1(n12014), .A2(n12001), .ZN(n12007) );
  NAND2_X1 U14564 ( .A1(n12097), .A2(n12707), .ZN(n12002) );
  OAI21_X1 U14565 ( .B1(n14245), .B2(n12017), .A(n12002), .ZN(n12003) );
  NOR2_X1 U14566 ( .A1(n12004), .A2(n12003), .ZN(n12005) );
  AOI22_X1 U14567 ( .A1(n12007), .A2(n11967), .B1(n12006), .B2(n12005), .ZN(
        n12011) );
  NAND2_X1 U14568 ( .A1(n12013), .A2(n12008), .ZN(n12009) );
  NAND2_X1 U14569 ( .A1(n12009), .A2(n12097), .ZN(n12010) );
  MUX2_X1 U14570 ( .A(n12014), .B(n12013), .S(n11967), .Z(n12015) );
  MUX2_X1 U14571 ( .A(n14431), .B(n14940), .S(n12017), .Z(n12034) );
  NAND2_X1 U14572 ( .A1(n12034), .A2(n14435), .ZN(n12016) );
  OR2_X1 U14573 ( .A1(n14431), .A2(n11967), .ZN(n12019) );
  AOI21_X1 U14574 ( .B1(n12016), .B2(n12019), .A(n14961), .ZN(n12023) );
  NAND2_X1 U14575 ( .A1(n12034), .A2(n12737), .ZN(n12018) );
  OR2_X1 U14576 ( .A1(n14940), .A2(n12097), .ZN(n12026) );
  AOI21_X1 U14577 ( .B1(n12018), .B2(n12026), .A(n14652), .ZN(n12022) );
  NAND2_X1 U14578 ( .A1(n14435), .A2(n11967), .ZN(n12027) );
  OR2_X1 U14579 ( .A1(n14940), .A2(n12027), .ZN(n12021) );
  INV_X1 U14580 ( .A(n12019), .ZN(n12030) );
  NAND2_X1 U14581 ( .A1(n12030), .A2(n12737), .ZN(n12020) );
  NAND2_X1 U14582 ( .A1(n12021), .A2(n12020), .ZN(n12033) );
  OR3_X1 U14583 ( .A1(n12023), .A2(n12022), .A3(n12033), .ZN(n12024) );
  NAND2_X1 U14584 ( .A1(n12025), .A2(n12024), .ZN(n12040) );
  INV_X1 U14585 ( .A(n12026), .ZN(n12029) );
  INV_X1 U14586 ( .A(n12027), .ZN(n12028) );
  AOI21_X1 U14587 ( .B1(n12034), .B2(n12029), .A(n12028), .ZN(n12037) );
  NAND2_X1 U14588 ( .A1(n12034), .A2(n12030), .ZN(n12031) );
  OAI21_X1 U14589 ( .B1(n11967), .B2(n14435), .A(n12031), .ZN(n12032) );
  NAND2_X1 U14590 ( .A1(n12032), .A2(n14652), .ZN(n12036) );
  NAND2_X1 U14591 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  OAI211_X1 U14592 ( .C1(n12037), .C2(n14652), .A(n12036), .B(n12035), .ZN(
        n12038) );
  NOR2_X1 U14593 ( .A1(n14629), .A2(n12038), .ZN(n12039) );
  NAND3_X1 U14594 ( .A1(n14638), .A2(n14416), .A3(n11967), .ZN(n12042) );
  OR3_X1 U14595 ( .A1(n14638), .A2(n14416), .A3(n11967), .ZN(n12041) );
  NAND2_X1 U14596 ( .A1(n12042), .A2(n12041), .ZN(n12043) );
  NAND2_X1 U14597 ( .A1(n14617), .A2(n12043), .ZN(n12047) );
  INV_X1 U14598 ( .A(n14417), .ZN(n12044) );
  OR2_X1 U14599 ( .A1(n14728), .A2(n12044), .ZN(n12045) );
  NAND2_X1 U14600 ( .A1(n14728), .A2(n12044), .ZN(n14439) );
  MUX2_X1 U14601 ( .A(n12045), .B(n14439), .S(n11967), .Z(n12046) );
  MUX2_X1 U14602 ( .A(n14441), .B(n14722), .S(n12017), .Z(n12049) );
  MUX2_X1 U14603 ( .A(n14418), .B(n14440), .S(n11967), .Z(n12048) );
  MUX2_X1 U14604 ( .A(n14564), .B(n14590), .S(n11967), .Z(n12053) );
  NAND2_X1 U14605 ( .A1(n12052), .A2(n12053), .ZN(n12051) );
  MUX2_X1 U14606 ( .A(n14564), .B(n14590), .S(n12017), .Z(n12050) );
  NAND2_X1 U14607 ( .A1(n12051), .A2(n12050), .ZN(n12057) );
  INV_X1 U14608 ( .A(n12053), .ZN(n12054) );
  NAND2_X1 U14609 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  MUX2_X1 U14610 ( .A(n14420), .B(n14711), .S(n12017), .Z(n12061) );
  NAND2_X1 U14611 ( .A1(n12060), .A2(n12061), .ZN(n12059) );
  MUX2_X1 U14612 ( .A(n14420), .B(n14711), .S(n11967), .Z(n12058) );
  NAND2_X1 U14613 ( .A1(n12059), .A2(n12058), .ZN(n12065) );
  INV_X1 U14614 ( .A(n12060), .ZN(n12063) );
  INV_X1 U14615 ( .A(n12061), .ZN(n12062) );
  MUX2_X1 U14616 ( .A(n14566), .B(n14557), .S(n11967), .Z(n12067) );
  MUX2_X1 U14617 ( .A(n14566), .B(n14557), .S(n12097), .Z(n12066) );
  MUX2_X1 U14618 ( .A(n14303), .B(n6677), .S(n12097), .Z(n12071) );
  NAND2_X1 U14619 ( .A1(n12070), .A2(n12071), .ZN(n12069) );
  MUX2_X1 U14620 ( .A(n14303), .B(n6677), .S(n11967), .Z(n12068) );
  NAND2_X1 U14621 ( .A1(n12069), .A2(n12068), .ZN(n12075) );
  INV_X1 U14622 ( .A(n12070), .ZN(n12073) );
  INV_X1 U14623 ( .A(n12071), .ZN(n12072) );
  NAND2_X1 U14624 ( .A1(n12075), .A2(n12074), .ZN(n12078) );
  MUX2_X1 U14625 ( .A(n14445), .B(n14694), .S(n11967), .Z(n12079) );
  NAND2_X1 U14626 ( .A1(n12078), .A2(n12079), .ZN(n12077) );
  MUX2_X1 U14627 ( .A(n14445), .B(n14694), .S(n12017), .Z(n12076) );
  NAND2_X1 U14628 ( .A1(n12077), .A2(n12076), .ZN(n12083) );
  INV_X1 U14629 ( .A(n12078), .ZN(n12081) );
  INV_X1 U14630 ( .A(n12079), .ZN(n12080) );
  NAND2_X1 U14631 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  MUX2_X1 U14632 ( .A(n14424), .B(n14688), .S(n12097), .Z(n12084) );
  MUX2_X1 U14633 ( .A(n14688), .B(n14424), .S(n12017), .Z(n12085) );
  INV_X1 U14634 ( .A(n14495), .ZN(n14681) );
  MUX2_X1 U14635 ( .A(n14426), .B(n14681), .S(n12097), .Z(n12086) );
  INV_X1 U14636 ( .A(n12100), .ZN(n12104) );
  INV_X1 U14637 ( .A(n14461), .ZN(n14427) );
  MUX2_X1 U14638 ( .A(n14427), .B(n14674), .S(n12017), .Z(n12099) );
  INV_X1 U14639 ( .A(n12099), .ZN(n12103) );
  OAI21_X1 U14640 ( .B1(n14402), .B2(n12089), .A(n14457), .ZN(n12090) );
  MUX2_X1 U14641 ( .A(n12090), .B(n14663), .S(n11935), .Z(n12107) );
  NAND2_X1 U14642 ( .A1(n14396), .A2(n12097), .ZN(n12096) );
  OAI22_X1 U14643 ( .A1(n12017), .A2(n12093), .B1(n12092), .B2(n12091), .ZN(
        n12094) );
  NAND2_X1 U14644 ( .A1(n12094), .A2(n14457), .ZN(n12095) );
  NAND2_X1 U14645 ( .A1(n12096), .A2(n12095), .ZN(n12112) );
  MUX2_X1 U14646 ( .A(n12831), .B(n14666), .S(n11967), .Z(n12106) );
  INV_X1 U14647 ( .A(n14666), .ZN(n14455) );
  MUX2_X1 U14648 ( .A(n14302), .B(n14455), .S(n12097), .Z(n12105) );
  MUX2_X1 U14649 ( .A(n14479), .B(n14461), .S(n12097), .Z(n12098) );
  AOI21_X1 U14650 ( .B1(n12100), .B2(n12099), .A(n12098), .ZN(n12101) );
  INV_X1 U14651 ( .A(n12112), .ZN(n12109) );
  NAND2_X1 U14652 ( .A1(n12106), .A2(n12105), .ZN(n12111) );
  INV_X1 U14653 ( .A(n12107), .ZN(n12108) );
  AOI21_X1 U14654 ( .B1(n12109), .B2(n12111), .A(n12108), .ZN(n12110) );
  INV_X1 U14655 ( .A(n12111), .ZN(n12113) );
  NOR2_X1 U14656 ( .A1(n12116), .A2(n14402), .ZN(n12117) );
  AOI211_X1 U14657 ( .C1(n12119), .C2(n14402), .A(n12118), .B(n12117), .ZN(
        n12120) );
  NOR2_X1 U14658 ( .A1(n12122), .A2(n12121), .ZN(n12123) );
  NAND3_X1 U14659 ( .A1(n12129), .A2(n12128), .A3(n14563), .ZN(n12130) );
  OAI211_X1 U14660 ( .C1(n14773), .C2(n12132), .A(n12130), .B(P1_B_REG_SCAN_IN), .ZN(n12131) );
  INV_X1 U14661 ( .A(n12133), .ZN(n14142) );
  OAI222_X1 U14662 ( .A1(n14771), .A2(n12134), .B1(n14768), .B2(n14142), .C1(
        P1_U3086), .C2(n6679), .ZN(P1_U3328) );
  NAND3_X1 U14663 ( .A1(n12135), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n12139) );
  NAND2_X1 U14664 ( .A1(n14759), .A2(n12136), .ZN(n12138) );
  NAND2_X1 U14665 ( .A1(n14138), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12137) );
  OAI211_X1 U14666 ( .C1(n12140), .C2(n12139), .A(n12138), .B(n12137), .ZN(
        P2_U3296) );
  INV_X1 U14667 ( .A(n12141), .ZN(n12142) );
  INV_X1 U14668 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12683) );
  OAI22_X1 U14669 ( .A1(n12143), .A2(n12142), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n12683), .ZN(n12149) );
  XNOR2_X1 U14670 ( .A(n12144), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12148) );
  XNOR2_X1 U14671 ( .A(n12149), .B(n12148), .ZN(n13458) );
  NAND2_X1 U14672 ( .A1(n13458), .A2(n7160), .ZN(n12146) );
  OR2_X1 U14673 ( .A1(n12152), .A2(n13460), .ZN(n12145) );
  INV_X1 U14674 ( .A(n12156), .ZN(n13396) );
  AND2_X1 U14675 ( .A1(n13396), .A2(n12147), .ZN(n12161) );
  OAI22_X1 U14676 ( .A1(n12149), .A2(n12148), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14761), .ZN(n12151) );
  XNOR2_X1 U14677 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12150) );
  XNOR2_X1 U14678 ( .A(n12151), .B(n12150), .ZN(n13456) );
  INV_X1 U14679 ( .A(SI_31_), .ZN(n13451) );
  NOR2_X1 U14680 ( .A1(n12152), .A2(n13451), .ZN(n12153) );
  INV_X1 U14681 ( .A(n13393), .ZN(n12160) );
  INV_X1 U14682 ( .A(n13116), .ZN(n12155) );
  AND2_X1 U14683 ( .A1(n13393), .A2(n13116), .ZN(n12351) );
  NAND2_X1 U14684 ( .A1(n12156), .A2(n12154), .ZN(n12317) );
  NAND2_X1 U14685 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  NAND3_X1 U14686 ( .A1(n12317), .A2(n12310), .A3(n12157), .ZN(n12158) );
  INV_X1 U14687 ( .A(n12161), .ZN(n12318) );
  NAND2_X1 U14688 ( .A1(n12318), .A2(n12317), .ZN(n12348) );
  INV_X1 U14689 ( .A(n12348), .ZN(n12305) );
  NOR2_X1 U14690 ( .A1(n12313), .A2(n12922), .ZN(n12347) );
  MUX2_X1 U14691 ( .A(n12163), .B(n12162), .S(n12320), .Z(n12164) );
  NAND2_X1 U14692 ( .A1(n13247), .A2(n13257), .ZN(n12166) );
  MUX2_X1 U14693 ( .A(n12166), .B(n12165), .S(n12292), .Z(n12167) );
  INV_X1 U14694 ( .A(n12167), .ZN(n12280) );
  NAND2_X1 U14695 ( .A1(n12210), .A2(n12168), .ZN(n12169) );
  NAND2_X1 U14696 ( .A1(n12169), .A2(n12320), .ZN(n12203) );
  INV_X1 U14697 ( .A(n12203), .ZN(n12211) );
  AND2_X1 U14698 ( .A1(n15652), .A2(n12170), .ZN(n12325) );
  INV_X1 U14699 ( .A(n12325), .ZN(n12172) );
  NAND2_X1 U14700 ( .A1(n12172), .A2(n12359), .ZN(n12175) );
  NAND2_X1 U14701 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  NAND3_X1 U14702 ( .A1(n12179), .A2(n12292), .A3(n12173), .ZN(n12174) );
  OAI21_X1 U14703 ( .B1(n15658), .B2(n12175), .A(n12174), .ZN(n12178) );
  NAND2_X1 U14704 ( .A1(n15651), .A2(n12176), .ZN(n12177) );
  NAND2_X1 U14705 ( .A1(n12178), .A2(n12177), .ZN(n12182) );
  MUX2_X1 U14706 ( .A(n12180), .B(n12179), .S(n12320), .Z(n12181) );
  NAND3_X1 U14707 ( .A1(n12182), .A2(n15640), .A3(n12181), .ZN(n12189) );
  NAND2_X1 U14708 ( .A1(n12191), .A2(n12183), .ZN(n12186) );
  NAND2_X1 U14709 ( .A1(n12190), .A2(n12184), .ZN(n12185) );
  MUX2_X1 U14710 ( .A(n12186), .B(n12185), .S(n12292), .Z(n12187) );
  INV_X1 U14711 ( .A(n12187), .ZN(n12188) );
  NAND2_X1 U14712 ( .A1(n12189), .A2(n12188), .ZN(n12193) );
  MUX2_X1 U14713 ( .A(n12191), .B(n12190), .S(n12320), .Z(n12192) );
  NAND3_X1 U14714 ( .A1(n12193), .A2(n12328), .A3(n12192), .ZN(n12197) );
  MUX2_X1 U14715 ( .A(n12195), .B(n12194), .S(n12292), .Z(n12196) );
  NAND3_X1 U14716 ( .A1(n12197), .A2(n15607), .A3(n12196), .ZN(n12204) );
  NAND2_X1 U14717 ( .A1(n12199), .A2(n12198), .ZN(n12200) );
  NAND2_X1 U14718 ( .A1(n12205), .A2(n12200), .ZN(n12201) );
  NAND2_X1 U14719 ( .A1(n12201), .A2(n12292), .ZN(n12202) );
  NAND3_X1 U14720 ( .A1(n12204), .A2(n12203), .A3(n12202), .ZN(n12209) );
  NOR2_X1 U14721 ( .A1(n12205), .A2(n12292), .ZN(n12206) );
  NOR2_X1 U14722 ( .A1(n12207), .A2(n12206), .ZN(n12208) );
  OAI211_X1 U14723 ( .C1(n12211), .C2(n12210), .A(n12209), .B(n12208), .ZN(
        n12215) );
  MUX2_X1 U14724 ( .A(n12213), .B(n12212), .S(n12320), .Z(n12214) );
  NAND3_X1 U14725 ( .A1(n12215), .A2(n15601), .A3(n12214), .ZN(n12222) );
  NAND2_X1 U14726 ( .A1(n12216), .A2(n12320), .ZN(n12220) );
  NAND2_X1 U14727 ( .A1(n12217), .A2(n12292), .ZN(n12219) );
  MUX2_X1 U14728 ( .A(n12220), .B(n12219), .S(n12218), .Z(n12221) );
  NAND3_X1 U14729 ( .A1(n12222), .A2(n12332), .A3(n12221), .ZN(n12228) );
  INV_X1 U14730 ( .A(n12223), .ZN(n12224) );
  MUX2_X1 U14731 ( .A(n12225), .B(n12224), .S(n12320), .Z(n12227) );
  AOI21_X1 U14732 ( .B1(n12228), .B2(n12227), .A(n12226), .ZN(n12235) );
  MUX2_X1 U14733 ( .A(n12230), .B(n12229), .S(n12320), .Z(n12231) );
  NAND2_X1 U14734 ( .A1(n12231), .A2(n12335), .ZN(n12234) );
  AND2_X1 U14735 ( .A1(n12240), .A2(n12232), .ZN(n12233) );
  OAI22_X1 U14736 ( .A1(n12235), .A2(n12234), .B1(n12320), .B2(n12233), .ZN(
        n12239) );
  AOI21_X1 U14737 ( .B1(n12238), .B2(n12236), .A(n12292), .ZN(n12237) );
  AOI21_X1 U14738 ( .B1(n12239), .B2(n12238), .A(n12237), .ZN(n12242) );
  NOR2_X1 U14739 ( .A1(n12240), .A2(n12292), .ZN(n12241) );
  OAI211_X1 U14740 ( .C1(n12242), .C2(n12241), .A(n12340), .B(n6705), .ZN(
        n12256) );
  NAND2_X1 U14741 ( .A1(n12259), .A2(n12243), .ZN(n12247) );
  OR2_X1 U14742 ( .A1(n12247), .A2(n12244), .ZN(n12245) );
  MUX2_X1 U14743 ( .A(n12246), .B(n12245), .S(n12320), .Z(n12253) );
  NAND2_X1 U14744 ( .A1(n12247), .A2(n12320), .ZN(n12254) );
  MUX2_X1 U14745 ( .A(n12249), .B(n12248), .S(n12292), .Z(n12250) );
  INV_X1 U14746 ( .A(n12250), .ZN(n12251) );
  NAND3_X1 U14747 ( .A1(n12254), .A2(n12340), .A3(n12251), .ZN(n12252) );
  NAND2_X1 U14748 ( .A1(n12253), .A2(n12252), .ZN(n12255) );
  INV_X1 U14749 ( .A(n13316), .ZN(n13312) );
  AOI22_X1 U14750 ( .A1(n12256), .A2(n12255), .B1(n13312), .B2(n12254), .ZN(
        n12262) );
  AOI21_X1 U14751 ( .B1(n12258), .B2(n12257), .A(n12320), .ZN(n12261) );
  MUX2_X1 U14752 ( .A(n12259), .B(n12258), .S(n12320), .Z(n12260) );
  OAI21_X1 U14753 ( .B1(n12262), .B2(n12261), .A(n12260), .ZN(n12263) );
  NAND3_X1 U14754 ( .A1(n12263), .A2(n13276), .A3(n13291), .ZN(n12274) );
  INV_X1 U14755 ( .A(n12268), .ZN(n12266) );
  OAI211_X1 U14756 ( .C1(n12266), .C2(n12265), .A(n12275), .B(n12264), .ZN(
        n12271) );
  NAND2_X1 U14757 ( .A1(n13276), .A2(n12267), .ZN(n12269) );
  NAND3_X1 U14758 ( .A1(n12269), .A2(n12276), .A3(n12268), .ZN(n12270) );
  MUX2_X1 U14759 ( .A(n12271), .B(n12270), .S(n12292), .Z(n12272) );
  INV_X1 U14760 ( .A(n12272), .ZN(n12273) );
  NAND2_X1 U14761 ( .A1(n12274), .A2(n12273), .ZN(n12278) );
  MUX2_X1 U14762 ( .A(n12276), .B(n12275), .S(n12292), .Z(n12277) );
  AOI21_X1 U14763 ( .B1(n12278), .B2(n12277), .A(n13241), .ZN(n12279) );
  OR3_X1 U14764 ( .A1(n12280), .A2(n13231), .A3(n12279), .ZN(n12284) );
  MUX2_X1 U14765 ( .A(n12282), .B(n12281), .S(n12320), .Z(n12283) );
  NAND2_X1 U14766 ( .A1(n12284), .A2(n12283), .ZN(n12288) );
  INV_X1 U14767 ( .A(n13214), .ZN(n13218) );
  MUX2_X1 U14768 ( .A(n12286), .B(n12285), .S(n12292), .Z(n12287) );
  OAI21_X1 U14769 ( .B1(n12288), .B2(n13218), .A(n12287), .ZN(n12290) );
  AND2_X1 U14770 ( .A1(n13217), .A2(n12320), .ZN(n12289) );
  AOI22_X1 U14771 ( .A1(n13204), .A2(n12290), .B1(n12289), .B2(n13209), .ZN(
        n12297) );
  INV_X1 U14772 ( .A(n12291), .ZN(n12295) );
  XNOR2_X1 U14773 ( .A(n12293), .B(n12292), .ZN(n12294) );
  OAI21_X1 U14774 ( .B1(n13184), .B2(n12295), .A(n12294), .ZN(n12296) );
  OAI211_X1 U14775 ( .C1(n13184), .C2(n12297), .A(n13173), .B(n12296), .ZN(
        n12298) );
  INV_X1 U14776 ( .A(n12299), .ZN(n12300) );
  MUX2_X1 U14777 ( .A(n12301), .B(n12300), .S(n12320), .Z(n12302) );
  INV_X1 U14778 ( .A(n12302), .ZN(n12303) );
  OR2_X1 U14779 ( .A1(n12307), .A2(n12306), .ZN(n12308) );
  OAI21_X1 U14780 ( .B1(n13141), .B2(n12922), .A(n12308), .ZN(n12309) );
  MUX2_X1 U14781 ( .A(n12309), .B(n12308), .S(n12320), .Z(n12314) );
  MUX2_X1 U14782 ( .A(n12311), .B(n12310), .S(n12320), .Z(n12312) );
  NAND2_X1 U14783 ( .A1(n12324), .A2(n12323), .ZN(n12356) );
  NOR2_X1 U14784 ( .A1(n15651), .A2(n12325), .ZN(n15428) );
  NAND4_X1 U14785 ( .A1(n15428), .A2(n12327), .A3(n15628), .A4(n12326), .ZN(
        n12331) );
  INV_X1 U14786 ( .A(n15658), .ZN(n12329) );
  NAND3_X1 U14787 ( .A1(n15640), .A2(n12329), .A3(n12328), .ZN(n12330) );
  NOR2_X1 U14788 ( .A1(n12331), .A2(n12330), .ZN(n12336) );
  AND3_X1 U14789 ( .A1(n15607), .A2(n12332), .A3(n15601), .ZN(n12333) );
  NAND4_X1 U14790 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12338) );
  NOR2_X1 U14791 ( .A1(n12338), .A2(n12337), .ZN(n12339) );
  NAND3_X1 U14792 ( .A1(n12340), .A2(n6705), .A3(n12339), .ZN(n12341) );
  NOR2_X1 U14793 ( .A1(n13298), .A2(n12341), .ZN(n12342) );
  NAND4_X1 U14794 ( .A1(n13276), .A2(n13316), .A3(n13291), .A4(n12342), .ZN(
        n12343) );
  NOR4_X1 U14795 ( .A1(n13231), .A2(n13241), .A3(n13261), .A4(n12343), .ZN(
        n12344) );
  NAND4_X1 U14796 ( .A1(n13173), .A2(n13204), .A3(n13214), .A4(n12344), .ZN(
        n12345) );
  NOR4_X1 U14797 ( .A1(n13141), .A2(n13155), .A3(n12345), .A4(n13184), .ZN(
        n12346) );
  NAND2_X1 U14798 ( .A1(n12347), .A2(n12346), .ZN(n12349) );
  NOR4_X1 U14799 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  XNOR2_X1 U14800 ( .A(n12352), .B(n13058), .ZN(n12354) );
  NOR2_X1 U14801 ( .A1(n12358), .A2(n13469), .ZN(n12361) );
  OAI21_X1 U14802 ( .B1(n12362), .B2(n12359), .A(P3_B_REG_SCAN_IN), .ZN(n12360) );
  OAI22_X1 U14803 ( .A1(n13842), .A2(n12655), .B1(n13664), .B2(n12584), .ZN(
        n12548) );
  NAND2_X1 U14804 ( .A1(n13704), .A2(n12368), .ZN(n12364) );
  NAND2_X1 U14805 ( .A1(n12368), .A2(n13705), .ZN(n12366) );
  OAI21_X1 U14806 ( .B1(n13705), .B2(n12367), .A(n12366), .ZN(n12373) );
  AND2_X1 U14807 ( .A1(n13705), .A2(n15291), .ZN(n12371) );
  INV_X1 U14808 ( .A(n7652), .ZN(n12369) );
  OAI21_X1 U14809 ( .B1(n7651), .B2(n13759), .A(n12369), .ZN(n12370) );
  INV_X1 U14810 ( .A(n12375), .ZN(n12378) );
  NAND2_X1 U14811 ( .A1(n12378), .A2(n12377), .ZN(n12379) );
  NAND2_X1 U14812 ( .A1(n12383), .A2(n13703), .ZN(n12382) );
  NAND2_X1 U14813 ( .A1(n12580), .A2(n15282), .ZN(n12381) );
  NAND2_X1 U14814 ( .A1(n12382), .A2(n12381), .ZN(n12385) );
  AOI22_X1 U14815 ( .A1(n12383), .A2(n15282), .B1(n13703), .B2(n12655), .ZN(
        n12384) );
  NAND2_X1 U14816 ( .A1(n12560), .A2(n12387), .ZN(n12389) );
  NAND2_X1 U14817 ( .A1(n13702), .A2(n6673), .ZN(n12388) );
  NAND2_X1 U14818 ( .A1(n12389), .A2(n12388), .ZN(n12394) );
  NAND2_X1 U14819 ( .A1(n12393), .A2(n12394), .ZN(n12392) );
  NAND2_X1 U14820 ( .A1(n12392), .A2(n12391), .ZN(n12398) );
  INV_X1 U14821 ( .A(n12393), .ZN(n12396) );
  INV_X1 U14822 ( .A(n12394), .ZN(n12395) );
  NAND2_X1 U14823 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  NAND2_X1 U14824 ( .A1(n12401), .A2(n6673), .ZN(n12400) );
  NAND2_X1 U14825 ( .A1(n12585), .A2(n13701), .ZN(n12399) );
  NAND2_X1 U14826 ( .A1(n12400), .A2(n12399), .ZN(n12403) );
  AOI22_X1 U14827 ( .A1(n12401), .A2(n12560), .B1(n13701), .B2(n6673), .ZN(
        n12402) );
  NAND2_X1 U14828 ( .A1(n15377), .A2(n12584), .ZN(n12406) );
  NAND2_X1 U14829 ( .A1(n13700), .A2(n6673), .ZN(n12405) );
  NAND2_X1 U14830 ( .A1(n12406), .A2(n12405), .ZN(n12408) );
  AOI22_X1 U14831 ( .A1(n15377), .A2(n6673), .B1(n12584), .B2(n13700), .ZN(
        n12407) );
  NAND2_X1 U14832 ( .A1(n12411), .A2(n12575), .ZN(n12410) );
  NAND2_X1 U14833 ( .A1(n12584), .A2(n13699), .ZN(n12409) );
  NAND2_X1 U14834 ( .A1(n12410), .A2(n12409), .ZN(n12417) );
  NAND2_X1 U14835 ( .A1(n12411), .A2(n12584), .ZN(n12412) );
  OAI21_X1 U14836 ( .B1(n12413), .B2(n12584), .A(n12412), .ZN(n12414) );
  NAND2_X1 U14837 ( .A1(n12415), .A2(n12414), .ZN(n12421) );
  NAND2_X1 U14838 ( .A1(n12419), .A2(n12418), .ZN(n12420) );
  NAND2_X1 U14839 ( .A1(n12424), .A2(n12584), .ZN(n12423) );
  NAND2_X1 U14840 ( .A1(n13698), .A2(n12575), .ZN(n12422) );
  AOI22_X1 U14841 ( .A1(n12424), .A2(n12575), .B1(n12584), .B2(n13698), .ZN(
        n12425) );
  NAND2_X1 U14842 ( .A1(n12428), .A2(n12655), .ZN(n12427) );
  NAND2_X1 U14843 ( .A1(n12584), .A2(n13697), .ZN(n12426) );
  NAND2_X1 U14844 ( .A1(n12427), .A2(n12426), .ZN(n12434) );
  NAND2_X1 U14845 ( .A1(n12428), .A2(n12584), .ZN(n12429) );
  OAI21_X1 U14846 ( .B1(n12430), .B2(n12585), .A(n12429), .ZN(n12431) );
  NAND2_X1 U14847 ( .A1(n12432), .A2(n12431), .ZN(n12438) );
  NAND2_X1 U14848 ( .A1(n12436), .A2(n12435), .ZN(n12437) );
  NAND2_X1 U14849 ( .A1(n12441), .A2(n12584), .ZN(n12440) );
  NAND2_X1 U14850 ( .A1(n13695), .A2(n6673), .ZN(n12439) );
  NAND2_X1 U14851 ( .A1(n12440), .A2(n12439), .ZN(n12446) );
  NAND2_X1 U14852 ( .A1(n12445), .A2(n12446), .ZN(n12444) );
  AOI22_X1 U14853 ( .A1(n12441), .A2(n12575), .B1(n12584), .B2(n13695), .ZN(
        n12442) );
  INV_X1 U14854 ( .A(n12442), .ZN(n12443) );
  NAND2_X1 U14855 ( .A1(n12444), .A2(n12443), .ZN(n12450) );
  INV_X1 U14856 ( .A(n12445), .ZN(n12448) );
  INV_X1 U14857 ( .A(n12446), .ZN(n12447) );
  NAND2_X1 U14858 ( .A1(n12448), .A2(n12447), .ZN(n12449) );
  NAND2_X1 U14859 ( .A1(n15393), .A2(n12655), .ZN(n12452) );
  NAND2_X1 U14860 ( .A1(n12584), .A2(n13694), .ZN(n12451) );
  NAND2_X1 U14861 ( .A1(n12452), .A2(n12451), .ZN(n12456) );
  NAND2_X1 U14862 ( .A1(n15393), .A2(n12584), .ZN(n12453) );
  OAI21_X1 U14863 ( .B1(n12454), .B2(n12560), .A(n12453), .ZN(n12455) );
  NAND2_X1 U14864 ( .A1(n12459), .A2(n12584), .ZN(n12458) );
  NAND2_X1 U14865 ( .A1(n13693), .A2(n12575), .ZN(n12457) );
  NAND2_X1 U14866 ( .A1(n12458), .A2(n12457), .ZN(n12462) );
  AOI22_X1 U14867 ( .A1(n12459), .A2(n12575), .B1(n12584), .B2(n13693), .ZN(
        n12460) );
  NAND2_X1 U14868 ( .A1(n14912), .A2(n12655), .ZN(n12465) );
  NAND2_X1 U14869 ( .A1(n12584), .A2(n13692), .ZN(n12464) );
  NAND2_X1 U14870 ( .A1(n12465), .A2(n12464), .ZN(n12467) );
  AOI22_X1 U14871 ( .A1(n14912), .A2(n12584), .B1(n13692), .B2(n12575), .ZN(
        n12466) );
  NAND2_X1 U14872 ( .A1(n12470), .A2(n12585), .ZN(n12469) );
  NAND2_X1 U14873 ( .A1(n13691), .A2(n6673), .ZN(n12468) );
  NAND2_X1 U14874 ( .A1(n12469), .A2(n12468), .ZN(n12476) );
  NAND2_X1 U14875 ( .A1(n12475), .A2(n12476), .ZN(n12474) );
  NAND2_X1 U14876 ( .A1(n12470), .A2(n6673), .ZN(n12471) );
  NAND2_X1 U14877 ( .A1(n12474), .A2(n12473), .ZN(n12480) );
  NAND2_X1 U14878 ( .A1(n12478), .A2(n12477), .ZN(n12479) );
  NAND2_X1 U14879 ( .A1(n12483), .A2(n12655), .ZN(n12482) );
  NAND2_X1 U14880 ( .A1(n12584), .A2(n13690), .ZN(n12481) );
  NAND2_X1 U14881 ( .A1(n12482), .A2(n12481), .ZN(n12486) );
  AOI22_X1 U14882 ( .A1(n12483), .A2(n12585), .B1(n13690), .B2(n12575), .ZN(
        n12484) );
  NAND2_X1 U14883 ( .A1(n14089), .A2(n12584), .ZN(n12489) );
  NAND2_X1 U14884 ( .A1(n13992), .A2(n12575), .ZN(n12488) );
  NAND2_X1 U14885 ( .A1(n12489), .A2(n12488), .ZN(n12494) );
  AND2_X1 U14886 ( .A1(n13689), .A2(n12584), .ZN(n12490) );
  AOI21_X1 U14887 ( .B1(n14084), .B2(n12575), .A(n12490), .ZN(n12498) );
  NAND2_X1 U14888 ( .A1(n14084), .A2(n12585), .ZN(n12492) );
  NAND2_X1 U14889 ( .A1(n13689), .A2(n6673), .ZN(n12491) );
  NAND2_X1 U14890 ( .A1(n12492), .A2(n12491), .ZN(n12497) );
  AOI22_X1 U14891 ( .A1(n14089), .A2(n12575), .B1(n12584), .B2(n13992), .ZN(
        n12493) );
  AOI22_X1 U14892 ( .A1(n14079), .A2(n12575), .B1(n12585), .B2(n13989), .ZN(
        n12499) );
  NAND2_X1 U14893 ( .A1(n14079), .A2(n12584), .ZN(n12496) );
  NAND2_X1 U14894 ( .A1(n13989), .A2(n12575), .ZN(n12495) );
  NAND2_X1 U14895 ( .A1(n12496), .A2(n12495), .ZN(n12502) );
  AOI22_X1 U14896 ( .A1(n12499), .A2(n12502), .B1(n12498), .B2(n12497), .ZN(
        n12500) );
  NOR2_X1 U14897 ( .A1(n14079), .A2(n13989), .ZN(n12501) );
  OR2_X1 U14898 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  NAND2_X1 U14899 ( .A1(n13961), .A2(n12575), .ZN(n12505) );
  NAND2_X1 U14900 ( .A1(n13939), .A2(n12560), .ZN(n12504) );
  NAND2_X1 U14901 ( .A1(n12505), .A2(n12504), .ZN(n12507) );
  AOI22_X1 U14902 ( .A1(n13961), .A2(n12584), .B1(n13939), .B2(n12575), .ZN(
        n12506) );
  NAND2_X1 U14903 ( .A1(n13934), .A2(n12585), .ZN(n12510) );
  NAND2_X1 U14904 ( .A1(n13920), .A2(n6673), .ZN(n12509) );
  NAND2_X1 U14905 ( .A1(n12510), .A2(n12509), .ZN(n12512) );
  AOI22_X1 U14906 ( .A1(n13934), .A2(n12575), .B1(n12584), .B2(n13920), .ZN(
        n12511) );
  NAND2_X1 U14907 ( .A1(n14063), .A2(n12575), .ZN(n12515) );
  NAND2_X1 U14908 ( .A1(n13940), .A2(n12585), .ZN(n12514) );
  NAND2_X1 U14909 ( .A1(n12515), .A2(n12514), .ZN(n12517) );
  AOI22_X1 U14910 ( .A1(n14063), .A2(n12584), .B1(n13940), .B2(n12575), .ZN(
        n12516) );
  NOR2_X1 U14911 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  NAND2_X1 U14912 ( .A1(n14120), .A2(n12584), .ZN(n12521) );
  NAND2_X1 U14913 ( .A1(n13919), .A2(n12575), .ZN(n12520) );
  NAND2_X1 U14914 ( .A1(n12521), .A2(n12520), .ZN(n12523) );
  AOI22_X1 U14915 ( .A1(n14120), .A2(n12575), .B1(n12560), .B2(n13919), .ZN(
        n12522) );
  NAND2_X1 U14916 ( .A1(n14118), .A2(n6673), .ZN(n12526) );
  NAND2_X1 U14917 ( .A1(n13688), .A2(n12585), .ZN(n12525) );
  NAND2_X1 U14918 ( .A1(n12526), .A2(n12525), .ZN(n12529) );
  NAND2_X1 U14919 ( .A1(n14118), .A2(n12560), .ZN(n12527) );
  OAI21_X1 U14920 ( .B1(n13534), .B2(n12584), .A(n12527), .ZN(n12528) );
  INV_X1 U14921 ( .A(n12528), .ZN(n12532) );
  NAND2_X1 U14922 ( .A1(n14045), .A2(n12585), .ZN(n12535) );
  NAND2_X1 U14923 ( .A1(n13687), .A2(n6673), .ZN(n12534) );
  NAND2_X1 U14924 ( .A1(n12535), .A2(n12534), .ZN(n12537) );
  NOR2_X1 U14925 ( .A1(n12538), .A2(n12537), .ZN(n12540) );
  AOI22_X1 U14926 ( .A1(n14045), .A2(n12575), .B1(n12584), .B2(n13687), .ZN(
        n12536) );
  AOI21_X1 U14927 ( .B1(n12538), .B2(n12537), .A(n12536), .ZN(n12539) );
  AOI22_X1 U14928 ( .A1(n14039), .A2(n12575), .B1(n12585), .B2(n13686), .ZN(
        n12543) );
  AOI22_X1 U14929 ( .A1(n14039), .A2(n12584), .B1(n13686), .B2(n12575), .ZN(
        n12541) );
  INV_X1 U14930 ( .A(n12541), .ZN(n12542) );
  AOI22_X1 U14931 ( .A1(n14034), .A2(n12575), .B1(n12585), .B2(n13685), .ZN(
        n12547) );
  AOI22_X1 U14932 ( .A1(n14111), .A2(n12575), .B1(n12560), .B2(n13684), .ZN(
        n12550) );
  AOI22_X1 U14933 ( .A1(n14111), .A2(n12560), .B1(n13684), .B2(n12575), .ZN(
        n12551) );
  NAND2_X1 U14934 ( .A1(n14759), .A2(n12576), .ZN(n12553) );
  NAND2_X1 U14935 ( .A1(n6687), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12552) );
  INV_X1 U14936 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14095) );
  NAND2_X1 U14937 ( .A1(n12554), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U14938 ( .A1(n8204), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12555) );
  OAI211_X1 U14939 ( .C1(n12557), .C2(n14095), .A(n12556), .B(n12555), .ZN(
        n13680) );
  XNOR2_X1 U14940 ( .A(n13765), .B(n13680), .ZN(n12645) );
  AND2_X1 U14941 ( .A1(n13682), .A2(n12575), .ZN(n12558) );
  AOI21_X1 U14942 ( .B1(n12559), .B2(n12585), .A(n12558), .ZN(n12589) );
  NAND2_X1 U14943 ( .A1(n12559), .A2(n12575), .ZN(n12562) );
  NAND2_X1 U14944 ( .A1(n13682), .A2(n12560), .ZN(n12561) );
  NAND2_X1 U14945 ( .A1(n12562), .A2(n12561), .ZN(n12588) );
  NAND2_X1 U14946 ( .A1(n12589), .A2(n12588), .ZN(n12596) );
  AND2_X1 U14947 ( .A1(n13806), .A2(n12575), .ZN(n12563) );
  AOI21_X1 U14948 ( .B1(n13797), .B2(n12584), .A(n12563), .ZN(n12594) );
  NAND2_X1 U14949 ( .A1(n13797), .A2(n6673), .ZN(n12565) );
  NAND2_X1 U14950 ( .A1(n13806), .A2(n12584), .ZN(n12564) );
  NAND2_X1 U14951 ( .A1(n12565), .A2(n12564), .ZN(n12593) );
  NAND2_X1 U14952 ( .A1(n12594), .A2(n12593), .ZN(n12566) );
  AND2_X1 U14953 ( .A1(n12596), .A2(n12566), .ZN(n12567) );
  NAND2_X1 U14954 ( .A1(n14107), .A2(n12584), .ZN(n12569) );
  NAND2_X1 U14955 ( .A1(n13683), .A2(n12575), .ZN(n12568) );
  AND2_X1 U14956 ( .A1(n13683), .A2(n12584), .ZN(n12570) );
  AOI21_X1 U14957 ( .B1(n14107), .B2(n12575), .A(n12570), .ZN(n12601) );
  NAND2_X1 U14958 ( .A1(n7613), .A2(n12571), .ZN(n12572) );
  NAND2_X1 U14959 ( .A1(n12574), .A2(n12573), .ZN(n12604) );
  INV_X1 U14960 ( .A(n13680), .ZN(n13767) );
  MUX2_X1 U14961 ( .A(n13767), .B(n12575), .S(n13765), .Z(n12592) );
  NOR2_X1 U14962 ( .A1(n12655), .A2(n13767), .ZN(n12591) );
  NAND2_X1 U14963 ( .A1(n12577), .A2(n12576), .ZN(n12579) );
  NAND2_X1 U14964 ( .A1(n7760), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12578) );
  NAND2_X1 U14965 ( .A1(n13680), .A2(n12575), .ZN(n12581) );
  NAND2_X1 U14966 ( .A1(n7651), .A2(n12666), .ZN(n12649) );
  NAND4_X1 U14967 ( .A1(n12581), .A2(n12646), .A3(n12657), .A4(n12649), .ZN(
        n12582) );
  AND2_X1 U14968 ( .A1(n12582), .A2(n13681), .ZN(n12583) );
  AOI21_X1 U14969 ( .B1(n13764), .B2(n12584), .A(n12583), .ZN(n12606) );
  NAND2_X1 U14970 ( .A1(n13764), .A2(n12655), .ZN(n12587) );
  NAND2_X1 U14971 ( .A1(n12585), .A2(n13681), .ZN(n12586) );
  NAND2_X1 U14972 ( .A1(n12587), .A2(n12586), .ZN(n12605) );
  OAI22_X1 U14973 ( .A1(n12606), .A2(n12605), .B1(n12589), .B2(n12588), .ZN(
        n12590) );
  OAI21_X1 U14974 ( .B1(n12592), .B2(n12591), .A(n12590), .ZN(n12599) );
  INV_X1 U14975 ( .A(n12593), .ZN(n12597) );
  INV_X1 U14976 ( .A(n12594), .ZN(n12595) );
  NAND4_X1 U14977 ( .A1(n12645), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12598) );
  INV_X1 U14978 ( .A(n12600), .ZN(n12602) );
  NOR2_X1 U14979 ( .A1(n7619), .A2(n7616), .ZN(n12603) );
  NAND2_X1 U14980 ( .A1(n12604), .A2(n12603), .ZN(n12608) );
  NAND2_X1 U14981 ( .A1(n12608), .A2(n12607), .ZN(n12680) );
  XNOR2_X1 U14982 ( .A(n13764), .B(n13681), .ZN(n12643) );
  XNOR2_X1 U14983 ( .A(n14120), .B(n13919), .ZN(n13910) );
  OAI21_X1 U14984 ( .B1(n13705), .B2(n12367), .A(n12609), .ZN(n15344) );
  NAND4_X1 U14985 ( .A1(n12612), .A2(n12611), .A3(n15344), .A4(n12610), .ZN(
        n12614) );
  NOR2_X1 U14986 ( .A1(n12614), .A2(n12613), .ZN(n12617) );
  NAND4_X1 U14987 ( .A1(n12618), .A2(n12617), .A3(n12616), .A4(n12615), .ZN(
        n12619) );
  NOR4_X1 U14988 ( .A1(n12622), .A2(n12621), .A3(n12620), .A4(n12619), .ZN(
        n12623) );
  NAND3_X1 U14989 ( .A1(n12625), .A2(n12624), .A3(n12623), .ZN(n12626) );
  OR4_X1 U14990 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12626), .ZN(
        n12630) );
  OR4_X1 U14991 ( .A1(n13979), .A2(n13986), .A3(n12631), .A4(n12630), .ZN(
        n12632) );
  NOR2_X1 U14992 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  NAND4_X1 U14993 ( .A1(n13910), .A2(n12634), .A3(n13917), .A4(n13956), .ZN(
        n12635) );
  OR4_X1 U14994 ( .A1(n13860), .A2(n13870), .A3(n13881), .A4(n12635), .ZN(
        n12639) );
  NAND2_X1 U14995 ( .A1(n12637), .A2(n12636), .ZN(n13823) );
  OR3_X1 U14996 ( .A1(n12639), .A2(n13823), .A3(n12638), .ZN(n12640) );
  NOR2_X1 U14997 ( .A1(n13800), .A2(n12640), .ZN(n12642) );
  AND4_X1 U14998 ( .A1(n12643), .A2(n12642), .A3(n12641), .A4(n13811), .ZN(
        n12644) );
  NOR2_X1 U14999 ( .A1(n12647), .A2(n12660), .ZN(n12665) );
  AOI21_X1 U15000 ( .B1(n12647), .B2(n12660), .A(n12646), .ZN(n12675) );
  INV_X1 U15001 ( .A(n12675), .ZN(n12648) );
  INV_X1 U15002 ( .A(n12661), .ZN(n12670) );
  NOR3_X1 U15003 ( .A1(n12665), .A2(n12648), .A3(n12670), .ZN(n12653) );
  OAI21_X1 U15004 ( .B1(n12650), .B2(n13759), .A(n12649), .ZN(n12651) );
  NAND2_X1 U15005 ( .A1(n12661), .A2(n12651), .ZN(n12672) );
  INV_X1 U15006 ( .A(n12672), .ZN(n12652) );
  NOR2_X1 U15007 ( .A1(n12653), .A2(n12652), .ZN(n12679) );
  MUX2_X1 U15008 ( .A(n13765), .B(n12560), .S(n13680), .Z(n12654) );
  OAI21_X1 U15009 ( .B1(n14097), .B2(n12655), .A(n12654), .ZN(n12673) );
  INV_X1 U15010 ( .A(n12656), .ZN(n12658) );
  OAI211_X1 U15011 ( .C1(n12660), .C2(n12659), .A(n12658), .B(n12657), .ZN(
        n12662) );
  AND2_X1 U15012 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  AND2_X1 U15013 ( .A1(n12673), .A2(n12663), .ZN(n12664) );
  NAND2_X1 U15014 ( .A1(n12680), .A2(n12664), .ZN(n12678) );
  AOI211_X1 U15015 ( .C1(n12666), .C2(n12673), .A(n12670), .B(n12665), .ZN(
        n12676) );
  NAND4_X1 U15016 ( .A1(n15343), .A2(n13991), .A3(n12668), .A4(n12667), .ZN(
        n12669) );
  OAI211_X1 U15017 ( .C1(n7651), .C2(n12670), .A(n12669), .B(P2_B_REG_SCAN_IN), 
        .ZN(n12671) );
  OAI21_X1 U15018 ( .B1(n12673), .B2(n12672), .A(n12671), .ZN(n12674) );
  AOI21_X1 U15019 ( .B1(n12676), .B2(n12675), .A(n12674), .ZN(n12677) );
  OAI211_X1 U15020 ( .C1(n12680), .C2(n12679), .A(n12678), .B(n12677), .ZN(
        P2_U3328) );
  INV_X1 U15021 ( .A(n12681), .ZN(n14766) );
  OAI222_X1 U15022 ( .A1(n14152), .A2(n12683), .B1(n14150), .B2(n14766), .C1(
        n12682), .C2(P2_U3088), .ZN(P2_U3298) );
  NAND2_X1 U15023 ( .A1(n14986), .A2(n12804), .ZN(n12685) );
  NAND2_X1 U15024 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  XNOR2_X1 U15025 ( .A(n12686), .B(n12824), .ZN(n12695) );
  NOR2_X1 U15026 ( .A1(n12687), .A2(n12826), .ZN(n12688) );
  AOI21_X1 U15027 ( .B1(n14986), .B2(n7074), .A(n12688), .ZN(n12693) );
  XNOR2_X1 U15028 ( .A(n12695), .B(n12693), .ZN(n14948) );
  INV_X1 U15029 ( .A(n12689), .ZN(n12691) );
  OR2_X1 U15030 ( .A1(n12691), .A2(n12690), .ZN(n14946) );
  INV_X1 U15031 ( .A(n12693), .ZN(n12694) );
  OR2_X1 U15032 ( .A1(n12695), .A2(n12694), .ZN(n12696) );
  NOR2_X1 U15033 ( .A1(n12697), .A2(n12826), .ZN(n12698) );
  AOI21_X1 U15034 ( .B1(n14801), .B2(n7074), .A(n12698), .ZN(n12704) );
  NAND2_X1 U15035 ( .A1(n14801), .A2(n12804), .ZN(n12700) );
  NAND2_X1 U15036 ( .A1(n14307), .A2(n7074), .ZN(n12699) );
  NAND2_X1 U15037 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  XNOR2_X1 U15038 ( .A(n12701), .B(n12824), .ZN(n12703) );
  XOR2_X1 U15039 ( .A(n12704), .B(n12703), .Z(n14201) );
  INV_X1 U15040 ( .A(n14201), .ZN(n12702) );
  INV_X1 U15041 ( .A(n12703), .ZN(n12705) );
  OR2_X1 U15042 ( .A1(n12705), .A2(n12704), .ZN(n12706) );
  NOR2_X1 U15043 ( .A1(n12707), .A2(n12826), .ZN(n12708) );
  AOI21_X1 U15044 ( .B1(n14245), .B2(n7074), .A(n12708), .ZN(n12715) );
  AOI22_X1 U15045 ( .A1(n14245), .A2(n12804), .B1(n7074), .B2(n14306), .ZN(
        n12709) );
  XNOR2_X1 U15046 ( .A(n12709), .B(n12824), .ZN(n12716) );
  XOR2_X1 U15047 ( .A(n12715), .B(n12716), .Z(n14247) );
  NAND2_X1 U15048 ( .A1(n14929), .A2(n12804), .ZN(n12711) );
  OR2_X1 U15049 ( .A1(n12713), .A2(n6686), .ZN(n12710) );
  NAND2_X1 U15050 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  XNOR2_X1 U15051 ( .A(n12712), .B(n12807), .ZN(n12719) );
  NOR2_X1 U15052 ( .A1(n12713), .A2(n12826), .ZN(n12714) );
  AOI21_X1 U15053 ( .B1(n14929), .B2(n7074), .A(n12714), .ZN(n12718) );
  XNOR2_X1 U15054 ( .A(n12719), .B(n12718), .ZN(n14924) );
  NOR2_X1 U15055 ( .A1(n12716), .A2(n12715), .ZN(n14925) );
  NOR2_X1 U15056 ( .A1(n14924), .A2(n14925), .ZN(n12717) );
  NAND2_X1 U15057 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  NAND2_X1 U15058 ( .A1(n12721), .A2(n12804), .ZN(n12723) );
  NAND2_X1 U15059 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  XNOR2_X1 U15060 ( .A(n12724), .B(n12807), .ZN(n12727) );
  INV_X1 U15061 ( .A(n12727), .ZN(n12725) );
  OAI22_X1 U15062 ( .A1(n14301), .A2(n6686), .B1(n12726), .B2(n12826), .ZN(
        n14290) );
  NOR2_X1 U15063 ( .A1(n12728), .A2(n12727), .ZN(n14936) );
  NAND2_X1 U15064 ( .A1(n14940), .A2(n12804), .ZN(n12730) );
  NAND2_X1 U15065 ( .A1(n14431), .A2(n7074), .ZN(n12729) );
  NAND2_X1 U15066 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  XNOR2_X1 U15067 ( .A(n12731), .B(n12807), .ZN(n12735) );
  AND2_X1 U15068 ( .A1(n14431), .A2(n12817), .ZN(n12732) );
  AOI21_X1 U15069 ( .B1(n14940), .B2(n7074), .A(n12732), .ZN(n12734) );
  XNOR2_X1 U15070 ( .A(n12735), .B(n12734), .ZN(n14935) );
  NOR2_X1 U15071 ( .A1(n14936), .A2(n14935), .ZN(n12733) );
  NAND2_X1 U15072 ( .A1(n12735), .A2(n12734), .ZN(n12736) );
  OAI22_X1 U15073 ( .A1(n14961), .A2(n12823), .B1(n12737), .B2(n6686), .ZN(
        n12738) );
  XNOR2_X1 U15074 ( .A(n12738), .B(n12824), .ZN(n14218) );
  OR2_X1 U15075 ( .A1(n14961), .A2(n6686), .ZN(n12740) );
  NAND2_X1 U15076 ( .A1(n14435), .A2(n12817), .ZN(n12739) );
  NAND2_X1 U15077 ( .A1(n12740), .A2(n12739), .ZN(n14217) );
  NAND2_X1 U15078 ( .A1(n14218), .A2(n14217), .ZN(n12741) );
  NAND2_X1 U15079 ( .A1(n12742), .A2(n12741), .ZN(n14268) );
  OAI22_X1 U15080 ( .A1(n14735), .A2(n12823), .B1(n14416), .B2(n6686), .ZN(
        n12743) );
  XNOR2_X1 U15081 ( .A(n12743), .B(n12824), .ZN(n12749) );
  OAI22_X1 U15082 ( .A1(n14735), .A2(n6686), .B1(n14416), .B2(n12826), .ZN(
        n12748) );
  XNOR2_X1 U15083 ( .A(n12749), .B(n12748), .ZN(n14271) );
  INV_X1 U15084 ( .A(n14271), .ZN(n12744) );
  AOI22_X1 U15085 ( .A1(n14728), .A2(n12804), .B1(n7074), .B2(n14417), .ZN(
        n12746) );
  XNOR2_X1 U15086 ( .A(n12746), .B(n12824), .ZN(n12751) );
  AND2_X1 U15087 ( .A1(n14417), .A2(n12817), .ZN(n12747) );
  AOI21_X1 U15088 ( .B1(n14728), .B2(n7074), .A(n12747), .ZN(n12752) );
  XNOR2_X1 U15089 ( .A(n12751), .B(n12752), .ZN(n14177) );
  NOR2_X1 U15090 ( .A1(n12749), .A2(n12748), .ZN(n14178) );
  NOR2_X1 U15091 ( .A1(n14177), .A2(n14178), .ZN(n12750) );
  INV_X1 U15092 ( .A(n12751), .ZN(n12754) );
  OAI22_X1 U15093 ( .A1(n14722), .A2(n6686), .B1(n14441), .B2(n12826), .ZN(
        n12756) );
  OAI22_X1 U15094 ( .A1(n14722), .A2(n12823), .B1(n14441), .B2(n6686), .ZN(
        n12755) );
  XNOR2_X1 U15095 ( .A(n12755), .B(n12824), .ZN(n12757) );
  XOR2_X1 U15096 ( .A(n12756), .B(n12757), .Z(n14237) );
  NAND2_X1 U15097 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  INV_X1 U15098 ( .A(n14188), .ZN(n12766) );
  NAND2_X1 U15099 ( .A1(n14590), .A2(n12804), .ZN(n12760) );
  NAND2_X1 U15100 ( .A1(n14564), .A2(n7074), .ZN(n12759) );
  NAND2_X1 U15101 ( .A1(n12760), .A2(n12759), .ZN(n12761) );
  XNOR2_X1 U15102 ( .A(n12761), .B(n12807), .ZN(n12764) );
  AND2_X1 U15103 ( .A1(n14564), .A2(n12817), .ZN(n12762) );
  AOI21_X1 U15104 ( .B1(n14590), .B2(n7074), .A(n12762), .ZN(n12763) );
  NAND2_X1 U15105 ( .A1(n12764), .A2(n12763), .ZN(n14255) );
  OAI21_X1 U15106 ( .B1(n12764), .B2(n12763), .A(n14255), .ZN(n14187) );
  INV_X1 U15107 ( .A(n14187), .ZN(n12765) );
  NAND2_X1 U15108 ( .A1(n14186), .A2(n14255), .ZN(n12774) );
  NAND2_X1 U15109 ( .A1(n14711), .A2(n12804), .ZN(n12768) );
  NAND2_X1 U15110 ( .A1(n12768), .A2(n12767), .ZN(n12769) );
  XNOR2_X1 U15111 ( .A(n12769), .B(n12807), .ZN(n12772) );
  NOR2_X1 U15112 ( .A1(n14443), .A2(n12826), .ZN(n12770) );
  AOI21_X1 U15113 ( .B1(n14711), .B2(n7074), .A(n12770), .ZN(n12771) );
  NAND2_X1 U15114 ( .A1(n12772), .A2(n12771), .ZN(n14164) );
  OR2_X1 U15115 ( .A1(n12772), .A2(n12771), .ZN(n12773) );
  NAND2_X1 U15116 ( .A1(n14557), .A2(n12804), .ZN(n12776) );
  NAND2_X1 U15117 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  XNOR2_X1 U15118 ( .A(n12777), .B(n12807), .ZN(n12779) );
  INV_X1 U15119 ( .A(n14566), .ZN(n14444) );
  NOR2_X1 U15120 ( .A1(n14444), .A2(n12826), .ZN(n12778) );
  AOI21_X1 U15121 ( .B1(n14557), .B2(n7074), .A(n12778), .ZN(n12780) );
  NAND2_X1 U15122 ( .A1(n12779), .A2(n12780), .ZN(n14231) );
  INV_X1 U15123 ( .A(n12779), .ZN(n12782) );
  INV_X1 U15124 ( .A(n12780), .ZN(n12781) );
  NAND2_X1 U15125 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  NAND2_X1 U15126 ( .A1(n6677), .A2(n12804), .ZN(n12786) );
  NAND2_X1 U15127 ( .A1(n12786), .A2(n12785), .ZN(n12787) );
  XNOR2_X1 U15128 ( .A(n12787), .B(n12807), .ZN(n12789) );
  NOR2_X1 U15129 ( .A1(n7399), .A2(n12826), .ZN(n12788) );
  AOI21_X1 U15130 ( .B1(n6677), .B2(n7074), .A(n12788), .ZN(n12790) );
  NAND2_X1 U15131 ( .A1(n12789), .A2(n12790), .ZN(n14210) );
  INV_X1 U15132 ( .A(n12789), .ZN(n12792) );
  INV_X1 U15133 ( .A(n12790), .ZN(n12791) );
  NAND2_X1 U15134 ( .A1(n12792), .A2(n12791), .ZN(n12793) );
  NAND2_X1 U15135 ( .A1(n14694), .A2(n12804), .ZN(n12795) );
  NAND2_X1 U15136 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  XNOR2_X1 U15137 ( .A(n12796), .B(n12807), .ZN(n12798) );
  INV_X1 U15138 ( .A(n14445), .ZN(n14227) );
  NOR2_X1 U15139 ( .A1(n14227), .A2(n12826), .ZN(n12797) );
  AOI21_X1 U15140 ( .B1(n14694), .B2(n7074), .A(n12797), .ZN(n12799) );
  NAND2_X1 U15141 ( .A1(n12798), .A2(n12799), .ZN(n12803) );
  INV_X1 U15142 ( .A(n12798), .ZN(n12801) );
  INV_X1 U15143 ( .A(n12799), .ZN(n12800) );
  NAND2_X1 U15144 ( .A1(n12801), .A2(n12800), .ZN(n12802) );
  NAND2_X1 U15145 ( .A1(n14688), .A2(n12804), .ZN(n12806) );
  NAND2_X1 U15146 ( .A1(n12806), .A2(n12805), .ZN(n12808) );
  XNOR2_X1 U15147 ( .A(n12808), .B(n12807), .ZN(n12811) );
  INV_X1 U15148 ( .A(n12811), .ZN(n12813) );
  NOR2_X1 U15149 ( .A1(n14205), .A2(n12826), .ZN(n12809) );
  AOI21_X1 U15150 ( .B1(n14688), .B2(n7074), .A(n12809), .ZN(n12810) );
  INV_X1 U15151 ( .A(n12810), .ZN(n12812) );
  AND2_X1 U15152 ( .A1(n12811), .A2(n12810), .ZN(n12814) );
  AOI21_X1 U15153 ( .B1(n12813), .B2(n12812), .A(n12814), .ZN(n14281) );
  NAND2_X1 U15154 ( .A1(n14280), .A2(n14281), .ZN(n14279) );
  INV_X1 U15155 ( .A(n12814), .ZN(n12815) );
  OAI22_X1 U15156 ( .A1(n14495), .A2(n12823), .B1(n12830), .B2(n6686), .ZN(
        n12816) );
  XNOR2_X1 U15157 ( .A(n12816), .B(n12824), .ZN(n12821) );
  OR2_X1 U15158 ( .A1(n14495), .A2(n6686), .ZN(n12819) );
  NAND2_X1 U15159 ( .A1(n14426), .A2(n12817), .ZN(n12818) );
  NAND2_X1 U15160 ( .A1(n12819), .A2(n12818), .ZN(n12820) );
  NOR2_X1 U15161 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  AOI21_X1 U15162 ( .B1(n12821), .B2(n12820), .A(n12822), .ZN(n14155) );
  OAI22_X1 U15163 ( .A1(n14479), .A2(n12823), .B1(n14461), .B2(n6686), .ZN(
        n12825) );
  XNOR2_X1 U15164 ( .A(n12825), .B(n12824), .ZN(n12828) );
  OAI22_X1 U15165 ( .A1(n14479), .A2(n6686), .B1(n14461), .B2(n12826), .ZN(
        n12827) );
  XNOR2_X1 U15166 ( .A(n12828), .B(n12827), .ZN(n12829) );
  OAI22_X1 U15167 ( .A1(n12831), .A2(n14401), .B1(n12830), .B2(n14460), .ZN(
        n14470) );
  AOI22_X1 U15168 ( .A1(n14953), .A2(n14470), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12832) );
  OAI21_X1 U15169 ( .B1(n14958), .B2(n14475), .A(n12832), .ZN(n12833) );
  AOI21_X1 U15170 ( .B1(n14674), .B2(n14950), .A(n12833), .ZN(n12834) );
  OAI21_X1 U15171 ( .B1(n12835), .B2(n14277), .A(n12834), .ZN(P1_U3220) );
  INV_X1 U15172 ( .A(n12836), .ZN(n14149) );
  OAI222_X1 U15173 ( .A1(n14771), .A2(n12839), .B1(n14768), .B2(n14149), .C1(
        n12838), .C2(P1_U3086), .ZN(P1_U3330) );
  XNOR2_X1 U15174 ( .A(n13148), .B(n12848), .ZN(n12918) );
  XNOR2_X1 U15175 ( .A(n12918), .B(n12925), .ZN(n12919) );
  XNOR2_X1 U15176 ( .A(n13220), .B(n12921), .ZN(n12899) );
  INV_X1 U15177 ( .A(n12899), .ZN(n12900) );
  XNOR2_X1 U15178 ( .A(n12976), .B(n12921), .ZN(n12970) );
  OR2_X1 U15179 ( .A1(n12970), .A2(n13200), .ZN(n12841) );
  XNOR2_X1 U15180 ( .A(n13209), .B(n12921), .ZN(n12966) );
  OR2_X1 U15181 ( .A1(n12966), .A2(n13217), .ZN(n12840) );
  NAND2_X1 U15182 ( .A1(n12841), .A2(n12840), .ZN(n12874) );
  NAND2_X1 U15183 ( .A1(n12844), .A2(n12994), .ZN(n12842) );
  NAND2_X1 U15184 ( .A1(n12843), .A2(n12842), .ZN(n12847) );
  INV_X1 U15185 ( .A(n12844), .ZN(n12845) );
  NAND2_X1 U15186 ( .A1(n12845), .A2(n13043), .ZN(n12846) );
  NAND2_X1 U15187 ( .A1(n12847), .A2(n12846), .ZN(n12989) );
  XNOR2_X1 U15188 ( .A(n12995), .B(n12848), .ZN(n12850) );
  NAND2_X1 U15189 ( .A1(n12850), .A2(n12849), .ZN(n12987) );
  NAND2_X1 U15190 ( .A1(n12989), .A2(n12987), .ZN(n12852) );
  INV_X1 U15191 ( .A(n12850), .ZN(n12851) );
  NAND2_X1 U15192 ( .A1(n12851), .A2(n12893), .ZN(n12988) );
  XNOR2_X1 U15193 ( .A(n13448), .B(n12921), .ZN(n12853) );
  XNOR2_X1 U15194 ( .A(n12853), .B(n13314), .ZN(n12890) );
  NAND2_X1 U15195 ( .A1(n12853), .A2(n12992), .ZN(n12854) );
  XNOR2_X1 U15196 ( .A(n13029), .B(n12921), .ZN(n12855) );
  XNOR2_X1 U15197 ( .A(n12855), .B(n13042), .ZN(n13031) );
  INV_X1 U15198 ( .A(n12855), .ZN(n12856) );
  NAND2_X1 U15199 ( .A1(n12856), .A2(n13042), .ZN(n12857) );
  XNOR2_X1 U15200 ( .A(n12949), .B(n12921), .ZN(n12858) );
  XNOR2_X1 U15201 ( .A(n12858), .B(n13287), .ZN(n12951) );
  NAND2_X1 U15202 ( .A1(n12952), .A2(n12951), .ZN(n12950) );
  INV_X1 U15203 ( .A(n12858), .ZN(n12859) );
  NAND2_X1 U15204 ( .A1(n12859), .A2(n13287), .ZN(n12860) );
  NAND2_X1 U15205 ( .A1(n12950), .A2(n12860), .ZN(n12961) );
  XNOR2_X1 U15206 ( .A(n13373), .B(n12921), .ZN(n12861) );
  XNOR2_X1 U15207 ( .A(n12861), .B(n12954), .ZN(n12960) );
  NAND2_X1 U15208 ( .A1(n12961), .A2(n12960), .ZN(n12959) );
  INV_X1 U15209 ( .A(n12861), .ZN(n12862) );
  NAND2_X1 U15210 ( .A1(n12862), .A2(n12954), .ZN(n12863) );
  XNOR2_X1 U15211 ( .A(n13278), .B(n12921), .ZN(n12864) );
  XNOR2_X1 U15212 ( .A(n12864), .B(n13256), .ZN(n13011) );
  NAND2_X1 U15213 ( .A1(n12864), .A2(n13256), .ZN(n12865) );
  XNOR2_X1 U15214 ( .A(n12909), .B(n12921), .ZN(n12866) );
  XNOR2_X1 U15215 ( .A(n12866), .B(n13274), .ZN(n12910) );
  INV_X1 U15216 ( .A(n12866), .ZN(n12867) );
  XNOR2_X1 U15217 ( .A(n13247), .B(n12921), .ZN(n12868) );
  XNOR2_X1 U15218 ( .A(n12868), .B(n13228), .ZN(n12980) );
  NAND2_X1 U15219 ( .A1(n12981), .A2(n12980), .ZN(n12979) );
  INV_X1 U15220 ( .A(n12868), .ZN(n12869) );
  NAND2_X1 U15221 ( .A1(n12869), .A2(n13228), .ZN(n12870) );
  NAND2_X1 U15222 ( .A1(n12979), .A2(n12870), .ZN(n12936) );
  XNOR2_X1 U15223 ( .A(n12933), .B(n12921), .ZN(n12871) );
  XNOR2_X1 U15224 ( .A(n12871), .B(n13002), .ZN(n12935) );
  NAND2_X1 U15225 ( .A1(n12936), .A2(n12935), .ZN(n12934) );
  INV_X1 U15226 ( .A(n12871), .ZN(n12872) );
  NAND2_X1 U15227 ( .A1(n12872), .A2(n13002), .ZN(n12873) );
  INV_X1 U15228 ( .A(n12970), .ZN(n12878) );
  AOI21_X1 U15229 ( .B1(n12966), .B2(n13217), .A(n13200), .ZN(n12877) );
  OR3_X1 U15230 ( .A1(n12874), .A2(n12900), .A3(n13229), .ZN(n12876) );
  NAND3_X1 U15231 ( .A1(n12966), .A2(n13217), .A3(n13200), .ZN(n12875) );
  OAI211_X1 U15232 ( .C1(n12878), .C2(n12877), .A(n12876), .B(n12875), .ZN(
        n12879) );
  XNOR2_X1 U15233 ( .A(n13335), .B(n12921), .ZN(n12881) );
  XNOR2_X1 U15234 ( .A(n12881), .B(n13157), .ZN(n12942) );
  XNOR2_X1 U15235 ( .A(n13407), .B(n12921), .ZN(n12882) );
  XNOR2_X1 U15236 ( .A(n12882), .B(n13169), .ZN(n13019) );
  INV_X1 U15237 ( .A(n12882), .ZN(n12883) );
  XOR2_X1 U15238 ( .A(n12919), .B(n12920), .Z(n12888) );
  AOI22_X1 U15239 ( .A1(n13149), .A2(n13037), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12885) );
  NAND2_X1 U15240 ( .A1(n13143), .A2(n13020), .ZN(n12884) );
  OAI211_X1 U15241 ( .C1(n13041), .C2(n13023), .A(n12885), .B(n12884), .ZN(
        n12886) );
  AOI21_X1 U15242 ( .B1(n13148), .B2(n15429), .A(n12886), .ZN(n12887) );
  OAI21_X1 U15243 ( .B1(n12888), .B2(n13027), .A(n12887), .ZN(P3_U3154) );
  OAI211_X1 U15244 ( .C1(n12891), .C2(n12890), .A(n12889), .B(n15432), .ZN(
        n12898) );
  INV_X1 U15245 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12892) );
  NOR2_X1 U15246 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12892), .ZN(n15580) );
  AOI21_X1 U15247 ( .B1(n12893), .B2(n13020), .A(n15580), .ZN(n12894) );
  OAI21_X1 U15248 ( .B1(n13302), .B2(n13023), .A(n12894), .ZN(n12895) );
  AOI21_X1 U15249 ( .B1(n12896), .B2(n13037), .A(n12895), .ZN(n12897) );
  OAI211_X1 U15250 ( .C1(n13040), .C2(n13448), .A(n12898), .B(n12897), .ZN(
        P3_U3155) );
  XNOR2_X1 U15251 ( .A(n12901), .B(n12899), .ZN(n13001) );
  NOR2_X1 U15252 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  AOI21_X1 U15253 ( .B1(n13001), .B2(n13199), .A(n12902), .ZN(n12967) );
  INV_X1 U15254 ( .A(n12967), .ZN(n12903) );
  XNOR2_X1 U15255 ( .A(n12969), .B(n13217), .ZN(n12908) );
  AOI22_X1 U15256 ( .A1(n13229), .A2(n13020), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12905) );
  NAND2_X1 U15257 ( .A1(n13208), .A2(n13037), .ZN(n12904) );
  OAI211_X1 U15258 ( .C1(n13200), .C2(n13023), .A(n12905), .B(n12904), .ZN(
        n12906) );
  AOI21_X1 U15259 ( .B1(n13209), .B2(n15429), .A(n12906), .ZN(n12907) );
  OAI21_X1 U15260 ( .B1(n12908), .B2(n13027), .A(n12907), .ZN(P3_U3156) );
  INV_X1 U15261 ( .A(n12909), .ZN(n13431) );
  AOI21_X1 U15262 ( .B1(n12911), .B2(n12910), .A(n13027), .ZN(n12913) );
  NAND2_X1 U15263 ( .A1(n12913), .A2(n12912), .ZN(n12917) );
  NAND2_X1 U15264 ( .A1(n13288), .A2(n13020), .ZN(n12914) );
  NAND2_X1 U15265 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13088)
         );
  OAI211_X1 U15266 ( .C1(n13257), .C2(n13023), .A(n12914), .B(n13088), .ZN(
        n12915) );
  AOI21_X1 U15267 ( .B1(n13263), .B2(n13037), .A(n12915), .ZN(n12916) );
  OAI211_X1 U15268 ( .C1(n13431), .C2(n13040), .A(n12917), .B(n12916), .ZN(
        P3_U3159) );
  XNOR2_X1 U15269 ( .A(n12922), .B(n12921), .ZN(n12923) );
  XNOR2_X1 U15270 ( .A(n12924), .B(n12923), .ZN(n12932) );
  AOI22_X1 U15271 ( .A1(n13130), .A2(n13037), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12927) );
  NAND2_X1 U15272 ( .A1(n12925), .A2(n13020), .ZN(n12926) );
  OAI211_X1 U15273 ( .C1(n12928), .C2(n13023), .A(n12927), .B(n12926), .ZN(
        n12929) );
  AOI21_X1 U15274 ( .B1(n12930), .B2(n15429), .A(n12929), .ZN(n12931) );
  OAI21_X1 U15275 ( .B1(n12932), .B2(n13027), .A(n12931), .ZN(P3_U3160) );
  INV_X1 U15276 ( .A(n12933), .ZN(n13423) );
  OAI211_X1 U15277 ( .C1(n12936), .C2(n12935), .A(n12934), .B(n15432), .ZN(
        n12940) );
  AOI22_X1 U15278 ( .A1(n13228), .A2(n13020), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12937) );
  OAI21_X1 U15279 ( .B1(n13199), .B2(n13023), .A(n12937), .ZN(n12938) );
  AOI21_X1 U15280 ( .B1(n13233), .B2(n13037), .A(n12938), .ZN(n12939) );
  OAI211_X1 U15281 ( .C1(n13423), .C2(n13040), .A(n12940), .B(n12939), .ZN(
        P3_U3163) );
  XOR2_X1 U15282 ( .A(n12942), .B(n12941), .Z(n12948) );
  OAI22_X1 U15283 ( .A1(n13200), .A2(n13035), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12943), .ZN(n12944) );
  AOI21_X1 U15284 ( .B1(n13175), .B2(n13037), .A(n12944), .ZN(n12945) );
  OAI21_X1 U15285 ( .B1(n13169), .B2(n13023), .A(n12945), .ZN(n12946) );
  AOI21_X1 U15286 ( .B1(n13335), .B2(n15429), .A(n12946), .ZN(n12947) );
  OAI21_X1 U15287 ( .B1(n12948), .B2(n13027), .A(n12947), .ZN(P3_U3165) );
  INV_X1 U15288 ( .A(n12949), .ZN(n13440) );
  OAI211_X1 U15289 ( .C1(n12952), .C2(n12951), .A(n12950), .B(n15432), .ZN(
        n12958) );
  NOR2_X1 U15290 ( .A1(n12953), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14838) );
  AOI21_X1 U15291 ( .B1(n12954), .B2(n15430), .A(n14838), .ZN(n12955) );
  OAI21_X1 U15292 ( .B1(n13302), .B2(n13035), .A(n12955), .ZN(n12956) );
  AOI21_X1 U15293 ( .B1(n13306), .B2(n13037), .A(n12956), .ZN(n12957) );
  OAI211_X1 U15294 ( .C1(n13440), .C2(n13040), .A(n12958), .B(n12957), .ZN(
        P3_U3166) );
  INV_X1 U15295 ( .A(n13373), .ZN(n13295) );
  OAI211_X1 U15296 ( .C1(n12961), .C2(n12960), .A(n12959), .B(n15432), .ZN(
        n12965) );
  AND2_X1 U15297 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14866) );
  AOI21_X1 U15298 ( .B1(n13288), .B2(n15430), .A(n14866), .ZN(n12962) );
  OAI21_X1 U15299 ( .B1(n13315), .B2(n13035), .A(n12962), .ZN(n12963) );
  AOI21_X1 U15300 ( .B1(n13293), .B2(n13037), .A(n12963), .ZN(n12964) );
  OAI211_X1 U15301 ( .C1(n13295), .C2(n13040), .A(n12965), .B(n12964), .ZN(
        P3_U3168) );
  INV_X1 U15302 ( .A(n12966), .ZN(n12968) );
  XNOR2_X1 U15303 ( .A(n12970), .B(n13200), .ZN(n12971) );
  XNOR2_X1 U15304 ( .A(n12972), .B(n12971), .ZN(n12978) );
  AOI22_X1 U15305 ( .A1(n13186), .A2(n13020), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12974) );
  NAND2_X1 U15306 ( .A1(n13191), .A2(n13037), .ZN(n12973) );
  OAI211_X1 U15307 ( .C1(n13157), .C2(n13023), .A(n12974), .B(n12973), .ZN(
        n12975) );
  AOI21_X1 U15308 ( .B1(n12976), .B2(n15429), .A(n12975), .ZN(n12977) );
  OAI21_X1 U15309 ( .B1(n12978), .B2(n13027), .A(n12977), .ZN(P3_U3169) );
  INV_X1 U15310 ( .A(n13247), .ZN(n13427) );
  OAI211_X1 U15311 ( .C1(n12981), .C2(n12980), .A(n12979), .B(n15432), .ZN(
        n12986) );
  AOI22_X1 U15312 ( .A1(n12982), .A2(n13020), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12983) );
  OAI21_X1 U15313 ( .B1(n13238), .B2(n13023), .A(n12983), .ZN(n12984) );
  AOI21_X1 U15314 ( .B1(n13245), .B2(n13037), .A(n12984), .ZN(n12985) );
  OAI211_X1 U15315 ( .C1(n13427), .C2(n13040), .A(n12986), .B(n12985), .ZN(
        P3_U3173) );
  NAND2_X1 U15316 ( .A1(n12988), .A2(n12987), .ZN(n12990) );
  XOR2_X1 U15317 ( .A(n12990), .B(n12989), .Z(n13000) );
  NOR2_X1 U15318 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12991), .ZN(n15562) );
  AOI21_X1 U15319 ( .B1(n15430), .B2(n12992), .A(n15562), .ZN(n12993) );
  OAI21_X1 U15320 ( .B1(n13035), .B2(n12994), .A(n12993), .ZN(n12997) );
  NOR2_X1 U15321 ( .A1(n12995), .A2(n13040), .ZN(n12996) );
  AOI211_X1 U15322 ( .C1(n12998), .C2(n13037), .A(n12997), .B(n12996), .ZN(
        n12999) );
  OAI21_X1 U15323 ( .B1(n13000), .B2(n13027), .A(n12999), .ZN(P3_U3174) );
  XNOR2_X1 U15324 ( .A(n13001), .B(n13229), .ZN(n13007) );
  AOI22_X1 U15325 ( .A1(n13002), .A2(n13020), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13004) );
  NAND2_X1 U15326 ( .A1(n13221), .A2(n13037), .ZN(n13003) );
  OAI211_X1 U15327 ( .C1(n13217), .C2(n13023), .A(n13004), .B(n13003), .ZN(
        n13005) );
  AOI21_X1 U15328 ( .B1(n13220), .B2(n15429), .A(n13005), .ZN(n13006) );
  OAI21_X1 U15329 ( .B1(n13007), .B2(n13027), .A(n13006), .ZN(P3_U3175) );
  INV_X1 U15330 ( .A(n13008), .ZN(n13009) );
  AOI21_X1 U15331 ( .B1(n13011), .B2(n13010), .A(n13009), .ZN(n13017) );
  NOR2_X1 U15332 ( .A1(n13301), .A2(n13035), .ZN(n13014) );
  OAI22_X1 U15333 ( .A1(n13274), .A2(n13023), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13012), .ZN(n13013) );
  AOI211_X1 U15334 ( .C1(n13279), .C2(n13037), .A(n13014), .B(n13013), .ZN(
        n13016) );
  NAND2_X1 U15335 ( .A1(n13278), .A2(n15429), .ZN(n13015) );
  OAI211_X1 U15336 ( .C1(n13017), .C2(n13027), .A(n13016), .B(n13015), .ZN(
        P3_U3178) );
  XOR2_X1 U15337 ( .A(n13019), .B(n13018), .Z(n13028) );
  AOI22_X1 U15338 ( .A1(n13162), .A2(n13037), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13022) );
  NAND2_X1 U15339 ( .A1(n13187), .A2(n13020), .ZN(n13021) );
  OAI211_X1 U15340 ( .C1(n13158), .C2(n13023), .A(n13022), .B(n13021), .ZN(
        n13024) );
  AOI21_X1 U15341 ( .B1(n13025), .B2(n15429), .A(n13024), .ZN(n13026) );
  OAI21_X1 U15342 ( .B1(n13028), .B2(n13027), .A(n13026), .ZN(P3_U3180) );
  INV_X1 U15343 ( .A(n13029), .ZN(n13444) );
  OAI211_X1 U15344 ( .C1(n13032), .C2(n13031), .A(n13030), .B(n15432), .ZN(
        n13039) );
  NOR2_X1 U15345 ( .A1(n13033), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14820) );
  AOI21_X1 U15346 ( .B1(n13287), .B2(n15430), .A(n14820), .ZN(n13034) );
  OAI21_X1 U15347 ( .B1(n13314), .B2(n13035), .A(n13034), .ZN(n13036) );
  AOI21_X1 U15348 ( .B1(n13318), .B2(n13037), .A(n13036), .ZN(n13038) );
  OAI211_X1 U15349 ( .C1(n13444), .C2(n13040), .A(n13039), .B(n13038), .ZN(
        P3_U3181) );
  INV_X1 U15350 ( .A(n13041), .ZN(n13144) );
  MUX2_X1 U15351 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13144), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15352 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13228), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15353 ( .A(n13042), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13044), .Z(
        P3_U3506) );
  MUX2_X1 U15354 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13043), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15355 ( .A(n15598), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13044), .Z(
        P3_U3500) );
  INV_X1 U15356 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14817) );
  NOR2_X1 U15357 ( .A1(n13047), .A2(n13048), .ZN(n13049) );
  AOI22_X1 U15358 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n13096), .B1(n15546), 
        .B2(n11525), .ZN(n15539) );
  INV_X1 U15359 ( .A(n15564), .ZN(n13069) );
  XNOR2_X1 U15360 ( .A(n13050), .B(n13069), .ZN(n15558) );
  NOR2_X1 U15361 ( .A1(n13069), .A2(n13050), .ZN(n13051) );
  XNOR2_X1 U15362 ( .A(n15583), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n15575) );
  INV_X1 U15363 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U15364 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13103), .B1(n14840), 
        .B2(n13053), .ZN(n14833) );
  NOR2_X1 U15365 ( .A1(n13054), .A2(n13055), .ZN(n13056) );
  INV_X1 U15366 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14854) );
  NOR2_X2 U15367 ( .A1(n14853), .A2(n14854), .ZN(n14852) );
  INV_X1 U15368 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U15369 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14869), .B1(n13090), 
        .B2(n13057), .ZN(n14880) );
  XNOR2_X1 U15370 ( .A(n13089), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13106) );
  MUX2_X1 U15371 ( .A(n6815), .B(n13106), .S(n6678), .Z(n13086) );
  INV_X1 U15372 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13371) );
  MUX2_X1 U15373 ( .A(n13057), .B(n13371), .S(n13078), .Z(n14875) );
  INV_X1 U15374 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13059) );
  MUX2_X1 U15375 ( .A(n14854), .B(n13059), .S(n6678), .Z(n13080) );
  NOR2_X1 U15376 ( .A1(n13080), .A2(n13054), .ZN(n13082) );
  OR2_X1 U15377 ( .A1(n13060), .A2(n13091), .ZN(n13061) );
  NAND2_X1 U15378 ( .A1(n13062), .A2(n13061), .ZN(n15533) );
  MUX2_X1 U15379 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6678), .Z(n13063) );
  XNOR2_X1 U15380 ( .A(n13063), .B(n13047), .ZN(n15532) );
  NAND2_X1 U15381 ( .A1(n15533), .A2(n15532), .ZN(n15531) );
  INV_X1 U15382 ( .A(n13063), .ZN(n13064) );
  NAND2_X1 U15383 ( .A1(n13064), .A2(n13047), .ZN(n13065) );
  NAND2_X1 U15384 ( .A1(n15531), .A2(n13065), .ZN(n15551) );
  MUX2_X1 U15385 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6678), .Z(n13066) );
  XNOR2_X1 U15386 ( .A(n13066), .B(n15546), .ZN(n15550) );
  NAND2_X1 U15387 ( .A1(n13066), .A2(n15546), .ZN(n13067) );
  MUX2_X1 U15388 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6678), .Z(n13068) );
  XNOR2_X1 U15389 ( .A(n13068), .B(n13069), .ZN(n15568) );
  NAND2_X1 U15390 ( .A1(n15569), .A2(n15568), .ZN(n15567) );
  INV_X1 U15391 ( .A(n13068), .ZN(n13070) );
  NAND2_X1 U15392 ( .A1(n13070), .A2(n13069), .ZN(n13071) );
  INV_X1 U15393 ( .A(n15575), .ZN(n13073) );
  NAND2_X1 U15394 ( .A1(n15583), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13099) );
  OR2_X1 U15395 ( .A1(n15583), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13072) );
  AND2_X1 U15396 ( .A1(n13099), .A2(n13072), .ZN(n15579) );
  MUX2_X1 U15397 ( .A(n13073), .B(n15579), .S(n6678), .Z(n15590) );
  NAND2_X1 U15398 ( .A1(n15591), .A2(n15590), .ZN(n15589) );
  NAND2_X1 U15399 ( .A1(n15583), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13074) );
  MUX2_X1 U15400 ( .A(n13074), .B(n13099), .S(n6678), .Z(n13075) );
  NAND2_X1 U15401 ( .A1(n15589), .A2(n13075), .ZN(n13076) );
  INV_X1 U15402 ( .A(n13076), .ZN(n13077) );
  XNOR2_X1 U15403 ( .A(n13076), .B(n14822), .ZN(n14826) );
  MUX2_X1 U15404 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6678), .Z(n14827) );
  NOR2_X1 U15405 ( .A1(n14826), .A2(n14827), .ZN(n14825) );
  AOI21_X1 U15406 ( .B1(n13077), .B2(n13101), .A(n14825), .ZN(n14848) );
  INV_X1 U15407 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13379) );
  MUX2_X1 U15408 ( .A(n13053), .B(n13379), .S(n13078), .Z(n13079) );
  NOR2_X1 U15409 ( .A1(n13079), .A2(n13103), .ZN(n14845) );
  NAND2_X1 U15410 ( .A1(n13079), .A2(n13103), .ZN(n14843) );
  OAI21_X1 U15411 ( .B1(n14848), .B2(n14845), .A(n14843), .ZN(n14859) );
  AOI21_X1 U15412 ( .B1(n13054), .B2(n13080), .A(n13082), .ZN(n13081) );
  INV_X1 U15413 ( .A(n13081), .ZN(n14860) );
  NOR2_X1 U15414 ( .A1(n14859), .A2(n14860), .ZN(n14858) );
  NOR2_X1 U15415 ( .A1(n13082), .A2(n14858), .ZN(n13083) );
  XNOR2_X1 U15416 ( .A(n13090), .B(n13083), .ZN(n14876) );
  NAND2_X1 U15417 ( .A1(n14875), .A2(n14876), .ZN(n14874) );
  NAND2_X1 U15418 ( .A1(n14869), .A2(n13083), .ZN(n13084) );
  NAND2_X1 U15419 ( .A1(n14874), .A2(n13084), .ZN(n13085) );
  XOR2_X1 U15420 ( .A(n13086), .B(n13085), .Z(n13111) );
  NAND2_X1 U15421 ( .A1(n15581), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13087) );
  OAI211_X1 U15422 ( .C1(n15584), .C2(n13089), .A(n13088), .B(n13087), .ZN(
        n13110) );
  AOI22_X1 U15423 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n13090), .B1(n14869), 
        .B2(n13371), .ZN(n14873) );
  AOI22_X1 U15424 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14840), .B1(n13103), 
        .B2(n13379), .ZN(n14837) );
  INV_X1 U15425 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14895) );
  AOI22_X1 U15426 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15546), .B1(n13096), 
        .B2(n14895), .ZN(n15543) );
  NAND2_X1 U15427 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n13091), .ZN(n13093) );
  NAND2_X1 U15428 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  NAND2_X1 U15429 ( .A1(n15528), .A2(n13094), .ZN(n13095) );
  XNOR2_X1 U15430 ( .A(n13047), .B(n13094), .ZN(n15525) );
  NAND2_X1 U15431 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15525), .ZN(n15524) );
  NAND2_X1 U15432 ( .A1(n13095), .A2(n15524), .ZN(n15542) );
  NAND2_X1 U15433 ( .A1(n15543), .A2(n15542), .ZN(n15541) );
  NAND2_X1 U15434 ( .A1(n15564), .A2(n13097), .ZN(n13098) );
  NAND2_X1 U15435 ( .A1(n13098), .A2(n15560), .ZN(n15578) );
  NAND2_X1 U15436 ( .A1(n15579), .A2(n15578), .ZN(n15577) );
  NAND2_X1 U15437 ( .A1(n13099), .A2(n15577), .ZN(n13100) );
  NAND2_X1 U15438 ( .A1(n14822), .A2(n13100), .ZN(n13102) );
  XNOR2_X1 U15439 ( .A(n13101), .B(n13100), .ZN(n14819) );
  NAND2_X1 U15440 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14819), .ZN(n14818) );
  NAND2_X1 U15441 ( .A1(n13102), .A2(n14818), .ZN(n14836) );
  NAND2_X1 U15442 ( .A1(n14837), .A2(n14836), .ZN(n14835) );
  NAND2_X1 U15443 ( .A1(n14862), .A2(n13104), .ZN(n13105) );
  NAND2_X1 U15444 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14856), .ZN(n14855) );
  NAND2_X1 U15445 ( .A1(n13105), .A2(n14855), .ZN(n14872) );
  XNOR2_X1 U15446 ( .A(n13107), .B(n13106), .ZN(n13108) );
  NOR2_X1 U15447 ( .A1(n13108), .A2(n15488), .ZN(n13109) );
  OAI21_X1 U15448 ( .B1(n13113), .B2(n15594), .A(n13112), .ZN(P3_U3201) );
  NAND2_X1 U15449 ( .A1(n15649), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13118) );
  INV_X1 U15450 ( .A(n13114), .ZN(n13115) );
  NOR2_X1 U15451 ( .A1(n13117), .A2(n15676), .ZN(n13122) );
  OAI21_X1 U15452 ( .B1(n13391), .B2(n13122), .A(n15682), .ZN(n13119) );
  OAI211_X1 U15453 ( .C1(n13393), .C2(n13320), .A(n13118), .B(n13119), .ZN(
        P3_U3202) );
  NAND2_X1 U15454 ( .A1(n15649), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13120) );
  OAI211_X1 U15455 ( .C1(n13396), .C2(n13320), .A(n13120), .B(n13119), .ZN(
        P3_U3203) );
  INV_X1 U15456 ( .A(n13121), .ZN(n13128) );
  AOI21_X1 U15457 ( .B1(n15649), .B2(P3_REG2_REG_29__SCAN_IN), .A(n13122), 
        .ZN(n13123) );
  OAI21_X1 U15458 ( .B1(n13124), .B2(n13320), .A(n13123), .ZN(n13125) );
  AOI21_X1 U15459 ( .B1(n13126), .B2(n15631), .A(n13125), .ZN(n13127) );
  OAI21_X1 U15460 ( .B1(n13128), .B2(n15649), .A(n13127), .ZN(P3_U3204) );
  INV_X1 U15461 ( .A(n13129), .ZN(n13135) );
  AOI22_X1 U15462 ( .A1(n13130), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13131) );
  OAI21_X1 U15463 ( .B1(n13400), .B2(n13320), .A(n13131), .ZN(n13132) );
  AOI21_X1 U15464 ( .B1(n13133), .B2(n15631), .A(n13132), .ZN(n13134) );
  OAI21_X1 U15465 ( .B1(n13135), .B2(n15649), .A(n13134), .ZN(P3_U3205) );
  INV_X1 U15466 ( .A(n13136), .ZN(n13138) );
  NAND2_X1 U15467 ( .A1(n13142), .A2(n15671), .ZN(n13146) );
  AOI22_X1 U15468 ( .A1(n13144), .A2(n15654), .B1(n15653), .B2(n13143), .ZN(
        n13145) );
  INV_X1 U15469 ( .A(n13327), .ZN(n13153) );
  INV_X1 U15470 ( .A(n13147), .ZN(n13328) );
  AOI22_X1 U15471 ( .A1(n13149), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13150) );
  OAI21_X1 U15472 ( .B1(n8883), .B2(n13320), .A(n13150), .ZN(n13151) );
  AOI21_X1 U15473 ( .B1(n13328), .B2(n15666), .A(n13151), .ZN(n13152) );
  OAI21_X1 U15474 ( .B1(n13153), .B2(n15649), .A(n13152), .ZN(P3_U3206) );
  XNOR2_X1 U15475 ( .A(n13154), .B(n13155), .ZN(n13161) );
  XNOR2_X1 U15476 ( .A(n13156), .B(n13155), .ZN(n13332) );
  OAI22_X1 U15477 ( .A1(n13158), .A2(n15673), .B1(n13157), .B2(n15637), .ZN(
        n13159) );
  AOI21_X1 U15478 ( .B1(n13332), .B2(n15645), .A(n13159), .ZN(n13160) );
  OAI21_X1 U15479 ( .B1(n13161), .B2(n15641), .A(n13160), .ZN(n13331) );
  INV_X1 U15480 ( .A(n13331), .ZN(n13166) );
  AOI22_X1 U15481 ( .A1(n13162), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13163) );
  OAI21_X1 U15482 ( .B1(n13407), .B2(n13320), .A(n13163), .ZN(n13164) );
  AOI21_X1 U15483 ( .B1(n13332), .B2(n15666), .A(n13164), .ZN(n13165) );
  OAI21_X1 U15484 ( .B1(n13166), .B2(n15649), .A(n13165), .ZN(P3_U3207) );
  INV_X1 U15485 ( .A(n13167), .ZN(n13168) );
  AOI21_X1 U15486 ( .B1(n13168), .B2(n13173), .A(n15641), .ZN(n13172) );
  OAI22_X1 U15487 ( .A1(n13169), .A2(n15673), .B1(n13200), .B2(n15637), .ZN(
        n13170) );
  AOI21_X1 U15488 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(n13338) );
  XNOR2_X1 U15489 ( .A(n13174), .B(n13173), .ZN(n13336) );
  NAND2_X1 U15490 ( .A1(n13335), .A2(n13246), .ZN(n13177) );
  AOI22_X1 U15491 ( .A1(n13175), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U15492 ( .A1(n13177), .A2(n13176), .ZN(n13178) );
  AOI21_X1 U15493 ( .B1(n13336), .B2(n15631), .A(n13178), .ZN(n13179) );
  OAI21_X1 U15494 ( .B1(n13338), .B2(n15649), .A(n13179), .ZN(P3_U3208) );
  INV_X1 U15495 ( .A(n13180), .ZN(n13181) );
  AOI21_X1 U15496 ( .B1(n13184), .B2(n13182), .A(n13181), .ZN(n13190) );
  OAI211_X1 U15497 ( .C1(n13185), .C2(n13184), .A(n13183), .B(n15671), .ZN(
        n13189) );
  AOI22_X1 U15498 ( .A1(n13187), .A2(n15654), .B1(n15653), .B2(n13186), .ZN(
        n13188) );
  OAI211_X1 U15499 ( .C1(n15662), .C2(n13190), .A(n13189), .B(n13188), .ZN(
        n13339) );
  INV_X1 U15500 ( .A(n13339), .ZN(n13195) );
  INV_X1 U15501 ( .A(n13190), .ZN(n13340) );
  AOI22_X1 U15502 ( .A1(n13191), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13192) );
  OAI21_X1 U15503 ( .B1(n13412), .B2(n13320), .A(n13192), .ZN(n13193) );
  AOI21_X1 U15504 ( .B1(n13340), .B2(n15666), .A(n13193), .ZN(n13194) );
  OAI21_X1 U15505 ( .B1(n13195), .B2(n15649), .A(n13194), .ZN(P3_U3209) );
  NAND2_X1 U15506 ( .A1(n13196), .A2(n13204), .ZN(n13197) );
  NAND3_X1 U15507 ( .A1(n13198), .A2(n15671), .A3(n13197), .ZN(n13203) );
  OAI22_X1 U15508 ( .A1(n13200), .A2(n15673), .B1(n13199), .B2(n15637), .ZN(
        n13201) );
  INV_X1 U15509 ( .A(n13201), .ZN(n13202) );
  NAND2_X1 U15510 ( .A1(n13203), .A2(n13202), .ZN(n13346) );
  OR2_X1 U15511 ( .A1(n13205), .A2(n13204), .ZN(n13206) );
  NAND2_X1 U15512 ( .A1(n13207), .A2(n13206), .ZN(n13344) );
  AOI22_X1 U15513 ( .A1(n13208), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U15514 ( .A1(n13209), .A2(n13246), .ZN(n13210) );
  OAI211_X1 U15515 ( .C1(n13344), .C2(n13250), .A(n13211), .B(n13210), .ZN(
        n13212) );
  AOI21_X1 U15516 ( .B1(n13346), .B2(n15682), .A(n13212), .ZN(n13213) );
  INV_X1 U15517 ( .A(n13213), .ZN(P3_U3210) );
  XNOR2_X1 U15518 ( .A(n13215), .B(n13214), .ZN(n13216) );
  OAI222_X1 U15519 ( .A1(n15673), .A2(n13217), .B1(n15637), .B2(n13238), .C1(
        n15641), .C2(n13216), .ZN(n13349) );
  INV_X1 U15520 ( .A(n13349), .ZN(n13225) );
  XNOR2_X1 U15521 ( .A(n13219), .B(n13218), .ZN(n13350) );
  INV_X1 U15522 ( .A(n13220), .ZN(n13419) );
  AOI22_X1 U15523 ( .A1(n13221), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13222) );
  OAI21_X1 U15524 ( .B1(n13419), .B2(n13320), .A(n13222), .ZN(n13223) );
  AOI21_X1 U15525 ( .B1(n13350), .B2(n15631), .A(n13223), .ZN(n13224) );
  OAI21_X1 U15526 ( .B1(n13225), .B2(n15649), .A(n13224), .ZN(P3_U3211) );
  OAI21_X1 U15527 ( .B1(n13227), .B2(n13231), .A(n13226), .ZN(n13230) );
  AOI222_X1 U15528 ( .A1(n15671), .A2(n13230), .B1(n13229), .B2(n15654), .C1(
        n13228), .C2(n15653), .ZN(n13353) );
  XNOR2_X1 U15529 ( .A(n13232), .B(n13231), .ZN(n13355) );
  AOI22_X1 U15530 ( .A1(n13233), .A2(n6668), .B1(n15649), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n13234) );
  OAI21_X1 U15531 ( .B1(n13423), .B2(n13320), .A(n13234), .ZN(n13235) );
  AOI21_X1 U15532 ( .B1(n13355), .B2(n15631), .A(n13235), .ZN(n13236) );
  OAI21_X1 U15533 ( .B1(n13353), .B2(n15649), .A(n13236), .ZN(P3_U3212) );
  XNOR2_X1 U15534 ( .A(n13237), .B(n8744), .ZN(n13240) );
  OAI22_X1 U15535 ( .A1(n13238), .A2(n15673), .B1(n13274), .B2(n15637), .ZN(
        n13239) );
  AOI21_X1 U15536 ( .B1(n13240), .B2(n15671), .A(n13239), .ZN(n13361) );
  NAND2_X1 U15537 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  NAND2_X1 U15538 ( .A1(n13244), .A2(n13243), .ZN(n13359) );
  AOI22_X1 U15539 ( .A1(n15649), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13245), 
        .B2(n6668), .ZN(n13249) );
  NAND2_X1 U15540 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  OAI211_X1 U15541 ( .C1(n13359), .C2(n13250), .A(n13249), .B(n13248), .ZN(
        n13251) );
  INV_X1 U15542 ( .A(n13251), .ZN(n13252) );
  OAI21_X1 U15543 ( .B1(n13361), .B2(n15649), .A(n13252), .ZN(P3_U3213) );
  NAND2_X1 U15544 ( .A1(n13271), .A2(n13253), .ZN(n13255) );
  AOI21_X1 U15545 ( .B1(n13255), .B2(n13254), .A(n15641), .ZN(n13260) );
  OAI22_X1 U15546 ( .A1(n13257), .A2(n15673), .B1(n13256), .B2(n15637), .ZN(
        n13258) );
  AOI21_X1 U15547 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(n13366) );
  XNOR2_X1 U15548 ( .A(n13262), .B(n13261), .ZN(n13364) );
  AOI22_X1 U15549 ( .A1(n15649), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n6668), 
        .B2(n13263), .ZN(n13264) );
  OAI21_X1 U15550 ( .B1(n13431), .B2(n13320), .A(n13264), .ZN(n13265) );
  AOI21_X1 U15551 ( .B1(n13364), .B2(n15631), .A(n13265), .ZN(n13266) );
  OAI21_X1 U15552 ( .B1(n13366), .B2(n15649), .A(n13266), .ZN(P3_U3214) );
  NAND2_X1 U15553 ( .A1(n13285), .A2(n13267), .ZN(n13269) );
  AND2_X1 U15554 ( .A1(n13269), .A2(n13268), .ZN(n13272) );
  AOI21_X1 U15555 ( .B1(n13276), .B2(n13272), .A(n7627), .ZN(n13273) );
  OAI222_X1 U15556 ( .A1(n15673), .A2(n13274), .B1(n15637), .B2(n13301), .C1(
        n15641), .C2(n13273), .ZN(n13369) );
  INV_X1 U15557 ( .A(n13369), .ZN(n13283) );
  NAND2_X1 U15558 ( .A1(n13290), .A2(n13275), .ZN(n13277) );
  XNOR2_X1 U15559 ( .A(n13277), .B(n13276), .ZN(n13370) );
  INV_X1 U15560 ( .A(n13278), .ZN(n13435) );
  AOI22_X1 U15561 ( .A1(n15649), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n6668), 
        .B2(n13279), .ZN(n13280) );
  OAI21_X1 U15562 ( .B1(n13435), .B2(n13320), .A(n13280), .ZN(n13281) );
  AOI21_X1 U15563 ( .B1(n13370), .B2(n15631), .A(n13281), .ZN(n13282) );
  OAI21_X1 U15564 ( .B1(n13283), .B2(n15649), .A(n13282), .ZN(P3_U3215) );
  NAND2_X1 U15565 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  XNOR2_X1 U15566 ( .A(n13286), .B(n13291), .ZN(n13289) );
  AOI222_X1 U15567 ( .A1(n15671), .A2(n13289), .B1(n13288), .B2(n15654), .C1(
        n13287), .C2(n15653), .ZN(n13376) );
  OAI21_X1 U15568 ( .B1(n13292), .B2(n13291), .A(n13290), .ZN(n13374) );
  AOI22_X1 U15569 ( .A1(n15649), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n6668), 
        .B2(n13293), .ZN(n13294) );
  OAI21_X1 U15570 ( .B1(n13295), .B2(n13320), .A(n13294), .ZN(n13296) );
  AOI21_X1 U15571 ( .B1(n13374), .B2(n15631), .A(n13296), .ZN(n13297) );
  OAI21_X1 U15572 ( .B1(n13376), .B2(n15649), .A(n13297), .ZN(P3_U3216) );
  XNOR2_X1 U15573 ( .A(n13299), .B(n13298), .ZN(n13300) );
  OAI222_X1 U15574 ( .A1(n15637), .A2(n13302), .B1(n15673), .B2(n13301), .C1(
        n13300), .C2(n15641), .ZN(n13377) );
  INV_X1 U15575 ( .A(n13377), .ZN(n13310) );
  OAI21_X1 U15576 ( .B1(n13305), .B2(n13304), .A(n13303), .ZN(n13378) );
  AOI22_X1 U15577 ( .A1(n15649), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n6668), 
        .B2(n13306), .ZN(n13307) );
  OAI21_X1 U15578 ( .B1(n13440), .B2(n13320), .A(n13307), .ZN(n13308) );
  AOI21_X1 U15579 ( .B1(n13378), .B2(n15631), .A(n13308), .ZN(n13309) );
  OAI21_X1 U15580 ( .B1(n13310), .B2(n15649), .A(n13309), .ZN(P3_U3217) );
  XNOR2_X1 U15581 ( .A(n13311), .B(n13312), .ZN(n13313) );
  OAI222_X1 U15582 ( .A1(n15673), .A2(n13315), .B1(n15637), .B2(n13314), .C1(
        n13313), .C2(n15641), .ZN(n13381) );
  INV_X1 U15583 ( .A(n13381), .ZN(n13323) );
  XNOR2_X1 U15584 ( .A(n13317), .B(n13316), .ZN(n13382) );
  AOI22_X1 U15585 ( .A1(n15649), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n6668), 
        .B2(n13318), .ZN(n13319) );
  OAI21_X1 U15586 ( .B1(n13444), .B2(n13320), .A(n13319), .ZN(n13321) );
  AOI21_X1 U15587 ( .B1(n13382), .B2(n15631), .A(n13321), .ZN(n13322) );
  OAI21_X1 U15588 ( .B1(n13323), .B2(n15649), .A(n13322), .ZN(P3_U3218) );
  NAND2_X1 U15589 ( .A1(n15761), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U15590 ( .A1(n13391), .A2(n15764), .ZN(n13326) );
  OAI211_X1 U15591 ( .C1(n13393), .C2(n13390), .A(n13324), .B(n13326), .ZN(
        P3_U3490) );
  NAND2_X1 U15592 ( .A1(n15761), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13325) );
  OAI211_X1 U15593 ( .C1(n13396), .C2(n13390), .A(n13326), .B(n13325), .ZN(
        P3_U3489) );
  INV_X1 U15594 ( .A(n15719), .ZN(n15739) );
  MUX2_X1 U15595 ( .A(n13329), .B(n13401), .S(n15764), .Z(n13330) );
  AOI21_X1 U15596 ( .B1(n15739), .B2(n13332), .A(n13331), .ZN(n13404) );
  MUX2_X1 U15597 ( .A(n13333), .B(n13404), .S(n15764), .Z(n13334) );
  OAI21_X1 U15598 ( .B1(n13407), .B2(n13390), .A(n13334), .ZN(P3_U3485) );
  AOI22_X1 U15599 ( .A1(n13336), .A2(n15732), .B1(n15677), .B2(n13335), .ZN(
        n13337) );
  NAND2_X1 U15600 ( .A1(n13338), .A2(n13337), .ZN(n13408) );
  MUX2_X1 U15601 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13408), .S(n15764), .Z(
        P3_U3484) );
  AOI21_X1 U15602 ( .B1(n15739), .B2(n13340), .A(n13339), .ZN(n13409) );
  MUX2_X1 U15603 ( .A(n13341), .B(n13409), .S(n15764), .Z(n13342) );
  OAI21_X1 U15604 ( .B1(n13412), .B2(n13390), .A(n13342), .ZN(P3_U3483) );
  INV_X1 U15605 ( .A(n15732), .ZN(n13358) );
  OAI22_X1 U15606 ( .A1(n13344), .A2(n13358), .B1(n13343), .B2(n15718), .ZN(
        n13345) );
  NOR2_X1 U15607 ( .A1(n13346), .A2(n13345), .ZN(n13413) );
  MUX2_X1 U15608 ( .A(n13347), .B(n13413), .S(n15764), .Z(n13348) );
  INV_X1 U15609 ( .A(n13348), .ZN(P3_U3482) );
  AOI21_X1 U15610 ( .B1(n15732), .B2(n13350), .A(n13349), .ZN(n13416) );
  MUX2_X1 U15611 ( .A(n13351), .B(n13416), .S(n15764), .Z(n13352) );
  OAI21_X1 U15612 ( .B1(n13419), .B2(n13390), .A(n13352), .ZN(P3_U3481) );
  INV_X1 U15613 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13356) );
  INV_X1 U15614 ( .A(n13353), .ZN(n13354) );
  AOI21_X1 U15615 ( .B1(n15732), .B2(n13355), .A(n13354), .ZN(n13420) );
  MUX2_X1 U15616 ( .A(n13356), .B(n13420), .S(n15764), .Z(n13357) );
  OAI21_X1 U15617 ( .B1(n13423), .B2(n13390), .A(n13357), .ZN(P3_U3480) );
  NAND2_X1 U15618 ( .A1(n13361), .A2(n13360), .ZN(n13424) );
  MUX2_X1 U15619 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13424), .S(n15764), .Z(
        n13362) );
  INV_X1 U15620 ( .A(n13362), .ZN(n13363) );
  OAI21_X1 U15621 ( .B1(n13427), .B2(n13390), .A(n13363), .ZN(P3_U3479) );
  NAND2_X1 U15622 ( .A1(n13364), .A2(n15732), .ZN(n13365) );
  NAND2_X1 U15623 ( .A1(n13366), .A2(n13365), .ZN(n13428) );
  MUX2_X1 U15624 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13428), .S(n15764), .Z(
        n13367) );
  INV_X1 U15625 ( .A(n13367), .ZN(n13368) );
  OAI21_X1 U15626 ( .B1(n13431), .B2(n13390), .A(n13368), .ZN(P3_U3478) );
  AOI21_X1 U15627 ( .B1(n13370), .B2(n15732), .A(n13369), .ZN(n13432) );
  MUX2_X1 U15628 ( .A(n13371), .B(n13432), .S(n15764), .Z(n13372) );
  OAI21_X1 U15629 ( .B1(n13435), .B2(n13390), .A(n13372), .ZN(P3_U3477) );
  AOI22_X1 U15630 ( .A1(n13374), .A2(n15732), .B1(n15677), .B2(n13373), .ZN(
        n13375) );
  NAND2_X1 U15631 ( .A1(n13376), .A2(n13375), .ZN(n13436) );
  MUX2_X1 U15632 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13436), .S(n15764), .Z(
        P3_U3476) );
  AOI21_X1 U15633 ( .B1(n15732), .B2(n13378), .A(n13377), .ZN(n13437) );
  MUX2_X1 U15634 ( .A(n13379), .B(n13437), .S(n15764), .Z(n13380) );
  OAI21_X1 U15635 ( .B1(n13440), .B2(n13390), .A(n13380), .ZN(P3_U3475) );
  INV_X1 U15636 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13383) );
  AOI21_X1 U15637 ( .B1(n13382), .B2(n15732), .A(n13381), .ZN(n13441) );
  MUX2_X1 U15638 ( .A(n13383), .B(n13441), .S(n15764), .Z(n13384) );
  OAI21_X1 U15639 ( .B1(n13444), .B2(n13390), .A(n13384), .ZN(P3_U3474) );
  NAND2_X1 U15640 ( .A1(n13385), .A2(n15732), .ZN(n13386) );
  NAND2_X1 U15641 ( .A1(n13387), .A2(n13386), .ZN(n13445) );
  MUX2_X1 U15642 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13445), .S(n15764), .Z(
        n13388) );
  INV_X1 U15643 ( .A(n13388), .ZN(n13389) );
  OAI21_X1 U15644 ( .B1(n13390), .B2(n13448), .A(n13389), .ZN(P3_U3473) );
  NAND2_X1 U15645 ( .A1(n15742), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13392) );
  NAND2_X1 U15646 ( .A1(n13391), .A2(n15740), .ZN(n13395) );
  OAI211_X1 U15647 ( .C1(n13393), .C2(n13449), .A(n13392), .B(n13395), .ZN(
        P3_U3458) );
  NAND2_X1 U15648 ( .A1(n15742), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13394) );
  OAI211_X1 U15649 ( .C1(n13396), .C2(n13449), .A(n13395), .B(n13394), .ZN(
        P3_U3457) );
  INV_X1 U15650 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13398) );
  MUX2_X1 U15651 ( .A(n13398), .B(n13397), .S(n15740), .Z(n13399) );
  OAI21_X1 U15652 ( .B1(n13400), .B2(n13449), .A(n13399), .ZN(P3_U3455) );
  INV_X1 U15653 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13402) );
  MUX2_X1 U15654 ( .A(n13402), .B(n13401), .S(n15740), .Z(n13403) );
  INV_X1 U15655 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13405) );
  MUX2_X1 U15656 ( .A(n13405), .B(n13404), .S(n15740), .Z(n13406) );
  OAI21_X1 U15657 ( .B1(n13407), .B2(n13449), .A(n13406), .ZN(P3_U3453) );
  MUX2_X1 U15658 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13408), .S(n15740), .Z(
        P3_U3452) );
  INV_X1 U15659 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13410) );
  MUX2_X1 U15660 ( .A(n13410), .B(n13409), .S(n15740), .Z(n13411) );
  OAI21_X1 U15661 ( .B1(n13412), .B2(n13449), .A(n13411), .ZN(P3_U3451) );
  INV_X1 U15662 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13414) );
  MUX2_X1 U15663 ( .A(n13414), .B(n13413), .S(n15740), .Z(n13415) );
  INV_X1 U15664 ( .A(n13415), .ZN(P3_U3450) );
  INV_X1 U15665 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13417) );
  MUX2_X1 U15666 ( .A(n13417), .B(n13416), .S(n15740), .Z(n13418) );
  OAI21_X1 U15667 ( .B1(n13419), .B2(n13449), .A(n13418), .ZN(P3_U3449) );
  INV_X1 U15668 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13421) );
  MUX2_X1 U15669 ( .A(n13421), .B(n13420), .S(n15740), .Z(n13422) );
  OAI21_X1 U15670 ( .B1(n13423), .B2(n13449), .A(n13422), .ZN(P3_U3448) );
  MUX2_X1 U15671 ( .A(n13424), .B(P3_REG0_REG_20__SCAN_IN), .S(n15742), .Z(
        n13425) );
  INV_X1 U15672 ( .A(n13425), .ZN(n13426) );
  OAI21_X1 U15673 ( .B1(n13427), .B2(n13449), .A(n13426), .ZN(P3_U3447) );
  MUX2_X1 U15674 ( .A(n13428), .B(P3_REG0_REG_19__SCAN_IN), .S(n15742), .Z(
        n13429) );
  INV_X1 U15675 ( .A(n13429), .ZN(n13430) );
  OAI21_X1 U15676 ( .B1(n13431), .B2(n13449), .A(n13430), .ZN(P3_U3446) );
  INV_X1 U15677 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13433) );
  MUX2_X1 U15678 ( .A(n13433), .B(n13432), .S(n15740), .Z(n13434) );
  OAI21_X1 U15679 ( .B1(n13435), .B2(n13449), .A(n13434), .ZN(P3_U3444) );
  MUX2_X1 U15680 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13436), .S(n15740), .Z(
        P3_U3441) );
  INV_X1 U15681 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13438) );
  MUX2_X1 U15682 ( .A(n13438), .B(n13437), .S(n15740), .Z(n13439) );
  OAI21_X1 U15683 ( .B1(n13440), .B2(n13449), .A(n13439), .ZN(P3_U3438) );
  INV_X1 U15684 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13442) );
  MUX2_X1 U15685 ( .A(n13442), .B(n13441), .S(n15740), .Z(n13443) );
  OAI21_X1 U15686 ( .B1(n13444), .B2(n13449), .A(n13443), .ZN(P3_U3435) );
  MUX2_X1 U15687 ( .A(n13445), .B(P3_REG0_REG_14__SCAN_IN), .S(n15742), .Z(
        n13446) );
  INV_X1 U15688 ( .A(n13446), .ZN(n13447) );
  OAI21_X1 U15689 ( .B1(n13449), .B2(n13448), .A(n13447), .ZN(P3_U3432) );
  INV_X1 U15690 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13450) );
  NAND3_X1 U15691 ( .A1(n13450), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13452) );
  OAI22_X1 U15692 ( .A1(n13453), .A2(n13452), .B1(n13451), .B2(n13471), .ZN(
        n13454) );
  AOI21_X1 U15693 ( .B1(n13456), .B2(n13455), .A(n13454), .ZN(n13457) );
  INV_X1 U15694 ( .A(n13457), .ZN(P3_U3264) );
  INV_X1 U15695 ( .A(n13458), .ZN(n13459) );
  OAI222_X1 U15696 ( .A1(n13461), .A2(P3_U3151), .B1(n13471), .B2(n13460), 
        .C1(n13468), .C2(n13459), .ZN(P3_U3265) );
  INV_X1 U15697 ( .A(n13462), .ZN(n13464) );
  OAI222_X1 U15698 ( .A1(n13471), .A2(n13465), .B1(n13468), .B2(n13464), .C1(
        P3_U3151), .C2(n13463), .ZN(P3_U3266) );
  INV_X1 U15699 ( .A(n13466), .ZN(n13467) );
  OAI222_X1 U15700 ( .A1(n13471), .A2(n13470), .B1(P3_U3151), .B2(n13469), 
        .C1(n13468), .C2(n13467), .ZN(P3_U3267) );
  MUX2_X1 U15701 ( .A(n13473), .B(n13472), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3295) );
  XNOR2_X1 U15702 ( .A(n14111), .B(n13525), .ZN(n13524) );
  NAND2_X1 U15703 ( .A1(n13684), .A2(n13922), .ZN(n13523) );
  NOR2_X1 U15704 ( .A1(n13540), .A2(n11160), .ZN(n13512) );
  XNOR2_X1 U15705 ( .A(n14045), .B(n13505), .ZN(n13511) );
  INV_X1 U15706 ( .A(n13474), .ZN(n13475) );
  OR2_X1 U15707 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  XNOR2_X1 U15708 ( .A(n14084), .B(n13525), .ZN(n13616) );
  NAND2_X1 U15709 ( .A1(n13689), .A2(n13922), .ZN(n13479) );
  XNOR2_X1 U15710 ( .A(n13616), .B(n13479), .ZN(n13604) );
  NAND2_X1 U15711 ( .A1(n13616), .A2(n13479), .ZN(n13480) );
  XNOR2_X1 U15712 ( .A(n14079), .B(n13493), .ZN(n13481) );
  NAND2_X1 U15713 ( .A1(n13989), .A2(n13922), .ZN(n13482) );
  XNOR2_X1 U15714 ( .A(n13481), .B(n13482), .ZN(n13614) );
  INV_X1 U15715 ( .A(n13481), .ZN(n13483) );
  NAND2_X1 U15716 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  XNOR2_X1 U15717 ( .A(n13961), .B(n13505), .ZN(n13485) );
  AND2_X1 U15718 ( .A1(n13939), .A2(n13509), .ZN(n13486) );
  NAND2_X1 U15719 ( .A1(n13485), .A2(n13486), .ZN(n13489) );
  INV_X1 U15720 ( .A(n13485), .ZN(n13552) );
  INV_X1 U15721 ( .A(n13486), .ZN(n13487) );
  NAND2_X1 U15722 ( .A1(n13552), .A2(n13487), .ZN(n13488) );
  NAND2_X1 U15723 ( .A1(n13489), .A2(n13488), .ZN(n13654) );
  XNOR2_X1 U15724 ( .A(n13934), .B(n13505), .ZN(n13491) );
  NAND2_X1 U15725 ( .A1(n13920), .A2(n13922), .ZN(n13492) );
  XNOR2_X1 U15726 ( .A(n13491), .B(n13492), .ZN(n13553) );
  AND2_X1 U15727 ( .A1(n13553), .A2(n13489), .ZN(n13490) );
  INV_X1 U15728 ( .A(n13491), .ZN(n13635) );
  XNOR2_X1 U15729 ( .A(n14063), .B(n13493), .ZN(n13494) );
  NAND2_X1 U15730 ( .A1(n13940), .A2(n13922), .ZN(n13495) );
  INV_X1 U15731 ( .A(n13494), .ZN(n13496) );
  NAND2_X1 U15732 ( .A1(n13496), .A2(n13495), .ZN(n13497) );
  NAND2_X1 U15733 ( .A1(n13640), .A2(n13497), .ZN(n13587) );
  INV_X1 U15734 ( .A(n13587), .ZN(n13499) );
  XNOR2_X1 U15735 ( .A(n14120), .B(n13525), .ZN(n13500) );
  NAND2_X1 U15736 ( .A1(n13919), .A2(n13922), .ZN(n13501) );
  XNOR2_X1 U15737 ( .A(n13500), .B(n13501), .ZN(n13588) );
  NAND2_X1 U15738 ( .A1(n13499), .A2(n13498), .ZN(n13585) );
  INV_X1 U15739 ( .A(n13500), .ZN(n13503) );
  INV_X1 U15740 ( .A(n13501), .ZN(n13502) );
  NAND2_X1 U15741 ( .A1(n13503), .A2(n13502), .ZN(n13504) );
  XNOR2_X1 U15742 ( .A(n14118), .B(n13505), .ZN(n13506) );
  AND2_X1 U15743 ( .A1(n13508), .A2(n13506), .ZN(n13536) );
  AOI21_X1 U15744 ( .B1(n13512), .B2(n13511), .A(n13536), .ZN(n13513) );
  INV_X1 U15745 ( .A(n13506), .ZN(n13507) );
  AND2_X1 U15746 ( .A1(n13688), .A2(n13509), .ZN(n13510) );
  INV_X1 U15747 ( .A(n13511), .ZN(n13538) );
  INV_X1 U15748 ( .A(n13512), .ZN(n13543) );
  XNOR2_X1 U15749 ( .A(n14039), .B(n13525), .ZN(n13593) );
  NAND2_X1 U15750 ( .A1(n13686), .A2(n13922), .ZN(n13514) );
  NOR2_X1 U15751 ( .A1(n13593), .A2(n13514), .ZN(n13515) );
  AOI21_X1 U15752 ( .B1(n13593), .B2(n13514), .A(n13515), .ZN(n13623) );
  INV_X1 U15753 ( .A(n13515), .ZN(n13520) );
  XNOR2_X1 U15754 ( .A(n13842), .B(n13525), .ZN(n13516) );
  NOR2_X1 U15755 ( .A1(n13664), .A2(n11160), .ZN(n13517) );
  NAND2_X1 U15756 ( .A1(n13516), .A2(n13517), .ZN(n13521) );
  INV_X1 U15757 ( .A(n13516), .ZN(n13665) );
  INV_X1 U15758 ( .A(n13517), .ZN(n13518) );
  NAND2_X1 U15759 ( .A1(n13665), .A2(n13518), .ZN(n13519) );
  NAND2_X1 U15760 ( .A1(n13521), .A2(n13519), .ZN(n13594) );
  INV_X1 U15761 ( .A(n13521), .ZN(n13522) );
  XNOR2_X1 U15762 ( .A(n13524), .B(n13523), .ZN(n13667) );
  XNOR2_X1 U15763 ( .A(n14107), .B(n13525), .ZN(n13527) );
  NAND2_X1 U15764 ( .A1(n13683), .A2(n13922), .ZN(n13526) );
  NOR2_X1 U15765 ( .A1(n13527), .A2(n13526), .ZN(n13558) );
  AOI21_X1 U15766 ( .B1(n13527), .B2(n13526), .A(n13558), .ZN(n13528) );
  OAI211_X1 U15767 ( .C1(n13529), .C2(n13528), .A(n13560), .B(n13676), .ZN(
        n13533) );
  AOI22_X1 U15768 ( .A1(n13684), .A2(n13659), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13532) );
  AOI22_X1 U15769 ( .A1(n13806), .A2(n13549), .B1(n13649), .B2(n13814), .ZN(
        n13531) );
  NAND2_X1 U15770 ( .A1(n14107), .A2(n13668), .ZN(n13530) );
  NAND4_X1 U15771 ( .A1(n13533), .A2(n13532), .A3(n13531), .A4(n13530), .ZN(
        P2_U3186) );
  OAI22_X1 U15772 ( .A1(n13592), .A2(n15294), .B1(n13534), .B2(n13953), .ZN(
        n13867) );
  AOI22_X1 U15773 ( .A1(n13867), .A2(n13671), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13535) );
  OAI21_X1 U15774 ( .B1(n13874), .B2(n13674), .A(n13535), .ZN(n13542) );
  INV_X1 U15775 ( .A(n13536), .ZN(n13537) );
  NAND2_X1 U15776 ( .A1(n13643), .A2(n13537), .ZN(n13539) );
  XNOR2_X1 U15777 ( .A(n13539), .B(n13538), .ZN(n13544) );
  NOR3_X1 U15778 ( .A1(n13544), .A2(n13540), .A3(n13663), .ZN(n13541) );
  AOI211_X1 U15779 ( .C1(n14045), .C2(n13668), .A(n13542), .B(n13541), .ZN(
        n13546) );
  NAND3_X1 U15780 ( .A1(n13544), .A2(n13676), .A3(n13543), .ZN(n13545) );
  NAND2_X1 U15781 ( .A1(n13546), .A2(n13545), .ZN(P2_U3188) );
  OAI21_X1 U15782 ( .B1(n13553), .B2(n13547), .A(n13637), .ZN(n13548) );
  NAND2_X1 U15783 ( .A1(n13548), .A2(n13676), .ZN(n13557) );
  NAND2_X1 U15784 ( .A1(n13549), .A2(n13940), .ZN(n13550) );
  NAND2_X1 U15785 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13762)
         );
  OAI211_X1 U15786 ( .C1(n13674), .C2(n13935), .A(n13550), .B(n13762), .ZN(
        n13551) );
  AOI21_X1 U15787 ( .B1(n13934), .B2(n13668), .A(n13551), .ZN(n13556) );
  NOR3_X1 U15788 ( .A1(n13553), .A2(n13552), .A3(n13663), .ZN(n13554) );
  OAI21_X1 U15789 ( .B1(n13554), .B2(n13659), .A(n13939), .ZN(n13555) );
  NAND3_X1 U15790 ( .A1(n13557), .A2(n13556), .A3(n13555), .ZN(P2_U3191) );
  INV_X1 U15791 ( .A(n13558), .ZN(n13559) );
  NAND2_X1 U15792 ( .A1(n13560), .A2(n13559), .ZN(n13564) );
  NAND2_X1 U15793 ( .A1(n13806), .A2(n13509), .ZN(n13561) );
  XNOR2_X1 U15794 ( .A(n13561), .B(n13493), .ZN(n13562) );
  XNOR2_X1 U15795 ( .A(n13797), .B(n13562), .ZN(n13563) );
  XNOR2_X1 U15796 ( .A(n13564), .B(n13563), .ZN(n13570) );
  NAND2_X1 U15797 ( .A1(n13682), .A2(n13988), .ZN(n13566) );
  NAND2_X1 U15798 ( .A1(n13683), .A2(n13991), .ZN(n13565) );
  NAND2_X1 U15799 ( .A1(n13566), .A2(n13565), .ZN(n13791) );
  AOI22_X1 U15800 ( .A1(n13791), .A2(n13671), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13567) );
  OAI21_X1 U15801 ( .B1(n13787), .B2(n13674), .A(n13567), .ZN(n13568) );
  AOI21_X1 U15802 ( .B1(n13797), .B2(n13668), .A(n13568), .ZN(n13569) );
  OAI21_X1 U15803 ( .B1(n13570), .B2(n13653), .A(n13569), .ZN(P2_U3192) );
  INV_X1 U15804 ( .A(n13575), .ZN(n13571) );
  NAND3_X1 U15805 ( .A1(n13641), .A2(n13572), .A3(n13571), .ZN(n13581) );
  AOI22_X1 U15806 ( .A1(n13671), .A2(n13573), .B1(n13668), .B2(n12363), .ZN(
        n13580) );
  OAI21_X1 U15807 ( .B1(n13576), .B2(n13575), .A(n13574), .ZN(n13577) );
  AOI22_X1 U15808 ( .A1(n13578), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n13676), 
        .B2(n13577), .ZN(n13579) );
  NAND3_X1 U15809 ( .A1(n13581), .A2(n13580), .A3(n13579), .ZN(P2_U3194) );
  NAND2_X1 U15810 ( .A1(n13688), .A2(n13988), .ZN(n13583) );
  NAND2_X1 U15811 ( .A1(n13940), .A2(n13991), .ZN(n13582) );
  NAND2_X1 U15812 ( .A1(n13583), .A2(n13582), .ZN(n13900) );
  AOI22_X1 U15813 ( .A1(n13900), .A2(n13671), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13584) );
  OAI21_X1 U15814 ( .B1(n13902), .B2(n13674), .A(n13584), .ZN(n13590) );
  INV_X1 U15815 ( .A(n13585), .ZN(n13586) );
  AOI211_X1 U15816 ( .C1(n13588), .C2(n13587), .A(n13653), .B(n13586), .ZN(
        n13589) );
  AOI211_X1 U15817 ( .C1(n14120), .C2(n13668), .A(n13590), .B(n13589), .ZN(
        n13591) );
  INV_X1 U15818 ( .A(n13591), .ZN(P2_U3195) );
  NOR3_X1 U15819 ( .A1(n13593), .A2(n13592), .A3(n13663), .ZN(n13598) );
  AOI21_X1 U15820 ( .B1(n13622), .B2(n13594), .A(n13653), .ZN(n13597) );
  INV_X1 U15821 ( .A(n13595), .ZN(n13596) );
  OAI21_X1 U15822 ( .B1(n13598), .B2(n13597), .A(n13596), .ZN(n13602) );
  AOI22_X1 U15823 ( .A1(n13684), .A2(n13988), .B1(n13991), .B2(n13686), .ZN(
        n13834) );
  OAI22_X1 U15824 ( .A1(n13834), .A2(n13646), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13599), .ZN(n13600) );
  AOI21_X1 U15825 ( .B1(n13840), .B2(n13649), .A(n13600), .ZN(n13601) );
  OAI211_X1 U15826 ( .C1(n13842), .C2(n13662), .A(n13602), .B(n13601), .ZN(
        P2_U3197) );
  AOI21_X1 U15827 ( .B1(n13604), .B2(n13603), .A(n6983), .ZN(n13609) );
  NAND2_X1 U15828 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15257)
         );
  OAI21_X1 U15829 ( .B1(n13630), .B2(n13605), .A(n15257), .ZN(n13607) );
  OAI22_X1 U15830 ( .A1(n13657), .A2(n13952), .B1(n13674), .B2(n13995), .ZN(
        n13606) );
  AOI211_X1 U15831 ( .C1(n14084), .C2(n13668), .A(n13607), .B(n13606), .ZN(
        n13608) );
  OAI21_X1 U15832 ( .B1(n13609), .B2(n13653), .A(n13608), .ZN(P2_U3198) );
  NAND2_X1 U15833 ( .A1(n13939), .A2(n13988), .ZN(n13611) );
  NAND2_X1 U15834 ( .A1(n13689), .A2(n13991), .ZN(n13610) );
  NAND2_X1 U15835 ( .A1(n13611), .A2(n13610), .ZN(n13970) );
  AOI22_X1 U15836 ( .A1(n13671), .A2(n13970), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13612) );
  OAI21_X1 U15837 ( .B1(n13975), .B2(n13674), .A(n13612), .ZN(n13613) );
  AOI21_X1 U15838 ( .B1(n14079), .B2(n13668), .A(n13613), .ZN(n13620) );
  OAI22_X1 U15839 ( .A1(n13616), .A2(n13653), .B1(n13615), .B2(n13663), .ZN(
        n13617) );
  NAND3_X1 U15840 ( .A1(n13618), .A2(n6988), .A3(n13617), .ZN(n13619) );
  OAI211_X1 U15841 ( .C1(n13621), .C2(n13653), .A(n13620), .B(n13619), .ZN(
        P2_U3200) );
  INV_X1 U15842 ( .A(n14039), .ZN(n13858) );
  OAI211_X1 U15843 ( .C1(n13624), .C2(n13623), .A(n13622), .B(n13676), .ZN(
        n13628) );
  AOI22_X1 U15844 ( .A1(n13685), .A2(n13988), .B1(n13991), .B2(n13687), .ZN(
        n13852) );
  OAI22_X1 U15845 ( .A1(n13852), .A2(n13646), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13625), .ZN(n13626) );
  AOI21_X1 U15846 ( .B1(n13856), .B2(n13649), .A(n13626), .ZN(n13627) );
  OAI211_X1 U15847 ( .C1(n13858), .C2(n13662), .A(n13628), .B(n13627), .ZN(
        P2_U3201) );
  OAI22_X1 U15848 ( .A1(n13630), .A2(n13954), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13629), .ZN(n13634) );
  INV_X1 U15849 ( .A(n13924), .ZN(n13631) );
  OAI22_X1 U15850 ( .A1(n13657), .A2(n13632), .B1(n13631), .B2(n13674), .ZN(
        n13633) );
  AOI211_X1 U15851 ( .C1(n14063), .C2(n13668), .A(n13634), .B(n13633), .ZN(
        n13639) );
  OAI22_X1 U15852 ( .A1(n13635), .A2(n13653), .B1(n13954), .B2(n13663), .ZN(
        n13636) );
  NAND3_X1 U15853 ( .A1(n13637), .A2(n6794), .A3(n13636), .ZN(n13638) );
  OAI211_X1 U15854 ( .C1(n13640), .C2(n13653), .A(n13639), .B(n13638), .ZN(
        P2_U3205) );
  AOI22_X1 U15855 ( .A1(n13642), .A2(n13676), .B1(n13641), .B2(n13688), .ZN(
        n13652) );
  INV_X1 U15856 ( .A(n13643), .ZN(n13651) );
  AND2_X1 U15857 ( .A1(n13919), .A2(n13991), .ZN(n13644) );
  AOI21_X1 U15858 ( .B1(n13687), .B2(n13988), .A(n13644), .ZN(n13885) );
  OAI22_X1 U15859 ( .A1(n13885), .A2(n13646), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13645), .ZN(n13648) );
  NOR2_X1 U15860 ( .A1(n13892), .A2(n13662), .ZN(n13647) );
  AOI211_X1 U15861 ( .C1(n13649), .C2(n13893), .A(n13648), .B(n13647), .ZN(
        n13650) );
  OAI21_X1 U15862 ( .B1(n13652), .B2(n13651), .A(n13650), .ZN(P2_U3207) );
  INV_X1 U15863 ( .A(n13961), .ZN(n14133) );
  AOI21_X1 U15864 ( .B1(n13655), .B2(n13654), .A(n13653), .ZN(n13656) );
  NAND2_X1 U15865 ( .A1(n13656), .A2(n13547), .ZN(n13661) );
  AND2_X1 U15866 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13741) );
  OAI22_X1 U15867 ( .A1(n13657), .A2(n13954), .B1(n13674), .B2(n13962), .ZN(
        n13658) );
  AOI211_X1 U15868 ( .C1(n13659), .C2(n13989), .A(n13741), .B(n13658), .ZN(
        n13660) );
  OAI211_X1 U15869 ( .C1(n14133), .C2(n13662), .A(n13661), .B(n13660), .ZN(
        P2_U3210) );
  NOR3_X1 U15870 ( .A1(n13665), .A2(n13664), .A3(n13663), .ZN(n13666) );
  AOI21_X1 U15871 ( .B1(n13595), .B2(n13676), .A(n13666), .ZN(n13679) );
  INV_X1 U15872 ( .A(n13667), .ZN(n13678) );
  NAND2_X1 U15873 ( .A1(n14111), .A2(n13668), .ZN(n13673) );
  NAND2_X1 U15874 ( .A1(n13683), .A2(n13988), .ZN(n13670) );
  NAND2_X1 U15875 ( .A1(n13685), .A2(n13991), .ZN(n13669) );
  NAND2_X1 U15876 ( .A1(n13670), .A2(n13669), .ZN(n13821) );
  AOI22_X1 U15877 ( .A1(n13821), .A2(n13671), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13672) );
  OAI211_X1 U15878 ( .C1(n13674), .C2(n13827), .A(n13673), .B(n13672), .ZN(
        n13675) );
  OAI21_X1 U15879 ( .B1(n13679), .B2(n13678), .A(n13677), .ZN(P2_U3212) );
  INV_X2 U15880 ( .A(P2_U3947), .ZN(n13696) );
  MUX2_X1 U15881 ( .A(n13680), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13696), .Z(
        P2_U3562) );
  MUX2_X1 U15882 ( .A(n13681), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13696), .Z(
        P2_U3561) );
  MUX2_X1 U15883 ( .A(n13682), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13696), .Z(
        P2_U3560) );
  MUX2_X1 U15884 ( .A(n13806), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13696), .Z(
        P2_U3559) );
  MUX2_X1 U15885 ( .A(n13683), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13696), .Z(
        P2_U3558) );
  MUX2_X1 U15886 ( .A(n13684), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13696), .Z(
        P2_U3557) );
  MUX2_X1 U15887 ( .A(n13685), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13696), .Z(
        P2_U3556) );
  MUX2_X1 U15888 ( .A(n13686), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13696), .Z(
        P2_U3555) );
  MUX2_X1 U15889 ( .A(n13687), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13696), .Z(
        P2_U3554) );
  MUX2_X1 U15890 ( .A(n13688), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13696), .Z(
        P2_U3553) );
  MUX2_X1 U15891 ( .A(n13919), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13696), .Z(
        P2_U3552) );
  MUX2_X1 U15892 ( .A(n13940), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13696), .Z(
        P2_U3551) );
  MUX2_X1 U15893 ( .A(n13920), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13696), .Z(
        P2_U3550) );
  MUX2_X1 U15894 ( .A(n13939), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13696), .Z(
        P2_U3549) );
  MUX2_X1 U15895 ( .A(n13989), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13696), .Z(
        P2_U3548) );
  MUX2_X1 U15896 ( .A(n13689), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13696), .Z(
        P2_U3547) );
  MUX2_X1 U15897 ( .A(n13992), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13696), .Z(
        P2_U3546) );
  MUX2_X1 U15898 ( .A(n13690), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13696), .Z(
        P2_U3545) );
  MUX2_X1 U15899 ( .A(n13691), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13696), .Z(
        P2_U3544) );
  MUX2_X1 U15900 ( .A(n13692), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13696), .Z(
        P2_U3543) );
  MUX2_X1 U15901 ( .A(n13693), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13696), .Z(
        P2_U3542) );
  MUX2_X1 U15902 ( .A(n13694), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13696), .Z(
        P2_U3541) );
  MUX2_X1 U15903 ( .A(n13695), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13696), .Z(
        P2_U3540) );
  MUX2_X1 U15904 ( .A(n13697), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13696), .Z(
        P2_U3539) );
  MUX2_X1 U15905 ( .A(n13698), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13696), .Z(
        P2_U3538) );
  MUX2_X1 U15906 ( .A(n13699), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13696), .Z(
        P2_U3537) );
  MUX2_X1 U15907 ( .A(n13700), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13696), .Z(
        P2_U3536) );
  MUX2_X1 U15908 ( .A(n13701), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13696), .Z(
        P2_U3535) );
  MUX2_X1 U15909 ( .A(n13702), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13696), .Z(
        P2_U3534) );
  MUX2_X1 U15910 ( .A(n13703), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13696), .Z(
        P2_U3533) );
  MUX2_X1 U15911 ( .A(n6854), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13696), .Z(
        P2_U3532) );
  MUX2_X1 U15912 ( .A(n13705), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13696), .Z(
        P2_U3531) );
  AOI21_X1 U15913 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(P2_REG2_REG_0__SCAN_IN), 
        .A(n13706), .ZN(n13707) );
  NOR3_X1 U15914 ( .A1(n15221), .A2(n13708), .A3(n13707), .ZN(n13709) );
  AOI21_X1 U15915 ( .B1(n15268), .B2(n13710), .A(n13709), .ZN(n13718) );
  AOI22_X1 U15916 ( .A1(n15266), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n13717) );
  INV_X1 U15917 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15410) );
  MUX2_X1 U15918 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n15412), .S(n13711), .Z(
        n13712) );
  OAI21_X1 U15919 ( .B1(n15410), .B2(n13713), .A(n13712), .ZN(n13714) );
  NAND3_X1 U15920 ( .A1(n15270), .A2(n13715), .A3(n13714), .ZN(n13716) );
  NAND3_X1 U15921 ( .A1(n13718), .A2(n13717), .A3(n13716), .ZN(P2_U3215) );
  NAND2_X1 U15922 ( .A1(n15267), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13729) );
  INV_X1 U15923 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U15924 ( .A1(n13739), .A2(n13720), .ZN(n13719) );
  OAI21_X1 U15925 ( .B1(n13739), .B2(n13720), .A(n13719), .ZN(n13721) );
  INV_X1 U15926 ( .A(n13721), .ZN(n15276) );
  INV_X1 U15927 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13728) );
  XNOR2_X1 U15928 ( .A(n15264), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U15929 ( .A1(n13723), .A2(n13722), .ZN(n13725) );
  NAND2_X1 U15930 ( .A1(n15244), .A2(n13726), .ZN(n13727) );
  NAND2_X1 U15931 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15246), .ZN(n15245) );
  NAND2_X1 U15932 ( .A1(n13727), .A2(n15245), .ZN(n15261) );
  NAND2_X1 U15933 ( .A1(n15260), .A2(n15261), .ZN(n15259) );
  NAND2_X1 U15934 ( .A1(n13729), .A2(n15273), .ZN(n13730) );
  AOI21_X1 U15935 ( .B1(n13731), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13749), 
        .ZN(n13747) );
  INV_X1 U15936 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13738) );
  XNOR2_X1 U15937 ( .A(n13739), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15272) );
  INV_X1 U15938 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13737) );
  XNOR2_X1 U15939 ( .A(n15264), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15254) );
  INV_X1 U15940 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14911) );
  OAI21_X1 U15941 ( .B1(n14911), .B2(n13733), .A(n13732), .ZN(n13734) );
  NAND2_X1 U15942 ( .A1(n15244), .A2(n13734), .ZN(n13736) );
  XNOR2_X1 U15943 ( .A(n13735), .B(n13734), .ZN(n15248) );
  NAND2_X1 U15944 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15248), .ZN(n15247) );
  NAND2_X1 U15945 ( .A1(n13736), .A2(n15247), .ZN(n15255) );
  NAND2_X1 U15946 ( .A1(n15254), .A2(n15255), .ZN(n15253) );
  OAI21_X1 U15947 ( .B1(n15264), .B2(n13737), .A(n15253), .ZN(n15271) );
  NAND2_X1 U15948 ( .A1(n15272), .A2(n15271), .ZN(n15269) );
  OAI21_X1 U15949 ( .B1(n13739), .B2(n13738), .A(n15269), .ZN(n13751) );
  XNOR2_X1 U15950 ( .A(n13744), .B(n13751), .ZN(n13740) );
  NAND2_X1 U15951 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n13740), .ZN(n13753) );
  OAI211_X1 U15952 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13740), .A(n15270), 
        .B(n13753), .ZN(n13743) );
  AOI21_X1 U15953 ( .B1(n15266), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13741), 
        .ZN(n13742) );
  OAI211_X1 U15954 ( .C1(n15265), .C2(n13744), .A(n13743), .B(n13742), .ZN(
        n13745) );
  INV_X1 U15955 ( .A(n13745), .ZN(n13746) );
  OAI21_X1 U15956 ( .B1(n13747), .B2(n15221), .A(n13746), .ZN(P2_U3232) );
  INV_X1 U15957 ( .A(n13758), .ZN(n13756) );
  NAND2_X1 U15958 ( .A1(n13751), .A2(n13750), .ZN(n13752) );
  NAND2_X1 U15959 ( .A1(n13753), .A2(n13752), .ZN(n13754) );
  XOR2_X1 U15960 ( .A(n13754), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13757) );
  OAI21_X1 U15961 ( .B1(n13757), .B2(n15214), .A(n15265), .ZN(n13755) );
  AOI21_X1 U15962 ( .B1(n13756), .B2(n15274), .A(n13755), .ZN(n13761) );
  AOI22_X1 U15963 ( .A1(n13758), .A2(n15274), .B1(n15270), .B2(n13757), .ZN(
        n13760) );
  OAI211_X1 U15964 ( .C1(n7685), .C2(n15231), .A(n13763), .B(n13762), .ZN(
        P2_U3233) );
  NAND2_X1 U15965 ( .A1(n14101), .A2(n13772), .ZN(n13771) );
  XNOR2_X1 U15966 ( .A(n13771), .B(n13765), .ZN(n13766) );
  NAND2_X1 U15967 ( .A1(n14009), .A2(n15285), .ZN(n13770) );
  NOR2_X1 U15968 ( .A1(n13768), .A2(n13767), .ZN(n14008) );
  INV_X1 U15969 ( .A(n14008), .ZN(n14012) );
  NOR2_X1 U15970 ( .A1(n15305), .A2(n14012), .ZN(n13774) );
  AOI21_X1 U15971 ( .B1(n15305), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13774), 
        .ZN(n13769) );
  OAI211_X1 U15972 ( .C1(n14097), .C2(n13998), .A(n13770), .B(n13769), .ZN(
        P2_U3234) );
  OAI211_X1 U15973 ( .C1(n14101), .C2(n13772), .A(n11160), .B(n13771), .ZN(
        n14013) );
  NOR2_X1 U15974 ( .A1(n14101), .A2(n13998), .ZN(n13773) );
  AOI211_X1 U15975 ( .C1(n15305), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13774), 
        .B(n13773), .ZN(n13775) );
  OAI21_X1 U15976 ( .B1(n13907), .B2(n14013), .A(n13775), .ZN(P2_U3235) );
  INV_X1 U15977 ( .A(n13776), .ZN(n13786) );
  NAND2_X1 U15978 ( .A1(n13777), .A2(n15285), .ZN(n13781) );
  INV_X1 U15979 ( .A(n13778), .ZN(n13779) );
  AOI22_X1 U15980 ( .A1(n13779), .A2(n15283), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15305), .ZN(n13780) );
  OAI211_X1 U15981 ( .C1(n13782), .C2(n13998), .A(n13781), .B(n13780), .ZN(
        n13783) );
  AOI21_X1 U15982 ( .B1(n15287), .B2(n13784), .A(n13783), .ZN(n13785) );
  OAI21_X1 U15983 ( .B1(n13786), .B2(n15305), .A(n13785), .ZN(P2_U3236) );
  INV_X1 U15984 ( .A(n13787), .ZN(n13794) );
  OAI211_X1 U15985 ( .C1(n13790), .C2(n13789), .A(n13788), .B(n15293), .ZN(
        n13793) );
  INV_X1 U15986 ( .A(n13791), .ZN(n13792) );
  NAND2_X1 U15987 ( .A1(n13793), .A2(n13792), .ZN(n14016) );
  AOI21_X1 U15988 ( .B1(n13794), .B2(n15283), .A(n14016), .ZN(n13804) );
  INV_X1 U15989 ( .A(n13795), .ZN(n13796) );
  AOI211_X1 U15990 ( .C1(n13797), .C2(n6726), .A(n13922), .B(n13796), .ZN(
        n14017) );
  INV_X1 U15991 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13798) );
  OAI22_X1 U15992 ( .A1(n8246), .A2(n13998), .B1(n15303), .B2(n13798), .ZN(
        n13799) );
  AOI21_X1 U15993 ( .B1(n14017), .B2(n15285), .A(n13799), .ZN(n13803) );
  XNOR2_X1 U15994 ( .A(n13801), .B(n13800), .ZN(n14018) );
  NAND2_X1 U15995 ( .A1(n14018), .A2(n15287), .ZN(n13802) );
  OAI211_X1 U15996 ( .C1(n13804), .C2(n15305), .A(n13803), .B(n13802), .ZN(
        P2_U3237) );
  XNOR2_X1 U15997 ( .A(n13805), .B(n13811), .ZN(n13810) );
  NAND2_X1 U15998 ( .A1(n13806), .A2(n13988), .ZN(n13807) );
  OAI21_X1 U15999 ( .B1(n13808), .B2(n13953), .A(n13807), .ZN(n13809) );
  XNOR2_X1 U16000 ( .A(n13812), .B(n13811), .ZN(n14021) );
  AOI21_X1 U16001 ( .B1(n14107), .B2(n13825), .A(n13922), .ZN(n13813) );
  NAND2_X1 U16002 ( .A1(n13813), .A2(n6726), .ZN(n14022) );
  AOI22_X1 U16003 ( .A1(n13814), .A2(n15283), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15305), .ZN(n13816) );
  NAND2_X1 U16004 ( .A1(n14107), .A2(n15281), .ZN(n13815) );
  OAI211_X1 U16005 ( .C1(n14022), .C2(n13907), .A(n13816), .B(n13815), .ZN(
        n13817) );
  AOI21_X1 U16006 ( .B1(n14021), .B2(n15287), .A(n13817), .ZN(n13818) );
  OAI21_X1 U16007 ( .B1(n14023), .B2(n15305), .A(n13818), .ZN(P2_U3238) );
  INV_X1 U16008 ( .A(n13823), .ZN(n13820) );
  XNOR2_X1 U16009 ( .A(n13819), .B(n13820), .ZN(n13822) );
  XNOR2_X1 U16010 ( .A(n13824), .B(n13823), .ZN(n14027) );
  AOI21_X1 U16011 ( .B1(n14111), .B2(n13837), .A(n13922), .ZN(n13826) );
  NAND2_X1 U16012 ( .A1(n13826), .A2(n13825), .ZN(n14028) );
  INV_X1 U16013 ( .A(n13827), .ZN(n13828) );
  AOI22_X1 U16014 ( .A1(n13828), .A2(n15283), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15305), .ZN(n13830) );
  NAND2_X1 U16015 ( .A1(n14111), .A2(n15281), .ZN(n13829) );
  OAI211_X1 U16016 ( .C1(n14028), .C2(n13907), .A(n13830), .B(n13829), .ZN(
        n13831) );
  AOI21_X1 U16017 ( .B1(n14027), .B2(n15287), .A(n13831), .ZN(n13832) );
  OAI21_X1 U16018 ( .B1(n14030), .B2(n15305), .A(n13832), .ZN(P2_U3239) );
  XNOR2_X1 U16019 ( .A(n13833), .B(n13846), .ZN(n13836) );
  INV_X1 U16020 ( .A(n13834), .ZN(n13835) );
  AOI21_X1 U16021 ( .B1(n13836), .B2(n15293), .A(n13835), .ZN(n14036) );
  INV_X1 U16022 ( .A(n13855), .ZN(n13839) );
  INV_X1 U16023 ( .A(n13837), .ZN(n13838) );
  AOI211_X1 U16024 ( .C1(n14034), .C2(n13839), .A(n13922), .B(n13838), .ZN(
        n14033) );
  AOI22_X1 U16025 ( .A1(n13840), .A2(n15283), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15305), .ZN(n13841) );
  OAI21_X1 U16026 ( .B1(n13842), .B2(n13998), .A(n13841), .ZN(n13848) );
  INV_X1 U16027 ( .A(n13843), .ZN(n13844) );
  AOI21_X1 U16028 ( .B1(n13846), .B2(n13845), .A(n13844), .ZN(n14037) );
  NOR2_X1 U16029 ( .A1(n14037), .A2(n14004), .ZN(n13847) );
  AOI211_X1 U16030 ( .C1(n14033), .C2(n15285), .A(n13848), .B(n13847), .ZN(
        n13849) );
  OAI21_X1 U16031 ( .B1(n15305), .B2(n14036), .A(n13849), .ZN(P2_U3240) );
  XNOR2_X1 U16032 ( .A(n13851), .B(n13850), .ZN(n13854) );
  INV_X1 U16033 ( .A(n13852), .ZN(n13853) );
  AOI21_X1 U16034 ( .B1(n13854), .B2(n15293), .A(n13853), .ZN(n14040) );
  AOI211_X1 U16035 ( .C1(n14039), .C2(n13872), .A(n13922), .B(n13855), .ZN(
        n14038) );
  AOI22_X1 U16036 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(n15305), .B1(n13856), 
        .B2(n15283), .ZN(n13857) );
  OAI21_X1 U16037 ( .B1(n13858), .B2(n13998), .A(n13857), .ZN(n13863) );
  OAI21_X1 U16038 ( .B1(n13861), .B2(n13860), .A(n13859), .ZN(n14042) );
  NOR2_X1 U16039 ( .A1(n14042), .A2(n14004), .ZN(n13862) );
  AOI211_X1 U16040 ( .C1(n14038), .C2(n15285), .A(n13863), .B(n13862), .ZN(
        n13864) );
  OAI21_X1 U16041 ( .B1(n15305), .B2(n14040), .A(n13864), .ZN(P2_U3241) );
  OAI21_X1 U16042 ( .B1(n6778), .B2(n13866), .A(n13865), .ZN(n13868) );
  AOI21_X1 U16043 ( .B1(n13868), .B2(n15293), .A(n13867), .ZN(n14047) );
  OAI21_X1 U16044 ( .B1(n13871), .B2(n13870), .A(n13869), .ZN(n14043) );
  INV_X1 U16045 ( .A(n14045), .ZN(n13878) );
  INV_X1 U16046 ( .A(n13872), .ZN(n13873) );
  AOI211_X1 U16047 ( .C1(n14045), .C2(n13891), .A(n13922), .B(n13873), .ZN(
        n14044) );
  NAND2_X1 U16048 ( .A1(n14044), .A2(n15285), .ZN(n13877) );
  INV_X1 U16049 ( .A(n13874), .ZN(n13875) );
  AOI22_X1 U16050 ( .A1(n15305), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13875), 
        .B2(n15283), .ZN(n13876) );
  OAI211_X1 U16051 ( .C1(n13878), .C2(n13998), .A(n13877), .B(n13876), .ZN(
        n13879) );
  AOI21_X1 U16052 ( .B1(n15287), .B2(n14043), .A(n13879), .ZN(n13880) );
  OAI21_X1 U16053 ( .B1(n14047), .B2(n15305), .A(n13880), .ZN(P2_U3242) );
  NAND2_X1 U16054 ( .A1(n13882), .A2(n13881), .ZN(n13883) );
  NAND3_X1 U16055 ( .A1(n13884), .A2(n15293), .A3(n13883), .ZN(n13886) );
  INV_X1 U16056 ( .A(n13887), .ZN(n13890) );
  NAND2_X1 U16057 ( .A1(n13888), .A2(n8283), .ZN(n13889) );
  NAND2_X1 U16058 ( .A1(n13890), .A2(n13889), .ZN(n14051) );
  INV_X1 U16059 ( .A(n14051), .ZN(n13897) );
  OAI211_X1 U16060 ( .C1(n13906), .C2(n13892), .A(n11160), .B(n13891), .ZN(
        n14049) );
  AOI22_X1 U16061 ( .A1(n15305), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13893), 
        .B2(n15283), .ZN(n13895) );
  NAND2_X1 U16062 ( .A1(n14118), .A2(n15281), .ZN(n13894) );
  OAI211_X1 U16063 ( .C1(n14049), .C2(n13907), .A(n13895), .B(n13894), .ZN(
        n13896) );
  AOI21_X1 U16064 ( .B1(n13897), .B2(n15287), .A(n13896), .ZN(n13898) );
  OAI21_X1 U16065 ( .B1(n14050), .B2(n15305), .A(n13898), .ZN(P2_U3243) );
  XNOR2_X1 U16066 ( .A(n13899), .B(n13910), .ZN(n13901) );
  AOI21_X1 U16067 ( .B1(n13901), .B2(n15293), .A(n13900), .ZN(n14057) );
  INV_X1 U16068 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13903) );
  OAI22_X1 U16069 ( .A1(n15303), .A2(n13903), .B1(n13902), .B2(n15298), .ZN(
        n13909) );
  NAND2_X1 U16070 ( .A1(n6706), .A2(n14120), .ZN(n13904) );
  NAND2_X1 U16071 ( .A1(n13904), .A2(n11160), .ZN(n13905) );
  OR2_X1 U16072 ( .A1(n13906), .A2(n13905), .ZN(n14055) );
  NOR2_X1 U16073 ( .A1(n14055), .A2(n13907), .ZN(n13908) );
  AOI211_X1 U16074 ( .C1(n15281), .C2(n14120), .A(n13909), .B(n13908), .ZN(
        n13913) );
  XNOR2_X1 U16075 ( .A(n13911), .B(n13910), .ZN(n14054) );
  NAND2_X1 U16076 ( .A1(n14054), .A2(n15287), .ZN(n13912) );
  OAI211_X1 U16077 ( .C1(n14057), .C2(n15305), .A(n13913), .B(n13912), .ZN(
        P2_U3244) );
  XNOR2_X1 U16078 ( .A(n13915), .B(n13914), .ZN(n14066) );
  OAI21_X1 U16079 ( .B1(n13918), .B2(n13917), .A(n13916), .ZN(n13921) );
  AOI222_X1 U16080 ( .A1(n13921), .A2(n15293), .B1(n13920), .B2(n13991), .C1(
        n13919), .C2(n13988), .ZN(n14065) );
  INV_X1 U16081 ( .A(n14065), .ZN(n13929) );
  INV_X1 U16082 ( .A(n14063), .ZN(n13927) );
  AOI21_X1 U16083 ( .B1(n13932), .B2(n14063), .A(n13922), .ZN(n13923) );
  AND2_X1 U16084 ( .A1(n13923), .A2(n6706), .ZN(n14062) );
  NAND2_X1 U16085 ( .A1(n14062), .A2(n15285), .ZN(n13926) );
  AOI22_X1 U16086 ( .A1(n15305), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13924), 
        .B2(n15283), .ZN(n13925) );
  OAI211_X1 U16087 ( .C1(n13927), .C2(n13998), .A(n13926), .B(n13925), .ZN(
        n13928) );
  AOI21_X1 U16088 ( .B1(n13929), .B2(n15303), .A(n13928), .ZN(n13930) );
  OAI21_X1 U16089 ( .B1(n14066), .B2(n14004), .A(n13930), .ZN(P2_U3245) );
  XNOR2_X1 U16090 ( .A(n13931), .B(n13943), .ZN(n14067) );
  INV_X1 U16091 ( .A(n13932), .ZN(n13933) );
  AOI211_X1 U16092 ( .C1(n13934), .C2(n13960), .A(n13922), .B(n13933), .ZN(
        n14069) );
  NOR2_X1 U16093 ( .A1(n7200), .A2(n13998), .ZN(n13938) );
  OAI22_X1 U16094 ( .A1(n15303), .A2(n13936), .B1(n13935), .B2(n15298), .ZN(
        n13937) );
  AOI211_X1 U16095 ( .C1(n14069), .C2(n15285), .A(n13938), .B(n13937), .ZN(
        n13948) );
  AOI22_X1 U16096 ( .A1(n13940), .A2(n13988), .B1(n13991), .B2(n13939), .ZN(
        n13946) );
  OAI21_X1 U16097 ( .B1(n13943), .B2(n13942), .A(n13941), .ZN(n13944) );
  NAND2_X1 U16098 ( .A1(n13944), .A2(n15293), .ZN(n13945) );
  NAND2_X1 U16099 ( .A1(n14068), .A2(n15303), .ZN(n13947) );
  OAI211_X1 U16100 ( .C1(n14067), .C2(n15300), .A(n13948), .B(n13947), .ZN(
        P2_U3246) );
  XOR2_X1 U16101 ( .A(n13956), .B(n13949), .Z(n13951) );
  OAI222_X1 U16102 ( .A1(n15294), .A2(n13954), .B1(n13953), .B2(n13952), .C1(
        n13951), .C2(n13950), .ZN(n14072) );
  INV_X1 U16103 ( .A(n14072), .ZN(n13968) );
  INV_X1 U16104 ( .A(n13955), .ZN(n13959) );
  INV_X1 U16105 ( .A(n13956), .ZN(n13958) );
  OAI21_X1 U16106 ( .B1(n13959), .B2(n13958), .A(n13957), .ZN(n14074) );
  AOI211_X1 U16107 ( .C1(n13961), .C2(n13972), .A(n13922), .B(n7201), .ZN(
        n14073) );
  NAND2_X1 U16108 ( .A1(n14073), .A2(n15285), .ZN(n13965) );
  INV_X1 U16109 ( .A(n13962), .ZN(n13963) );
  AOI22_X1 U16110 ( .A1(n15305), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13963), 
        .B2(n15283), .ZN(n13964) );
  OAI211_X1 U16111 ( .C1(n14133), .C2(n13998), .A(n13965), .B(n13964), .ZN(
        n13966) );
  AOI21_X1 U16112 ( .B1(n15287), .B2(n14074), .A(n13966), .ZN(n13967) );
  OAI21_X1 U16113 ( .B1(n13968), .B2(n15305), .A(n13967), .ZN(P2_U3247) );
  XNOR2_X1 U16114 ( .A(n13969), .B(n13979), .ZN(n13971) );
  AOI21_X1 U16115 ( .B1(n13971), .B2(n15293), .A(n13970), .ZN(n14081) );
  INV_X1 U16116 ( .A(n13993), .ZN(n13974) );
  INV_X1 U16117 ( .A(n13972), .ZN(n13973) );
  AOI211_X1 U16118 ( .C1(n14079), .C2(n13974), .A(n13922), .B(n13973), .ZN(
        n14078) );
  INV_X1 U16119 ( .A(n13975), .ZN(n13976) );
  AOI22_X1 U16120 ( .A1(n15305), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13976), 
        .B2(n15283), .ZN(n13977) );
  OAI21_X1 U16121 ( .B1(n13978), .B2(n13998), .A(n13977), .ZN(n13984) );
  OR2_X1 U16122 ( .A1(n13980), .A2(n13979), .ZN(n13981) );
  NAND2_X1 U16123 ( .A1(n13982), .A2(n13981), .ZN(n14082) );
  NOR2_X1 U16124 ( .A1(n14082), .A2(n14004), .ZN(n13983) );
  AOI211_X1 U16125 ( .C1(n14078), .C2(n15285), .A(n13984), .B(n13983), .ZN(
        n13985) );
  OAI21_X1 U16126 ( .B1(n15305), .B2(n14081), .A(n13985), .ZN(P2_U3248) );
  XNOR2_X1 U16127 ( .A(n13987), .B(n13986), .ZN(n13990) );
  AOI222_X1 U16128 ( .A1(n13992), .A2(n13991), .B1(n15293), .B2(n13990), .C1(
        n13989), .C2(n13988), .ZN(n14086) );
  AOI211_X1 U16129 ( .C1(n14084), .C2(n13994), .A(n13922), .B(n13993), .ZN(
        n14083) );
  INV_X1 U16130 ( .A(n14084), .ZN(n13999) );
  INV_X1 U16131 ( .A(n13995), .ZN(n13996) );
  AOI22_X1 U16132 ( .A1(n15305), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13996), 
        .B2(n15283), .ZN(n13997) );
  OAI21_X1 U16133 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n14006) );
  NAND2_X1 U16134 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  NAND2_X1 U16135 ( .A1(n14003), .A2(n14002), .ZN(n14087) );
  NOR2_X1 U16136 ( .A1(n14087), .A2(n14004), .ZN(n14005) );
  AOI211_X1 U16137 ( .C1(n14083), .C2(n15285), .A(n14006), .B(n14005), .ZN(
        n14007) );
  OAI21_X1 U16138 ( .B1(n14086), .B2(n15305), .A(n14007), .ZN(P2_U3249) );
  INV_X1 U16139 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14010) );
  NOR2_X1 U16140 ( .A1(n14009), .A2(n14008), .ZN(n14094) );
  MUX2_X1 U16141 ( .A(n14010), .B(n14094), .S(n15427), .Z(n14011) );
  OAI21_X1 U16142 ( .B1(n14097), .B2(n14077), .A(n14011), .ZN(P2_U3530) );
  INV_X1 U16143 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14014) );
  AND2_X1 U16144 ( .A1(n14013), .A2(n14012), .ZN(n14098) );
  MUX2_X1 U16145 ( .A(n14014), .B(n14098), .S(n15427), .Z(n14015) );
  OAI21_X1 U16146 ( .B1(n14101), .B2(n14077), .A(n14015), .ZN(P2_U3529) );
  INV_X1 U16147 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n14019) );
  MUX2_X1 U16148 ( .A(n14019), .B(n14102), .S(n15427), .Z(n14020) );
  OAI21_X1 U16149 ( .B1(n8246), .B2(n14077), .A(n14020), .ZN(P2_U3527) );
  NAND2_X1 U16150 ( .A1(n14021), .A2(n15390), .ZN(n14024) );
  NAND3_X1 U16151 ( .A1(n14024), .A2(n14023), .A3(n14022), .ZN(n14105) );
  MUX2_X1 U16152 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14105), .S(n15427), .Z(
        n14025) );
  AOI21_X1 U16153 ( .B1(n14059), .B2(n14107), .A(n14025), .ZN(n14026) );
  INV_X1 U16154 ( .A(n14026), .ZN(P2_U3526) );
  NAND2_X1 U16155 ( .A1(n14027), .A2(n15390), .ZN(n14029) );
  NAND3_X1 U16156 ( .A1(n14030), .A2(n14029), .A3(n14028), .ZN(n14109) );
  MUX2_X1 U16157 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14109), .S(n15427), .Z(
        n14031) );
  AOI21_X1 U16158 ( .B1(n14059), .B2(n14111), .A(n14031), .ZN(n14032) );
  INV_X1 U16159 ( .A(n14032), .ZN(P2_U3525) );
  AOI21_X1 U16160 ( .B1(n15392), .B2(n14034), .A(n14033), .ZN(n14035) );
  OAI211_X1 U16161 ( .C1(n14037), .C2(n14093), .A(n14036), .B(n14035), .ZN(
        n14113) );
  MUX2_X1 U16162 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14113), .S(n15427), .Z(
        P2_U3524) );
  AOI21_X1 U16163 ( .B1(n15392), .B2(n14039), .A(n14038), .ZN(n14041) );
  OAI211_X1 U16164 ( .C1(n14093), .C2(n14042), .A(n14041), .B(n14040), .ZN(
        n14114) );
  MUX2_X1 U16165 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14114), .S(n15427), .Z(
        P2_U3523) );
  INV_X1 U16166 ( .A(n14043), .ZN(n14048) );
  AOI21_X1 U16167 ( .B1(n15392), .B2(n14045), .A(n14044), .ZN(n14046) );
  OAI211_X1 U16168 ( .C1(n14093), .C2(n14048), .A(n14047), .B(n14046), .ZN(
        n14115) );
  MUX2_X1 U16169 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14115), .S(n15427), .Z(
        P2_U3522) );
  OAI211_X1 U16170 ( .C1(n14093), .C2(n14051), .A(n14050), .B(n14049), .ZN(
        n14116) );
  MUX2_X1 U16171 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14116), .S(n15427), .Z(
        n14052) );
  AOI21_X1 U16172 ( .B1(n14059), .B2(n14118), .A(n14052), .ZN(n14053) );
  INV_X1 U16173 ( .A(n14053), .ZN(P2_U3521) );
  NAND2_X1 U16174 ( .A1(n14054), .A2(n15390), .ZN(n14056) );
  NAND3_X1 U16175 ( .A1(n14057), .A2(n14056), .A3(n14055), .ZN(n14121) );
  MUX2_X1 U16176 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14121), .S(n15427), .Z(
        n14058) );
  INV_X1 U16177 ( .A(n14058), .ZN(n14061) );
  NAND2_X1 U16178 ( .A1(n14120), .A2(n14059), .ZN(n14060) );
  NAND2_X1 U16179 ( .A1(n14061), .A2(n14060), .ZN(P2_U3520) );
  AOI21_X1 U16180 ( .B1(n15392), .B2(n14063), .A(n14062), .ZN(n14064) );
  OAI211_X1 U16181 ( .C1(n14093), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        n14125) );
  MUX2_X1 U16182 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14125), .S(n15427), .Z(
        P2_U3519) );
  INV_X1 U16183 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14070) );
  AOI211_X1 U16184 ( .C1(n15399), .C2(n6975), .A(n14069), .B(n14068), .ZN(
        n14126) );
  MUX2_X1 U16185 ( .A(n14070), .B(n14126), .S(n15427), .Z(n14071) );
  OAI21_X1 U16186 ( .B1(n7200), .B2(n14077), .A(n14071), .ZN(P2_U3518) );
  AOI211_X1 U16187 ( .C1(n15390), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        n14129) );
  MUX2_X1 U16188 ( .A(n14075), .B(n14129), .S(n15427), .Z(n14076) );
  OAI21_X1 U16189 ( .B1(n14133), .B2(n14077), .A(n14076), .ZN(P2_U3517) );
  AOI21_X1 U16190 ( .B1(n15392), .B2(n14079), .A(n14078), .ZN(n14080) );
  OAI211_X1 U16191 ( .C1(n14082), .C2(n14093), .A(n14081), .B(n14080), .ZN(
        n14134) );
  MUX2_X1 U16192 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14134), .S(n15427), .Z(
        P2_U3516) );
  AOI21_X1 U16193 ( .B1(n15392), .B2(n14084), .A(n14083), .ZN(n14085) );
  OAI211_X1 U16194 ( .C1(n14093), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        n14135) );
  MUX2_X1 U16195 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14135), .S(n15427), .Z(
        P2_U3515) );
  AOI21_X1 U16196 ( .B1(n15392), .B2(n14089), .A(n14088), .ZN(n14090) );
  OAI211_X1 U16197 ( .C1(n14093), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14136) );
  MUX2_X1 U16198 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14136), .S(n15427), .Z(
        P2_U3514) );
  MUX2_X1 U16199 ( .A(n14095), .B(n14094), .S(n15409), .Z(n14096) );
  OAI21_X1 U16200 ( .B1(n14097), .B2(n14132), .A(n14096), .ZN(P2_U3498) );
  MUX2_X1 U16201 ( .A(n14099), .B(n14098), .S(n15409), .Z(n14100) );
  OAI21_X1 U16202 ( .B1(n14101), .B2(n14132), .A(n14100), .ZN(P2_U3497) );
  MUX2_X1 U16203 ( .A(n14103), .B(n14102), .S(n15409), .Z(n14104) );
  MUX2_X1 U16204 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14105), .S(n15409), .Z(
        n14106) );
  AOI21_X1 U16205 ( .B1(n8335), .B2(n14107), .A(n14106), .ZN(n14108) );
  INV_X1 U16206 ( .A(n14108), .ZN(P2_U3494) );
  MUX2_X1 U16207 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14109), .S(n15409), .Z(
        n14110) );
  AOI21_X1 U16208 ( .B1(n8335), .B2(n14111), .A(n14110), .ZN(n14112) );
  INV_X1 U16209 ( .A(n14112), .ZN(P2_U3493) );
  MUX2_X1 U16210 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14113), .S(n15409), .Z(
        P2_U3492) );
  MUX2_X1 U16211 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14114), .S(n15409), .Z(
        P2_U3491) );
  MUX2_X1 U16212 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14115), .S(n15409), .Z(
        P2_U3490) );
  MUX2_X1 U16213 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14116), .S(n15409), .Z(
        n14117) );
  AOI21_X1 U16214 ( .B1(n8335), .B2(n14118), .A(n14117), .ZN(n14119) );
  INV_X1 U16215 ( .A(n14119), .ZN(P2_U3489) );
  INV_X1 U16216 ( .A(n14120), .ZN(n14124) );
  MUX2_X1 U16217 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14121), .S(n15409), .Z(
        n14122) );
  INV_X1 U16218 ( .A(n14122), .ZN(n14123) );
  OAI21_X1 U16219 ( .B1(n14124), .B2(n14132), .A(n14123), .ZN(P2_U3488) );
  MUX2_X1 U16220 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14125), .S(n15409), .Z(
        P2_U3487) );
  INV_X1 U16221 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14127) );
  MUX2_X1 U16222 ( .A(n14127), .B(n14126), .S(n15409), .Z(n14128) );
  OAI21_X1 U16223 ( .B1(n7200), .B2(n14132), .A(n14128), .ZN(P2_U3486) );
  INV_X1 U16224 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14130) );
  MUX2_X1 U16225 ( .A(n14130), .B(n14129), .S(n15409), .Z(n14131) );
  OAI21_X1 U16226 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(P2_U3484) );
  MUX2_X1 U16227 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14134), .S(n15409), .Z(
        P2_U3481) );
  MUX2_X1 U16228 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14135), .S(n15409), .Z(
        P2_U3478) );
  MUX2_X1 U16229 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14136), .S(n15409), .Z(
        P2_U3475) );
  AOI21_X1 U16230 ( .B1(n14138), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14137), 
        .ZN(n14139) );
  OAI21_X1 U16231 ( .B1(n14140), .B2(n14150), .A(n14139), .ZN(P2_U3299) );
  OAI222_X1 U16232 ( .A1(n14152), .A2(n14143), .B1(n14150), .B2(n14142), .C1(
        P2_U3088), .C2(n14141), .ZN(P2_U3300) );
  INV_X1 U16233 ( .A(n14144), .ZN(n14767) );
  OAI222_X1 U16234 ( .A1(P2_U3088), .A2(n14146), .B1(n14150), .B2(n14767), 
        .C1(n14145), .C2(n14152), .ZN(P2_U3301) );
  OAI222_X1 U16235 ( .A1(n14152), .A2(n14151), .B1(n14150), .B2(n14149), .C1(
        P2_U3088), .C2(n14147), .ZN(P2_U3302) );
  INV_X1 U16236 ( .A(n14153), .ZN(n14154) );
  MUX2_X1 U16237 ( .A(n14154), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16238 ( .A(n14496), .ZN(n14158) );
  AOI22_X1 U16239 ( .A1(n14427), .A2(n14565), .B1(n14563), .B2(n14424), .ZN(
        n14486) );
  OAI22_X1 U16240 ( .A1(n14294), .A2(n14486), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14156), .ZN(n14157) );
  AOI21_X1 U16241 ( .B1(n14158), .B2(n14296), .A(n14157), .ZN(n14159) );
  OAI211_X1 U16242 ( .C1(n14495), .C2(n14300), .A(n14160), .B(n14159), .ZN(
        P1_U3214) );
  NAND2_X1 U16243 ( .A1(n14557), .A2(n15116), .ZN(n14705) );
  NAND2_X1 U16244 ( .A1(n14162), .A2(n14161), .ZN(n14190) );
  INV_X1 U16245 ( .A(n14163), .ZN(n14259) );
  INV_X1 U16246 ( .A(n14164), .ZN(n14166) );
  NOR3_X1 U16247 ( .A1(n14259), .A2(n14166), .A3(n14165), .ZN(n14168) );
  INV_X1 U16248 ( .A(n14232), .ZN(n14167) );
  OAI21_X1 U16249 ( .B1(n14168), .B2(n14167), .A(n14951), .ZN(n14175) );
  INV_X1 U16250 ( .A(n14554), .ZN(n14173) );
  NAND2_X1 U16251 ( .A1(n14420), .A2(n14563), .ZN(n14170) );
  NAND2_X1 U16252 ( .A1(n14303), .A2(n14565), .ZN(n14169) );
  AND2_X1 U16253 ( .A1(n14170), .A2(n14169), .ZN(n14706) );
  INV_X1 U16254 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14171) );
  OAI22_X1 U16255 ( .A1(n14294), .A2(n14706), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14171), .ZN(n14172) );
  AOI21_X1 U16256 ( .B1(n14173), .B2(n14296), .A(n14172), .ZN(n14174) );
  OAI211_X1 U16257 ( .C1(n14705), .C2(n14190), .A(n14175), .B(n14174), .ZN(
        P1_U3216) );
  INV_X1 U16258 ( .A(n14728), .ZN(n14615) );
  INV_X1 U16259 ( .A(n14176), .ZN(n14269) );
  OAI21_X1 U16260 ( .B1(n14269), .B2(n14178), .A(n14177), .ZN(n14180) );
  NAND3_X1 U16261 ( .A1(n14180), .A2(n14951), .A3(n14179), .ZN(n14185) );
  OR2_X1 U16262 ( .A1(n14441), .A2(n14401), .ZN(n14182) );
  OR2_X1 U16263 ( .A1(n14416), .A2(n14460), .ZN(n14181) );
  NAND2_X1 U16264 ( .A1(n14182), .A2(n14181), .ZN(n14619) );
  AND2_X1 U16265 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14393) );
  NOR2_X1 U16266 ( .A1(n14958), .A2(n14611), .ZN(n14183) );
  AOI211_X1 U16267 ( .C1(n14619), .C2(n14953), .A(n14393), .B(n14183), .ZN(
        n14184) );
  OAI211_X1 U16268 ( .C1(n14615), .C2(n14300), .A(n14185), .B(n14184), .ZN(
        P1_U3219) );
  INV_X1 U16269 ( .A(n14186), .ZN(n14258) );
  AOI21_X1 U16270 ( .B1(n14188), .B2(n14187), .A(n14258), .ZN(n14194) );
  AOI22_X1 U16271 ( .A1(n14418), .A2(n14563), .B1(n14565), .B2(n14420), .ZN(
        n14580) );
  INV_X1 U16272 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14189) );
  OAI22_X1 U16273 ( .A1(n14580), .A2(n14294), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14189), .ZN(n14192) );
  NAND2_X1 U16274 ( .A1(n14590), .A2(n15116), .ZN(n14717) );
  NOR2_X1 U16275 ( .A1(n14717), .A2(n14190), .ZN(n14191) );
  AOI211_X1 U16276 ( .C1(n14296), .C2(n14589), .A(n14192), .B(n14191), .ZN(
        n14193) );
  OAI21_X1 U16277 ( .B1(n14194), .B2(n14277), .A(n14193), .ZN(P1_U3223) );
  NAND2_X1 U16278 ( .A1(n14308), .A2(n14563), .ZN(n14196) );
  NAND2_X1 U16279 ( .A1(n14306), .A2(n14565), .ZN(n14195) );
  NAND2_X1 U16280 ( .A1(n14196), .A2(n14195), .ZN(n14798) );
  AOI22_X1 U16281 ( .A1(n14953), .A2(n14798), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14197) );
  OAI21_X1 U16282 ( .B1(n14958), .B2(n14799), .A(n14197), .ZN(n14203) );
  INV_X1 U16283 ( .A(n14198), .ZN(n14199) );
  AOI211_X1 U16284 ( .C1(n14201), .C2(n14200), .A(n14277), .B(n14199), .ZN(
        n14202) );
  AOI211_X1 U16285 ( .C1(n14950), .C2(n14801), .A(n14203), .B(n14202), .ZN(
        n14204) );
  INV_X1 U16286 ( .A(n14204), .ZN(P1_U3224) );
  OAI22_X1 U16287 ( .A1(n7399), .A2(n14460), .B1(n14205), .B2(n14401), .ZN(
        n14693) );
  AOI22_X1 U16288 ( .A1(n14953), .A2(n14693), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14206) );
  OAI21_X1 U16289 ( .B1(n14958), .B2(n14521), .A(n14206), .ZN(n14214) );
  INV_X1 U16290 ( .A(n14208), .ZN(n14209) );
  NAND3_X1 U16291 ( .A1(n14207), .A2(n14210), .A3(n14209), .ZN(n14211) );
  AOI21_X1 U16292 ( .B1(n14212), .B2(n14211), .A(n14277), .ZN(n14213) );
  AOI211_X1 U16293 ( .C1(n14950), .C2(n14694), .A(n14214), .B(n14213), .ZN(
        n14215) );
  INV_X1 U16294 ( .A(n14215), .ZN(P1_U3225) );
  XNOR2_X1 U16295 ( .A(n14218), .B(n14217), .ZN(n14219) );
  XNOR2_X1 U16296 ( .A(n14216), .B(n14219), .ZN(n14226) );
  OR2_X1 U16297 ( .A1(n14416), .A2(n14401), .ZN(n14221) );
  NAND2_X1 U16298 ( .A1(n14431), .A2(n14563), .ZN(n14220) );
  AND2_X1 U16299 ( .A1(n14221), .A2(n14220), .ZN(n14959) );
  NAND2_X1 U16300 ( .A1(n14296), .A2(n14647), .ZN(n14222) );
  OAI211_X1 U16301 ( .C1(n14959), .C2(n14294), .A(n14223), .B(n14222), .ZN(
        n14224) );
  AOI21_X1 U16302 ( .B1(n14652), .B2(n14950), .A(n14224), .ZN(n14225) );
  OAI21_X1 U16303 ( .B1(n14226), .B2(n14277), .A(n14225), .ZN(P1_U3228) );
  OAI22_X1 U16304 ( .A1(n14444), .A2(n14460), .B1(n14227), .B2(n14401), .ZN(
        n14534) );
  AOI22_X1 U16305 ( .A1(n14953), .A2(n14534), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14228) );
  OAI21_X1 U16306 ( .B1(n14958), .B2(n14537), .A(n14228), .ZN(n14235) );
  INV_X1 U16307 ( .A(n14229), .ZN(n14230) );
  NAND3_X1 U16308 ( .A1(n14232), .A2(n14231), .A3(n14230), .ZN(n14233) );
  AOI21_X1 U16309 ( .B1(n14207), .B2(n14233), .A(n14277), .ZN(n14234) );
  AOI211_X1 U16310 ( .C1(n14950), .C2(n6677), .A(n14235), .B(n14234), .ZN(
        n14236) );
  INV_X1 U16311 ( .A(n14236), .ZN(P1_U3229) );
  XNOR2_X1 U16312 ( .A(n14238), .B(n14237), .ZN(n14244) );
  AND2_X1 U16313 ( .A1(n14417), .A2(n14563), .ZN(n14239) );
  AOI21_X1 U16314 ( .B1(n14564), .B2(n14565), .A(n14239), .ZN(n14720) );
  AOI22_X1 U16315 ( .A1(n14296), .A2(n14240), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14241) );
  OAI21_X1 U16316 ( .B1(n14720), .B2(n14294), .A(n14241), .ZN(n14242) );
  AOI21_X1 U16317 ( .B1(n14440), .B2(n14950), .A(n14242), .ZN(n14243) );
  OAI21_X1 U16318 ( .B1(n14244), .B2(n14277), .A(n14243), .ZN(P1_U3233) );
  OAI211_X1 U16319 ( .C1(n14247), .C2(n14246), .A(n14923), .B(n14951), .ZN(
        n14254) );
  INV_X1 U16320 ( .A(n14248), .ZN(n14251) );
  NOR2_X1 U16321 ( .A1(n14958), .A2(n14249), .ZN(n14250) );
  AOI211_X1 U16322 ( .C1(n14953), .C2(n14252), .A(n14251), .B(n14250), .ZN(
        n14253) );
  OAI211_X1 U16323 ( .C1(n11302), .C2(n14300), .A(n14254), .B(n14253), .ZN(
        P1_U3234) );
  INV_X1 U16324 ( .A(n14255), .ZN(n14257) );
  NOR3_X1 U16325 ( .A1(n14258), .A2(n14257), .A3(n14256), .ZN(n14260) );
  OAI21_X1 U16326 ( .B1(n14260), .B2(n14259), .A(n14951), .ZN(n14267) );
  NOR2_X1 U16327 ( .A1(n14958), .A2(n14571), .ZN(n14264) );
  OAI22_X1 U16328 ( .A1(n14262), .A2(n14444), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14261), .ZN(n14263) );
  AOI211_X1 U16329 ( .C1(n14265), .C2(n14564), .A(n14264), .B(n14263), .ZN(
        n14266) );
  OAI211_X1 U16330 ( .C1(n14300), .C2(n7346), .A(n14267), .B(n14266), .ZN(
        P1_U3235) );
  AOI21_X1 U16331 ( .B1(n14271), .B2(n14270), .A(n14269), .ZN(n14278) );
  AND2_X1 U16332 ( .A1(n14435), .A2(n14563), .ZN(n14272) );
  AOI21_X1 U16333 ( .B1(n14417), .B2(n14565), .A(n14272), .ZN(n14626) );
  NAND2_X1 U16334 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15040)
         );
  NAND2_X1 U16335 ( .A1(n14296), .A2(n14273), .ZN(n14274) );
  OAI211_X1 U16336 ( .C1(n14626), .C2(n14294), .A(n15040), .B(n14274), .ZN(
        n14275) );
  AOI21_X1 U16337 ( .B1(n14638), .B2(n14950), .A(n14275), .ZN(n14276) );
  OAI21_X1 U16338 ( .B1(n14278), .B2(n14277), .A(n14276), .ZN(P1_U3238) );
  INV_X1 U16339 ( .A(n14688), .ZN(n14288) );
  OAI21_X1 U16340 ( .B1(n14281), .B2(n14280), .A(n14279), .ZN(n14282) );
  NAND2_X1 U16341 ( .A1(n14282), .A2(n14951), .ZN(n14287) );
  INV_X1 U16342 ( .A(n14505), .ZN(n14285) );
  AOI22_X1 U16343 ( .A1(n14426), .A2(n14565), .B1(n14563), .B2(n14445), .ZN(
        n14685) );
  OAI22_X1 U16344 ( .A1(n14294), .A2(n14685), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14283), .ZN(n14284) );
  AOI21_X1 U16345 ( .B1(n14285), .B2(n14296), .A(n14284), .ZN(n14286) );
  OAI211_X1 U16346 ( .C1(n14288), .C2(n14300), .A(n14287), .B(n14286), .ZN(
        P1_U3240) );
  OAI211_X1 U16347 ( .C1(n14291), .C2(n14290), .A(n14289), .B(n14951), .ZN(
        n14299) );
  INV_X1 U16348 ( .A(n14292), .ZN(n14297) );
  NAND2_X1 U16349 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15026)
         );
  OAI21_X1 U16350 ( .B1(n14294), .B2(n14293), .A(n15026), .ZN(n14295) );
  AOI21_X1 U16351 ( .B1(n14297), .B2(n14296), .A(n14295), .ZN(n14298) );
  OAI211_X1 U16352 ( .C1(n14301), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        P1_U3241) );
  MUX2_X1 U16353 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14402), .S(n14319), .Z(
        P1_U3591) );
  MUX2_X1 U16354 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14457), .S(n14319), .Z(
        P1_U3590) );
  MUX2_X1 U16355 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14302), .S(n14319), .Z(
        P1_U3589) );
  MUX2_X1 U16356 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14427), .S(n14319), .Z(
        P1_U3588) );
  MUX2_X1 U16357 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14426), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16358 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14424), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16359 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14445), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16360 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14303), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16361 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14566), .S(n14319), .Z(
        P1_U3583) );
  MUX2_X1 U16362 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14420), .S(n14319), .Z(
        P1_U3582) );
  MUX2_X1 U16363 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14564), .S(n14319), .Z(
        P1_U3581) );
  MUX2_X1 U16364 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14418), .S(n14319), .Z(
        P1_U3580) );
  MUX2_X1 U16365 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14417), .S(n14319), .Z(
        P1_U3579) );
  INV_X1 U16366 ( .A(n14416), .ZN(n14437) );
  MUX2_X1 U16367 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14437), .S(n14319), .Z(
        P1_U3578) );
  MUX2_X1 U16368 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14435), .S(n14319), .Z(
        P1_U3577) );
  MUX2_X1 U16369 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14431), .S(n14319), .Z(
        P1_U3576) );
  MUX2_X1 U16370 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14304), .S(n14319), .Z(
        P1_U3575) );
  MUX2_X1 U16371 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14305), .S(n14319), .Z(
        P1_U3574) );
  MUX2_X1 U16372 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14306), .S(n14319), .Z(
        P1_U3573) );
  MUX2_X1 U16373 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14307), .S(n14319), .Z(
        P1_U3572) );
  MUX2_X1 U16374 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14308), .S(n14319), .Z(
        P1_U3571) );
  MUX2_X1 U16375 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14309), .S(n14319), .Z(
        P1_U3570) );
  MUX2_X1 U16376 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14310), .S(n14319), .Z(
        P1_U3569) );
  MUX2_X1 U16377 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14311), .S(n14319), .Z(
        P1_U3568) );
  MUX2_X1 U16378 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14312), .S(n14319), .Z(
        P1_U3567) );
  MUX2_X1 U16379 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14313), .S(n14319), .Z(
        P1_U3566) );
  MUX2_X1 U16380 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14314), .S(n14319), .Z(
        P1_U3565) );
  MUX2_X1 U16381 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14315), .S(n14319), .Z(
        P1_U3564) );
  MUX2_X1 U16382 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14316), .S(n14319), .Z(
        P1_U3563) );
  MUX2_X1 U16383 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14317), .S(n14319), .Z(
        P1_U3562) );
  MUX2_X1 U16384 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14318), .S(n14319), .Z(
        P1_U3561) );
  MUX2_X1 U16385 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14320), .S(n14319), .Z(
        P1_U3560) );
  INV_X1 U16386 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14322) );
  OAI21_X1 U16387 ( .B1(n15042), .B2(n14322), .A(n14321), .ZN(n14323) );
  AOI21_X1 U16388 ( .B1(n14324), .B2(n14387), .A(n14323), .ZN(n14335) );
  MUX2_X1 U16389 ( .A(n10121), .B(P1_REG1_REG_3__SCAN_IN), .S(n14324), .Z(
        n14327) );
  NAND3_X1 U16390 ( .A1(n14327), .A2(n14326), .A3(n14325), .ZN(n14328) );
  NAND3_X1 U16391 ( .A1(n14383), .A2(n14347), .A3(n14328), .ZN(n14334) );
  OR3_X1 U16392 ( .A1(n14331), .A2(n14330), .A3(n14329), .ZN(n14332) );
  NAND3_X1 U16393 ( .A1(n14389), .A2(n14338), .A3(n14332), .ZN(n14333) );
  NAND3_X1 U16394 ( .A1(n14335), .A2(n14334), .A3(n14333), .ZN(P1_U3246) );
  AND3_X1 U16395 ( .A1(n14338), .A2(n14337), .A3(n14336), .ZN(n14339) );
  NOR3_X1 U16396 ( .A1(n15034), .A2(n14340), .A3(n14339), .ZN(n14341) );
  AOI211_X1 U16397 ( .C1(n14343), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n14342), .B(
        n14341), .ZN(n14353) );
  NAND2_X1 U16398 ( .A1(n14387), .A2(n14344), .ZN(n14352) );
  INV_X1 U16399 ( .A(n14345), .ZN(n14350) );
  NAND3_X1 U16400 ( .A1(n14348), .A2(n14347), .A3(n14346), .ZN(n14349) );
  NAND3_X1 U16401 ( .A1(n14383), .A2(n14350), .A3(n14349), .ZN(n14351) );
  NAND4_X1 U16402 ( .A1(n14354), .A2(n14353), .A3(n14352), .A4(n14351), .ZN(
        P1_U3247) );
  OAI21_X1 U16403 ( .B1(n14357), .B2(n14356), .A(n14355), .ZN(n14358) );
  NAND2_X1 U16404 ( .A1(n14358), .A2(n14383), .ZN(n14371) );
  NAND2_X1 U16405 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14932)
         );
  OAI21_X1 U16406 ( .B1(n15042), .B2(n14359), .A(n14932), .ZN(n14360) );
  AOI21_X1 U16407 ( .B1(n14361), .B2(n14387), .A(n14360), .ZN(n14370) );
  MUX2_X1 U16408 ( .A(n14362), .B(P1_REG2_REG_14__SCAN_IN), .S(n14361), .Z(
        n14365) );
  INV_X1 U16409 ( .A(n14363), .ZN(n14364) );
  NAND2_X1 U16410 ( .A1(n14365), .A2(n14364), .ZN(n14367) );
  OAI211_X1 U16411 ( .C1(n14368), .C2(n14367), .A(n14366), .B(n14389), .ZN(
        n14369) );
  NAND3_X1 U16412 ( .A1(n14371), .A2(n14370), .A3(n14369), .ZN(P1_U3257) );
  INV_X1 U16413 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14965) );
  OAI21_X1 U16414 ( .B1(n14965), .B2(n14373), .A(n14372), .ZN(n14374) );
  XOR2_X1 U16415 ( .A(n14380), .B(n14374), .Z(n15030) );
  NAND2_X1 U16416 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n15030), .ZN(n15029) );
  NAND2_X1 U16417 ( .A1(n14380), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U16418 ( .A1(n14376), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14378) );
  NAND2_X1 U16419 ( .A1(n14378), .A2(n14377), .ZN(n14379) );
  XOR2_X1 U16420 ( .A(n14380), .B(n14379), .Z(n15032) );
  NAND2_X1 U16421 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15032), .ZN(n15031) );
  NAND2_X1 U16422 ( .A1(n14380), .A2(n14379), .ZN(n14381) );
  NAND2_X1 U16423 ( .A1(n15031), .A2(n14381), .ZN(n14382) );
  XOR2_X1 U16424 ( .A(n14382), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14384) );
  AOI22_X1 U16425 ( .A1(n14385), .A2(n14383), .B1(n14389), .B2(n14384), .ZN(
        n14392) );
  INV_X1 U16426 ( .A(n14384), .ZN(n14388) );
  NOR2_X1 U16427 ( .A1(n14385), .A2(n15036), .ZN(n14386) );
  AOI211_X1 U16428 ( .C1(n14389), .C2(n14388), .A(n14387), .B(n14386), .ZN(
        n14391) );
  MUX2_X1 U16429 ( .A(n14392), .B(n14391), .S(n14390), .Z(n14395) );
  INV_X1 U16430 ( .A(n14393), .ZN(n14394) );
  OAI211_X1 U16431 ( .C1(n7683), .C2(n15042), .A(n14395), .B(n14394), .ZN(
        P1_U3262) );
  NOR2_X2 U16432 ( .A1(n14600), .A2(n14590), .ZN(n14568) );
  NAND2_X1 U16433 ( .A1(n14452), .A2(n14666), .ZN(n14405) );
  NOR2_X1 U16434 ( .A1(n14396), .A2(n14405), .ZN(n14406) );
  XNOR2_X1 U16435 ( .A(n14406), .B(n14397), .ZN(n14398) );
  NAND2_X1 U16436 ( .A1(n14398), .A2(n15055), .ZN(n14659) );
  NOR2_X1 U16437 ( .A1(n6679), .A2(n14399), .ZN(n14400) );
  NOR2_X1 U16438 ( .A1(n14401), .A2(n14400), .ZN(n14456) );
  NAND2_X1 U16439 ( .A1(n14456), .A2(n14402), .ZN(n14661) );
  NOR2_X1 U16440 ( .A1(n15074), .A2(n14661), .ZN(n14409) );
  NOR2_X1 U16441 ( .A1(n14660), .A2(n14614), .ZN(n14403) );
  AOI211_X1 U16442 ( .C1(n15074), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14409), 
        .B(n14403), .ZN(n14404) );
  OAI21_X1 U16443 ( .B1(n14659), .B2(n14654), .A(n14404), .ZN(P1_U3263) );
  INV_X1 U16444 ( .A(n14405), .ZN(n14453) );
  INV_X1 U16445 ( .A(n14406), .ZN(n14407) );
  OAI211_X1 U16446 ( .C1(n14663), .C2(n14453), .A(n14407), .B(n15055), .ZN(
        n14662) );
  NOR2_X1 U16447 ( .A1(n14663), .A2(n14614), .ZN(n14408) );
  AOI211_X1 U16448 ( .C1(n15074), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14409), 
        .B(n14408), .ZN(n14410) );
  OAI21_X1 U16449 ( .B1(n14662), .B2(n14654), .A(n14410), .ZN(P1_U3264) );
  INV_X1 U16450 ( .A(n6677), .ZN(n14540) );
  NOR2_X1 U16451 ( .A1(n14940), .A2(n14431), .ZN(n14411) );
  INV_X1 U16452 ( .A(n14413), .ZN(n14414) );
  INV_X1 U16453 ( .A(n14557), .ZN(n14421) );
  INV_X1 U16454 ( .A(n14485), .ZN(n14490) );
  INV_X1 U16455 ( .A(n14629), .ZN(n14438) );
  INV_X1 U16456 ( .A(n14431), .ZN(n14432) );
  NAND2_X1 U16457 ( .A1(n14940), .A2(n14432), .ZN(n14433) );
  NOR2_X1 U16458 ( .A1(n14961), .A2(n14435), .ZN(n14434) );
  NAND2_X1 U16459 ( .A1(n14961), .A2(n14435), .ZN(n14436) );
  INV_X1 U16460 ( .A(n14599), .ZN(n14595) );
  INV_X1 U16461 ( .A(n14584), .ZN(n14442) );
  INV_X1 U16462 ( .A(n14590), .ZN(n14587) );
  INV_X1 U16463 ( .A(n14548), .ZN(n14551) );
  OAI21_X1 U16464 ( .B1(n7399), .B2(n6677), .A(n14535), .ZN(n14527) );
  NAND2_X1 U16465 ( .A1(n14503), .A2(n14507), .ZN(n14502) );
  INV_X1 U16466 ( .A(n14447), .ZN(n14448) );
  INV_X1 U16467 ( .A(n14452), .ZN(n14454) );
  AOI211_X1 U16468 ( .C1(n14455), .C2(n14454), .A(n14630), .B(n14453), .ZN(
        n14668) );
  NAND2_X1 U16469 ( .A1(n14668), .A2(n15058), .ZN(n14465) );
  NAND2_X1 U16470 ( .A1(n14457), .A2(n14456), .ZN(n14664) );
  OAI22_X1 U16471 ( .A1(n14459), .A2(n14664), .B1(n14458), .B2(n14633), .ZN(
        n14463) );
  OR2_X1 U16472 ( .A1(n14461), .A2(n14460), .ZN(n14665) );
  NOR2_X1 U16473 ( .A1(n15074), .A2(n14665), .ZN(n14462) );
  AOI211_X1 U16474 ( .C1(n15074), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14463), 
        .B(n14462), .ZN(n14464) );
  OAI211_X1 U16475 ( .C1(n14666), .C2(n14614), .A(n14465), .B(n14464), .ZN(
        n14466) );
  AOI21_X1 U16476 ( .B1(n14669), .B2(n14528), .A(n14466), .ZN(n14467) );
  OAI21_X1 U16477 ( .B1(n14671), .B2(n15067), .A(n14467), .ZN(P1_U3356) );
  OAI21_X1 U16478 ( .B1(n14472), .B2(n14469), .A(n14468), .ZN(n14471) );
  NAND2_X1 U16479 ( .A1(n14473), .A2(n14472), .ZN(n14672) );
  NAND3_X1 U16480 ( .A1(n7121), .A2(n14656), .A3(n14672), .ZN(n14482) );
  XNOR2_X1 U16481 ( .A(n14479), .B(n14492), .ZN(n14474) );
  AND2_X1 U16482 ( .A1(n14474), .A2(n15055), .ZN(n14673) );
  OAI22_X1 U16483 ( .A1(n14636), .A2(n14476), .B1(n14475), .B2(n14633), .ZN(
        n14477) );
  INV_X1 U16484 ( .A(n14477), .ZN(n14478) );
  OAI21_X1 U16485 ( .B1(n14479), .B2(n14614), .A(n14478), .ZN(n14480) );
  AOI21_X1 U16486 ( .B1(n14673), .B2(n15058), .A(n14480), .ZN(n14481) );
  OAI211_X1 U16487 ( .C1(n15074), .C2(n14676), .A(n14482), .B(n14481), .ZN(
        P1_U3265) );
  OAI21_X1 U16488 ( .B1(n14485), .B2(n14484), .A(n14483), .ZN(n14488) );
  INV_X1 U16489 ( .A(n14486), .ZN(n14487) );
  OAI21_X1 U16490 ( .B1(n14491), .B2(n14490), .A(n14489), .ZN(n14679) );
  NAND2_X1 U16491 ( .A1(n14679), .A2(n14641), .ZN(n14501) );
  INV_X1 U16492 ( .A(n14513), .ZN(n14494) );
  INV_X1 U16493 ( .A(n14492), .ZN(n14493) );
  AOI211_X1 U16494 ( .C1(n14681), .C2(n14494), .A(n14630), .B(n14493), .ZN(
        n14680) );
  NOR2_X1 U16495 ( .A1(n14495), .A2(n14614), .ZN(n14499) );
  OAI22_X1 U16496 ( .A1(n14636), .A2(n14497), .B1(n14496), .B2(n14633), .ZN(
        n14498) );
  AOI211_X1 U16497 ( .C1(n14680), .C2(n15058), .A(n14499), .B(n14498), .ZN(
        n14500) );
  OAI211_X1 U16498 ( .C1(n15074), .C2(n14683), .A(n14501), .B(n14500), .ZN(
        P1_U3266) );
  OAI21_X1 U16499 ( .B1(n14507), .B2(n14503), .A(n14502), .ZN(n14504) );
  NAND2_X1 U16500 ( .A1(n14504), .A2(n14792), .ZN(n14689) );
  OAI211_X1 U16501 ( .C1(n14505), .C2(n14633), .A(n14689), .B(n14685), .ZN(
        n14517) );
  AOI21_X1 U16502 ( .B1(n14508), .B2(n14507), .A(n14506), .ZN(n14509) );
  INV_X1 U16503 ( .A(n14509), .ZN(n14691) );
  AOI22_X1 U16504 ( .A1(n14688), .A2(n15052), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15074), .ZN(n14515) );
  NAND2_X1 U16505 ( .A1(n14688), .A2(n14510), .ZN(n14511) );
  NAND2_X1 U16506 ( .A1(n14511), .A2(n15055), .ZN(n14512) );
  NOR2_X1 U16507 ( .A1(n14513), .A2(n14512), .ZN(n14686) );
  NAND2_X1 U16508 ( .A1(n14686), .A2(n15058), .ZN(n14514) );
  OAI211_X1 U16509 ( .C1(n14691), .C2(n15067), .A(n14515), .B(n14514), .ZN(
        n14516) );
  AOI21_X1 U16510 ( .B1(n14636), .B2(n14517), .A(n14516), .ZN(n14518) );
  INV_X1 U16511 ( .A(n14518), .ZN(P1_U3267) );
  XNOR2_X1 U16512 ( .A(n14519), .B(n14526), .ZN(n14698) );
  XNOR2_X1 U16513 ( .A(n14694), .B(n7179), .ZN(n14520) );
  AND2_X1 U16514 ( .A1(n14520), .A2(n15055), .ZN(n14692) );
  INV_X1 U16515 ( .A(n14693), .ZN(n14522) );
  OAI22_X1 U16516 ( .A1(n15074), .A2(n14522), .B1(n14521), .B2(n14633), .ZN(
        n14523) );
  AOI21_X1 U16517 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n15074), .A(n14523), 
        .ZN(n14524) );
  OAI21_X1 U16518 ( .B1(n7178), .B2(n14614), .A(n14524), .ZN(n14525) );
  AOI21_X1 U16519 ( .B1(n14692), .B2(n15058), .A(n14525), .ZN(n14530) );
  XNOR2_X1 U16520 ( .A(n14527), .B(n14526), .ZN(n14695) );
  NAND2_X1 U16521 ( .A1(n14695), .A2(n14528), .ZN(n14529) );
  OAI211_X1 U16522 ( .C1(n14698), .C2(n15067), .A(n14530), .B(n14529), .ZN(
        P1_U3268) );
  INV_X1 U16523 ( .A(n14531), .ZN(n14533) );
  AOI21_X1 U16524 ( .B1(n14533), .B2(n14532), .A(n15128), .ZN(n14536) );
  AOI21_X1 U16525 ( .B1(n14536), .B2(n14535), .A(n14534), .ZN(n14702) );
  AOI211_X1 U16526 ( .C1(n6677), .C2(n14556), .A(n14630), .B(n7179), .ZN(
        n14699) );
  INV_X1 U16527 ( .A(n14537), .ZN(n14538) );
  AOI22_X1 U16528 ( .A1(n15074), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14538), 
        .B2(n15070), .ZN(n14539) );
  OAI21_X1 U16529 ( .B1(n14540), .B2(n14614), .A(n14539), .ZN(n14546) );
  AOI21_X1 U16530 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14703) );
  NOR2_X1 U16531 ( .A1(n14703), .A2(n14544), .ZN(n14545) );
  AOI211_X1 U16532 ( .C1(n14699), .C2(n15058), .A(n14546), .B(n14545), .ZN(
        n14547) );
  OAI21_X1 U16533 ( .B1(n15074), .B2(n14702), .A(n14547), .ZN(P1_U3269) );
  XNOR2_X1 U16534 ( .A(n14549), .B(n14548), .ZN(n14709) );
  AOI21_X1 U16535 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14553) );
  OR2_X1 U16536 ( .A1(n14553), .A2(n15128), .ZN(n14707) );
  OAI211_X1 U16537 ( .C1(n14633), .C2(n14554), .A(n14707), .B(n14706), .ZN(
        n14560) );
  NAND2_X1 U16538 ( .A1(n14569), .A2(n14557), .ZN(n14555) );
  NAND3_X1 U16539 ( .A1(n14556), .A2(n15055), .A3(n14555), .ZN(n14704) );
  AOI22_X1 U16540 ( .A1(n14557), .A2(n15052), .B1(n15074), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n14558) );
  OAI21_X1 U16541 ( .B1(n14704), .B2(n14654), .A(n14558), .ZN(n14559) );
  AOI21_X1 U16542 ( .B1(n14560), .B2(n14636), .A(n14559), .ZN(n14561) );
  OAI21_X1 U16543 ( .B1(n15067), .B2(n14709), .A(n14561), .ZN(P1_U3270) );
  XNOR2_X1 U16544 ( .A(n14562), .B(n14575), .ZN(n14567) );
  AOI222_X1 U16545 ( .A1(n14792), .A2(n14567), .B1(n14566), .B2(n14565), .C1(
        n14564), .C2(n14563), .ZN(n14713) );
  INV_X1 U16546 ( .A(n14568), .ZN(n14586) );
  INV_X1 U16547 ( .A(n14569), .ZN(n14570) );
  AOI211_X1 U16548 ( .C1(n14711), .C2(n14586), .A(n14630), .B(n14570), .ZN(
        n14710) );
  INV_X1 U16549 ( .A(n14571), .ZN(n14572) );
  AOI22_X1 U16550 ( .A1(n15074), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14572), 
        .B2(n15070), .ZN(n14573) );
  OAI21_X1 U16551 ( .B1(n7346), .B2(n14614), .A(n14573), .ZN(n14577) );
  XOR2_X1 U16552 ( .A(n14575), .B(n14574), .Z(n14714) );
  NOR2_X1 U16553 ( .A1(n14714), .A2(n15067), .ZN(n14576) );
  AOI211_X1 U16554 ( .C1(n14710), .C2(n15058), .A(n14577), .B(n14576), .ZN(
        n14578) );
  OAI21_X1 U16555 ( .B1(n15074), .B2(n14713), .A(n14578), .ZN(P1_U3271) );
  XNOR2_X1 U16556 ( .A(n14579), .B(n14584), .ZN(n14582) );
  INV_X1 U16557 ( .A(n14580), .ZN(n14581) );
  AOI21_X1 U16558 ( .B1(n14582), .B2(n14792), .A(n14581), .ZN(n14718) );
  OAI21_X1 U16559 ( .B1(n14585), .B2(n14584), .A(n14583), .ZN(n14715) );
  INV_X1 U16560 ( .A(n14600), .ZN(n14588) );
  OAI211_X1 U16561 ( .C1(n14588), .C2(n14587), .A(n15055), .B(n14586), .ZN(
        n14716) );
  AOI22_X1 U16562 ( .A1(n14589), .A2(n15070), .B1(n15074), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U16563 ( .A1(n14590), .A2(n15052), .ZN(n14591) );
  OAI211_X1 U16564 ( .C1(n14716), .C2(n14654), .A(n14592), .B(n14591), .ZN(
        n14593) );
  AOI21_X1 U16565 ( .B1(n14715), .B2(n14656), .A(n14593), .ZN(n14594) );
  OAI21_X1 U16566 ( .B1(n15074), .B2(n14718), .A(n14594), .ZN(P1_U3272) );
  XNOR2_X1 U16567 ( .A(n14596), .B(n14595), .ZN(n14726) );
  AOI21_X1 U16568 ( .B1(n14599), .B2(n14598), .A(n14597), .ZN(n14724) );
  OAI211_X1 U16569 ( .C1(n6793), .C2(n14722), .A(n15055), .B(n14600), .ZN(
        n14721) );
  NOR2_X1 U16570 ( .A1(n14721), .A2(n14654), .ZN(n14607) );
  INV_X1 U16571 ( .A(n14720), .ZN(n14604) );
  INV_X1 U16572 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14601) );
  OAI22_X1 U16573 ( .A1(n14602), .A2(n14633), .B1(n14636), .B2(n14601), .ZN(
        n14603) );
  AOI21_X1 U16574 ( .B1(n14604), .B2(n14636), .A(n14603), .ZN(n14605) );
  OAI21_X1 U16575 ( .B1(n14722), .B2(n14614), .A(n14605), .ZN(n14606) );
  AOI211_X1 U16576 ( .C1(n14724), .C2(n14656), .A(n14607), .B(n14606), .ZN(
        n14608) );
  OAI21_X1 U16577 ( .B1(n14726), .B2(n15068), .A(n14608), .ZN(P1_U3273) );
  XNOR2_X1 U16578 ( .A(n14610), .B(n14609), .ZN(n14731) );
  AOI211_X1 U16579 ( .C1(n14728), .C2(n14631), .A(n14630), .B(n6793), .ZN(
        n14727) );
  INV_X1 U16580 ( .A(n14611), .ZN(n14612) );
  AOI22_X1 U16581 ( .A1(n15074), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14612), 
        .B2(n15070), .ZN(n14613) );
  OAI21_X1 U16582 ( .B1(n14615), .B2(n14614), .A(n14613), .ZN(n14622) );
  OAI21_X1 U16583 ( .B1(n14618), .B2(n14617), .A(n14616), .ZN(n14620) );
  AOI21_X1 U16584 ( .B1(n14620), .B2(n14792), .A(n14619), .ZN(n14729) );
  NOR2_X1 U16585 ( .A1(n14729), .A2(n15074), .ZN(n14621) );
  AOI211_X1 U16586 ( .C1(n14727), .C2(n15058), .A(n14622), .B(n14621), .ZN(
        n14623) );
  OAI21_X1 U16587 ( .B1(n15067), .B2(n14731), .A(n14623), .ZN(P1_U3274) );
  XNOR2_X1 U16588 ( .A(n14629), .B(n14624), .ZN(n14625) );
  NAND2_X1 U16589 ( .A1(n14625), .A2(n14792), .ZN(n14627) );
  NAND2_X1 U16590 ( .A1(n14627), .A2(n14626), .ZN(n14737) );
  INV_X1 U16591 ( .A(n14737), .ZN(n14643) );
  XNOR2_X1 U16592 ( .A(n14629), .B(n14628), .ZN(n14733) );
  AOI21_X1 U16593 ( .B1(n14638), .B2(n14650), .A(n14630), .ZN(n14632) );
  NAND2_X1 U16594 ( .A1(n14632), .A2(n14631), .ZN(n14734) );
  OAI22_X1 U16595 ( .A1(n14636), .A2(n14635), .B1(n14634), .B2(n14633), .ZN(
        n14637) );
  AOI21_X1 U16596 ( .B1(n14638), .B2(n15052), .A(n14637), .ZN(n14639) );
  OAI21_X1 U16597 ( .B1(n14734), .B2(n14654), .A(n14639), .ZN(n14640) );
  AOI21_X1 U16598 ( .B1(n14733), .B2(n14641), .A(n14640), .ZN(n14642) );
  OAI21_X1 U16599 ( .B1(n14643), .B2(n15074), .A(n14642), .ZN(P1_U3275) );
  INV_X1 U16600 ( .A(n14959), .ZN(n14646) );
  XOR2_X1 U16601 ( .A(n14644), .B(n14648), .Z(n14645) );
  NOR2_X1 U16602 ( .A1(n14645), .A2(n15128), .ZN(n14962) );
  AOI211_X1 U16603 ( .C1(n15070), .C2(n14647), .A(n14646), .B(n14962), .ZN(
        n14658) );
  XNOR2_X1 U16604 ( .A(n14649), .B(n14648), .ZN(n14964) );
  OAI211_X1 U16605 ( .C1(n14961), .C2(n14651), .A(n15055), .B(n14650), .ZN(
        n14960) );
  AOI22_X1 U16606 ( .A1(n14652), .A2(n15052), .B1(n15074), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n14653) );
  OAI21_X1 U16607 ( .B1(n14960), .B2(n14654), .A(n14653), .ZN(n14655) );
  AOI21_X1 U16608 ( .B1(n14964), .B2(n14656), .A(n14655), .ZN(n14657) );
  OAI21_X1 U16609 ( .B1(n14658), .B2(n15074), .A(n14657), .ZN(P1_U3276) );
  OAI211_X1 U16610 ( .C1(n14660), .C2(n15126), .A(n14659), .B(n14661), .ZN(
        n14739) );
  INV_X2 U16611 ( .A(n15148), .ZN(n15150) );
  MUX2_X1 U16612 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14739), .S(n15150), .Z(
        P1_U3559) );
  OAI211_X1 U16613 ( .C1(n14663), .C2(n15126), .A(n14662), .B(n14661), .ZN(
        n14740) );
  MUX2_X1 U16614 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14740), .S(n15150), .Z(
        P1_U3558) );
  OAI211_X1 U16615 ( .C1(n14666), .C2(n15126), .A(n14665), .B(n14664), .ZN(
        n14667) );
  NAND2_X1 U16616 ( .A1(n14672), .A2(n15134), .ZN(n14677) );
  AOI21_X1 U16617 ( .B1(n15116), .B2(n14674), .A(n14673), .ZN(n14675) );
  MUX2_X1 U16618 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14742), .S(n15150), .Z(
        P1_U3556) );
  INV_X1 U16619 ( .A(n14679), .ZN(n14684) );
  AOI21_X1 U16620 ( .B1(n15116), .B2(n14681), .A(n14680), .ZN(n14682) );
  OAI211_X1 U16621 ( .C1(n14684), .C2(n14732), .A(n14683), .B(n14682), .ZN(
        n14743) );
  MUX2_X1 U16622 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14743), .S(n15150), .Z(
        P1_U3555) );
  INV_X1 U16623 ( .A(n14685), .ZN(n14687) );
  AOI211_X1 U16624 ( .C1(n15116), .C2(n14688), .A(n14687), .B(n14686), .ZN(
        n14690) );
  OAI211_X1 U16625 ( .C1(n14691), .C2(n14732), .A(n14690), .B(n14689), .ZN(
        n14744) );
  MUX2_X1 U16626 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14744), .S(n15150), .Z(
        P1_U3554) );
  AOI211_X1 U16627 ( .C1(n15116), .C2(n14694), .A(n14693), .B(n14692), .ZN(
        n14697) );
  NAND2_X1 U16628 ( .A1(n14695), .A2(n14792), .ZN(n14696) );
  OAI211_X1 U16629 ( .C1(n14698), .C2(n14732), .A(n14697), .B(n14696), .ZN(
        n14745) );
  MUX2_X1 U16630 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14745), .S(n15150), .Z(
        P1_U3553) );
  AOI21_X1 U16631 ( .B1(n15116), .B2(n6677), .A(n14699), .ZN(n14701) );
  OAI211_X1 U16632 ( .C1(n14703), .C2(n14732), .A(n14702), .B(n14701), .ZN(
        n14746) );
  MUX2_X1 U16633 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14746), .S(n15150), .Z(
        P1_U3552) );
  AND4_X1 U16634 ( .A1(n14707), .A2(n14706), .A3(n14705), .A4(n14704), .ZN(
        n14708) );
  OAI21_X1 U16635 ( .B1(n14732), .B2(n14709), .A(n14708), .ZN(n14747) );
  MUX2_X1 U16636 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14747), .S(n15150), .Z(
        P1_U3551) );
  AOI21_X1 U16637 ( .B1(n15116), .B2(n14711), .A(n14710), .ZN(n14712) );
  OAI211_X1 U16638 ( .C1(n14714), .C2(n14732), .A(n14713), .B(n14712), .ZN(
        n14748) );
  MUX2_X1 U16639 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14748), .S(n15150), .Z(
        P1_U3550) );
  NAND2_X1 U16640 ( .A1(n14715), .A2(n15134), .ZN(n14719) );
  NAND4_X1 U16641 ( .A1(n14719), .A2(n14718), .A3(n14717), .A4(n14716), .ZN(
        n14749) );
  MUX2_X1 U16642 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14749), .S(n15150), .Z(
        P1_U3549) );
  OAI211_X1 U16643 ( .C1(n14722), .C2(n15126), .A(n14721), .B(n14720), .ZN(
        n14723) );
  AOI21_X1 U16644 ( .B1(n14724), .B2(n15134), .A(n14723), .ZN(n14725) );
  OAI21_X1 U16645 ( .B1(n15128), .B2(n14726), .A(n14725), .ZN(n14750) );
  MUX2_X1 U16646 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14750), .S(n15150), .Z(
        P1_U3548) );
  AOI21_X1 U16647 ( .B1(n15116), .B2(n14728), .A(n14727), .ZN(n14730) );
  OAI211_X1 U16648 ( .C1(n14732), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14751) );
  MUX2_X1 U16649 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14751), .S(n15150), .Z(
        P1_U3547) );
  AND2_X1 U16650 ( .A1(n14733), .A2(n15134), .ZN(n14738) );
  OAI21_X1 U16651 ( .B1(n14735), .B2(n15126), .A(n14734), .ZN(n14736) );
  MUX2_X1 U16652 ( .A(n14752), .B(P1_REG1_REG_18__SCAN_IN), .S(n15148), .Z(
        P1_U3546) );
  MUX2_X1 U16653 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14739), .S(n15113), .Z(
        P1_U3527) );
  MUX2_X1 U16654 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14740), .S(n15113), .Z(
        P1_U3526) );
  MUX2_X1 U16655 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14742), .S(n15113), .Z(
        P1_U3524) );
  MUX2_X1 U16656 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14743), .S(n15113), .Z(
        P1_U3523) );
  MUX2_X1 U16657 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14744), .S(n15113), .Z(
        P1_U3522) );
  MUX2_X1 U16658 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14745), .S(n15113), .Z(
        P1_U3521) );
  MUX2_X1 U16659 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14746), .S(n15113), .Z(
        P1_U3520) );
  MUX2_X1 U16660 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14747), .S(n15113), .Z(
        P1_U3519) );
  MUX2_X1 U16661 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14748), .S(n15113), .Z(
        P1_U3518) );
  MUX2_X1 U16662 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14749), .S(n15113), .Z(
        P1_U3517) );
  MUX2_X1 U16663 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14750), .S(n15113), .Z(
        P1_U3516) );
  MUX2_X1 U16664 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14751), .S(n15113), .Z(
        P1_U3515) );
  MUX2_X1 U16665 ( .A(n14752), .B(P1_REG0_REG_18__SCAN_IN), .S(n15135), .Z(
        P1_U3513) );
  INV_X1 U16666 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14753) );
  NAND3_X1 U16667 ( .A1(n14753), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14755) );
  OAI22_X1 U16668 ( .A1(n14756), .A2(n14755), .B1(n14754), .B2(n14764), .ZN(
        n14757) );
  AOI21_X1 U16669 ( .B1(n14759), .B2(n14758), .A(n14757), .ZN(n14760) );
  INV_X1 U16670 ( .A(n14760), .ZN(P1_U3324) );
  OAI222_X1 U16671 ( .A1(n14768), .A2(n14763), .B1(P1_U3086), .B2(n14762), 
        .C1(n14761), .C2(n14764), .ZN(P1_U3325) );
  OAI222_X1 U16672 ( .A1(n14768), .A2(n14766), .B1(P1_U3086), .B2(n9782), .C1(
        n14765), .C2(n14764), .ZN(P1_U3326) );
  OAI222_X1 U16673 ( .A1(n14771), .A2(n14770), .B1(P1_U3086), .B2(n14769), 
        .C1(n14768), .C2(n14767), .ZN(P1_U3329) );
  MUX2_X1 U16674 ( .A(n14773), .B(n14772), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16675 ( .A(n14774), .ZN(n14776) );
  MUX2_X1 U16676 ( .A(n14776), .B(n14775), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  XNOR2_X1 U16677 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14777), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16678 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14778) );
  OAI21_X1 U16679 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14778), 
        .ZN(U28) );
  OAI221_X1 U16680 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7686), .C2(n7684), .A(n14779), .ZN(U29) );
  XOR2_X1 U16681 ( .A(n14780), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16682 ( .A(n14782), .B(n14781), .Z(SUB_1596_U57) );
  XNOR2_X1 U16683 ( .A(n14783), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XNOR2_X1 U16684 ( .A(n14785), .B(n14784), .ZN(SUB_1596_U54) );
  AOI21_X1 U16685 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n14789) );
  XOR2_X1 U16686 ( .A(n14789), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16687 ( .A(n14790), .B(n14791), .ZN(n14811) );
  OAI211_X1 U16688 ( .C1(n14795), .C2(n14794), .A(n14793), .B(n14792), .ZN(
        n14796) );
  INV_X1 U16689 ( .A(n14796), .ZN(n14797) );
  AOI211_X1 U16690 ( .C1(n15123), .C2(n14811), .A(n14798), .B(n14797), .ZN(
        n14808) );
  INV_X1 U16691 ( .A(n14799), .ZN(n14800) );
  AOI222_X1 U16692 ( .A1(n14801), .A2(n15052), .B1(n14800), .B2(n15070), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n15074), .ZN(n14806) );
  INV_X1 U16693 ( .A(n14802), .ZN(n14803) );
  OAI211_X1 U16694 ( .C1(n7185), .C2(n14803), .A(n15055), .B(n6806), .ZN(
        n14807) );
  INV_X1 U16695 ( .A(n14807), .ZN(n14804) );
  AOI22_X1 U16696 ( .A1(n14811), .A2(n15059), .B1(n15058), .B2(n14804), .ZN(
        n14805) );
  OAI211_X1 U16697 ( .C1(n15074), .C2(n14808), .A(n14806), .B(n14805), .ZN(
        P1_U3281) );
  OAI21_X1 U16698 ( .B1(n7185), .B2(n15126), .A(n14807), .ZN(n14810) );
  INV_X1 U16699 ( .A(n14808), .ZN(n14809) );
  AOI211_X1 U16700 ( .C1(n15097), .C2(n14811), .A(n14810), .B(n14809), .ZN(
        n14813) );
  AOI22_X1 U16701 ( .A1(n15113), .A2(n14813), .B1(n10980), .B2(n15135), .ZN(
        P1_U3495) );
  AOI22_X1 U16702 ( .A1(n15150), .A2(n14813), .B1(n14812), .B2(n15148), .ZN(
        P1_U3540) );
  XNOR2_X1 U16703 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14814), .ZN(SUB_1596_U63)
         );
  AOI21_X1 U16704 ( .B1(n14817), .B2(n14816), .A(n14815), .ZN(n14831) );
  OAI21_X1 U16705 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14819), .A(n14818), 
        .ZN(n14824) );
  AOI21_X1 U16706 ( .B1(n15581), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14820), 
        .ZN(n14821) );
  OAI21_X1 U16707 ( .B1(n15584), .B2(n14822), .A(n14821), .ZN(n14823) );
  AOI21_X1 U16708 ( .B1(n14824), .B2(n15586), .A(n14823), .ZN(n14830) );
  AOI21_X1 U16709 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14828) );
  OR2_X1 U16710 ( .A1(n14828), .A2(n15549), .ZN(n14829) );
  OAI211_X1 U16711 ( .C1(n14831), .C2(n15594), .A(n14830), .B(n14829), .ZN(
        P3_U3197) );
  AOI21_X1 U16712 ( .B1(n14834), .B2(n14833), .A(n14832), .ZN(n14851) );
  OAI21_X1 U16713 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n14842) );
  AOI21_X1 U16714 ( .B1(n15581), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n14838), 
        .ZN(n14839) );
  OAI21_X1 U16715 ( .B1(n15584), .B2(n14840), .A(n14839), .ZN(n14841) );
  AOI21_X1 U16716 ( .B1(n14842), .B2(n15586), .A(n14841), .ZN(n14850) );
  INV_X1 U16717 ( .A(n14843), .ZN(n14844) );
  NOR2_X1 U16718 ( .A1(n14845), .A2(n14844), .ZN(n14847) );
  AOI21_X1 U16719 ( .B1(n14848), .B2(n14847), .A(n15549), .ZN(n14846) );
  OAI21_X1 U16720 ( .B1(n14848), .B2(n14847), .A(n14846), .ZN(n14849) );
  OAI211_X1 U16721 ( .C1(n14851), .C2(n15594), .A(n14850), .B(n14849), .ZN(
        P3_U3198) );
  AOI21_X1 U16722 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n14868) );
  OAI21_X1 U16723 ( .B1(n14856), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14855), 
        .ZN(n14857) );
  AND2_X1 U16724 ( .A1(n14857), .A2(n15586), .ZN(n14865) );
  AOI211_X1 U16725 ( .C1(n14860), .C2(n14859), .A(n15549), .B(n14858), .ZN(
        n14864) );
  OAI22_X1 U16726 ( .A1(n15584), .A2(n14862), .B1(n14861), .B2(n15519), .ZN(
        n14863) );
  NOR4_X1 U16727 ( .A1(n14866), .A2(n14865), .A3(n14864), .A4(n14863), .ZN(
        n14867) );
  OAI21_X1 U16728 ( .B1(n14868), .B2(n15594), .A(n14867), .ZN(P3_U3199) );
  AOI22_X1 U16729 ( .A1(n14870), .A2(n14869), .B1(n15581), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14885) );
  OAI21_X1 U16730 ( .B1(n14873), .B2(n14872), .A(n14871), .ZN(n14878) );
  OAI21_X1 U16731 ( .B1(n14876), .B2(n14875), .A(n14874), .ZN(n14877) );
  AOI22_X1 U16732 ( .A1(n14878), .A2(n15586), .B1(n15588), .B2(n14877), .ZN(
        n14884) );
  NAND2_X1 U16733 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14883)
         );
  AOI21_X1 U16734 ( .B1(n14887), .B2(n15732), .A(n14886), .ZN(n14888) );
  AND2_X1 U16735 ( .A1(n14889), .A2(n14888), .ZN(n14900) );
  INV_X1 U16736 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U16737 ( .A1(n15764), .A2(n14900), .B1(n14890), .B2(n15761), .ZN(
        P3_U3472) );
  AOI21_X1 U16738 ( .B1(n14892), .B2(n15732), .A(n14891), .ZN(n14893) );
  AND2_X1 U16739 ( .A1(n14894), .A2(n14893), .ZN(n14902) );
  AOI22_X1 U16740 ( .A1(n15764), .A2(n14902), .B1(n14895), .B2(n15761), .ZN(
        P3_U3471) );
  AOI211_X1 U16741 ( .C1(n14898), .C2(n15732), .A(n14897), .B(n14896), .ZN(
        n14904) );
  INV_X1 U16742 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U16743 ( .A1(n15764), .A2(n14904), .B1(n14899), .B2(n15761), .ZN(
        P3_U3470) );
  INV_X1 U16744 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14901) );
  AOI22_X1 U16745 ( .A1(n15742), .A2(n14901), .B1(n14900), .B2(n15740), .ZN(
        P3_U3429) );
  INV_X1 U16746 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14903) );
  AOI22_X1 U16747 ( .A1(n15742), .A2(n14903), .B1(n14902), .B2(n15740), .ZN(
        P3_U3426) );
  INV_X1 U16748 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U16749 ( .A1(n15742), .A2(n14905), .B1(n14904), .B2(n15740), .ZN(
        P3_U3423) );
  OAI21_X1 U16750 ( .B1(n14907), .B2(n15403), .A(n14906), .ZN(n14909) );
  AOI211_X1 U16751 ( .C1(n14910), .C2(n15390), .A(n14909), .B(n14908), .ZN(
        n14920) );
  AOI22_X1 U16752 ( .A1(n15427), .A2(n14920), .B1(n14911), .B2(n15424), .ZN(
        P2_U3513) );
  NAND2_X1 U16753 ( .A1(n14912), .A2(n15392), .ZN(n14913) );
  NAND2_X1 U16754 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  AOI21_X1 U16755 ( .B1(n14916), .B2(n15390), .A(n14915), .ZN(n14917) );
  AOI22_X1 U16756 ( .A1(n15427), .A2(n14922), .B1(n15211), .B2(n15424), .ZN(
        P2_U3511) );
  INV_X1 U16757 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14919) );
  AOI22_X1 U16758 ( .A1(n15409), .A2(n14920), .B1(n14919), .B2(n15407), .ZN(
        P2_U3472) );
  INV_X1 U16759 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U16760 ( .A1(n15409), .A2(n14922), .B1(n14921), .B2(n15407), .ZN(
        P2_U3466) );
  INV_X1 U16761 ( .A(n14923), .ZN(n14926) );
  OAI21_X1 U16762 ( .B1(n14926), .B2(n14925), .A(n14924), .ZN(n14928) );
  NAND2_X1 U16763 ( .A1(n14928), .A2(n14927), .ZN(n14930) );
  AOI222_X1 U16764 ( .A1(n14931), .A2(n14953), .B1(n14930), .B2(n14951), .C1(
        n14929), .C2(n14950), .ZN(n14933) );
  OAI211_X1 U16765 ( .C1(n14958), .C2(n14934), .A(n14933), .B(n14932), .ZN(
        P1_U3215) );
  INV_X1 U16766 ( .A(n14289), .ZN(n14937) );
  OAI21_X1 U16767 ( .B1(n14937), .B2(n14936), .A(n14935), .ZN(n14939) );
  NAND2_X1 U16768 ( .A1(n14939), .A2(n14938), .ZN(n14941) );
  AOI222_X1 U16769 ( .A1(n14942), .A2(n14953), .B1(n14941), .B2(n14951), .C1(
        n14940), .C2(n14950), .ZN(n14944) );
  OAI211_X1 U16770 ( .C1(n14958), .C2(n14945), .A(n14944), .B(n14943), .ZN(
        P1_U3226) );
  AND2_X1 U16771 ( .A1(n12692), .A2(n14946), .ZN(n14949) );
  OAI21_X1 U16772 ( .B1(n14949), .B2(n14948), .A(n14947), .ZN(n14952) );
  AOI222_X1 U16773 ( .A1(n14954), .A2(n14953), .B1(n14952), .B2(n14951), .C1(
        n14986), .C2(n14950), .ZN(n14956) );
  OAI211_X1 U16774 ( .C1(n14958), .C2(n14957), .A(n14956), .B(n14955), .ZN(
        P1_U3236) );
  OAI211_X1 U16775 ( .C1(n14961), .C2(n15126), .A(n14960), .B(n14959), .ZN(
        n14963) );
  AOI211_X1 U16776 ( .C1(n14964), .C2(n15134), .A(n14963), .B(n14962), .ZN(
        n14993) );
  AOI22_X1 U16777 ( .A1(n15150), .A2(n14993), .B1(n14965), .B2(n15148), .ZN(
        P1_U3545) );
  OAI21_X1 U16778 ( .B1(n14967), .B2(n15126), .A(n14966), .ZN(n14969) );
  AOI211_X1 U16779 ( .C1(n14970), .C2(n15134), .A(n14969), .B(n14968), .ZN(
        n14995) );
  AOI22_X1 U16780 ( .A1(n15150), .A2(n14995), .B1(n11172), .B2(n15148), .ZN(
        P1_U3544) );
  NAND3_X1 U16781 ( .A1(n14972), .A2(n14971), .A3(n15134), .ZN(n14974) );
  OAI211_X1 U16782 ( .C1(n14975), .C2(n15126), .A(n14974), .B(n14973), .ZN(
        n14976) );
  NOR2_X1 U16783 ( .A1(n14977), .A2(n14976), .ZN(n14997) );
  AOI22_X1 U16784 ( .A1(n15150), .A2(n14997), .B1(n14978), .B2(n15148), .ZN(
        P1_U3542) );
  AND2_X1 U16785 ( .A1(n14979), .A2(n15134), .ZN(n14982) );
  OAI21_X1 U16786 ( .B1(n11302), .B2(n15126), .A(n14980), .ZN(n14981) );
  NOR3_X1 U16787 ( .A1(n14983), .A2(n14982), .A3(n14981), .ZN(n14998) );
  AOI22_X1 U16788 ( .A1(n15150), .A2(n14998), .B1(n14984), .B2(n15148), .ZN(
        P1_U3541) );
  AND2_X1 U16789 ( .A1(n14985), .A2(n15134), .ZN(n14990) );
  INV_X1 U16790 ( .A(n14986), .ZN(n14988) );
  OAI21_X1 U16791 ( .B1(n14988), .B2(n15126), .A(n14987), .ZN(n14989) );
  NOR3_X1 U16792 ( .A1(n14991), .A2(n14990), .A3(n14989), .ZN(n14999) );
  AOI22_X1 U16793 ( .A1(n15150), .A2(n14999), .B1(n10956), .B2(n15148), .ZN(
        P1_U3539) );
  INV_X1 U16794 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16795 ( .A1(n15113), .A2(n14993), .B1(n14992), .B2(n15135), .ZN(
        P1_U3510) );
  INV_X1 U16796 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U16797 ( .A1(n15113), .A2(n14995), .B1(n14994), .B2(n15135), .ZN(
        P1_U3507) );
  INV_X1 U16798 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U16799 ( .A1(n15113), .A2(n14997), .B1(n14996), .B2(n15135), .ZN(
        P1_U3501) );
  AOI22_X1 U16800 ( .A1(n15113), .A2(n14998), .B1(n11284), .B2(n15135), .ZN(
        P1_U3498) );
  AOI22_X1 U16801 ( .A1(n15113), .A2(n14999), .B1(n10955), .B2(n15135), .ZN(
        P1_U3492) );
  NOR2_X1 U16802 ( .A1(n15001), .A2(n6683), .ZN(n15002) );
  XOR2_X1 U16803 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15002), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16804 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15006) );
  XOR2_X1 U16805 ( .A(n15006), .B(P2_ADDR_REG_12__SCAN_IN), .Z(SUB_1596_U68)
         );
  AOI21_X1 U16806 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15010) );
  XOR2_X1 U16807 ( .A(n15010), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16808 ( .A1(n15012), .A2(n15011), .ZN(n15013) );
  XOR2_X1 U16809 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n15013), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16810 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  XOR2_X1 U16811 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15016), .Z(SUB_1596_U65)
         );
  XOR2_X1 U16812 ( .A(n15017), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16813 ( .B1(n15019), .B2(P1_REG1_REG_15__SCAN_IN), .A(n15018), 
        .ZN(n15023) );
  AOI21_X1 U16814 ( .B1(n15021), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15020), 
        .ZN(n15022) );
  OAI222_X1 U16815 ( .A1(n15038), .A2(n15024), .B1(n15036), .B2(n15023), .C1(
        n15034), .C2(n15022), .ZN(n15025) );
  INV_X1 U16816 ( .A(n15025), .ZN(n15027) );
  OAI211_X1 U16817 ( .C1(n15028), .C2(n15042), .A(n15027), .B(n15026), .ZN(
        P1_U3258) );
  OAI21_X1 U16818 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n15030), .A(n15029), 
        .ZN(n15035) );
  OAI21_X1 U16819 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n15032), .A(n15031), 
        .ZN(n15033) );
  OAI222_X1 U16820 ( .A1(n15038), .A2(n15037), .B1(n15036), .B2(n15035), .C1(
        n15034), .C2(n15033), .ZN(n15039) );
  INV_X1 U16821 ( .A(n15039), .ZN(n15041) );
  OAI211_X1 U16822 ( .C1(n15043), .C2(n15042), .A(n15041), .B(n15040), .ZN(
        P1_U3261) );
  XNOR2_X1 U16823 ( .A(n15044), .B(n15045), .ZN(n15096) );
  XNOR2_X1 U16824 ( .A(n15046), .B(n15045), .ZN(n15047) );
  NOR2_X1 U16825 ( .A1(n15047), .A2(n15128), .ZN(n15048) );
  AOI211_X1 U16826 ( .C1(n15096), .C2(n15123), .A(n15049), .B(n15048), .ZN(
        n15093) );
  INV_X1 U16827 ( .A(n15050), .ZN(n15051) );
  AOI222_X1 U16828 ( .A1(n15053), .A2(n15052), .B1(n15051), .B2(n15070), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(n15074), .ZN(n15061) );
  OAI211_X1 U16829 ( .C1(n15092), .C2(n15056), .A(n15055), .B(n15054), .ZN(
        n15091) );
  INV_X1 U16830 ( .A(n15091), .ZN(n15057) );
  AOI22_X1 U16831 ( .A1(n15096), .A2(n15059), .B1(n15058), .B2(n15057), .ZN(
        n15060) );
  OAI211_X1 U16832 ( .C1(n15074), .C2(n15093), .A(n15061), .B(n15060), .ZN(
        P1_U3287) );
  INV_X1 U16833 ( .A(n15062), .ZN(n15065) );
  AOI21_X1 U16834 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15073) );
  AOI21_X1 U16835 ( .B1(n15068), .B2(n15067), .A(n15066), .ZN(n15069) );
  AOI21_X1 U16836 ( .B1(n15070), .B2(P1_REG3_REG_0__SCAN_IN), .A(n15069), .ZN(
        n15071) );
  OAI221_X1 U16837 ( .B1(n15074), .B2(n15073), .C1(n14636), .C2(n15072), .A(
        n15071), .ZN(P1_U3293) );
  AND2_X1 U16838 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15075), .ZN(P1_U3294) );
  AND2_X1 U16839 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15075), .ZN(P1_U3295) );
  AND2_X1 U16840 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15075), .ZN(P1_U3296) );
  AND2_X1 U16841 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15075), .ZN(P1_U3297) );
  AND2_X1 U16842 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15075), .ZN(P1_U3298) );
  AND2_X1 U16843 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15075), .ZN(P1_U3299) );
  AND2_X1 U16844 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15075), .ZN(P1_U3300) );
  AND2_X1 U16845 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15075), .ZN(P1_U3301) );
  AND2_X1 U16846 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15075), .ZN(P1_U3302) );
  AND2_X1 U16847 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15075), .ZN(P1_U3303) );
  AND2_X1 U16848 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15075), .ZN(P1_U3304) );
  AND2_X1 U16849 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15075), .ZN(P1_U3305) );
  AND2_X1 U16850 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15075), .ZN(P1_U3306) );
  AND2_X1 U16851 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15075), .ZN(P1_U3307) );
  AND2_X1 U16852 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15075), .ZN(P1_U3308) );
  AND2_X1 U16853 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15075), .ZN(P1_U3309) );
  AND2_X1 U16854 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15075), .ZN(P1_U3310) );
  AND2_X1 U16855 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15075), .ZN(P1_U3311) );
  AND2_X1 U16856 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15075), .ZN(P1_U3312) );
  AND2_X1 U16857 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15075), .ZN(P1_U3313) );
  AND2_X1 U16858 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15075), .ZN(P1_U3314) );
  AND2_X1 U16859 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15075), .ZN(P1_U3315) );
  AND2_X1 U16860 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15075), .ZN(P1_U3316) );
  AND2_X1 U16861 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15075), .ZN(P1_U3317) );
  AND2_X1 U16862 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15075), .ZN(P1_U3318) );
  AND2_X1 U16863 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15075), .ZN(P1_U3319) );
  AND2_X1 U16864 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15075), .ZN(P1_U3320) );
  AND2_X1 U16865 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15075), .ZN(P1_U3321) );
  AND2_X1 U16866 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15075), .ZN(P1_U3322) );
  AND2_X1 U16867 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15075), .ZN(P1_U3323) );
  AOI21_X1 U16868 ( .B1(n15077), .B2(n15116), .A(n15076), .ZN(n15079) );
  NAND3_X1 U16869 ( .A1(n15080), .A2(n15079), .A3(n15078), .ZN(n15081) );
  AOI21_X1 U16870 ( .B1(n15082), .B2(n15134), .A(n15081), .ZN(n15137) );
  INV_X1 U16871 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U16872 ( .A1(n15113), .A2(n15137), .B1(n15083), .B2(n15135), .ZN(
        P1_U3471) );
  NAND2_X1 U16873 ( .A1(n15090), .A2(n15097), .ZN(n15088) );
  NAND2_X1 U16874 ( .A1(n15084), .A2(n15116), .ZN(n15085) );
  NAND4_X1 U16875 ( .A1(n15088), .A2(n15087), .A3(n15086), .A4(n15085), .ZN(
        n15089) );
  AOI21_X1 U16876 ( .B1(n15123), .B2(n15090), .A(n15089), .ZN(n15139) );
  AOI22_X1 U16877 ( .A1(n15113), .A2(n15139), .B1(n10429), .B2(n15135), .ZN(
        P1_U3474) );
  OAI21_X1 U16878 ( .B1(n15092), .B2(n15126), .A(n15091), .ZN(n15095) );
  INV_X1 U16879 ( .A(n15093), .ZN(n15094) );
  AOI211_X1 U16880 ( .C1(n15097), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15141) );
  AOI22_X1 U16881 ( .A1(n15113), .A2(n15141), .B1(n10595), .B2(n15135), .ZN(
        P1_U3477) );
  NAND2_X1 U16882 ( .A1(n15098), .A2(n15123), .ZN(n15104) );
  NAND2_X1 U16883 ( .A1(n15098), .A2(n15097), .ZN(n15103) );
  OAI21_X1 U16884 ( .B1(n7176), .B2(n15126), .A(n15099), .ZN(n15100) );
  NOR2_X1 U16885 ( .A1(n15101), .A2(n15100), .ZN(n15102) );
  AOI22_X1 U16886 ( .A1(n15113), .A2(n15143), .B1(n10723), .B2(n15135), .ZN(
        P1_U3480) );
  AOI211_X1 U16887 ( .C1(n15116), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15108) );
  OAI21_X1 U16888 ( .B1(n15128), .B2(n15109), .A(n15108), .ZN(n15110) );
  AOI21_X1 U16889 ( .B1(n15111), .B2(n15134), .A(n15110), .ZN(n15145) );
  INV_X1 U16890 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U16891 ( .A1(n15113), .A2(n15145), .B1(n15112), .B2(n15135), .ZN(
        P1_U3483) );
  AOI21_X1 U16892 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(n15117) );
  OAI211_X1 U16893 ( .C1(n15120), .C2(n15119), .A(n15118), .B(n15117), .ZN(
        n15121) );
  AOI21_X1 U16894 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15147) );
  AOI22_X1 U16895 ( .A1(n15113), .A2(n15147), .B1(n10926), .B2(n15135), .ZN(
        P1_U3486) );
  OAI211_X1 U16896 ( .C1(n15127), .C2(n15126), .A(n15125), .B(n15124), .ZN(
        n15132) );
  NOR3_X1 U16897 ( .A1(n15130), .A2(n15129), .A3(n15128), .ZN(n15131) );
  AOI211_X1 U16898 ( .C1(n15134), .C2(n15133), .A(n15132), .B(n15131), .ZN(
        n15149) );
  AOI22_X1 U16899 ( .A1(n15113), .A2(n15149), .B1(n10941), .B2(n15135), .ZN(
        P1_U3489) );
  AOI22_X1 U16900 ( .A1(n15150), .A2(n15137), .B1(n15136), .B2(n15148), .ZN(
        P1_U3532) );
  AOI22_X1 U16901 ( .A1(n15150), .A2(n15139), .B1(n15138), .B2(n15148), .ZN(
        P1_U3533) );
  AOI22_X1 U16902 ( .A1(n15150), .A2(n15141), .B1(n15140), .B2(n15148), .ZN(
        P1_U3534) );
  AOI22_X1 U16903 ( .A1(n15150), .A2(n15143), .B1(n15142), .B2(n15148), .ZN(
        P1_U3535) );
  AOI22_X1 U16904 ( .A1(n15150), .A2(n15145), .B1(n15144), .B2(n15148), .ZN(
        P1_U3536) );
  AOI22_X1 U16905 ( .A1(n15150), .A2(n15147), .B1(n15146), .B2(n15148), .ZN(
        P1_U3537) );
  AOI22_X1 U16906 ( .A1(n15150), .A2(n15149), .B1(n9660), .B2(n15148), .ZN(
        P1_U3538) );
  NOR2_X1 U16907 ( .A1(n15266), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16908 ( .A(n15151), .ZN(n15166) );
  OAI21_X1 U16909 ( .B1(n15166), .B2(n15152), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15153) );
  OAI21_X1 U16910 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15153), .ZN(n15164) );
  XOR2_X1 U16911 ( .A(n15155), .B(n15154), .Z(n15156) );
  NAND2_X1 U16912 ( .A1(n15270), .A2(n15156), .ZN(n15163) );
  NAND2_X1 U16913 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n15266), .ZN(n15162) );
  AOI211_X1 U16914 ( .C1(n15159), .C2(n15158), .A(n15157), .B(n15221), .ZN(
        n15160) );
  INV_X1 U16915 ( .A(n15160), .ZN(n15161) );
  NAND4_X1 U16916 ( .A1(n15164), .A2(n15163), .A3(n15162), .A4(n15161), .ZN(
        P2_U3216) );
  OAI21_X1 U16917 ( .B1(n15166), .B2(n15165), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15167) );
  OAI21_X1 U16918 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15167), .ZN(n15179) );
  AOI211_X1 U16919 ( .C1(n15170), .C2(n15169), .A(n15168), .B(n15221), .ZN(
        n15171) );
  INV_X1 U16920 ( .A(n15171), .ZN(n15178) );
  NAND2_X1 U16921 ( .A1(n15173), .A2(n15172), .ZN(n15174) );
  NAND3_X1 U16922 ( .A1(n15270), .A2(n15175), .A3(n15174), .ZN(n15177) );
  NAND2_X1 U16923 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15266), .ZN(n15176) );
  NAND4_X1 U16924 ( .A1(n15179), .A2(n15178), .A3(n15177), .A4(n15176), .ZN(
        P2_U3217) );
  NAND2_X1 U16925 ( .A1(n15266), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n15180) );
  OAI211_X1 U16926 ( .C1(n15265), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15183) );
  INV_X1 U16927 ( .A(n15183), .ZN(n15194) );
  NAND2_X1 U16928 ( .A1(n15185), .A2(n15184), .ZN(n15186) );
  NAND3_X1 U16929 ( .A1(n15187), .A2(n15274), .A3(n15186), .ZN(n15193) );
  NAND2_X1 U16930 ( .A1(n15189), .A2(n15188), .ZN(n15190) );
  NAND3_X1 U16931 ( .A1(n15270), .A2(n15191), .A3(n15190), .ZN(n15192) );
  NAND3_X1 U16932 ( .A1(n15194), .A2(n15193), .A3(n15192), .ZN(P2_U3219) );
  NAND2_X1 U16933 ( .A1(n15266), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n15195) );
  OAI211_X1 U16934 ( .C1(n15265), .C2(n15197), .A(n15196), .B(n15195), .ZN(
        n15198) );
  INV_X1 U16935 ( .A(n15198), .ZN(n15209) );
  AOI211_X1 U16936 ( .C1(n15201), .C2(n15200), .A(n15199), .B(n15214), .ZN(
        n15202) );
  INV_X1 U16937 ( .A(n15202), .ZN(n15208) );
  AOI211_X1 U16938 ( .C1(n15205), .C2(n15204), .A(n15221), .B(n15203), .ZN(
        n15206) );
  INV_X1 U16939 ( .A(n15206), .ZN(n15207) );
  NAND3_X1 U16940 ( .A1(n15209), .A2(n15208), .A3(n15207), .ZN(P2_U3221) );
  INV_X1 U16941 ( .A(n15210), .ZN(n15213) );
  NAND2_X1 U16942 ( .A1(n15226), .A2(n15211), .ZN(n15212) );
  OAI211_X1 U16943 ( .C1(n15226), .C2(n15211), .A(n15213), .B(n15212), .ZN(
        n15215) );
  AOI21_X1 U16944 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15225) );
  INV_X1 U16945 ( .A(n15217), .ZN(n15223) );
  NAND3_X1 U16946 ( .A1(n15220), .A2(n15219), .A3(n15218), .ZN(n15222) );
  AOI21_X1 U16947 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15224) );
  AOI211_X1 U16948 ( .C1(n15268), .C2(n15226), .A(n15225), .B(n15224), .ZN(
        n15228) );
  OAI211_X1 U16949 ( .C1(n15229), .C2(n15231), .A(n15228), .B(n15227), .ZN(
        P2_U3226) );
  OAI22_X1 U16950 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15232), .B1(n15231), .B2(
        n15230), .ZN(n15233) );
  AOI21_X1 U16951 ( .B1(n15234), .B2(n15268), .A(n15233), .ZN(n15243) );
  OAI211_X1 U16952 ( .C1(n15237), .C2(n15236), .A(n15270), .B(n15235), .ZN(
        n15242) );
  OAI211_X1 U16953 ( .C1(n15240), .C2(n15239), .A(n15274), .B(n15238), .ZN(
        n15241) );
  NAND3_X1 U16954 ( .A1(n15243), .A2(n15242), .A3(n15241), .ZN(P2_U3227) );
  AOI22_X1 U16955 ( .A1(n15266), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15252) );
  NAND2_X1 U16956 ( .A1(n15268), .A2(n15244), .ZN(n15251) );
  OAI211_X1 U16957 ( .C1(n15246), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15274), 
        .B(n15245), .ZN(n15250) );
  OAI211_X1 U16958 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15248), .A(n15270), 
        .B(n15247), .ZN(n15249) );
  NAND4_X1 U16959 ( .A1(n15252), .A2(n15251), .A3(n15250), .A4(n15249), .ZN(
        P2_U3229) );
  OAI211_X1 U16960 ( .C1(n15255), .C2(n15254), .A(n15270), .B(n15253), .ZN(
        n15256) );
  NAND2_X1 U16961 ( .A1(n15257), .A2(n15256), .ZN(n15258) );
  AOI21_X1 U16962 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n15266), .A(n15258), 
        .ZN(n15263) );
  OAI211_X1 U16963 ( .C1(n15261), .C2(n15260), .A(n15274), .B(n15259), .ZN(
        n15262) );
  OAI211_X1 U16964 ( .C1(n15265), .C2(n15264), .A(n15263), .B(n15262), .ZN(
        P2_U3230) );
  AOI22_X1 U16965 ( .A1(n15266), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15280) );
  NAND2_X1 U16966 ( .A1(n15268), .A2(n15267), .ZN(n15279) );
  OAI211_X1 U16967 ( .C1(n15272), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        n15278) );
  OAI211_X1 U16968 ( .C1(n15276), .C2(n15275), .A(n15274), .B(n15273), .ZN(
        n15277) );
  NAND4_X1 U16969 ( .A1(n15280), .A2(n15279), .A3(n15278), .A4(n15277), .ZN(
        P2_U3231) );
  AOI222_X1 U16970 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n15305), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n15283), .C1(n15282), .C2(n15281), .ZN(
        n15289) );
  AOI22_X1 U16971 ( .A1(n15287), .A2(n15286), .B1(n15285), .B2(n15284), .ZN(
        n15288) );
  OAI211_X1 U16972 ( .C1(n15305), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        P2_U3263) );
  NOR2_X1 U16973 ( .A1(n15292), .A2(n15291), .ZN(n15346) );
  NOR2_X1 U16974 ( .A1(n15376), .A2(n15293), .ZN(n15296) );
  OAI22_X1 U16975 ( .A1(n15296), .A2(n15344), .B1(n15295), .B2(n15294), .ZN(
        n15345) );
  AOI21_X1 U16976 ( .B1(n15346), .B2(n15297), .A(n15345), .ZN(n15304) );
  INV_X1 U16977 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15299) );
  OAI22_X1 U16978 ( .A1(n15300), .A2(n15344), .B1(n15299), .B2(n15298), .ZN(
        n15301) );
  INV_X1 U16979 ( .A(n15301), .ZN(n15302) );
  OAI221_X1 U16980 ( .B1(n15305), .B2(n15304), .C1(n15303), .C2(n9746), .A(
        n15302), .ZN(P2_U3265) );
  INV_X1 U16981 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15307) );
  NOR2_X1 U16982 ( .A1(n15338), .A2(n15307), .ZN(P2_U3266) );
  INV_X1 U16983 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15308) );
  NOR2_X1 U16984 ( .A1(n15338), .A2(n15308), .ZN(P2_U3267) );
  INV_X1 U16985 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15309) );
  NOR2_X1 U16986 ( .A1(n15338), .A2(n15309), .ZN(P2_U3268) );
  INV_X1 U16987 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15310) );
  NOR2_X1 U16988 ( .A1(n15338), .A2(n15310), .ZN(P2_U3269) );
  INV_X1 U16989 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15311) );
  NOR2_X1 U16990 ( .A1(n15321), .A2(n15311), .ZN(P2_U3270) );
  INV_X1 U16991 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15312) );
  NOR2_X1 U16992 ( .A1(n15321), .A2(n15312), .ZN(P2_U3271) );
  INV_X1 U16993 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15313) );
  NOR2_X1 U16994 ( .A1(n15321), .A2(n15313), .ZN(P2_U3272) );
  INV_X1 U16995 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15314) );
  NOR2_X1 U16996 ( .A1(n15321), .A2(n15314), .ZN(P2_U3273) );
  INV_X1 U16997 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15315) );
  NOR2_X1 U16998 ( .A1(n15321), .A2(n15315), .ZN(P2_U3274) );
  INV_X1 U16999 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15316) );
  NOR2_X1 U17000 ( .A1(n15321), .A2(n15316), .ZN(P2_U3275) );
  INV_X1 U17001 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15317) );
  NOR2_X1 U17002 ( .A1(n15321), .A2(n15317), .ZN(P2_U3276) );
  INV_X1 U17003 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15318) );
  NOR2_X1 U17004 ( .A1(n15321), .A2(n15318), .ZN(P2_U3277) );
  INV_X1 U17005 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15319) );
  NOR2_X1 U17006 ( .A1(n15321), .A2(n15319), .ZN(P2_U3278) );
  INV_X1 U17007 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15320) );
  NOR2_X1 U17008 ( .A1(n15321), .A2(n15320), .ZN(P2_U3279) );
  INV_X1 U17009 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15322) );
  NOR2_X1 U17010 ( .A1(n15338), .A2(n15322), .ZN(P2_U3280) );
  INV_X1 U17011 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15323) );
  NOR2_X1 U17012 ( .A1(n15338), .A2(n15323), .ZN(P2_U3281) );
  INV_X1 U17013 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15324) );
  NOR2_X1 U17014 ( .A1(n15338), .A2(n15324), .ZN(P2_U3282) );
  INV_X1 U17015 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15325) );
  NOR2_X1 U17016 ( .A1(n15338), .A2(n15325), .ZN(P2_U3283) );
  INV_X1 U17017 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15326) );
  NOR2_X1 U17018 ( .A1(n15338), .A2(n15326), .ZN(P2_U3284) );
  INV_X1 U17019 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15327) );
  NOR2_X1 U17020 ( .A1(n15338), .A2(n15327), .ZN(P2_U3285) );
  INV_X1 U17021 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15328) );
  NOR2_X1 U17022 ( .A1(n15338), .A2(n15328), .ZN(P2_U3286) );
  INV_X1 U17023 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U17024 ( .A1(n15338), .A2(n15329), .ZN(P2_U3287) );
  INV_X1 U17025 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15330) );
  NOR2_X1 U17026 ( .A1(n15338), .A2(n15330), .ZN(P2_U3288) );
  INV_X1 U17027 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15331) );
  NOR2_X1 U17028 ( .A1(n15338), .A2(n15331), .ZN(P2_U3289) );
  INV_X1 U17029 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U17030 ( .A1(n15338), .A2(n15332), .ZN(P2_U3290) );
  INV_X1 U17031 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U17032 ( .A1(n15338), .A2(n15333), .ZN(P2_U3291) );
  INV_X1 U17033 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15334) );
  NOR2_X1 U17034 ( .A1(n15338), .A2(n15334), .ZN(P2_U3292) );
  INV_X1 U17035 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U17036 ( .A1(n15338), .A2(n15335), .ZN(P2_U3293) );
  INV_X1 U17037 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U17038 ( .A1(n15338), .A2(n15336), .ZN(P2_U3294) );
  INV_X1 U17039 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U17040 ( .A1(n15338), .A2(n15337), .ZN(P2_U3295) );
  MUX2_X1 U17041 ( .A(P2_D_REG_0__SCAN_IN), .B(n15339), .S(n15338), .Z(
        P2_U3416) );
  AOI22_X1 U17042 ( .A1(n15343), .A2(n15342), .B1(n15341), .B2(n15340), .ZN(
        P2_U3417) );
  INV_X1 U17043 ( .A(n15344), .ZN(n15347) );
  AOI211_X1 U17044 ( .C1(n15347), .C2(n15399), .A(n15346), .B(n15345), .ZN(
        n15411) );
  INV_X1 U17045 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15348) );
  AOI22_X1 U17046 ( .A1(n15409), .A2(n15411), .B1(n15348), .B2(n15407), .ZN(
        P2_U3430) );
  INV_X1 U17047 ( .A(n15354), .ZN(n15352) );
  AOI211_X1 U17048 ( .C1(n15392), .C2(n12363), .A(n15350), .B(n15349), .ZN(
        n15351) );
  OAI21_X1 U17049 ( .B1(n15359), .B2(n15352), .A(n15351), .ZN(n15353) );
  AOI21_X1 U17050 ( .B1(n15376), .B2(n15354), .A(n15353), .ZN(n15413) );
  INV_X1 U17051 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U17052 ( .A1(n15409), .A2(n15413), .B1(n15355), .B2(n15407), .ZN(
        P2_U3433) );
  INV_X1 U17053 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U17054 ( .A1(n15409), .A2(n15357), .B1(n15356), .B2(n15407), .ZN(
        P2_U3436) );
  INV_X1 U17055 ( .A(n15360), .ZN(n15361) );
  OAI211_X1 U17056 ( .C1(n15363), .C2(n15403), .A(n15362), .B(n15361), .ZN(
        n15364) );
  NOR2_X1 U17057 ( .A1(n15365), .A2(n15364), .ZN(n15415) );
  INV_X1 U17058 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U17059 ( .A1(n15409), .A2(n15415), .B1(n15366), .B2(n15407), .ZN(
        P2_U3439) );
  OAI21_X1 U17060 ( .B1(n15368), .B2(n15403), .A(n15367), .ZN(n15371) );
  INV_X1 U17061 ( .A(n15369), .ZN(n15370) );
  AOI211_X1 U17062 ( .C1(n15399), .C2(n15372), .A(n15371), .B(n15370), .ZN(
        n15417) );
  INV_X1 U17063 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U17064 ( .A1(n15409), .A2(n15417), .B1(n15373), .B2(n15407), .ZN(
        P2_U3442) );
  INV_X1 U17065 ( .A(n15374), .ZN(n15375) );
  OAI21_X1 U17066 ( .B1(n15399), .B2(n15376), .A(n15375), .ZN(n15382) );
  AND2_X1 U17067 ( .A1(n15377), .A2(n15392), .ZN(n15378) );
  NOR2_X1 U17068 ( .A1(n15379), .A2(n15378), .ZN(n15380) );
  AND3_X1 U17069 ( .A1(n15382), .A2(n15381), .A3(n15380), .ZN(n15419) );
  INV_X1 U17070 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U17071 ( .A1(n15409), .A2(n15419), .B1(n15383), .B2(n15407), .ZN(
        P2_U3445) );
  OAI21_X1 U17072 ( .B1(n15385), .B2(n15403), .A(n15384), .ZN(n15387) );
  AOI211_X1 U17073 ( .C1(n15399), .C2(n15388), .A(n15387), .B(n15386), .ZN(
        n15421) );
  INV_X1 U17074 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U17075 ( .A1(n15409), .A2(n15421), .B1(n15389), .B2(n15407), .ZN(
        P2_U3454) );
  AND2_X1 U17076 ( .A1(n15391), .A2(n15390), .ZN(n15396) );
  AND2_X1 U17077 ( .A1(n15393), .A2(n15392), .ZN(n15394) );
  NOR4_X1 U17078 ( .A1(n15397), .A2(n15396), .A3(n15395), .A4(n15394), .ZN(
        n15423) );
  INV_X1 U17079 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15398) );
  AOI22_X1 U17080 ( .A1(n15409), .A2(n15423), .B1(n15398), .B2(n15407), .ZN(
        P2_U3460) );
  NAND2_X1 U17081 ( .A1(n15400), .A2(n15399), .ZN(n15402) );
  OAI211_X1 U17082 ( .C1(n15404), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        n15405) );
  NOR2_X1 U17083 ( .A1(n15406), .A2(n15405), .ZN(n15426) );
  INV_X1 U17084 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U17085 ( .A1(n15409), .A2(n15426), .B1(n15408), .B2(n15407), .ZN(
        P2_U3463) );
  AOI22_X1 U17086 ( .A1(n15427), .A2(n15411), .B1(n15410), .B2(n15424), .ZN(
        P2_U3499) );
  AOI22_X1 U17087 ( .A1(n15427), .A2(n15413), .B1(n15412), .B2(n15424), .ZN(
        P2_U3500) );
  AOI22_X1 U17088 ( .A1(n15427), .A2(n15415), .B1(n15414), .B2(n15424), .ZN(
        P2_U3502) );
  AOI22_X1 U17089 ( .A1(n15427), .A2(n15417), .B1(n15416), .B2(n15424), .ZN(
        P2_U3503) );
  AOI22_X1 U17090 ( .A1(n15427), .A2(n15419), .B1(n15418), .B2(n15424), .ZN(
        P2_U3504) );
  AOI22_X1 U17091 ( .A1(n15427), .A2(n15421), .B1(n15420), .B2(n15424), .ZN(
        P2_U3507) );
  AOI22_X1 U17092 ( .A1(n15427), .A2(n15423), .B1(n15422), .B2(n15424), .ZN(
        P2_U3509) );
  AOI22_X1 U17093 ( .A1(n15427), .A2(n15426), .B1(n15425), .B2(n15424), .ZN(
        P2_U3510) );
  NOR2_X1 U17094 ( .A1(P3_U3897), .A2(n15581), .ZN(P3_U3150) );
  INV_X1 U17095 ( .A(n15428), .ZN(n15670) );
  AOI222_X1 U17096 ( .A1(n15670), .A2(n15432), .B1(n15431), .B2(n15430), .C1(
        n15678), .C2(n15429), .ZN(n15433) );
  OAI21_X1 U17097 ( .B1(n15434), .B2(n15675), .A(n15433), .ZN(P3_U3172) );
  XNOR2_X1 U17098 ( .A(n15436), .B(n15435), .ZN(n15447) );
  NOR2_X1 U17099 ( .A1(n15584), .A2(n15437), .ZN(n15446) );
  AOI21_X1 U17100 ( .B1(n15440), .B2(n15439), .A(n15438), .ZN(n15444) );
  XOR2_X1 U17101 ( .A(n15442), .B(n15441), .Z(n15443) );
  OAI22_X1 U17102 ( .A1(n15594), .A2(n15444), .B1(n15443), .B2(n15488), .ZN(
        n15445) );
  AOI211_X1 U17103 ( .C1(n15447), .C2(n15588), .A(n15446), .B(n15445), .ZN(
        n15449) );
  OAI211_X1 U17104 ( .C1(n15450), .C2(n15519), .A(n15449), .B(n15448), .ZN(
        P3_U3186) );
  XNOR2_X1 U17105 ( .A(n15452), .B(n15451), .ZN(n15463) );
  AOI21_X1 U17106 ( .B1(n15455), .B2(n15454), .A(n15453), .ZN(n15456) );
  NOR2_X1 U17107 ( .A1(n15456), .A2(n15594), .ZN(n15462) );
  XOR2_X1 U17108 ( .A(n15458), .B(n15457), .Z(n15460) );
  OAI22_X1 U17109 ( .A1(n15460), .A2(n15488), .B1(n15584), .B2(n15459), .ZN(
        n15461) );
  AOI211_X1 U17110 ( .C1(n15463), .C2(n15588), .A(n15462), .B(n15461), .ZN(
        n15465) );
  OAI211_X1 U17111 ( .C1(n15466), .C2(n15519), .A(n15465), .B(n15464), .ZN(
        P3_U3188) );
  XNOR2_X1 U17112 ( .A(n15468), .B(n15467), .ZN(n15478) );
  XOR2_X1 U17113 ( .A(n15469), .B(P3_REG1_REG_7__SCAN_IN), .Z(n15471) );
  OAI22_X1 U17114 ( .A1(n15471), .A2(n15488), .B1(n15470), .B2(n15584), .ZN(
        n15477) );
  AOI21_X1 U17115 ( .B1(n15474), .B2(n15473), .A(n15472), .ZN(n15475) );
  NOR2_X1 U17116 ( .A1(n15475), .A2(n15594), .ZN(n15476) );
  AOI211_X1 U17117 ( .C1(n15588), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15480) );
  OAI211_X1 U17118 ( .C1(n15481), .C2(n15519), .A(n15480), .B(n15479), .ZN(
        P3_U3189) );
  OAI21_X1 U17119 ( .B1(n15484), .B2(n15483), .A(n15482), .ZN(n15496) );
  XOR2_X1 U17120 ( .A(n15486), .B(n15485), .Z(n15489) );
  OAI22_X1 U17121 ( .A1(n15489), .A2(n15488), .B1(n15487), .B2(n15584), .ZN(
        n15495) );
  AOI21_X1 U17122 ( .B1(n15492), .B2(n15491), .A(n15490), .ZN(n15493) );
  NOR2_X1 U17123 ( .A1(n15493), .A2(n15594), .ZN(n15494) );
  AOI211_X1 U17124 ( .C1(n15588), .C2(n15496), .A(n15495), .B(n15494), .ZN(
        n15498) );
  OAI211_X1 U17125 ( .C1(n15499), .C2(n15519), .A(n15498), .B(n15497), .ZN(
        P3_U3190) );
  NAND2_X1 U17126 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  XNOR2_X1 U17127 ( .A(n15503), .B(n15502), .ZN(n15515) );
  AOI21_X1 U17128 ( .B1(n15506), .B2(n15505), .A(n6874), .ZN(n15507) );
  OR2_X1 U17129 ( .A1(n15507), .A2(n15594), .ZN(n15514) );
  OAI21_X1 U17130 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15509), .A(n15508), .ZN(
        n15512) );
  NOR2_X1 U17131 ( .A1(n15584), .A2(n15510), .ZN(n15511) );
  AOI21_X1 U17132 ( .B1(n15512), .B2(n15586), .A(n15511), .ZN(n15513) );
  OAI211_X1 U17133 ( .C1(n15515), .C2(n15549), .A(n15514), .B(n15513), .ZN(
        n15516) );
  INV_X1 U17134 ( .A(n15516), .ZN(n15518) );
  OAI211_X1 U17135 ( .C1(n15520), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        P3_U3191) );
  AOI21_X1 U17136 ( .B1(n15523), .B2(n15522), .A(n15521), .ZN(n15537) );
  OAI21_X1 U17137 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15525), .A(n15524), 
        .ZN(n15530) );
  AOI21_X1 U17138 ( .B1(n15581), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15526), 
        .ZN(n15527) );
  OAI21_X1 U17139 ( .B1(n15584), .B2(n15528), .A(n15527), .ZN(n15529) );
  AOI21_X1 U17140 ( .B1(n15530), .B2(n15586), .A(n15529), .ZN(n15536) );
  OAI21_X1 U17141 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15534) );
  NAND2_X1 U17142 ( .A1(n15534), .A2(n15588), .ZN(n15535) );
  OAI211_X1 U17143 ( .C1(n15537), .C2(n15594), .A(n15536), .B(n15535), .ZN(
        P3_U3193) );
  AOI21_X1 U17144 ( .B1(n15540), .B2(n15539), .A(n15538), .ZN(n15556) );
  OAI21_X1 U17145 ( .B1(n15543), .B2(n15542), .A(n15541), .ZN(n15548) );
  AOI21_X1 U17146 ( .B1(n15581), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15544), 
        .ZN(n15545) );
  OAI21_X1 U17147 ( .B1(n15584), .B2(n15546), .A(n15545), .ZN(n15547) );
  AOI21_X1 U17148 ( .B1(n15548), .B2(n15586), .A(n15547), .ZN(n15555) );
  AOI21_X1 U17149 ( .B1(n15551), .B2(n15550), .A(n15549), .ZN(n15553) );
  NAND2_X1 U17150 ( .A1(n15553), .A2(n15552), .ZN(n15554) );
  OAI211_X1 U17151 ( .C1(n15556), .C2(n15594), .A(n15555), .B(n15554), .ZN(
        P3_U3194) );
  AOI21_X1 U17152 ( .B1(n15559), .B2(n15558), .A(n15557), .ZN(n15573) );
  OAI21_X1 U17153 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15561), .A(n15560), 
        .ZN(n15566) );
  AOI21_X1 U17154 ( .B1(n15581), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15562), 
        .ZN(n15563) );
  OAI21_X1 U17155 ( .B1(n15584), .B2(n15564), .A(n15563), .ZN(n15565) );
  AOI21_X1 U17156 ( .B1(n15566), .B2(n15586), .A(n15565), .ZN(n15572) );
  OAI21_X1 U17157 ( .B1(n15569), .B2(n15568), .A(n15567), .ZN(n15570) );
  NAND2_X1 U17158 ( .A1(n15570), .A2(n15588), .ZN(n15571) );
  OAI211_X1 U17159 ( .C1(n15573), .C2(n15594), .A(n15572), .B(n15571), .ZN(
        P3_U3195) );
  AOI21_X1 U17160 ( .B1(n15576), .B2(n15575), .A(n15574), .ZN(n15595) );
  OAI21_X1 U17161 ( .B1(n15579), .B2(n15578), .A(n15577), .ZN(n15587) );
  AOI21_X1 U17162 ( .B1(n15581), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n15580), 
        .ZN(n15582) );
  OAI21_X1 U17163 ( .B1(n15584), .B2(n15583), .A(n15582), .ZN(n15585) );
  AOI21_X1 U17164 ( .B1(n15587), .B2(n15586), .A(n15585), .ZN(n15593) );
  OAI211_X1 U17165 ( .C1(n15591), .C2(n15590), .A(n15589), .B(n15588), .ZN(
        n15592) );
  OAI211_X1 U17166 ( .C1(n15595), .C2(n15594), .A(n15593), .B(n15592), .ZN(
        P3_U3196) );
  XNOR2_X1 U17167 ( .A(n15596), .B(n15601), .ZN(n15599) );
  AOI222_X1 U17168 ( .A1(n15671), .A2(n15599), .B1(n15598), .B2(n15654), .C1(
        n15597), .C2(n15653), .ZN(n15724) );
  AOI22_X1 U17169 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15649), .B1(n6668), .B2(
        n15600), .ZN(n15605) );
  XNOR2_X1 U17170 ( .A(n15602), .B(n15601), .ZN(n15727) );
  NOR2_X1 U17171 ( .A1(n15603), .A2(n15718), .ZN(n15726) );
  AOI22_X1 U17172 ( .A1(n15727), .A2(n15631), .B1(n15726), .B2(n15679), .ZN(
        n15604) );
  OAI211_X1 U17173 ( .C1(n15649), .C2(n15724), .A(n15605), .B(n15604), .ZN(
        P3_U3225) );
  XOR2_X1 U17174 ( .A(n15607), .B(n15606), .Z(n15615) );
  INV_X1 U17175 ( .A(n15615), .ZN(n15710) );
  INV_X1 U17176 ( .A(n15607), .ZN(n15609) );
  OAI21_X1 U17177 ( .B1(n15610), .B2(n15609), .A(n15608), .ZN(n15613) );
  OAI22_X1 U17178 ( .A1(n15623), .A2(n15637), .B1(n15611), .B2(n15673), .ZN(
        n15612) );
  AOI21_X1 U17179 ( .B1(n15613), .B2(n15671), .A(n15612), .ZN(n15614) );
  OAI21_X1 U17180 ( .B1(n15615), .B2(n15662), .A(n15614), .ZN(n15708) );
  AOI21_X1 U17181 ( .B1(n15616), .B2(n15710), .A(n15708), .ZN(n15621) );
  AND2_X1 U17182 ( .A1(n15617), .A2(n15677), .ZN(n15709) );
  AOI22_X1 U17183 ( .A1(n15679), .A2(n15709), .B1(n6668), .B2(n15618), .ZN(
        n15619) );
  OAI221_X1 U17184 ( .B1(n15649), .B2(n15621), .C1(n15682), .C2(n15620), .A(
        n15619), .ZN(P3_U3228) );
  AOI21_X1 U17185 ( .B1(n15622), .B2(n15628), .A(n15641), .ZN(n15627) );
  OAI22_X1 U17186 ( .A1(n15624), .A2(n15637), .B1(n15623), .B2(n15673), .ZN(
        n15625) );
  AOI21_X1 U17187 ( .B1(n15627), .B2(n15626), .A(n15625), .ZN(n15698) );
  AOI22_X1 U17188 ( .A1(n15649), .A2(P3_REG2_REG_3__SCAN_IN), .B1(n6668), .B2(
        n8475), .ZN(n15633) );
  XNOR2_X1 U17189 ( .A(n15629), .B(n15628), .ZN(n15701) );
  NOR2_X1 U17190 ( .A1(n15630), .A2(n15718), .ZN(n15700) );
  AOI22_X1 U17191 ( .A1(n15701), .A2(n15631), .B1(n15700), .B2(n15679), .ZN(
        n15632) );
  OAI211_X1 U17192 ( .C1(n15649), .C2(n15698), .A(n15633), .B(n15632), .ZN(
        P3_U3230) );
  OAI21_X1 U17193 ( .B1(n15635), .B2(n15640), .A(n15634), .ZN(n15696) );
  OAI22_X1 U17194 ( .A1(n15674), .A2(n15637), .B1(n15636), .B2(n15673), .ZN(
        n15644) );
  NAND3_X1 U17195 ( .A1(n15656), .A2(n15640), .A3(n15639), .ZN(n15642) );
  AOI21_X1 U17196 ( .B1(n15638), .B2(n15642), .A(n15641), .ZN(n15643) );
  AOI211_X1 U17197 ( .C1(n15645), .C2(n15696), .A(n15644), .B(n15643), .ZN(
        n15693) );
  NOR2_X1 U17198 ( .A1(n15646), .A2(n15718), .ZN(n15695) );
  AOI22_X1 U17199 ( .A1(n15695), .A2(n15663), .B1(n6668), .B2(
        P3_REG3_REG_2__SCAN_IN), .ZN(n15648) );
  AOI22_X1 U17200 ( .A1(n15696), .A2(n15666), .B1(P3_REG2_REG_2__SCAN_IN), 
        .B2(n15649), .ZN(n15647) );
  OAI221_X1 U17201 ( .B1(n15649), .B2(n15693), .C1(n15649), .C2(n15648), .A(
        n15647), .ZN(P3_U3231) );
  NOR2_X1 U17202 ( .A1(n15650), .A2(n15718), .ZN(n15690) );
  XNOR2_X1 U17203 ( .A(n15658), .B(n15651), .ZN(n15664) );
  AOI22_X1 U17204 ( .A1(n15655), .A2(n15654), .B1(n15653), .B2(n15652), .ZN(
        n15661) );
  OAI21_X1 U17205 ( .B1(n15658), .B2(n15657), .A(n15656), .ZN(n15659) );
  NAND2_X1 U17206 ( .A1(n15659), .A2(n15671), .ZN(n15660) );
  OAI211_X1 U17207 ( .C1(n15664), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        n15689) );
  AOI21_X1 U17208 ( .B1(n15690), .B2(n15663), .A(n15689), .ZN(n15669) );
  INV_X1 U17209 ( .A(n15664), .ZN(n15691) );
  AOI22_X1 U17210 ( .A1(n15691), .A2(n15666), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n6668), .ZN(n15667) );
  OAI221_X1 U17211 ( .B1(n15649), .B2(n15669), .C1(n15682), .C2(n15668), .A(
        n15667), .ZN(P3_U3232) );
  OAI21_X1 U17212 ( .B1(n15672), .B2(n15671), .A(n15670), .ZN(n15687) );
  OR2_X1 U17213 ( .A1(n15674), .A2(n15673), .ZN(n15685) );
  OAI211_X1 U17214 ( .C1(n15676), .C2(n15675), .A(n15687), .B(n15685), .ZN(
        n15680) );
  AND2_X1 U17215 ( .A1(n15678), .A2(n15677), .ZN(n15684) );
  AOI22_X1 U17216 ( .A1(n15680), .A2(n15682), .B1(n15684), .B2(n15679), .ZN(
        n15681) );
  OAI21_X1 U17217 ( .B1(n15683), .B2(n15682), .A(n15681), .ZN(P3_U3233) );
  INV_X1 U17218 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n15688) );
  INV_X1 U17219 ( .A(n15684), .ZN(n15686) );
  AND3_X1 U17220 ( .A1(n15687), .A2(n15686), .A3(n15685), .ZN(n15744) );
  AOI22_X1 U17221 ( .A1(n15742), .A2(n15688), .B1(n15744), .B2(n15740), .ZN(
        P3_U3390) );
  INV_X1 U17222 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15692) );
  AOI211_X1 U17223 ( .C1(n15739), .C2(n15691), .A(n15690), .B(n15689), .ZN(
        n15745) );
  AOI22_X1 U17224 ( .A1(n15742), .A2(n15692), .B1(n15745), .B2(n15740), .ZN(
        P3_U3393) );
  INV_X1 U17225 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15697) );
  INV_X1 U17226 ( .A(n15693), .ZN(n15694) );
  AOI211_X1 U17227 ( .C1(n15739), .C2(n15696), .A(n15695), .B(n15694), .ZN(
        n15746) );
  AOI22_X1 U17228 ( .A1(n15742), .A2(n15697), .B1(n15746), .B2(n15740), .ZN(
        P3_U3396) );
  INV_X1 U17229 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15702) );
  INV_X1 U17230 ( .A(n15698), .ZN(n15699) );
  AOI211_X1 U17231 ( .C1(n15701), .C2(n15732), .A(n15700), .B(n15699), .ZN(
        n15748) );
  AOI22_X1 U17232 ( .A1(n15742), .A2(n15702), .B1(n15748), .B2(n15740), .ZN(
        P3_U3399) );
  INV_X1 U17233 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15707) );
  OAI22_X1 U17234 ( .A1(n15704), .A2(n15719), .B1(n15718), .B2(n15703), .ZN(
        n15705) );
  NOR2_X1 U17235 ( .A1(n15706), .A2(n15705), .ZN(n15750) );
  AOI22_X1 U17236 ( .A1(n15742), .A2(n15707), .B1(n15750), .B2(n15740), .ZN(
        P3_U3402) );
  INV_X1 U17237 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15711) );
  AOI211_X1 U17238 ( .C1(n15710), .C2(n15739), .A(n15709), .B(n15708), .ZN(
        n15752) );
  AOI22_X1 U17239 ( .A1(n15742), .A2(n15711), .B1(n15752), .B2(n15740), .ZN(
        P3_U3405) );
  INV_X1 U17240 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15716) );
  NOR2_X1 U17241 ( .A1(n15712), .A2(n15718), .ZN(n15714) );
  AOI211_X1 U17242 ( .C1(n15715), .C2(n15732), .A(n15714), .B(n15713), .ZN(
        n15754) );
  AOI22_X1 U17243 ( .A1(n15742), .A2(n15716), .B1(n15754), .B2(n15740), .ZN(
        P3_U3408) );
  INV_X1 U17244 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15723) );
  OAI22_X1 U17245 ( .A1(n15720), .A2(n15719), .B1(n15718), .B2(n15717), .ZN(
        n15721) );
  NOR2_X1 U17246 ( .A1(n15722), .A2(n15721), .ZN(n15756) );
  AOI22_X1 U17247 ( .A1(n15742), .A2(n15723), .B1(n15756), .B2(n15740), .ZN(
        P3_U3411) );
  INV_X1 U17248 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15728) );
  INV_X1 U17249 ( .A(n15724), .ZN(n15725) );
  AOI211_X1 U17250 ( .C1(n15732), .C2(n15727), .A(n15726), .B(n15725), .ZN(
        n15758) );
  AOI22_X1 U17251 ( .A1(n15742), .A2(n15728), .B1(n15758), .B2(n15740), .ZN(
        P3_U3414) );
  INV_X1 U17252 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15734) );
  INV_X1 U17253 ( .A(n15729), .ZN(n15730) );
  AOI211_X1 U17254 ( .C1(n15733), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        n15760) );
  AOI22_X1 U17255 ( .A1(n15742), .A2(n15734), .B1(n15760), .B2(n15740), .ZN(
        P3_U3417) );
  INV_X1 U17256 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15741) );
  INV_X1 U17257 ( .A(n15735), .ZN(n15738) );
  AOI211_X1 U17258 ( .C1(n15739), .C2(n15738), .A(n15737), .B(n15736), .ZN(
        n15763) );
  AOI22_X1 U17259 ( .A1(n15742), .A2(n15741), .B1(n15763), .B2(n15740), .ZN(
        P3_U3420) );
  AOI22_X1 U17260 ( .A1(n15764), .A2(n15744), .B1(n15743), .B2(n15761), .ZN(
        P3_U3459) );
  AOI22_X1 U17261 ( .A1(n15764), .A2(n15745), .B1(n10012), .B2(n15761), .ZN(
        P3_U3460) );
  AOI22_X1 U17262 ( .A1(n15764), .A2(n15746), .B1(n9873), .B2(n15761), .ZN(
        P3_U3461) );
  INV_X1 U17263 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15747) );
  AOI22_X1 U17264 ( .A1(n15764), .A2(n15748), .B1(n15747), .B2(n15761), .ZN(
        P3_U3462) );
  AOI22_X1 U17265 ( .A1(n15764), .A2(n15750), .B1(n15749), .B2(n15761), .ZN(
        P3_U3463) );
  INV_X1 U17266 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U17267 ( .A1(n15764), .A2(n15752), .B1(n15751), .B2(n15761), .ZN(
        P3_U3464) );
  AOI22_X1 U17268 ( .A1(n15764), .A2(n15754), .B1(n15753), .B2(n15761), .ZN(
        P3_U3465) );
  INV_X1 U17269 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U17270 ( .A1(n15764), .A2(n15756), .B1(n15755), .B2(n15761), .ZN(
        P3_U3466) );
  AOI22_X1 U17271 ( .A1(n15764), .A2(n15758), .B1(n15757), .B2(n15761), .ZN(
        P3_U3467) );
  AOI22_X1 U17272 ( .A1(n15764), .A2(n15760), .B1(n15759), .B2(n15761), .ZN(
        P3_U3468) );
  AOI22_X1 U17273 ( .A1(n15764), .A2(n15763), .B1(n15762), .B2(n15761), .ZN(
        P3_U3469) );
  XOR2_X1 U17274 ( .A(n15766), .B(n15765), .Z(SUB_1596_U59) );
  XNOR2_X1 U17275 ( .A(n15767), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17276 ( .B1(n15769), .B2(n15768), .A(n15777), .ZN(SUB_1596_U53) );
  XOR2_X1 U17277 ( .A(n15770), .B(n15771), .Z(SUB_1596_U56) );
  AOI21_X1 U17278 ( .B1(n15774), .B2(n15773), .A(n15772), .ZN(n15775) );
  XOR2_X1 U17279 ( .A(n15775), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  XOR2_X1 U17280 ( .A(n15777), .B(n15776), .Z(SUB_1596_U5) );
  INV_X1 U7549 ( .A(n12655), .ZN(n12585) );
  INV_X2 U7550 ( .A(n12655), .ZN(n12584) );
  CLKBUF_X1 U7440 ( .A(n12580), .Z(n6673) );
  INV_X1 U7548 ( .A(n12655), .ZN(n12560) );
  NAND2_X2 U7556 ( .A1(n13469), .A2(n13078), .ZN(n9868) );
  BUF_X1 U7660 ( .A(n7669), .Z(n12140) );
endmodule

