

module b17_C_SARLock_k_128_9 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407;

  NAND2_X1 U11154 ( .A1(n15691), .A2(n10250), .ZN(n15679) );
  AND2_X1 U11155 ( .A1(n10159), .A2(n10157), .ZN(n15619) );
  AOI21_X1 U11156 ( .B1(n10211), .B2(n10209), .A(n10208), .ZN(n10207) );
  INV_X2 U11157 ( .A(n19024), .ZN(n19036) );
  INV_X1 U11158 ( .A(n19020), .ZN(n19038) );
  AND2_X1 U11159 ( .A1(n9885), .A2(n9757), .ZN(n10212) );
  INV_X1 U11160 ( .A(n21407), .ZN(n15063) );
  NAND2_X1 U11161 ( .A1(n13121), .A2(n9828), .ZN(n15466) );
  INV_X1 U11162 ( .A(n19037), .ZN(n16209) );
  NOR3_X1 U11163 ( .A1(n17575), .A2(n11746), .A3(n14440), .ZN(n10393) );
  NOR2_X1 U11164 ( .A1(n17575), .A2(n18574), .ZN(n19037) );
  OR2_X1 U11165 ( .A1(n10628), .A2(n16001), .ZN(n20010) );
  AND2_X1 U11166 ( .A1(n10989), .A2(n9736), .ZN(n11195) );
  INV_X1 U11167 ( .A(n10631), .ZN(n9904) );
  CLKBUF_X2 U11168 ( .A(n10331), .Z(n17533) );
  AND3_X1 U11169 ( .A1(n10574), .A2(n10573), .A3(n10572), .ZN(n10605) );
  OR2_X1 U11170 ( .A1(n9741), .A2(n10577), .ZN(n10580) );
  INV_X4 U11171 ( .A(n10449), .ZN(n11455) );
  CLKBUF_X1 U11172 ( .A(n11624), .Z(n17510) );
  OR2_X1 U11173 ( .A1(n10590), .A2(n16014), .ZN(n10574) );
  INV_X1 U11174 ( .A(n14458), .ZN(n17522) );
  BUF_X1 U11175 ( .A(n10567), .Z(n13841) );
  CLKBUF_X1 U11176 ( .A(n11661), .Z(n17521) );
  INV_X1 U11177 ( .A(n11074), .ZN(n13307) );
  INV_X2 U11178 ( .A(n13826), .ZN(n13298) );
  CLKBUF_X2 U11179 ( .A(n11844), .Z(n12958) );
  CLKBUF_X1 U11180 ( .A(n12798), .Z(n12959) );
  CLKBUF_X2 U11181 ( .A(n9747), .Z(n9735) );
  CLKBUF_X1 U11182 ( .A(n11983), .Z(n14024) );
  AND2_X1 U11184 ( .A1(n10656), .A2(n10429), .ZN(n13202) );
  INV_X1 U11185 ( .A(n10669), .ZN(n13296) );
  INV_X1 U11186 ( .A(n10739), .ZN(n11121) );
  BUF_X1 U11187 ( .A(n11969), .Z(n14621) );
  INV_X2 U11188 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19175) );
  CLKBUF_X2 U11189 ( .A(n14136), .Z(n9728) );
  INV_X1 U11191 ( .A(n12138), .ZN(n13934) );
  NOR2_X2 U11192 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13268) );
  INV_X1 U11193 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10429) );
  AND2_X2 U11194 ( .A1(n10638), .A2(n13819), .ZN(n9715) );
  AND2_X1 U11195 ( .A1(n11848), .A2(n11847), .ZN(n12004) );
  AND2_X2 U11196 ( .A1(n13638), .A2(n11846), .ZN(n12951) );
  NOR2_X2 U11197 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10645) );
  CLKBUF_X1 U11198 ( .A(n18722), .Z(n9709) );
  NOR2_X1 U11199 ( .A1(n19042), .A2(n18681), .ZN(n18722) );
  CLKBUF_X1 U11200 ( .A(n12976), .Z(n9710) );
  NOR2_X1 U11201 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12976) );
  CLKBUF_X1 U11202 ( .A(n18989), .Z(n9711) );
  NOR2_X1 U11203 ( .A1(n18877), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18989) );
  OAI22_X1 U11204 ( .A1(n13944), .A2(n14022), .B1(n16832), .B2(n14021), .ZN(
        n20932) );
  NAND2_X2 U11205 ( .A1(n20477), .A2(n14918), .ZN(n14021) );
  NAND2_X2 U11206 ( .A1(n20477), .A2(n14634), .ZN(n14022) );
  OAI22_X1 U11207 ( .A1(n13143), .A2(n19905), .B1(n16078), .B2(n10621), .ZN(
        n10625) );
  NOR2_X1 U11208 ( .A1(n12064), .A2(n9919), .ZN(n12292) );
  AND4_X1 U11209 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n10272) );
  NAND2_X1 U11210 ( .A1(n10661), .A2(n10429), .ZN(n13292) );
  INV_X1 U11211 ( .A(n11036), .ZN(n13304) );
  XNOR2_X1 U11212 ( .A(n10879), .B(n10878), .ZN(n11434) );
  OR3_X1 U11213 ( .A1(n10631), .A2(n19629), .A3(n10611), .ZN(n14139) );
  NAND2_X1 U11214 ( .A1(n11978), .A2(n11977), .ZN(n12049) );
  NAND2_X2 U11215 ( .A1(n11881), .A2(n10272), .ZN(n11957) );
  AND2_X2 U11216 ( .A1(n9717), .A2(n14156), .ZN(n14155) );
  OR2_X1 U11217 ( .A1(n15419), .A2(n15418), .ZN(n10219) );
  INV_X1 U11218 ( .A(n13287), .ZN(n13201) );
  NAND2_X1 U11219 ( .A1(n9742), .A2(n10488), .ZN(n10991) );
  OR2_X1 U11220 ( .A1(n10879), .A2(n10874), .ZN(n10905) );
  XNOR2_X1 U11221 ( .A(n10833), .B(n10834), .ZN(n11426) );
  INV_X1 U11222 ( .A(n9728), .ZN(n13873) );
  OR3_X1 U11223 ( .A1(n10631), .A2(n9750), .A3(n10629), .ZN(n19773) );
  INV_X1 U11225 ( .A(n10245), .ZN(n17511) );
  NOR2_X1 U11226 ( .A1(n17863), .A2(n11744), .ZN(n11745) );
  OR2_X1 U11227 ( .A1(n14749), .A2(n14736), .ZN(n14734) );
  NAND2_X1 U11228 ( .A1(n11957), .A2(n11958), .ZN(n14637) );
  NAND2_X1 U11229 ( .A1(n11557), .A2(n11482), .ZN(n11518) );
  XNOR2_X1 U11230 ( .A(n13317), .B(n13337), .ZN(n15439) );
  NAND2_X1 U11231 ( .A1(n10143), .A2(n10144), .ZN(n15595) );
  AND2_X1 U11232 ( .A1(n15624), .A2(n10908), .ZN(n15609) );
  NOR2_X2 U11233 ( .A1(n15679), .A2(n10096), .ZN(n15624) );
  NAND2_X1 U11234 ( .A1(n10529), .A2(n10528), .ZN(n10551) );
  NOR4_X1 U11235 ( .A1(n18458), .A2(n18476), .A3(n18244), .A4(n18243), .ZN(
        n18247) );
  NAND2_X1 U11236 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19033) );
  XNOR2_X1 U11238 ( .A(n12149), .B(n12148), .ZN(n14668) );
  BUF_X1 U11239 ( .A(n12495), .Z(n9729) );
  OAI21_X1 U11240 ( .B1(n15671), .B2(n9993), .A(n9992), .ZN(n15687) );
  NAND2_X1 U11241 ( .A1(n15929), .A2(n15886), .ZN(n16583) );
  NAND2_X1 U11242 ( .A1(n10088), .A2(n10907), .ZN(n15717) );
  INV_X1 U11243 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n21192) );
  NOR2_X1 U11244 ( .A1(n11821), .A2(n18348), .ZN(n18240) );
  INV_X1 U11245 ( .A(n18035), .ZN(n18050) );
  INV_X1 U11246 ( .A(n20341), .ZN(n21398) );
  OR2_X1 U11248 ( .A1(n15623), .A2(n15622), .ZN(n15822) );
  INV_X1 U11249 ( .A(n18196), .ZN(n18187) );
  AOI211_X1 U11250 ( .C1(n18110), .C2(n16787), .A(n16786), .B(n16785), .ZN(
        n16793) );
  NOR2_X1 U11251 ( .A1(n17980), .A2(n18050), .ZN(n18194) );
  AND2_X1 U11252 ( .A1(n11434), .A2(n15761), .ZN(n9712) );
  AND2_X1 U11253 ( .A1(n13848), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10638) );
  OAI21_X2 U11254 ( .B1(n11772), .B2(n11810), .A(n18107), .ZN(n11728) );
  BUF_X2 U11255 ( .A(n10489), .Z(n10488) );
  AND2_X2 U11256 ( .A1(n12093), .A2(n12092), .ZN(n14284) );
  AOI21_X2 U11258 ( .B1(n10587), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10569), .ZN(n10604) );
  AND2_X1 U11259 ( .A1(n13638), .A2(n11846), .ZN(n9713) );
  AND2_X2 U11260 ( .A1(n10638), .A2(n13819), .ZN(n9714) );
  AND2_X1 U11261 ( .A1(n10638), .A2(n13819), .ZN(n13266) );
  INV_X1 U11262 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9716) );
  NAND4_X1 U11263 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n9717) );
  NOR2_X2 U11264 ( .A1(n16670), .A2(n16660), .ZN(n16659) );
  NOR2_X1 U11266 ( .A1(n10296), .A2(n10298), .ZN(n11645) );
  OAI21_X2 U11267 ( .B1(n13620), .B2(n13621), .A(n13112), .ZN(n13692) );
  NOR2_X2 U11268 ( .A1(n18157), .A2(n11723), .ZN(n18138) );
  XNOR2_X2 U11269 ( .A(n11418), .B(n11406), .ZN(n14321) );
  AND2_X2 U11271 ( .A1(n14756), .A2(n9831), .ZN(n14640) );
  AND3_X1 U11272 ( .A1(n11591), .A2(n9760), .A3(n10147), .ZN(n15612) );
  AND2_X1 U11273 ( .A1(n12674), .A2(n10164), .ZN(n14861) );
  NAND2_X1 U11274 ( .A1(n10903), .A2(n10902), .ZN(n16623) );
  NOR2_X1 U11275 ( .A1(n16188), .A2(n16783), .ZN(n16746) );
  AND2_X1 U11276 ( .A1(n14774), .A2(n14759), .ZN(n14761) );
  NOR2_X1 U11277 ( .A1(n15538), .A2(n15529), .ZN(n15523) );
  OR2_X1 U11278 ( .A1(n14845), .A2(n14804), .ZN(n14806) );
  NOR3_X1 U11279 ( .A1(n17649), .A2(n17617), .A3(n17574), .ZN(n17614) );
  INV_X1 U11281 ( .A(n11475), .ZN(n11477) );
  AND2_X1 U11282 ( .A1(n11557), .A2(n11478), .ZN(n11475) );
  NOR2_X2 U11283 ( .A1(n18413), .A2(n19036), .ZN(n18335) );
  OR2_X1 U11285 ( .A1(n14258), .A2(n14409), .ZN(n14423) );
  AOI21_X2 U11286 ( .B1(n19015), .B2(n19022), .A(n19014), .ZN(n19024) );
  NAND2_X1 U11287 ( .A1(n9899), .A2(n10581), .ZN(n10583) );
  NOR2_X1 U11288 ( .A1(n11803), .A2(n19025), .ZN(n19028) );
  AND2_X1 U11289 ( .A1(n14059), .A2(n14058), .ZN(n14061) );
  INV_X2 U11290 ( .A(n18109), .ZN(n18107) );
  OR2_X1 U11291 ( .A1(n13632), .A2(n14637), .ZN(n12431) );
  NAND2_X1 U11292 ( .A1(n17575), .A2(n17578), .ZN(n10390) );
  BUF_X1 U11293 ( .A(n10494), .Z(n16038) );
  INV_X2 U11294 ( .A(n12327), .ZN(n12337) );
  OAI21_X2 U11295 ( .B1(n14195), .B2(n9728), .A(n13059), .ZN(n11239) );
  INV_X1 U11296 ( .A(n10489), .ZN(n13113) );
  AND2_X1 U11297 ( .A1(n10517), .A2(n10516), .ZN(n14136) );
  INV_X2 U11298 ( .A(n14157), .ZN(n9720) );
  AND4_X1 U11299 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11954) );
  CLKBUF_X2 U11300 ( .A(n12004), .Z(n12613) );
  CLKBUF_X2 U11301 ( .A(n11902), .Z(n12811) );
  INV_X2 U11302 ( .A(n11704), .ZN(n10374) );
  INV_X4 U11303 ( .A(n17476), .ZN(n11673) );
  CLKBUF_X2 U11304 ( .A(n12009), .Z(n12960) );
  AND2_X2 U11305 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10475) );
  CLKBUF_X2 U11307 ( .A(n14480), .Z(n9732) );
  BUF_X2 U11308 ( .A(n11889), .Z(n12928) );
  CLKBUF_X2 U11309 ( .A(n14480), .Z(n9731) );
  CLKBUF_X2 U11310 ( .A(n11944), .Z(n12934) );
  CLKBUF_X2 U11311 ( .A(n11993), .Z(n12873) );
  AND2_X2 U11312 ( .A1(n13644), .A2(n11848), .ZN(n11844) );
  OR2_X1 U11313 ( .A1(n10298), .A2(n17252), .ZN(n17525) );
  NAND2_X4 U11314 ( .A1(n19192), .A2(n19198), .ZN(n17252) );
  AND2_X2 U11315 ( .A1(n13821), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10663) );
  INV_X2 U11316 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12237) );
  INV_X1 U11317 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13819) );
  AOI21_X1 U11318 ( .B1(n15001), .B2(n20477), .A(n15000), .ZN(n15002) );
  OAI21_X1 U11319 ( .B1(n14640), .B2(n14642), .A(n14641), .ZN(n14996) );
  XNOR2_X1 U11320 ( .A(n14641), .B(n12981), .ZN(n14710) );
  AND2_X1 U11321 ( .A1(n11393), .A2(n11392), .ZN(n11589) );
  OAI21_X1 U11322 ( .B1(n14732), .B2(n14733), .A(n14723), .ZN(n15018) );
  NAND2_X1 U11323 ( .A1(n14640), .A2(n14642), .ZN(n14641) );
  AOI21_X1 U11324 ( .B1(n14724), .B2(n14723), .A(n14640), .ZN(n15010) );
  NAND2_X1 U11325 ( .A1(n9892), .A2(n9889), .ZN(n15004) );
  NOR2_X1 U11326 ( .A1(n16583), .A2(n11507), .ZN(n16579) );
  OR2_X1 U11327 ( .A1(n11594), .A2(n11593), .ZN(n10263) );
  NAND2_X1 U11328 ( .A1(n15588), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10909) );
  NAND2_X1 U11329 ( .A1(n9890), .A2(n12228), .ZN(n9889) );
  NAND2_X1 U11330 ( .A1(n9796), .A2(n12228), .ZN(n12229) );
  INV_X1 U11331 ( .A(n16617), .ZN(n15929) );
  NAND2_X1 U11332 ( .A1(n15717), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15743) );
  NAND2_X1 U11333 ( .A1(n15717), .A2(n9849), .ZN(n16617) );
  NAND2_X1 U11334 ( .A1(n10206), .A2(n10211), .ZN(n15105) );
  NOR2_X1 U11335 ( .A1(n11391), .A2(n11390), .ZN(n11392) );
  XNOR2_X1 U11336 ( .A(n10901), .B(n10899), .ZN(n15752) );
  XNOR2_X1 U11337 ( .A(n15325), .B(n13058), .ZN(n15773) );
  XNOR2_X1 U11338 ( .A(n10139), .B(n10138), .ZN(n16489) );
  NAND2_X1 U11339 ( .A1(n17836), .A2(n17837), .ZN(n17835) );
  NAND2_X1 U11340 ( .A1(n17855), .A2(n11834), .ZN(n17836) );
  AND2_X1 U11341 ( .A1(n9887), .A2(n9886), .ZN(n10211) );
  AND2_X1 U11342 ( .A1(n10201), .A2(n9799), .ZN(n10199) );
  AND2_X1 U11343 ( .A1(n15451), .A2(n13337), .ZN(n13318) );
  OR2_X1 U11344 ( .A1(n12176), .A2(n12168), .ZN(n10252) );
  AND2_X1 U11345 ( .A1(n10154), .A2(n15650), .ZN(n10153) );
  OAI21_X1 U11346 ( .B1(n10060), .B2(n10058), .A(n10057), .ZN(n16493) );
  NAND2_X1 U11347 ( .A1(n14427), .A2(n14429), .ZN(n14428) );
  OAI21_X1 U11348 ( .B1(n11419), .B2(n9877), .A(n11425), .ZN(n9875) );
  OR2_X1 U11349 ( .A1(n12193), .A2(n15301), .ZN(n12194) );
  NAND2_X1 U11350 ( .A1(n10832), .A2(n15987), .ZN(n15760) );
  NAND2_X1 U11351 ( .A1(n11426), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15761) );
  AND2_X1 U11352 ( .A1(n12521), .A2(n12520), .ZN(n14007) );
  INV_X1 U11353 ( .A(n20166), .ZN(n20173) );
  NOR2_X1 U11354 ( .A1(n14245), .A2(n14244), .ZN(n14251) );
  NOR2_X1 U11355 ( .A1(n19866), .A2(n20257), .ZN(n19922) );
  XNOR2_X1 U11356 ( .A(n12178), .B(n12177), .ZN(n12530) );
  NAND2_X1 U11357 ( .A1(n14120), .A2(n9793), .ZN(n14244) );
  NAND2_X1 U11358 ( .A1(n12170), .A2(n12161), .ZN(n20515) );
  AND2_X1 U11359 ( .A1(n10831), .A2(n10830), .ZN(n10834) );
  AND2_X1 U11360 ( .A1(n13992), .A2(n13983), .ZN(n14120) );
  CLKBUF_X1 U11361 ( .A(n12481), .Z(n20652) );
  NOR2_X1 U11362 ( .A1(n13981), .A2(n13982), .ZN(n13983) );
  OAI211_X1 U11363 ( .C1(n11798), .C2(n11797), .A(n18114), .B(n11796), .ZN(
        n18100) );
  AOI22_X1 U11364 ( .A1(n19740), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n19776), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U11365 ( .A1(n13907), .A2(n13895), .ZN(n13981) );
  AND2_X1 U11366 ( .A1(n11500), .A2(n11505), .ZN(n19322) );
  AND2_X1 U11367 ( .A1(n13905), .A2(n13904), .ZN(n13907) );
  AND2_X1 U11368 ( .A1(n13095), .A2(n13775), .ZN(n13691) );
  NOR2_X1 U11369 ( .A1(n16710), .A2(n15954), .ZN(n16683) );
  OAI22_X1 U11370 ( .A1(n14139), .A2(n10676), .B1(n10797), .B2(n10677), .ZN(
        n10612) );
  OR2_X1 U11371 ( .A1(n10628), .A2(n15396), .ZN(n20076) );
  NAND2_X1 U11372 ( .A1(n9904), .A2(n10607), .ZN(n10845) );
  NAND2_X1 U11373 ( .A1(n9904), .A2(n10608), .ZN(n10801) );
  CLKBUF_X2 U11374 ( .A(n13630), .Z(n9749) );
  OR2_X1 U11375 ( .A1(n13115), .A2(n13094), .ZN(n13095) );
  CLKBUF_X1 U11376 ( .A(n13678), .Z(n9748) );
  NAND2_X1 U11377 ( .A1(n9986), .A2(n9904), .ZN(n16055) );
  AND2_X1 U11378 ( .A1(n13887), .A2(n13781), .ZN(n13905) );
  NAND2_X2 U11379 ( .A1(n14985), .A2(n13963), .ZN(n14990) );
  NOR2_X2 U11380 ( .A1(n19215), .A2(n16915), .ZN(n18143) );
  NOR2_X2 U11381 ( .A1(n18552), .A2(n16915), .ZN(n18191) );
  AND2_X1 U11382 ( .A1(n18106), .A2(n9801), .ZN(n18016) );
  NOR2_X1 U11383 ( .A1(n13779), .A2(n13780), .ZN(n13781) );
  OR2_X1 U11384 ( .A1(n12044), .A2(n12043), .ZN(n10179) );
  OR2_X2 U11385 ( .A1(n20474), .A2(n13617), .ZN(n20482) );
  NAND2_X1 U11386 ( .A1(n9917), .A2(n12051), .ZN(n12490) );
  NOR2_X1 U11387 ( .A1(n16001), .A2(n10630), .ZN(n9986) );
  NAND2_X1 U11388 ( .A1(n13961), .A2(n13960), .ZN(n14985) );
  NAND2_X1 U11389 ( .A1(n12056), .A2(n12055), .ZN(n9884) );
  CLKBUF_X3 U11390 ( .A(n14555), .Z(n19410) );
  AND3_X1 U11391 ( .A1(n10053), .A2(n15714), .A3(n10052), .ZN(n19269) );
  INV_X2 U11392 ( .A(n13768), .ZN(n20470) );
  OR2_X2 U11393 ( .A1(n11461), .A2(n11455), .ZN(n11557) );
  NAND2_X1 U11394 ( .A1(n13098), .A2(n13097), .ZN(n16010) );
  AND2_X1 U11395 ( .A1(n10610), .A2(n13096), .ZN(n10622) );
  AND2_X1 U11396 ( .A1(n10982), .A2(n13899), .ZN(n11587) );
  CLKBUF_X1 U11397 ( .A(n16568), .Z(n16632) );
  XNOR2_X1 U11398 ( .A(n10603), .B(n10609), .ZN(n13099) );
  NAND2_X1 U11399 ( .A1(n10068), .A2(n9788), .ZN(n11729) );
  NOR2_X2 U11400 ( .A1(n19532), .A2(n19874), .ZN(n14194) );
  NOR2_X2 U11401 ( .A1(n14144), .A2(n19874), .ZN(n14145) );
  XNOR2_X1 U11402 ( .A(n11289), .B(n11290), .ZN(n11287) );
  AND2_X1 U11403 ( .A1(n11286), .A2(n11285), .ZN(n13779) );
  INV_X2 U11404 ( .A(n17569), .ZN(n17556) );
  XNOR2_X1 U11405 ( .A(n10606), .B(n10605), .ZN(n10609) );
  OAI21_X1 U11406 ( .B1(n10601), .B2(n10604), .A(n10605), .ZN(n10576) );
  OR2_X1 U11407 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  AND3_X1 U11408 ( .A1(n10594), .A2(n10593), .A3(n10592), .ZN(n11290) );
  NAND2_X1 U11409 ( .A1(n10589), .A2(n10588), .ZN(n11289) );
  NOR2_X1 U11410 ( .A1(n11001), .A2(n11000), .ZN(n11010) );
  NAND2_X1 U11411 ( .A1(n12046), .A2(n11976), .ZN(n12057) );
  OAI21_X1 U11412 ( .B1(n14609), .B2(n11771), .A(n19213), .ZN(n18530) );
  OAI22_X1 U11413 ( .A1(n10566), .A2(n10541), .B1(n9752), .B2(n10540), .ZN(
        n10550) );
  OR2_X1 U11414 ( .A1(n11805), .A2(n9867), .ZN(n19025) );
  AND3_X1 U11415 ( .A1(n11992), .A2(n11991), .A3(n11990), .ZN(n12047) );
  NAND2_X1 U11416 ( .A1(n9780), .A2(n10559), .ZN(n10566) );
  NOR2_X1 U11417 ( .A1(n13510), .A2(n13883), .ZN(n19379) );
  AND3_X1 U11418 ( .A1(n10538), .A2(n10537), .A3(n11244), .ZN(n10559) );
  INV_X2 U11419 ( .A(n10571), .ZN(n11367) );
  AOI21_X1 U11420 ( .B1(n11717), .B2(n18178), .A(n11716), .ZN(n11719) );
  AND2_X2 U11421 ( .A1(n11253), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U11422 ( .A1(n12309), .A2(n14621), .ZN(n11988) );
  NOR2_X1 U11423 ( .A1(n18186), .A2(n11714), .ZN(n18180) );
  NAND2_X1 U11424 ( .A1(n10532), .A2(n19696), .ZN(n11238) );
  AND3_X2 U11425 ( .A1(n9935), .A2(n11239), .A3(n10542), .ZN(n11226) );
  OR2_X1 U11426 ( .A1(n11984), .A2(n11968), .ZN(n12309) );
  AND2_X1 U11427 ( .A1(n10708), .A2(n10707), .ZN(n11004) );
  INV_X1 U11428 ( .A(n10551), .ZN(n10552) );
  AND3_X1 U11429 ( .A1(n10214), .A2(n10495), .A3(n10213), .ZN(n11249) );
  AND2_X1 U11430 ( .A1(n10214), .A2(n10495), .ZN(n10532) );
  NAND2_X1 U11431 ( .A1(n14155), .A2(n12398), .ZN(n12419) );
  NAND2_X1 U11432 ( .A1(n11971), .A2(n9912), .ZN(n13631) );
  NAND2_X1 U11433 ( .A1(n12337), .A2(n14155), .ZN(n12422) );
  NOR2_X1 U11434 ( .A1(n17875), .A2(n17884), .ZN(n17866) );
  NAND4_X1 U11435 ( .A1(n10689), .A2(n10688), .A3(n10687), .A4(n10686), .ZN(
        n11395) );
  INV_X1 U11436 ( .A(n18589), .ZN(n17659) );
  CLKBUF_X1 U11437 ( .A(n11962), .Z(n14016) );
  CLKBUF_X3 U11438 ( .A(n13071), .Z(n9736) );
  NAND3_X1 U11439 ( .A1(n10330), .A2(n10329), .A3(n10328), .ZN(n17206) );
  NOR2_X1 U11440 ( .A1(n13034), .A2(n10045), .ZN(n13031) );
  NAND2_X2 U11441 ( .A1(n10562), .A2(n14136), .ZN(n13059) );
  NAND2_X1 U11442 ( .A1(n10083), .A2(n10078), .ZN(n17709) );
  CLKBUF_X1 U11443 ( .A(n12017), .Z(n13954) );
  AOI211_X1 U11444 ( .C1(n17477), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n10327), .B(n10326), .ZN(n10328) );
  INV_X2 U11445 ( .A(n12017), .ZN(n11967) );
  NAND2_X1 U11446 ( .A1(n10490), .A2(n10489), .ZN(n10543) );
  INV_X1 U11447 ( .A(n11245), .ZN(n10494) );
  AND4_X1 U11448 ( .A1(n10079), .A2(n9800), .A3(n11675), .A4(n11676), .ZN(
        n10078) );
  CLKBUF_X3 U11449 ( .A(n10562), .Z(n14195) );
  OR2_X2 U11450 ( .A1(n16863), .A2(n16809), .ZN(n16866) );
  OR2_X1 U11451 ( .A1(n12003), .A2(n12002), .ZN(n12142) );
  OR2_X2 U11452 ( .A1(n11864), .A2(n11863), .ZN(n14661) );
  NAND2_X1 U11453 ( .A1(n9882), .A2(n9881), .ZN(n10562) );
  NAND2_X1 U11454 ( .A1(n10461), .A2(n10460), .ZN(n11245) );
  NAND2_X1 U11455 ( .A1(n10472), .A2(n10471), .ZN(n10493) );
  NAND2_X1 U11456 ( .A1(n10437), .A2(n10436), .ZN(n10489) );
  OR2_X2 U11457 ( .A1(n11895), .A2(n11894), .ZN(n11958) );
  INV_X2 U11458 ( .A(U214), .ZN(n16863) );
  NAND2_X1 U11459 ( .A1(n10119), .A2(n10118), .ZN(n19682) );
  NAND2_X1 U11460 ( .A1(n9778), .A2(n10429), .ZN(n10516) );
  NAND2_X1 U11461 ( .A1(n10511), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10517) );
  NAND2_X1 U11462 ( .A1(n10251), .A2(n10459), .ZN(n10460) );
  NAND2_X1 U11463 ( .A1(n10254), .A2(n10470), .ZN(n10471) );
  AND4_X1 U11464 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11953) );
  AND4_X1 U11465 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11931) );
  AND4_X1 U11466 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n11930) );
  AND4_X1 U11467 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11932) );
  AND4_X1 U11468 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11881) );
  AND4_X1 U11469 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11956) );
  AND4_X1 U11470 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11929) );
  AND2_X1 U11471 ( .A1(n10469), .A2(n10468), .ZN(n10470) );
  AND2_X1 U11472 ( .A1(n10423), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10427) );
  AND3_X1 U11473 ( .A1(n10439), .A2(n10438), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10442) );
  AND4_X1 U11474 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10511) );
  CLKBUF_X2 U11475 ( .A(n11924), .Z(n9737) );
  BUF_X2 U11476 ( .A(n11671), .Z(n17477) );
  NAND2_X1 U11477 ( .A1(n9745), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13287) );
  INV_X4 U11478 ( .A(n17525), .ZN(n17325) );
  BUF_X2 U11479 ( .A(n11924), .Z(n9738) );
  BUF_X2 U11480 ( .A(n12032), .Z(n12912) );
  AND2_X1 U11481 ( .A1(n10450), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10454) );
  AND2_X1 U11482 ( .A1(n10522), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10121) );
  AND2_X1 U11483 ( .A1(n9871), .A2(n9870), .ZN(n10501) );
  NAND2_X2 U11484 ( .A1(n20314), .A2(n20200), .ZN(n20249) );
  NAND2_X2 U11485 ( .A1(n19225), .A2(n19098), .ZN(n19155) );
  NOR2_X1 U11486 ( .A1(n13041), .A2(n19625), .ZN(n13042) );
  NOR2_X4 U11487 ( .A1(n10299), .A2(n10300), .ZN(n10331) );
  NAND2_X1 U11488 ( .A1(n9866), .A2(n9865), .ZN(n14469) );
  NOR2_X4 U11489 ( .A1(n10301), .A2(n17252), .ZN(n14480) );
  OR2_X1 U11490 ( .A1(n10299), .A2(n17252), .ZN(n14458) );
  OR2_X1 U11491 ( .A1(n19033), .A2(n10298), .ZN(n10309) );
  NOR2_X2 U11492 ( .A1(n19045), .A2(n18703), .ZN(n18740) );
  AND2_X2 U11493 ( .A1(n10637), .A2(n13819), .ZN(n10523) );
  AND2_X2 U11494 ( .A1(n10637), .A2(n13819), .ZN(n9744) );
  AND2_X2 U11495 ( .A1(n11849), .A2(n11847), .ZN(n11902) );
  AND2_X1 U11496 ( .A1(n11848), .A2(n11846), .ZN(n12032) );
  NOR2_X1 U11497 ( .A1(n19186), .A2(n19192), .ZN(n19012) );
  NAND2_X1 U11498 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19175), .ZN(
        n10299) );
  AND2_X2 U11499 ( .A1(n13638), .A2(n11846), .ZN(n9727) );
  NAND2_X1 U11500 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19198), .ZN(
        n10300) );
  AND2_X1 U11501 ( .A1(n11838), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11848) );
  NAND2_X1 U11502 ( .A1(n19186), .A2(n19175), .ZN(n10298) );
  NAND2_X2 U11503 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19192), .ZN(
        n10296) );
  AND2_X1 U11504 ( .A1(n11839), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11850) );
  AND2_X1 U11505 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10655) );
  INV_X2 U11506 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19198) );
  INV_X2 U11507 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19192) );
  INV_X2 U11508 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19186) );
  NOR2_X2 U11509 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11847) );
  AND2_X1 U11510 ( .A1(n9721), .A2(n10022), .ZN(n14897) );
  NOR2_X1 U11511 ( .A1(n14895), .A2(n14901), .ZN(n9721) );
  NOR2_X1 U11512 ( .A1(n14110), .A2(n10009), .ZN(n9722) );
  NOR2_X1 U11513 ( .A1(n14110), .A2(n10009), .ZN(n14268) );
  NAND2_X1 U11514 ( .A1(n14061), .A2(n14012), .ZN(n14110) );
  XNOR2_X1 U11515 ( .A(n12335), .B(n13787), .ZN(n14166) );
  OAI21_X1 U11516 ( .B1(n9758), .B2(n9880), .A(n10003), .ZN(n9879) );
  NAND2_X1 U11517 ( .A1(n10198), .A2(n9794), .ZN(n15144) );
  NAND2_X1 U11518 ( .A1(n16364), .A2(n16363), .ZN(n16362) );
  NAND2_X1 U11519 ( .A1(n14428), .A2(n10252), .ZN(n16364) );
  NAND2_X1 U11520 ( .A1(n10117), .A2(n13816), .ZN(n9723) );
  NAND2_X1 U11521 ( .A1(n10117), .A2(n13816), .ZN(n11376) );
  NAND2_X2 U11522 ( .A1(n10480), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10487) );
  NOR2_X2 U11523 ( .A1(n11448), .A2(n11447), .ZN(n11460) );
  NAND2_X2 U11524 ( .A1(n14596), .A2(n12610), .ZN(n14605) );
  NAND2_X1 U11525 ( .A1(n9884), .A2(n12063), .ZN(n14034) );
  BUF_X4 U11526 ( .A(n12111), .Z(n12950) );
  BUF_X2 U11527 ( .A(n11934), .Z(n12779) );
  NAND2_X1 U11528 ( .A1(n9914), .A2(n9913), .ZN(n12056) );
  XNOR2_X1 U11529 ( .A(n9888), .B(n12054), .ZN(n9914) );
  NOR2_X2 U11530 ( .A1(n18204), .A2(n17879), .ZN(n18211) );
  NOR2_X2 U11531 ( .A1(n17607), .A2(n17732), .ZN(n17603) );
  AOI221_X1 U11532 ( .B1(n18552), .B2(n14608), .C1(n17781), .C2(n14608), .A(
        n14612), .ZN(n16206) );
  NOR2_X2 U11533 ( .A1(n14600), .A2(n14601), .ZN(n10022) );
  AND2_X1 U11534 ( .A1(n15624), .A2(n9724), .ZN(n15588) );
  AND2_X1 U11535 ( .A1(n10908), .A2(n10093), .ZN(n9724) );
  NAND2_X1 U11536 ( .A1(n11226), .A2(n10547), .ZN(n9725) );
  NAND2_X1 U11537 ( .A1(n11226), .A2(n10547), .ZN(n13816) );
  INV_X2 U11538 ( .A(n14240), .ZN(n13121) );
  AND2_X2 U11539 ( .A1(n10539), .A2(n11249), .ZN(n11253) );
  OAI21_X2 U11540 ( .B1(n13053), .B2(n10042), .A(n10041), .ZN(n15358) );
  NOR2_X2 U11541 ( .A1(n13021), .A2(n16523), .ZN(n13020) );
  AOI21_X1 U11542 ( .B1(n12057), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12045), .ZN(n9888) );
  NOR2_X2 U11543 ( .A1(n11979), .A2(n11933), .ZN(n12311) );
  AOI21_X1 U11544 ( .B1(n15671), .B2(n15670), .A(n15722), .ZN(n15713) );
  OAI21_X2 U11545 ( .B1(n16597), .B2(n15665), .A(n16594), .ZN(n16586) );
  NOR2_X2 U11547 ( .A1(n11567), .A2(n11593), .ZN(n11590) );
  XNOR2_X1 U11548 ( .A(n13621), .B(n13620), .ZN(n20271) );
  NAND2_X1 U11549 ( .A1(n9750), .A2(n13625), .ZN(n10630) );
  XNOR2_X1 U11550 ( .A(n12137), .B(n12136), .ZN(n12495) );
  BUF_X4 U11551 ( .A(n12111), .Z(n12935) );
  NAND2_X1 U11552 ( .A1(n15765), .A2(n9712), .ZN(n9903) );
  NAND2_X1 U11553 ( .A1(n15760), .A2(n15762), .ZN(n9726) );
  NAND2_X1 U11554 ( .A1(n15760), .A2(n15762), .ZN(n15765) );
  INV_X2 U11555 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11845) );
  AND3_X2 U11556 ( .A1(n10544), .A2(n19682), .A3(n11245), .ZN(n10528) );
  NAND2_X2 U11557 ( .A1(n10553), .A2(n13873), .ZN(n10951) );
  OAI21_X1 U11558 ( .B1(n10488), .B2(n10490), .A(n10543), .ZN(n10950) );
  AOI211_X2 U11559 ( .C1(n15166), .C2(n20486), .A(n15165), .B(n15164), .ZN(
        n15167) );
  NAND2_X2 U11560 ( .A1(n16362), .A2(n12185), .ZN(n14584) );
  AND3_X1 U11561 ( .A1(n10431), .A2(n10430), .A3(n10429), .ZN(n10435) );
  INV_X2 U11562 ( .A(n13665), .ZN(n12302) );
  INV_X2 U11563 ( .A(n19682), .ZN(n10533) );
  NOR2_X2 U11564 ( .A1(n13017), .A2(n10051), .ZN(n13012) );
  AOI21_X1 U11565 ( .B1(n13011), .B2(n21192), .A(n10055), .ZN(n14555) );
  XNOR2_X2 U11566 ( .A(n12175), .B(n12168), .ZN(n14427) );
  AOI21_X1 U11567 ( .B1(n10644), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n10475), .ZN(n10476) );
  OAI211_X2 U11568 ( .C1(n9741), .C2(n13532), .A(n10565), .B(n10564), .ZN(
        n10598) );
  NOR2_X1 U11569 ( .A1(n16513), .A2(n19410), .ZN(n15348) );
  AND2_X4 U11570 ( .A1(n14769), .A2(n12863), .ZN(n14756) );
  NOR2_X2 U11571 ( .A1(n14783), .A2(n14785), .ZN(n14769) );
  XNOR2_X2 U11572 ( .A(n13382), .B(n10265), .ZN(n15419) );
  NAND2_X2 U11573 ( .A1(n15422), .A2(n9789), .ZN(n13382) );
  AND2_X2 U11574 ( .A1(n10790), .A2(n10789), .ZN(n15762) );
  BUF_X1 U11575 ( .A(n14721), .Z(n9730) );
  NOR2_X2 U11576 ( .A1(n14668), .A2(n20498), .ZN(n14667) );
  XNOR2_X1 U11577 ( .A(n10596), .B(n10595), .ZN(n13104) );
  NAND3_X2 U11578 ( .A1(n9869), .A2(n10748), .A3(n10151), .ZN(n10784) );
  AOI21_X2 U11579 ( .B1(n15063), .B2(n15198), .A(n15012), .ZN(n15014) );
  INV_X2 U11580 ( .A(n15033), .ZN(n15012) );
  NAND2_X2 U11581 ( .A1(n14323), .A2(n10760), .ZN(n19618) );
  NAND3_X2 U11582 ( .A1(n10092), .A2(n10758), .A3(n10784), .ZN(n14323) );
  NAND2_X4 U11583 ( .A1(n10487), .A2(n10486), .ZN(n10544) );
  NOR2_X2 U11584 ( .A1(n14006), .A2(n14234), .ZN(n14233) );
  INV_X1 U11585 ( .A(n15690), .ZN(n15691) );
  AND2_X1 U11586 ( .A1(n11849), .A2(n11846), .ZN(n9747) );
  AND2_X1 U11587 ( .A1(n11849), .A2(n11846), .ZN(n12957) );
  OAI21_X2 U11588 ( .B1(n16623), .B2(n10091), .A(n10089), .ZN(n15690) );
  AND2_X2 U11589 ( .A1(n11253), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9752) );
  AND2_X2 U11590 ( .A1(n10527), .A2(n13113), .ZN(n9756) );
  INV_X2 U11591 ( .A(n10493), .ZN(n10527) );
  BUF_X4 U11592 ( .A(n10650), .Z(n9739) );
  BUF_X4 U11593 ( .A(n10650), .Z(n9740) );
  NAND2_X1 U11594 ( .A1(n9723), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9741) );
  NOR2_X2 U11595 ( .A1(n13772), .A2(n13117), .ZN(n13894) );
  OAI21_X2 U11596 ( .B1(n13777), .B2(n13116), .A(n13773), .ZN(n13772) );
  INV_X1 U11597 ( .A(n10490), .ZN(n9742) );
  NAND2_X2 U11598 ( .A1(n10448), .A2(n10447), .ZN(n10490) );
  INV_X1 U11599 ( .A(n14156), .ZN(n9743) );
  AND2_X2 U11600 ( .A1(n10637), .A2(n13819), .ZN(n9745) );
  INV_X2 U11601 ( .A(n10544), .ZN(n11241) );
  AND3_X1 U11602 ( .A1(n13848), .A2(n10087), .A3(n9716), .ZN(n10650) );
  INV_X2 U11603 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13848) );
  AND2_X1 U11604 ( .A1(n11849), .A2(n11846), .ZN(n9746) );
  AND3_X2 U11605 ( .A1(n10534), .A2(n9756), .A3(n10449), .ZN(n10553) );
  OAI21_X2 U11606 ( .B1(n12495), .B2(n12147), .A(n12140), .ZN(n13611) );
  BUF_X4 U11607 ( .A(n13104), .Z(n9750) );
  AND2_X1 U11608 ( .A1(n11253), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9751) );
  NOR2_X1 U11609 ( .A1(n19061), .A2(n10414), .ZN(n17247) );
  NAND2_X1 U11610 ( .A1(n10492), .A2(n10491), .ZN(n10214) );
  AOI21_X1 U11611 ( .B1(n15105), .B2(n12232), .A(n9925), .ZN(n9924) );
  NAND2_X1 U11612 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  OR2_X1 U11613 ( .A1(n16537), .A2(n11444), .ZN(n11551) );
  NAND2_X1 U11614 ( .A1(n12300), .A2(n12299), .ZN(n13661) );
  NAND2_X1 U11615 ( .A1(n10938), .A2(n10937), .ZN(n20304) );
  NAND2_X1 U11616 ( .A1(n10936), .A2(n10935), .ZN(n10938) );
  AND2_X1 U11617 ( .A1(n9991), .A2(n14195), .ZN(n9990) );
  NOR2_X1 U11618 ( .A1(n10629), .A2(n13153), .ZN(n9988) );
  INV_X1 U11619 ( .A(n10212), .ZN(n10209) );
  AND2_X1 U11620 ( .A1(n12177), .A2(n12169), .ZN(n9896) );
  NAND2_X1 U11621 ( .A1(n9918), .A2(n12056), .ZN(n9917) );
  AND2_X1 U11622 ( .A1(n20548), .A2(n9919), .ZN(n9918) );
  INV_X1 U11623 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9919) );
  INV_X1 U11624 ( .A(n10075), .ZN(n10070) );
  NAND2_X1 U11625 ( .A1(n9898), .A2(n10189), .ZN(n12178) );
  NOR2_X1 U11626 ( .A1(n14284), .A2(n10190), .ZN(n9898) );
  NAND2_X1 U11627 ( .A1(n12220), .A2(n9757), .ZN(n9887) );
  INV_X1 U11628 ( .A(n9820), .ZN(n9886) );
  OR2_X1 U11629 ( .A1(n12015), .A2(n12014), .ZN(n12206) );
  NAND2_X1 U11630 ( .A1(n10189), .A2(n9897), .ZN(n12170) );
  AND2_X1 U11631 ( .A1(n15475), .A2(n15367), .ZN(n10124) );
  NAND2_X1 U11632 ( .A1(n15619), .A2(n15621), .ZN(n11567) );
  INV_X1 U11633 ( .A(n15861), .ZN(n10116) );
  AND2_X1 U11634 ( .A1(n9814), .A2(n15378), .ZN(n10113) );
  AND4_X1 U11635 ( .A1(n10259), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n11444) );
  NAND2_X1 U11636 ( .A1(n10506), .A2(n10429), .ZN(n9882) );
  NAND2_X1 U11637 ( .A1(n10505), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9881) );
  AND2_X1 U11638 ( .A1(n11420), .A2(n11399), .ZN(n10962) );
  INV_X1 U11639 ( .A(n17903), .ZN(n9972) );
  OR2_X1 U11640 ( .A1(n21064), .A2(n14152), .ZN(n20376) );
  OR2_X1 U11641 ( .A1(n15105), .A2(n9929), .ZN(n9923) );
  AND2_X1 U11642 ( .A1(n12315), .A2(n14709), .ZN(n12461) );
  INV_X1 U11643 ( .A(n10056), .ZN(n10055) );
  NAND2_X1 U11644 ( .A1(n10586), .A2(n10585), .ZN(n11288) );
  NAND2_X1 U11645 ( .A1(n10266), .A2(n10240), .ZN(n14240) );
  NOR2_X1 U11646 ( .A1(n10241), .A2(n9818), .ZN(n10240) );
  NAND2_X1 U11647 ( .A1(n10227), .A2(n13436), .ZN(n10229) );
  NAND2_X1 U11648 ( .A1(n13406), .A2(n10231), .ZN(n10230) );
  NAND2_X1 U11649 ( .A1(n16659), .A2(n9767), .ZN(n15893) );
  AOI22_X1 U11650 ( .A1(n13868), .A2(n13541), .B1(n13540), .B2(n13864), .ZN(
        n13573) );
  AND2_X1 U11651 ( .A1(n15523), .A2(n9774), .ZN(n15328) );
  NAND2_X1 U11652 ( .A1(n10435), .A2(n10434), .ZN(n10436) );
  NOR2_X2 U11653 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20259) );
  NOR2_X1 U11654 ( .A1(n20264), .A2(n20292), .ZN(n20048) );
  AND2_X1 U11655 ( .A1(n13536), .A2(n13661), .ZN(n13959) );
  AND2_X1 U11656 ( .A1(n19642), .A2(n13528), .ZN(n19613) );
  NAND2_X1 U11657 ( .A1(n12241), .A2(n12240), .ZN(n12245) );
  NAND2_X1 U11658 ( .A1(n12232), .A2(n9929), .ZN(n9926) );
  NAND2_X1 U11660 ( .A1(n11884), .A2(n11883), .ZN(n11911) );
  OAI22_X1 U11661 ( .A1(n10927), .A2(n10926), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20278), .ZN(n10933) );
  AND2_X1 U11662 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20278), .ZN(
        n10926) );
  OR2_X1 U11663 ( .A1(n10040), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10039) );
  INV_X1 U11664 ( .A(n11445), .ZN(n10040) );
  AND2_X1 U11665 ( .A1(n10644), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10739) );
  INV_X1 U11666 ( .A(n10833), .ZN(n10835) );
  OAI21_X1 U11667 ( .B1(n11234), .B2(n11241), .A(n10496), .ZN(n10555) );
  AND2_X1 U11668 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11726), .ZN(
        n11727) );
  INV_X1 U11669 ( .A(n17694), .ZN(n11776) );
  NOR2_X1 U11670 ( .A1(n17697), .A2(n11724), .ZN(n11725) );
  NOR2_X1 U11671 ( .A1(n17705), .A2(n11702), .ZN(n11721) );
  NAND2_X1 U11672 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19042), .ZN(
        n11757) );
  AND2_X1 U11673 ( .A1(n10187), .A2(n14733), .ZN(n10186) );
  NOR2_X1 U11674 ( .A1(n14746), .A2(n10188), .ZN(n10187) );
  INV_X1 U11675 ( .A(n14757), .ZN(n10188) );
  NOR2_X1 U11676 ( .A1(n14872), .A2(n10165), .ZN(n10164) );
  INV_X1 U11677 ( .A(n10166), .ZN(n10165) );
  NOR2_X1 U11678 ( .A1(n14621), .A2(n9919), .ZN(n12945) );
  NOR2_X1 U11679 ( .A1(n14893), .A2(n10175), .ZN(n10174) );
  INV_X1 U11680 ( .A(n14604), .ZN(n10175) );
  NAND2_X1 U11681 ( .A1(n12596), .A2(n12595), .ZN(n12610) );
  INV_X1 U11682 ( .A(n9710), .ZN(n12795) );
  NOR2_X2 U11683 ( .A1(n11957), .A2(n20913), .ZN(n12654) );
  NAND2_X1 U11684 ( .A1(n14000), .A2(n12158), .ZN(n12166) );
  AND2_X1 U11685 ( .A1(n12482), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12513) );
  OR2_X1 U11686 ( .A1(n11958), .A2(n20913), .ZN(n12943) );
  NOR2_X1 U11687 ( .A1(n9894), .A2(n15197), .ZN(n9891) );
  NOR2_X1 U11688 ( .A1(n12232), .A2(n12472), .ZN(n9894) );
  NAND2_X1 U11689 ( .A1(n15012), .A2(n10192), .ZN(n10191) );
  AND2_X1 U11690 ( .A1(n15035), .A2(n9848), .ZN(n10192) );
  INV_X1 U11691 ( .A(n10211), .ZN(n10210) );
  INV_X1 U11692 ( .A(n15107), .ZN(n10208) );
  NAND2_X1 U11693 ( .A1(n9920), .A2(n12146), .ZN(n12150) );
  NAND2_X1 U11694 ( .A1(n9917), .A2(n9915), .ZN(n9920) );
  NOR2_X1 U11695 ( .A1(n13954), .A2(n9919), .ZN(n12134) );
  NAND2_X1 U11696 ( .A1(n12044), .A2(n12043), .ZN(n10178) );
  INV_X1 U11697 ( .A(n12046), .ZN(n12054) );
  OAI21_X1 U11698 ( .B1(n13678), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12075), 
        .ZN(n12152) );
  INV_X1 U11699 ( .A(n20652), .ZN(n20516) );
  NOR2_X1 U11700 ( .A1(n11517), .A2(n10032), .ZN(n10031) );
  INV_X1 U11701 ( .A(n11490), .ZN(n10032) );
  AND2_X1 U11702 ( .A1(n10111), .A2(n15522), .ZN(n10110) );
  INV_X1 U11703 ( .A(n15341), .ZN(n10111) );
  NAND2_X1 U11704 ( .A1(n9832), .A2(n15430), .ZN(n10233) );
  AND2_X1 U11705 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  INV_X1 U11706 ( .A(n15452), .ZN(n10236) );
  INV_X1 U11707 ( .A(n15491), .ZN(n10239) );
  INV_X1 U11708 ( .A(n19424), .ZN(n10105) );
  INV_X1 U11709 ( .A(n14327), .ZN(n10107) );
  NAND2_X1 U11710 ( .A1(n10047), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10046) );
  INV_X1 U11711 ( .A(n10048), .ZN(n10047) );
  AND2_X1 U11712 ( .A1(n10709), .A2(n10747), .ZN(n10151) );
  NAND2_X1 U11713 ( .A1(n10133), .A2(n15426), .ZN(n10132) );
  INV_X1 U11714 ( .A(n15434), .ZN(n10133) );
  INV_X1 U11715 ( .A(n10007), .ZN(n9880) );
  NOR2_X1 U11716 ( .A1(n15711), .A2(n15721), .ZN(n9998) );
  INV_X1 U11717 ( .A(n15932), .ZN(n10005) );
  AND2_X1 U11718 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  INV_X1 U11719 ( .A(n14229), .ZN(n10126) );
  AND2_X1 U11720 ( .A1(n9783), .A2(n10008), .ZN(n10007) );
  INV_X1 U11721 ( .A(n16611), .ZN(n10008) );
  NAND2_X1 U11722 ( .A1(n10552), .A2(n9728), .ZN(n13069) );
  NOR2_X1 U11723 ( .A1(n19696), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10996) );
  NOR2_X1 U11724 ( .A1(n11455), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10989) );
  AND2_X1 U11725 ( .A1(n16038), .A2(n10527), .ZN(n10542) );
  AND2_X1 U11726 ( .A1(n10546), .A2(n10545), .ZN(n9935) );
  OAI21_X1 U11727 ( .B1(n10562), .B2(n10543), .A(n11241), .ZN(n10546) );
  INV_X1 U11728 ( .A(n10630), .ZN(n10613) );
  NAND2_X1 U11729 ( .A1(n21192), .A2(n10591), .ZN(n13511) );
  NOR2_X1 U11730 ( .A1(n9957), .A2(n9958), .ZN(n9953) );
  NOR2_X1 U11731 ( .A1(n10275), .A2(n9965), .ZN(n9957) );
  INV_X1 U11732 ( .A(n17853), .ZN(n9955) );
  NAND2_X1 U11733 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19186), .ZN(
        n10301) );
  INV_X1 U11734 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n21223) );
  OR2_X1 U11735 ( .A1(n17252), .A2(n10297), .ZN(n10245) );
  NOR2_X1 U11736 ( .A1(n18066), .A2(n9946), .ZN(n9945) );
  NOR2_X1 U11737 ( .A1(n18144), .A2(n9948), .ZN(n9947) );
  NAND2_X1 U11738 ( .A1(n10256), .A2(n11743), .ZN(n11744) );
  NAND2_X1 U11739 ( .A1(n18109), .A2(n18204), .ZN(n11743) );
  NAND2_X1 U11740 ( .A1(n11776), .A2(n11725), .ZN(n11815) );
  NOR2_X1 U11741 ( .A1(n18589), .A2(n18563), .ZN(n11804) );
  AND2_X1 U11742 ( .A1(n10395), .A2(n18552), .ZN(n9867) );
  NOR2_X1 U11743 ( .A1(n14438), .A2(n16741), .ZN(n14610) );
  AND2_X1 U11744 ( .A1(n20913), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12978) );
  XNOR2_X1 U11745 ( .A(n12166), .B(n12159), .ZN(n14218) );
  NAND2_X1 U11746 ( .A1(n15004), .A2(n12232), .ZN(n9911) );
  NAND2_X1 U11747 ( .A1(n15112), .A2(n10212), .ZN(n10206) );
  NAND2_X1 U11748 ( .A1(n12230), .A2(n12209), .ZN(n15151) );
  NAND2_X1 U11749 ( .A1(n12194), .A2(n9813), .ZN(n10202) );
  NAND2_X1 U11750 ( .A1(n10204), .A2(n9813), .ZN(n10201) );
  INV_X1 U11751 ( .A(n12194), .ZN(n10205) );
  NAND2_X1 U11752 ( .A1(n9749), .A2(n9919), .ZN(n12093) );
  NAND3_X1 U11753 ( .A1(n10528), .A2(n9756), .A3(n10449), .ZN(n13872) );
  NAND2_X1 U11754 ( .A1(n10576), .A2(n10575), .ZN(n10596) );
  NAND2_X1 U11755 ( .A1(n10242), .A2(n13119), .ZN(n10241) );
  INV_X1 U11756 ( .A(n10244), .ZN(n10242) );
  NOR2_X1 U11757 ( .A1(n10226), .A2(n10224), .ZN(n10223) );
  INV_X1 U11758 ( .A(n10231), .ZN(n10224) );
  INV_X1 U11759 ( .A(n10217), .ZN(n10216) );
  OAI21_X1 U11760 ( .B1(n13383), .B2(n10221), .A(n13403), .ZN(n10217) );
  INV_X1 U11761 ( .A(n15948), .ZN(n10114) );
  NAND2_X1 U11762 ( .A1(n9728), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19539) );
  AND2_X1 U11763 ( .A1(n9769), .A2(n13496), .ZN(n10122) );
  NOR2_X1 U11764 ( .A1(n15581), .A2(n10142), .ZN(n10141) );
  NOR2_X1 U11765 ( .A1(n10094), .A2(n15589), .ZN(n10093) );
  INV_X1 U11766 ( .A(n10095), .ZN(n10094) );
  NAND2_X1 U11767 ( .A1(n15609), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15611) );
  INV_X1 U11768 ( .A(n11567), .ZN(n15622) );
  OR3_X1 U11769 ( .A1(n16528), .A2(n11444), .A3(n15813), .ZN(n15630) );
  NAND2_X1 U11770 ( .A1(n15847), .A2(n10156), .ZN(n10159) );
  NOR2_X1 U11771 ( .A1(n15641), .A2(n10160), .ZN(n10156) );
  NAND2_X1 U11772 ( .A1(n15892), .A2(n9840), .ZN(n15538) );
  INV_X1 U11773 ( .A(n15535), .ZN(n10115) );
  NOR2_X2 U11774 ( .A1(n15893), .A2(n15894), .ZN(n15892) );
  NAND2_X1 U11775 ( .A1(n15671), .A2(n9998), .ZN(n9994) );
  AND2_X1 U11776 ( .A1(n15668), .A2(n16575), .ZN(n10000) );
  NAND2_X1 U11777 ( .A1(n16704), .A2(n10113), .ZN(n15936) );
  INV_X1 U11778 ( .A(n16684), .ZN(n9942) );
  AND2_X1 U11779 ( .A1(n10162), .A2(n11453), .ZN(n10161) );
  INV_X1 U11780 ( .A(n15745), .ZN(n10162) );
  NOR2_X1 U11781 ( .A1(n16705), .A2(n16706), .ZN(n16704) );
  NAND2_X1 U11782 ( .A1(n15958), .A2(n15957), .ZN(n16705) );
  NAND2_X1 U11783 ( .A1(n20264), .A2(n19453), .ZN(n19866) );
  AND2_X1 U11784 ( .A1(n20271), .A2(n20281), .ZN(n19931) );
  OAI22_X2 U11785 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16730), .B1(n20295), 
        .B2(n13515), .ZN(n20125) );
  INV_X1 U11786 ( .A(n20125), .ZN(n19874) );
  AND2_X1 U11787 ( .A1(n20304), .A2(n10948), .ZN(n13862) );
  INV_X1 U11788 ( .A(n18452), .ZN(n19004) );
  NOR2_X1 U11789 ( .A1(n16931), .A2(n16933), .ZN(n16932) );
  OAI21_X1 U11790 ( .B1(n9969), .B2(n9965), .A(n9970), .ZN(n9973) );
  NOR2_X1 U11791 ( .A1(n16992), .A2(n17903), .ZN(n16993) );
  INV_X1 U11792 ( .A(n10297), .ZN(n9865) );
  INV_X1 U11793 ( .A(n19033), .ZN(n9866) );
  CLKBUF_X2 U11794 ( .A(n11671), .Z(n17448) );
  CLKBUF_X2 U11795 ( .A(n11692), .Z(n14517) );
  INV_X1 U11796 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21174) );
  NOR2_X1 U11797 ( .A1(n10082), .A2(n10080), .ZN(n10079) );
  NAND2_X1 U11798 ( .A1(n11674), .A2(n10081), .ZN(n10080) );
  INV_X1 U11799 ( .A(n11677), .ZN(n10082) );
  NAND2_X1 U11800 ( .A1(n10342), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10081) );
  AOI22_X1 U11801 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11675) );
  NOR2_X2 U11802 ( .A1(n10298), .A2(n10300), .ZN(n11692) );
  CLKBUF_X1 U11803 ( .A(n9968), .Z(n9965) );
  NAND2_X1 U11804 ( .A1(n17112), .A2(n10261), .ZN(n17994) );
  NOR3_X1 U11805 ( .A1(n18109), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U11806 ( .A1(n18552), .A2(n18335), .ZN(n18397) );
  NAND2_X1 U11807 ( .A1(n10076), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10075) );
  INV_X1 U11808 ( .A(n10074), .ZN(n10072) );
  NAND2_X1 U11809 ( .A1(n18139), .A2(n10077), .ZN(n10074) );
  XNOR2_X1 U11810 ( .A(n11715), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18178) );
  INV_X1 U11811 ( .A(n13959), .ZN(n13554) );
  INV_X1 U11812 ( .A(n14969), .ZN(n14964) );
  INV_X2 U11813 ( .A(n15131), .ZN(n20474) );
  NAND2_X1 U11814 ( .A1(n10013), .A2(n10012), .ZN(n14829) );
  NAND2_X1 U11815 ( .A1(n9730), .A2(n10015), .ZN(n10013) );
  OR2_X1 U11816 ( .A1(n9730), .A2(n10014), .ZN(n10012) );
  XNOR2_X1 U11817 ( .A(n14644), .B(n12429), .ZN(n10015) );
  AND2_X1 U11818 ( .A1(n12461), .A2(n12432), .ZN(n20486) );
  NAND2_X1 U11819 ( .A1(n10059), .A2(n15604), .ZN(n10058) );
  AND2_X1 U11820 ( .A1(n13510), .A2(n13077), .ZN(n19431) );
  INV_X1 U11821 ( .A(n19447), .ZN(n19422) );
  INV_X1 U11822 ( .A(n19420), .ZN(n19454) );
  NOR2_X2 U11823 ( .A1(n15480), .A2(n19696), .ZN(n15492) );
  INV_X1 U11824 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19318) );
  NAND2_X1 U11825 ( .A1(n16580), .A2(n12997), .ZN(n9907) );
  NAND2_X1 U11826 ( .A1(n16650), .A2(n19622), .ZN(n9906) );
  NAND2_X1 U11827 ( .A1(n13524), .A2(n13001), .ZN(n19642) );
  NAND2_X1 U11828 ( .A1(n15778), .A2(n19669), .ZN(n10102) );
  OR2_X1 U11829 ( .A1(n15780), .A2(n15779), .ZN(n10101) );
  NAND2_X1 U11830 ( .A1(n15595), .A2(n15593), .ZN(n15580) );
  OR2_X1 U11831 ( .A1(n15328), .A2(n15327), .ZN(n15791) );
  AND2_X1 U11832 ( .A1(n16583), .A2(n11507), .ZN(n9908) );
  OR2_X1 U11833 ( .A1(n16010), .A2(n13578), .ZN(n20292) );
  INV_X1 U11834 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20288) );
  XNOR2_X1 U11835 ( .A(n13627), .B(n13628), .ZN(n20284) );
  INV_X1 U11836 ( .A(n20284), .ZN(n20281) );
  NAND2_X1 U11837 ( .A1(n13868), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16730) );
  INV_X1 U11838 ( .A(n19068), .ZN(n19213) );
  NOR2_X1 U11839 ( .A1(n16932), .A2(n19076), .ZN(n9983) );
  NAND2_X1 U11840 ( .A1(n16931), .A2(n16933), .ZN(n9984) );
  AND2_X1 U11841 ( .A1(n9981), .A2(n9822), .ZN(n9979) );
  OR2_X1 U11842 ( .A1(n16940), .A2(n19153), .ZN(n9981) );
  AND2_X1 U11843 ( .A1(n17266), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n9980) );
  INV_X1 U11844 ( .A(n17585), .ZN(n17580) );
  OR2_X2 U11845 ( .A1(n9863), .A2(n9862), .ZN(n17585) );
  INV_X1 U11846 ( .A(n17618), .ZN(n17647) );
  NOR2_X1 U11847 ( .A1(n16209), .A2(n16208), .ZN(n17716) );
  INV_X1 U11848 ( .A(n17716), .ZN(n17711) );
  NAND2_X1 U11849 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9871) );
  NAND2_X1 U11850 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9870) );
  OR2_X1 U11851 ( .A1(n12038), .A2(n12037), .ZN(n12141) );
  NAND2_X1 U11852 ( .A1(n9932), .A2(n12232), .ZN(n9927) );
  OR2_X1 U11853 ( .A1(n12117), .A2(n12116), .ZN(n12188) );
  NOR2_X1 U11854 ( .A1(n9916), .A2(n12147), .ZN(n9915) );
  INV_X1 U11855 ( .A(n12051), .ZN(n9916) );
  INV_X1 U11856 ( .A(n12435), .ZN(n12316) );
  NAND2_X1 U11857 ( .A1(n9739), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U11858 ( .A1(n9797), .A2(n9986), .ZN(n9989) );
  INV_X1 U11859 ( .A(n10668), .ZN(n10778) );
  NAND2_X1 U11860 ( .A1(n10667), .A2(n10666), .ZN(n10990) );
  OAI211_X1 U11861 ( .C1(n10950), .C2(n10494), .A(n10952), .B(n10527), .ZN(
        n11234) );
  AOI22_X1 U11862 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10497) );
  AND2_X1 U11863 ( .A1(n20298), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10913) );
  OAI21_X1 U11864 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19192), .A(
        n10396), .ZN(n10397) );
  AND2_X1 U11865 ( .A1(n12292), .A2(n12256), .ZN(n12287) );
  AND2_X1 U11866 ( .A1(n12243), .A2(n12244), .ZN(n12257) );
  OR2_X1 U11867 ( .A1(n12245), .A2(n12242), .ZN(n12243) );
  NAND2_X1 U11868 ( .A1(n12331), .A2(n10016), .ZN(n12335) );
  NAND2_X1 U11869 ( .A1(n12138), .A2(n14156), .ZN(n12327) );
  OR2_X1 U11870 ( .A1(n12845), .A2(n14791), .ZN(n12884) );
  INV_X1 U11871 ( .A(n14841), .ZN(n10167) );
  AND2_X1 U11872 ( .A1(n12774), .A2(n10170), .ZN(n10169) );
  INV_X1 U11873 ( .A(n14847), .ZN(n12774) );
  NOR2_X1 U11874 ( .A1(n14819), .A2(n10171), .ZN(n10170) );
  INV_X1 U11875 ( .A(n14855), .ZN(n10171) );
  INV_X1 U11876 ( .A(n12945), .ZN(n12972) );
  AND2_X1 U11877 ( .A1(n12691), .A2(n12673), .ZN(n10166) );
  NAND2_X1 U11878 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n12657), .ZN(
        n12675) );
  NOR2_X1 U11879 ( .A1(n14537), .A2(n10181), .ZN(n10180) );
  INV_X1 U11880 ( .A(n10182), .ZN(n10181) );
  NOR2_X1 U11881 ( .A1(n14421), .A2(n10183), .ZN(n10182) );
  INV_X1 U11882 ( .A(n14393), .ZN(n10183) );
  AND2_X1 U11883 ( .A1(n12525), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12532) );
  INV_X1 U11884 ( .A(n12654), .ZN(n12671) );
  OR2_X1 U11885 ( .A1(n12074), .A2(n12073), .ZN(n12162) );
  AOI21_X1 U11886 ( .B1(n15063), .B2(n12224), .A(n9933), .ZN(n9932) );
  NAND2_X1 U11887 ( .A1(n12226), .A2(n9934), .ZN(n9929) );
  NOR2_X1 U11888 ( .A1(n14874), .A2(n10020), .ZN(n10019) );
  INV_X1 U11889 ( .A(n14865), .ZN(n10020) );
  OR2_X1 U11890 ( .A1(n15113), .A2(n12220), .ZN(n9885) );
  NAND2_X1 U11891 ( .A1(n10199), .A2(n10202), .ZN(n10197) );
  OR2_X1 U11892 ( .A1(n12129), .A2(n12128), .ZN(n12200) );
  NAND2_X1 U11893 ( .A1(n12133), .A2(n12132), .ZN(n12198) );
  INV_X1 U11894 ( .A(n16460), .ZN(n10010) );
  NAND2_X1 U11895 ( .A1(n12166), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12167) );
  INV_X1 U11896 ( .A(n14109), .ZN(n12350) );
  INV_X1 U11897 ( .A(n14110), .ZN(n10011) );
  OR2_X1 U11898 ( .A1(n12462), .A2(n13789), .ZN(n14430) );
  NOR2_X1 U11899 ( .A1(n11965), .A2(n11960), .ZN(n11961) );
  OR2_X1 U11900 ( .A1(n13661), .A2(n12305), .ZN(n13667) );
  NAND2_X1 U11901 ( .A1(n10177), .A2(n10178), .ZN(n12076) );
  OR2_X1 U11902 ( .A1(n12091), .A2(n12090), .ZN(n12171) );
  AND2_X1 U11903 ( .A1(n12064), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12271) );
  NOR2_X1 U11904 ( .A1(n9717), .A2(n12138), .ZN(n10195) );
  NOR2_X1 U11905 ( .A1(n14156), .A2(n13665), .ZN(n10194) );
  OAI21_X1 U11906 ( .B1(n16184), .B2(n14048), .A(n13918), .ZN(n13919) );
  AND2_X1 U11907 ( .A1(n10929), .A2(n10928), .ZN(n10936) );
  NAND2_X1 U11908 ( .A1(n10026), .A2(n10025), .ZN(n11394) );
  NAND2_X1 U11909 ( .A1(n11004), .A2(n10027), .ZN(n10026) );
  NAND2_X1 U11910 ( .A1(n13059), .A2(n10960), .ZN(n10025) );
  NOR2_X1 U11911 ( .A1(n11570), .A2(n11571), .ZN(n11574) );
  OR2_X1 U11912 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n11558), .ZN(n11564) );
  NOR2_X1 U11913 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  INV_X1 U11914 ( .A(n11502), .ZN(n10030) );
  INV_X1 U11915 ( .A(n11476), .ZN(n10029) );
  NAND2_X1 U11916 ( .A1(n11477), .A2(n11476), .ZN(n11503) );
  NOR2_X1 U11917 ( .A1(n11448), .A2(n10036), .ZN(n11468) );
  INV_X1 U11918 ( .A(n10039), .ZN(n10038) );
  NOR3_X1 U11919 ( .A1(n11448), .A2(n11447), .A3(n10039), .ZN(n11467) );
  NOR3_X1 U11920 ( .A1(n11448), .A2(n11447), .A3(n10040), .ZN(n11456) );
  NAND2_X1 U11921 ( .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10056) );
  OR2_X1 U11922 ( .A1(n10745), .A2(n10744), .ZN(n11402) );
  NAND2_X1 U11923 ( .A1(n11405), .A2(n11410), .ZN(n11428) );
  NAND2_X1 U11924 ( .A1(n10024), .A2(n10023), .ZN(n11412) );
  NAND2_X1 U11925 ( .A1(n11455), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U11926 ( .A1(n11394), .A2(n10449), .ZN(n10024) );
  NAND2_X1 U11927 ( .A1(n10587), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9899) );
  INV_X1 U11928 ( .A(n11054), .ZN(n13303) );
  INV_X1 U11929 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9900) );
  AND2_X1 U11930 ( .A1(n13405), .A2(n13436), .ZN(n10231) );
  INV_X1 U11931 ( .A(n15418), .ZN(n10221) );
  AND2_X1 U11932 ( .A1(n13243), .A2(n15462), .ZN(n10237) );
  AND2_X1 U11933 ( .A1(n11241), .A2(n10493), .ZN(n10213) );
  AND2_X1 U11934 ( .A1(n11599), .A2(n15321), .ZN(n10137) );
  INV_X1 U11935 ( .A(n15464), .ZN(n10123) );
  AND2_X1 U11936 ( .A1(n14119), .A2(n14125), .ZN(n10127) );
  NAND2_X1 U11937 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10048) );
  INV_X1 U11938 ( .A(n11603), .ZN(n10109) );
  NOR2_X1 U11939 ( .A1(n11568), .A2(n11569), .ZN(n10095) );
  NOR2_X1 U11940 ( .A1(n10098), .A2(n15853), .ZN(n10097) );
  INV_X1 U11941 ( .A(n10099), .ZN(n10098) );
  INV_X1 U11942 ( .A(n16111), .ZN(n10108) );
  NAND2_X1 U11943 ( .A1(n10877), .A2(n10876), .ZN(n10901) );
  NAND2_X1 U11944 ( .A1(n9726), .A2(n15761), .ZN(n10875) );
  INV_X1 U11945 ( .A(n11434), .ZN(n9902) );
  NOR2_X1 U11946 ( .A1(n10878), .A2(n15987), .ZN(n9936) );
  AND2_X1 U11947 ( .A1(n10871), .A2(n10870), .ZN(n11437) );
  AND2_X1 U11948 ( .A1(n10151), .A2(n11016), .ZN(n9909) );
  AND3_X1 U11949 ( .A1(n11019), .A2(n11018), .A3(n11017), .ZN(n19424) );
  AND2_X1 U11950 ( .A1(n13580), .A2(n13579), .ZN(n13582) );
  NOR2_X1 U11951 ( .A1(n13376), .A2(n16037), .ZN(n13102) );
  AND2_X1 U11952 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10657), .ZN(
        n10965) );
  OR2_X1 U11953 ( .A1(n9750), .A2(n13096), .ZN(n10618) );
  NAND2_X1 U11954 ( .A1(n9987), .A2(n9904), .ZN(n19868) );
  NOR2_X1 U11955 ( .A1(n10629), .A2(n19629), .ZN(n9987) );
  AND2_X1 U11956 ( .A1(n10518), .A2(n10429), .ZN(n10120) );
  AOI22_X1 U11957 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10656), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U11958 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U11959 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10484) );
  AND2_X1 U11960 ( .A1(n10474), .A2(n10473), .ZN(n10479) );
  NAND2_X1 U11961 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10297) );
  NAND3_X1 U11962 ( .A1(n19012), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n19198), .ZN(n17476) );
  NOR2_X1 U11963 ( .A1(n10085), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10084) );
  INV_X1 U11964 ( .A(n10086), .ZN(n10085) );
  OR2_X1 U11965 ( .A1(n14607), .A2(n9868), .ZN(n11805) );
  NOR2_X1 U11966 ( .A1(n11727), .A2(n10070), .ZN(n10069) );
  AOI21_X1 U11967 ( .B1(n10409), .B2(n11757), .A(n10408), .ZN(n11758) );
  AOI211_X1 U11968 ( .C1(n11748), .C2(n10390), .A(n10389), .B(n11753), .ZN(
        n11809) );
  NOR2_X1 U11969 ( .A1(n19033), .A2(n10301), .ZN(n10342) );
  INV_X1 U11970 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16275) );
  AND2_X1 U11971 ( .A1(n12385), .A2(n12384), .ZN(n14883) );
  NAND2_X2 U11972 ( .A1(n12345), .A2(n12327), .ZN(n13786) );
  INV_X1 U11973 ( .A(n14155), .ZN(n14054) );
  AND2_X1 U11974 ( .A1(n12705), .A2(n12704), .ZN(n14872) );
  CLKBUF_X1 U11975 ( .A(n14861), .Z(n14862) );
  AND2_X1 U11976 ( .A1(n12488), .A2(n12505), .ZN(n10264) );
  NAND2_X1 U11977 ( .A1(n10264), .A2(n12504), .ZN(n13969) );
  AND2_X1 U11978 ( .A1(n13589), .A2(n13588), .ZN(n20414) );
  INV_X1 U11979 ( .A(n12943), .ZN(n12979) );
  INV_X1 U11980 ( .A(n14724), .ZN(n10185) );
  OR2_X1 U11981 ( .A1(n12923), .A2(n14737), .ZN(n12974) );
  NAND2_X1 U11982 ( .A1(n12793), .A2(n12792), .ZN(n12826) );
  INV_X1 U11983 ( .A(n12791), .ZN(n12793) );
  CLKBUF_X1 U11984 ( .A(n14797), .Z(n14798) );
  AND2_X1 U11985 ( .A1(n12757), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12758) );
  AND2_X1 U11986 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n12707), .ZN(
        n12757) );
  NOR2_X1 U11987 ( .A1(n12675), .A2(n16275), .ZN(n12676) );
  NOR2_X1 U11988 ( .A1(n10176), .A2(n10173), .ZN(n10172) );
  INV_X1 U11989 ( .A(n14888), .ZN(n10176) );
  INV_X1 U11990 ( .A(n10174), .ZN(n10173) );
  NOR2_X1 U11991 ( .A1(n12642), .A2(n16285), .ZN(n12657) );
  NAND2_X1 U11992 ( .A1(n12627), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12642) );
  INV_X1 U11993 ( .A(n12611), .ZN(n12627) );
  AND2_X1 U11994 ( .A1(n12592), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12593) );
  NAND2_X1 U11995 ( .A1(n12593), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12611) );
  NOR2_X1 U11996 ( .A1(n12577), .A2(n20344), .ZN(n12592) );
  INV_X1 U11997 ( .A(n12559), .ZN(n12562) );
  NAND2_X1 U11998 ( .A1(n12542), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12559) );
  AND2_X1 U11999 ( .A1(n12532), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12542) );
  AND2_X1 U12000 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12524), .ZN(
        n12525) );
  AOI21_X1 U12001 ( .B1(n12530), .B2(n12654), .A(n12529), .ZN(n14234) );
  INV_X1 U12002 ( .A(n14007), .ZN(n12522) );
  OR2_X1 U12003 ( .A1(n16179), .A2(n9919), .ZN(n13953) );
  XNOR2_X1 U12004 ( .A(n12429), .B(n12337), .ZN(n10014) );
  NAND2_X1 U12005 ( .A1(n9893), .A2(n12472), .ZN(n14993) );
  INV_X1 U12006 ( .A(n12229), .ZN(n9893) );
  INV_X1 U12007 ( .A(n10191), .ZN(n9895) );
  NAND2_X1 U12008 ( .A1(n10191), .A2(n12232), .ZN(n9892) );
  AND2_X1 U12009 ( .A1(n15044), .A2(n9891), .ZN(n9890) );
  NAND2_X1 U12010 ( .A1(n10019), .A2(n14857), .ZN(n10018) );
  NOR2_X1 U12011 ( .A1(n15105), .A2(n9930), .ZN(n15081) );
  NOR2_X1 U12012 ( .A1(n14885), .A2(n10017), .ZN(n14867) );
  INV_X1 U12013 ( .A(n10019), .ZN(n10017) );
  OR2_X1 U12014 ( .A1(n16269), .A2(n14883), .ZN(n14885) );
  NOR2_X1 U12015 ( .A1(n14885), .A2(n14874), .ZN(n14875) );
  XNOR2_X1 U12016 ( .A(n15063), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9883) );
  AND2_X1 U12017 ( .A1(n14897), .A2(n14889), .ZN(n16271) );
  NAND2_X1 U12018 ( .A1(n16271), .A2(n16270), .ZN(n16269) );
  NAND2_X1 U12019 ( .A1(n10022), .A2(n10021), .ZN(n14904) );
  INV_X1 U12020 ( .A(n14901), .ZN(n10021) );
  NOR2_X1 U12021 ( .A1(n15144), .A2(n9795), .ZN(n16347) );
  NAND2_X1 U12022 ( .A1(n9785), .A2(n14266), .ZN(n10009) );
  NAND2_X1 U12023 ( .A1(n10011), .A2(n12350), .ZN(n16461) );
  INV_X1 U12024 ( .A(n14433), .ZN(n20502) );
  AND2_X1 U12025 ( .A1(n16396), .A2(n16385), .ZN(n20495) );
  NAND2_X1 U12026 ( .A1(n20495), .A2(n20502), .ZN(n15300) );
  INV_X1 U12027 ( .A(n12050), .ZN(n9913) );
  NAND2_X1 U12028 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  NAND2_X1 U12029 ( .A1(n12081), .A2(n12080), .ZN(n14286) );
  NAND2_X1 U12030 ( .A1(n9919), .A2(n13919), .ZN(n14342) );
  CLKBUF_X1 U12031 ( .A(n12311), .Z(n12312) );
  NAND2_X1 U12032 ( .A1(n13661), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13918) );
  CLKBUF_X1 U12033 ( .A(n12319), .Z(n12320) );
  OR2_X1 U12034 ( .A1(n20650), .A2(n13917), .ZN(n20738) );
  INV_X1 U12035 ( .A(n20623), .ZN(n20615) );
  AND2_X1 U12036 ( .A1(n20652), .A2(n20651), .ZN(n20687) );
  INV_X1 U12037 ( .A(n20711), .ZN(n14293) );
  AND2_X1 U12038 ( .A1(n20650), .A2(n13917), .ZN(n20622) );
  NAND2_X1 U12039 ( .A1(n14065), .A2(n20516), .ZN(n20784) );
  NAND3_X1 U12040 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n9919), .A3(n13919), 
        .ZN(n14025) );
  OAI21_X1 U12041 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20817), .A(
        n20522), .ZN(n20910) );
  NOR2_X2 U12042 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20911) );
  AND2_X1 U12043 ( .A1(n20650), .A2(n9729), .ZN(n20574) );
  AND2_X1 U12044 ( .A1(n20652), .A2(n9897), .ZN(n20862) );
  INV_X1 U12045 ( .A(n10253), .ZN(n10059) );
  AND2_X1 U12046 ( .A1(n9736), .A2(n11455), .ZN(n10984) );
  OAI22_X1 U12047 ( .A1(n16521), .A2(n9838), .B1(n16514), .B2(n10049), .ZN(
        n16513) );
  OR2_X1 U12048 ( .A1(n16521), .A2(n16522), .ZN(n10050) );
  NOR2_X1 U12049 ( .A1(n11546), .A2(n10035), .ZN(n10034) );
  INV_X1 U12050 ( .A(n11537), .ZN(n10035) );
  NOR2_X1 U12051 ( .A1(n15358), .A2(n19410), .ZN(n16534) );
  OR2_X1 U12052 ( .A1(n19261), .A2(n19410), .ZN(n13491) );
  NOR2_X1 U12053 ( .A1(n19410), .A2(n15362), .ZN(n19262) );
  NOR2_X1 U12054 ( .A1(n19263), .A2(n19262), .ZN(n19261) );
  NAND2_X1 U12055 ( .A1(n11518), .A2(n10031), .ZN(n11521) );
  NAND2_X1 U12056 ( .A1(n10054), .A2(n13011), .ZN(n10053) );
  NOR2_X1 U12057 ( .A1(n13051), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10054) );
  OR2_X1 U12058 ( .A1(n13051), .A2(n10056), .ZN(n10052) );
  AND2_X1 U12059 ( .A1(n10137), .A2(n10136), .ZN(n10135) );
  INV_X1 U12060 ( .A(n13058), .ZN(n10136) );
  NAND2_X1 U12061 ( .A1(n15485), .A2(n10124), .ZN(n15463) );
  CLKBUF_X1 U12062 ( .A(n15460), .Z(n15461) );
  NAND2_X1 U12063 ( .A1(n13987), .A2(n9816), .ZN(n10244) );
  INV_X1 U12064 ( .A(n10266), .ZN(n10243) );
  NAND2_X1 U12065 ( .A1(n13092), .A2(n13091), .ZN(n13115) );
  NAND2_X1 U12066 ( .A1(n10227), .A2(n10225), .ZN(n10228) );
  NOR2_X1 U12067 ( .A1(n10226), .A2(n15407), .ZN(n10225) );
  NAND2_X1 U12068 ( .A1(n15523), .A2(n10110), .ZN(n15343) );
  NAND2_X1 U12069 ( .A1(n10218), .A2(n13407), .ZN(n15412) );
  NAND2_X1 U12070 ( .A1(n10219), .A2(n9759), .ZN(n10218) );
  XNOR2_X1 U12071 ( .A(n13360), .B(n13357), .ZN(n15424) );
  AND2_X1 U12072 ( .A1(n13265), .A2(n13264), .ZN(n15452) );
  AND2_X1 U12073 ( .A1(n11205), .A2(n11204), .ZN(n15894) );
  CLKBUF_X1 U12074 ( .A(n15466), .Z(n15467) );
  AND3_X1 U12075 ( .A1(n11176), .A2(n11175), .A3(n11174), .ZN(n16660) );
  NOR2_X1 U12076 ( .A1(n14558), .A2(n10104), .ZN(n19425) );
  NAND2_X1 U12077 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  OAI21_X1 U12078 ( .B1(n13489), .B2(n13488), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13715) );
  INV_X1 U12079 ( .A(n13715), .ZN(n14685) );
  OR2_X1 U12080 ( .A1(n10046), .A2(n21272), .ZN(n10045) );
  AND2_X1 U12081 ( .A1(n11317), .A2(n11316), .ZN(n14229) );
  NAND2_X1 U12082 ( .A1(n14120), .A2(n10127), .ZN(n14228) );
  AND2_X1 U12083 ( .A1(n11305), .A2(n11304), .ZN(n13982) );
  INV_X1 U12084 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13040) );
  NAND2_X1 U12085 ( .A1(n9869), .A2(n10709), .ZN(n10750) );
  NAND2_X1 U12086 ( .A1(n10748), .A2(n10747), .ZN(n10749) );
  NOR2_X1 U12087 ( .A1(n11578), .A2(n11579), .ZN(n10149) );
  INV_X1 U12088 ( .A(n15592), .ZN(n11578) );
  AND2_X1 U12089 ( .A1(n11576), .A2(n10150), .ZN(n11579) );
  NOR2_X1 U12090 ( .A1(n11444), .A2(n15779), .ZN(n10150) );
  AOI21_X1 U12091 ( .B1(n15622), .B2(n15788), .A(n10146), .ZN(n10144) );
  NAND2_X1 U12092 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  OAI21_X1 U12093 ( .B1(n11577), .B2(n11444), .A(n15589), .ZN(n15593) );
  NAND2_X1 U12094 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  INV_X1 U12095 ( .A(n15352), .ZN(n10131) );
  NOR2_X1 U12096 ( .A1(n10158), .A2(n15632), .ZN(n10157) );
  NOR3_X1 U12097 ( .A1(n15447), .A2(n15352), .A3(n15434), .ZN(n15433) );
  NAND2_X1 U12098 ( .A1(n10097), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10096) );
  NAND2_X1 U12099 ( .A1(n15692), .A2(n10097), .ZN(n15844) );
  NOR2_X1 U12100 ( .A1(n15881), .A2(n15864), .ZN(n10099) );
  AND2_X1 U12101 ( .A1(n15892), .A2(n9836), .ZN(n15859) );
  INV_X1 U12102 ( .A(n9879), .ZN(n9878) );
  NAND2_X1 U12103 ( .A1(n15892), .A2(n13497), .ZN(n15860) );
  OR2_X1 U12104 ( .A1(n15674), .A2(n9997), .ZN(n9993) );
  NAND2_X1 U12105 ( .A1(n9995), .A2(n15673), .ZN(n9992) );
  NAND2_X1 U12106 ( .A1(n15687), .A2(n15685), .ZN(n15689) );
  NAND2_X1 U12107 ( .A1(n16659), .A2(n9753), .ZN(n15565) );
  AND2_X1 U12108 ( .A1(n15485), .A2(n15475), .ZN(n15474) );
  NAND2_X1 U12109 ( .A1(n16124), .A2(n15669), .ZN(n15724) );
  NAND2_X1 U12110 ( .A1(n14251), .A2(n14250), .ZN(n15494) );
  AND2_X1 U12111 ( .A1(n11323), .A2(n11322), .ZN(n15495) );
  NAND2_X1 U12112 ( .A1(n16659), .A2(n16645), .ZN(n16644) );
  OAI21_X1 U12113 ( .B1(n10163), .B2(n10004), .A(n10001), .ZN(n16597) );
  INV_X1 U12114 ( .A(n10002), .ZN(n10001) );
  OAI21_X1 U12115 ( .B1(n10004), .B2(n10007), .A(n15931), .ZN(n10002) );
  AND2_X1 U12116 ( .A1(n16704), .A2(n9827), .ZN(n16672) );
  INV_X1 U12117 ( .A(n15935), .ZN(n10112) );
  NAND2_X1 U12118 ( .A1(n16672), .A2(n16671), .ZN(n16670) );
  NAND2_X1 U12119 ( .A1(n10163), .A2(n10007), .ZN(n10006) );
  INV_X1 U12120 ( .A(n16654), .ZN(n16669) );
  NAND2_X1 U12121 ( .A1(n10163), .A2(n9783), .ZN(n16609) );
  AND2_X1 U12122 ( .A1(n14120), .A2(n14119), .ZN(n14126) );
  NAND2_X1 U12123 ( .A1(n16704), .A2(n15948), .ZN(n16694) );
  NAND2_X1 U12124 ( .A1(n16623), .A2(n16624), .ZN(n10088) );
  AND2_X1 U12125 ( .A1(n19387), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16625) );
  NAND2_X1 U12126 ( .A1(n10530), .A2(n10551), .ZN(n11227) );
  INV_X1 U12127 ( .A(n9875), .ZN(n9874) );
  OR2_X1 U12128 ( .A1(n13872), .A2(n13062), .ZN(n20303) );
  NAND2_X1 U12129 ( .A1(n13101), .A2(n13100), .ZN(n13628) );
  AND2_X1 U12130 ( .A1(n21192), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13103) );
  OAI21_X1 U12131 ( .B1(n10489), .B2(n21192), .A(n19936), .ZN(n13105) );
  OAI22_X1 U12132 ( .A1(n13627), .A2(n13628), .B1(n13102), .B2(n16010), .ZN(
        n13620) );
  NAND2_X1 U12133 ( .A1(n10663), .A2(n10429), .ZN(n13826) );
  NAND2_X1 U12134 ( .A1(n10941), .A2(n10964), .ZN(n10942) );
  AND2_X1 U12135 ( .A1(n20271), .A2(n20284), .ZN(n19744) );
  INV_X1 U12136 ( .A(n19695), .ZN(n19686) );
  INV_X1 U12137 ( .A(n20257), .ZN(n20071) );
  NOR2_X1 U12138 ( .A1(n20264), .A2(n19453), .ZN(n20072) );
  NOR2_X2 U12139 ( .A1(n14685), .A2(n14135), .ZN(n19693) );
  NOR2_X2 U12140 ( .A1(n14688), .A2(n14135), .ZN(n19694) );
  INV_X1 U12141 ( .A(n19694), .ZN(n19701) );
  NAND2_X1 U12142 ( .A1(n19215), .A2(n18547), .ZN(n11801) );
  NOR2_X1 U12143 ( .A1(n19028), .A2(n11805), .ZN(n19000) );
  NOR2_X1 U12144 ( .A1(n9950), .A2(n9949), .ZN(n16944) );
  INV_X1 U12145 ( .A(n9952), .ZN(n9949) );
  AOI21_X1 U12146 ( .B1(n9953), .B2(n9955), .A(n9965), .ZN(n9952) );
  NAND2_X1 U12147 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  INV_X1 U12148 ( .A(n9957), .ZN(n9956) );
  NOR2_X1 U12149 ( .A1(n16963), .A2(n17867), .ZN(n16962) );
  NAND2_X1 U12150 ( .A1(n9971), .A2(n9958), .ZN(n9967) );
  NOR2_X1 U12152 ( .A1(n17877), .A2(n16971), .ZN(n16972) );
  OAI21_X1 U12153 ( .B1(n17055), .B2(n9963), .A(n9962), .ZN(n17046) );
  NAND2_X1 U12154 ( .A1(n9966), .A2(n9964), .ZN(n9963) );
  NAND2_X1 U12155 ( .A1(n9965), .A2(n9966), .ZN(n9962) );
  INV_X1 U12156 ( .A(n17984), .ZN(n9964) );
  NOR2_X1 U12157 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17082), .ZN(n17067) );
  AOI21_X1 U12158 ( .B1(n10289), .B2(n17256), .A(n9968), .ZN(n17066) );
  NOR2_X1 U12159 ( .A1(n18101), .A2(n18066), .ZN(n17125) );
  NOR2_X1 U12160 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17181), .ZN(n17162) );
  INV_X1 U12161 ( .A(n19231), .ZN(n17205) );
  NAND2_X1 U12162 ( .A1(n17595), .A2(n9861), .ZN(n9863) );
  NOR2_X1 U12163 ( .A1(n17727), .A2(n17799), .ZN(n9861) );
  NAND3_X1 U12164 ( .A1(n10352), .A2(n10351), .A3(n10350), .ZN(n17575) );
  AOI211_X1 U12165 ( .C1(n11704), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n10349), .B(n10348), .ZN(n10350) );
  NAND2_X1 U12166 ( .A1(n17720), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17658) );
  INV_X1 U12167 ( .A(n11664), .ZN(n11665) );
  AOI21_X1 U12168 ( .B1(n16206), .B2(n19213), .A(n16205), .ZN(n16208) );
  NAND4_X1 U12169 ( .A1(n11804), .A2(n18574), .A3(n10393), .A4(n17206), .ZN(
        n17781) );
  AND2_X1 U12170 ( .A1(n17866), .A2(n9829), .ZN(n10287) );
  NAND2_X1 U12171 ( .A1(n17866), .A2(n9763), .ZN(n16752) );
  NOR2_X1 U12172 ( .A1(n17843), .A2(n9960), .ZN(n9959) );
  INV_X1 U12173 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U12174 ( .A1(n17866), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17842) );
  NOR2_X1 U12175 ( .A1(n17884), .A2(n10277), .ZN(n17838) );
  NAND2_X1 U12176 ( .A1(n10281), .A2(n9810), .ZN(n17924) );
  NOR2_X1 U12177 ( .A1(n17963), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U12178 ( .A1(n18065), .A2(n9945), .ZN(n18014) );
  NOR2_X1 U12179 ( .A1(n18145), .A2(n18101), .ZN(n9943) );
  NAND2_X1 U12180 ( .A1(n9944), .A2(n9947), .ZN(n18064) );
  INV_X1 U12181 ( .A(n18145), .ZN(n9944) );
  NOR2_X1 U12182 ( .A1(n11819), .A2(n11818), .ZN(n11820) );
  NAND2_X1 U12183 ( .A1(n11816), .A2(n10067), .ZN(n17855) );
  NOR2_X1 U12184 ( .A1(n16190), .A2(n18107), .ZN(n10067) );
  NOR2_X1 U12185 ( .A1(n10066), .A2(n17904), .ZN(n17881) );
  NAND2_X1 U12186 ( .A1(n10065), .A2(n10064), .ZN(n17904) );
  INV_X1 U12187 ( .A(n11823), .ZN(n10064) );
  INV_X1 U12188 ( .A(n10065), .ZN(n17969) );
  NAND2_X1 U12189 ( .A1(n11739), .A2(n11738), .ZN(n17990) );
  NAND2_X1 U12190 ( .A1(n18106), .A2(n10084), .ZN(n18052) );
  NOR2_X1 U12191 ( .A1(n11746), .A2(n10391), .ZN(n19015) );
  NAND2_X1 U12192 ( .A1(n18106), .A2(n18107), .ZN(n18092) );
  NAND3_X1 U12193 ( .A1(n10320), .A2(n10319), .A3(n10318), .ZN(n14440) );
  AOI21_X1 U12194 ( .B1(n11766), .B2(n11765), .A(n11764), .ZN(n19003) );
  INV_X1 U12195 ( .A(n16913), .ZN(n19001) );
  INV_X1 U12196 ( .A(n19010), .ZN(n19031) );
  INV_X1 U12197 ( .A(n19025), .ZN(n19022) );
  INV_X1 U12198 ( .A(n19028), .ZN(n14608) );
  INV_X1 U12199 ( .A(n17578), .ZN(n18574) );
  INV_X1 U12200 ( .A(n17206), .ZN(n18547) );
  NAND2_X1 U12202 ( .A1(n19218), .A2(n18545), .ZN(n18657) );
  OAI22_X1 U12203 ( .A1(n18998), .A2(n19004), .B1(n18397), .B2(n16741), .ZN(
        n19059) );
  OR2_X1 U12204 ( .A1(n13568), .A2(n13953), .ZN(n13555) );
  AND2_X1 U12205 ( .A1(n16257), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16239) );
  INV_X1 U12206 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16285) );
  AND2_X1 U12207 ( .A1(n20376), .A2(n14168), .ZN(n20341) );
  AND2_X1 U12208 ( .A1(n20376), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21395) );
  INV_X1 U12209 ( .A(n21403), .ZN(n20368) );
  INV_X1 U12210 ( .A(n21395), .ZN(n20389) );
  INV_X1 U12211 ( .A(n20353), .ZN(n21391) );
  NAND2_X1 U12212 ( .A1(n14175), .A2(n14161), .ZN(n20373) );
  OR2_X1 U12213 ( .A1(n14722), .A2(n9730), .ZN(n15174) );
  INV_X1 U12214 ( .A(n14899), .ZN(n20405) );
  NAND2_X1 U12215 ( .A1(n14985), .A2(n14635), .ZN(n14969) );
  INV_X1 U12216 ( .A(n14985), .ZN(n14982) );
  INV_X1 U12217 ( .A(n14988), .ZN(n14983) );
  NAND2_X1 U12218 ( .A1(n13952), .A2(n14709), .ZN(n13961) );
  OR2_X1 U12219 ( .A1(n14982), .A2(n13963), .ZN(n14988) );
  NAND2_X1 U12220 ( .A1(n20321), .A2(n12984), .ZN(n15131) );
  NAND2_X1 U12221 ( .A1(n9922), .A2(n9921), .ZN(n15025) );
  NAND2_X1 U12222 ( .A1(n12229), .A2(n12230), .ZN(n9921) );
  NAND2_X1 U12223 ( .A1(n15024), .A2(n21407), .ZN(n9922) );
  NAND2_X1 U12224 ( .A1(n9923), .A2(n12232), .ZN(n15074) );
  NAND2_X1 U12225 ( .A1(n9931), .A2(n15063), .ZN(n15073) );
  NAND2_X1 U12226 ( .A1(n10200), .A2(n10201), .ZN(n15153) );
  OR2_X1 U12227 ( .A1(n14584), .A2(n10202), .ZN(n10200) );
  NAND2_X1 U12228 ( .A1(n10203), .A2(n12194), .ZN(n16358) );
  NAND2_X1 U12229 ( .A1(n14584), .A2(n10249), .ZN(n10203) );
  NOR2_X1 U12230 ( .A1(n20495), .A2(n14680), .ZN(n20493) );
  INV_X1 U12231 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20905) );
  CLKBUF_X1 U12232 ( .A(n13915), .Z(n20650) );
  INV_X1 U12233 ( .A(n20911), .ZN(n20915) );
  INV_X1 U12234 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14633) );
  NOR2_X1 U12235 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16471) );
  NOR2_X2 U12236 ( .A1(n20615), .A2(n20738), .ZN(n20570) );
  AND2_X1 U12237 ( .A1(n20623), .A2(n20622), .ZN(n20677) );
  AND2_X1 U12238 ( .A1(n20687), .A2(n13917), .ZN(n20732) );
  AND2_X1 U12239 ( .A1(n15315), .A2(n9729), .ZN(n20733) );
  OAI211_X1 U12240 ( .C1(n20817), .C2(n20771), .A(n20748), .B(n20814), .ZN(
        n20773) );
  NOR2_X1 U12241 ( .A1(n14291), .A2(n9729), .ZN(n20772) );
  AND2_X1 U12242 ( .A1(n20862), .A2(n20861), .ZN(n20972) );
  AND2_X1 U12243 ( .A1(n20862), .A2(n20547), .ZN(n20970) );
  NAND2_X1 U12244 ( .A1(n21247), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16179) );
  INV_X1 U12245 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21247) );
  NOR2_X1 U12246 ( .A1(n16500), .A2(n16501), .ZN(n16499) );
  NAND2_X1 U12247 ( .A1(n10043), .A2(n15654), .ZN(n10042) );
  NAND2_X1 U12248 ( .A1(n19410), .A2(n10043), .ZN(n10041) );
  INV_X1 U12249 ( .A(n16558), .ZN(n10043) );
  NOR2_X1 U12250 ( .A1(n16134), .A2(n16135), .ZN(n16133) );
  NOR2_X1 U12251 ( .A1(n13492), .A2(n19410), .ZN(n16134) );
  AND2_X1 U12252 ( .A1(n11518), .A2(n9811), .ZN(n11496) );
  NOR2_X1 U12253 ( .A1(n19269), .A2(n14555), .ZN(n15363) );
  NOR2_X1 U12254 ( .A1(n15364), .A2(n15363), .ZN(n15362) );
  NAND2_X1 U12255 ( .A1(n16486), .A2(n13075), .ZN(n19444) );
  OR2_X1 U12256 ( .A1(n19431), .A2(n19936), .ZN(n19420) );
  NOR2_X1 U12257 ( .A1(n14558), .A2(n11011), .ZN(n14328) );
  CLKBUF_X1 U12258 ( .A(n14240), .Z(n14241) );
  INV_X1 U12259 ( .A(n15492), .ZN(n15482) );
  NAND2_X1 U12260 ( .A1(n13121), .A2(n13120), .ZN(n15490) );
  AND2_X1 U12261 ( .A1(n14686), .A2(n14685), .ZN(n19461) );
  AND2_X1 U12262 ( .A1(n19489), .A2(n13575), .ZN(n19459) );
  AND2_X1 U12263 ( .A1(n16704), .A2(n9814), .ZN(n15379) );
  INV_X1 U12264 ( .A(n15576), .ZN(n19523) );
  INV_X1 U12265 ( .A(n19489), .ZN(n19522) );
  AND2_X1 U12266 ( .A1(n19489), .A2(n10992), .ZN(n19505) );
  INV_X1 U12267 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n21272) );
  INV_X1 U12268 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16637) );
  INV_X1 U12269 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19625) );
  INV_X1 U12270 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19641) );
  INV_X1 U12271 ( .A(n16568), .ZN(n19636) );
  INV_X1 U12272 ( .A(n13099), .ZN(n15396) );
  INV_X1 U12273 ( .A(n19613), .ZN(n19634) );
  NOR2_X1 U12274 ( .A1(n13524), .A2(n14195), .ZN(n16568) );
  XNOR2_X1 U12275 ( .A(n9872), .B(n11596), .ZN(n15608) );
  NAND2_X1 U12276 ( .A1(n15613), .A2(n10263), .ZN(n9872) );
  NAND2_X1 U12277 ( .A1(n10159), .A2(n15640), .ZN(n15633) );
  NAND2_X1 U12278 ( .A1(n15892), .A2(n9772), .ZN(n15536) );
  NAND2_X1 U12279 ( .A1(n9994), .A2(n9996), .ZN(n15702) );
  INV_X1 U12280 ( .A(n10090), .ZN(n10089) );
  OAI21_X1 U12281 ( .B1(n16624), .B2(n10091), .A(n15887), .ZN(n10090) );
  INV_X1 U12282 ( .A(n10907), .ZN(n10091) );
  NOR2_X1 U12283 ( .A1(n16144), .A2(n16145), .ZN(n9939) );
  NOR2_X1 U12284 ( .A1(n16726), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9941) );
  NAND2_X1 U12285 ( .A1(n15667), .A2(n16575), .ZN(n16122) );
  AND2_X1 U12286 ( .A1(n10163), .A2(n10161), .ZN(n15732) );
  NAND2_X1 U12287 ( .A1(n10163), .A2(n11453), .ZN(n15747) );
  INV_X1 U12288 ( .A(n15761), .ZN(n15764) );
  NAND2_X1 U12289 ( .A1(n14321), .A2(n14322), .ZN(n9876) );
  INV_X1 U12290 ( .A(n19667), .ZN(n19645) );
  INV_X1 U12291 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20298) );
  NOR2_X1 U12292 ( .A1(n13514), .A2(n10591), .ZN(n20295) );
  OR2_X1 U12293 ( .A1(n20271), .A2(n20281), .ZN(n20257) );
  INV_X1 U12294 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16203) );
  NOR2_X1 U12295 ( .A1(n19708), .A2(n19866), .ZN(n19762) );
  NOR2_X1 U12296 ( .A1(n19866), .A2(n20260), .ZN(n19801) );
  INV_X1 U12297 ( .A(n16055), .ZN(n16060) );
  OAI21_X1 U12298 ( .B1(n19909), .B2(n19908), .A(n19907), .ZN(n19926) );
  OAI22_X1 U12299 ( .A1(n19940), .A2(n19939), .B1(n19938), .B2(n13514), .ZN(
        n19958) );
  NOR2_X1 U12300 ( .A1(n20002), .A2(n20260), .ZN(n19992) );
  INV_X1 U12301 ( .A(n19992), .ZN(n20001) );
  OR2_X1 U12302 ( .A1(n20007), .A2(n20006), .ZN(n20035) );
  INV_X1 U12303 ( .A(n20130), .ZN(n20080) );
  INV_X1 U12304 ( .A(n20141), .ZN(n20092) );
  INV_X1 U12305 ( .A(n20147), .ZN(n20095) );
  OAI22_X1 U12306 ( .A1(n16825), .A2(n19701), .B1(n18581), .B2(n19699), .ZN(
        n20105) );
  AND2_X1 U12307 ( .A1(n20048), .A2(n20047), .ZN(n20109) );
  INV_X1 U12308 ( .A(n19881), .ZN(n20127) );
  INV_X1 U12309 ( .A(n20055), .ZN(n20138) );
  AND2_X1 U12310 ( .A1(n10544), .A2(n19686), .ZN(n20142) );
  INV_X1 U12311 ( .A(n19951), .ZN(n20150) );
  INV_X1 U12312 ( .A(n19725), .ZN(n20148) );
  INV_X1 U12313 ( .A(n19973), .ZN(n20156) );
  INV_X1 U12314 ( .A(n20177), .ZN(n20163) );
  INV_X1 U12315 ( .A(n19730), .ZN(n20160) );
  NAND2_X1 U12316 ( .A1(n20072), .A2(n20071), .ZN(n20177) );
  AND2_X1 U12317 ( .A1(n20294), .A2(n10971), .ZN(n20302) );
  NAND2_X1 U12318 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10981), .ZN(n19533) );
  AND2_X1 U12319 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n10591), .ZN(n10981) );
  INV_X1 U12320 ( .A(n19533), .ZN(n13899) );
  AND3_X1 U12321 ( .A1(n20189), .A2(n20247), .A3(n20194), .ZN(n20188) );
  INV_X2 U12322 ( .A(n20315), .ZN(n20314) );
  OR2_X1 U12323 ( .A1(n20182), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n20315) );
  AND2_X1 U12324 ( .A1(n17781), .A2(n11754), .ZN(n16914) );
  NAND2_X1 U12325 ( .A1(n19213), .A2(n19059), .ZN(n16915) );
  NOR2_X1 U12326 ( .A1(n16993), .A2(n9965), .ZN(n16985) );
  INV_X1 U12327 ( .A(n9973), .ZN(n16984) );
  NOR2_X1 U12328 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17014), .ZN(n17002) );
  NOR2_X1 U12329 ( .A1(n19136), .A2(n17021), .ZN(n17020) );
  NOR2_X1 U12330 ( .A1(n17065), .A2(n9968), .ZN(n17055) );
  NOR2_X1 U12331 ( .A1(n17055), .A2(n17984), .ZN(n17054) );
  NOR2_X1 U12332 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17128), .ZN(n17111) );
  INV_X1 U12333 ( .A(n17244), .ZN(n17254) );
  INV_X1 U12334 ( .A(n17247), .ZN(n17245) );
  INV_X1 U12335 ( .A(n17268), .ZN(n17246) );
  INV_X1 U12336 ( .A(n17266), .ZN(n17259) );
  NOR3_X1 U12337 ( .A1(n17274), .A2(n17333), .A3(n17332), .ZN(n17320) );
  NOR2_X1 U12338 ( .A1(n17659), .A2(n17374), .ZN(n17362) );
  INV_X1 U12339 ( .A(n17377), .ZN(n17375) );
  NAND2_X1 U12340 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17375), .ZN(n17374) );
  NAND2_X1 U12341 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17415), .ZN(n17402) );
  INV_X1 U12342 ( .A(n17432), .ZN(n17415) );
  NOR2_X1 U12343 ( .A1(n17560), .A2(n17537), .ZN(n17548) );
  INV_X1 U12344 ( .A(n17572), .ZN(n17560) );
  NOR3_X1 U12345 ( .A1(n18552), .A2(n18547), .A3(n16204), .ZN(n17572) );
  INV_X1 U12346 ( .A(n17598), .ZN(n17595) );
  NAND2_X1 U12347 ( .A1(n17595), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17594) );
  NAND2_X1 U12348 ( .A1(n17603), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17598) );
  NOR2_X1 U12349 ( .A1(n17613), .A2(n17659), .ZN(n17608) );
  NAND2_X1 U12350 ( .A1(n17608), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17607) );
  NAND2_X1 U12351 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17653), .ZN(n17649) );
  NOR2_X1 U12352 ( .A1(n17834), .A2(n17661), .ZN(n17653) );
  NOR2_X1 U12353 ( .A1(n17658), .A2(n17689), .ZN(n17686) );
  NOR2_X1 U12354 ( .A1(n11634), .A2(n11633), .ZN(n17694) );
  NOR2_X1 U12355 ( .A1(n11644), .A2(n11643), .ZN(n17697) );
  INV_X1 U12356 ( .A(n11678), .ZN(n10083) );
  INV_X1 U12357 ( .A(n17708), .ZN(n17718) );
  NOR2_X1 U12358 ( .A1(n17719), .A2(n19037), .ZN(n17717) );
  NOR2_X1 U12359 ( .A1(n16208), .A2(n21141), .ZN(n17720) );
  NOR2_X2 U12360 ( .A1(n10341), .A2(n10340), .ZN(n18589) );
  INV_X1 U12361 ( .A(n17717), .ZN(n17714) );
  NOR2_X1 U12362 ( .A1(n17784), .A2(n17723), .ZN(n17770) );
  NOR2_X1 U12363 ( .A1(n17778), .A2(n17770), .ZN(n17773) );
  CLKBUF_X1 U12364 ( .A(n17773), .Z(n17777) );
  NOR2_X1 U12365 ( .A1(n17784), .A2(n19062), .ZN(n17824) );
  NOR2_X1 U12366 ( .A1(n17830), .A2(n18552), .ZN(n17831) );
  AND2_X1 U12367 ( .A1(n10281), .A2(n9974), .ZN(n17902) );
  AND2_X1 U12368 ( .A1(n9810), .A2(n9975), .ZN(n9974) );
  INV_X1 U12369 ( .A(n17925), .ZN(n9975) );
  AND2_X1 U12370 ( .A1(n10281), .A2(n9976), .ZN(n17949) );
  NOR2_X1 U12371 ( .A1(n18046), .A2(n18036), .ZN(n18030) );
  INV_X1 U12372 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18036) );
  INV_X1 U12373 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18046) );
  INV_X1 U12374 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18118) );
  NOR2_X1 U12375 ( .A1(n18145), .A2(n18144), .ZN(n18129) );
  NAND2_X1 U12376 ( .A1(n17185), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18145) );
  INV_X1 U12377 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18184) );
  OAI21_X1 U12378 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19212), .A(n16915), 
        .ZN(n18197) );
  INV_X1 U12379 ( .A(n18143), .ZN(n18202) );
  INV_X1 U12380 ( .A(n18191), .ZN(n18201) );
  XNOR2_X1 U12381 ( .A(n16103), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16779) );
  NAND2_X1 U12382 ( .A1(n16188), .A2(n16102), .ZN(n16103) );
  NOR2_X1 U12383 ( .A1(n18523), .A2(n18512), .ZN(n18458) );
  AND2_X1 U12384 ( .A1(n18106), .A2(n10086), .ZN(n18061) );
  NAND2_X1 U12385 ( .A1(n19031), .A2(n19038), .ZN(n18413) );
  NOR2_X1 U12386 ( .A1(n18399), .A2(n18106), .ZN(n18443) );
  NAND2_X1 U12387 ( .A1(n18138), .A2(n10075), .ZN(n10073) );
  INV_X1 U12388 ( .A(n18530), .ZN(n18512) );
  NAND2_X1 U12389 ( .A1(n18999), .A2(n18512), .ZN(n18521) );
  CLKBUF_X1 U12390 ( .A(n18418), .Z(n18529) );
  INV_X1 U12391 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19042) );
  INV_X1 U12392 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19049) );
  INV_X1 U12393 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19053) );
  AOI211_X1 U12394 ( .C1(n19213), .C2(n19035), .A(n18546), .B(n14613), .ZN(
        n19199) );
  INV_X1 U12395 ( .A(n17229), .ZN(n19076) );
  INV_X1 U12396 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19169) );
  NAND2_X1 U12397 ( .A1(n19096), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19226) );
  AND2_X1 U12398 ( .A1(n13478), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14918)
         );
  CLKBUF_X1 U12399 ( .A(n16890), .Z(n16900) );
  AOI21_X1 U12400 ( .B1(n14829), .B2(n20486), .A(n12477), .ZN(n12478) );
  AOI21_X1 U12401 ( .B1(n15334), .B2(n15333), .A(n15332), .ZN(n15335) );
  OAI21_X1 U12402 ( .B1(n15773), .B2(n13461), .A(n13462), .ZN(n13463) );
  AOI21_X1 U12403 ( .B1(n9784), .B2(n16632), .A(n9905), .ZN(n16581) );
  NAND2_X1 U12404 ( .A1(n9907), .A2(n9906), .ZN(n9905) );
  OAI21_X1 U12405 ( .B1(n15777), .B2(n19667), .A(n9792), .ZN(n15781) );
  OAI21_X1 U12406 ( .B1(n9940), .B2(n16148), .A(n9937), .ZN(P2_U3029) );
  NOR2_X1 U12407 ( .A1(n9787), .A2(n9938), .ZN(n9937) );
  NOR2_X1 U12408 ( .A1(n16141), .A2(n9941), .ZN(n9940) );
  OAI21_X1 U12409 ( .B1(n16150), .B2(n16702), .A(n9939), .ZN(n9938) );
  NAND2_X1 U12410 ( .A1(n9982), .A2(n9978), .ZN(P3_U2642) );
  AND2_X1 U12411 ( .A1(n16939), .A2(n9979), .ZN(n9978) );
  NAND2_X1 U12412 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  NAND2_X1 U12413 ( .A1(n17581), .A2(n9864), .ZN(P3_U2705) );
  AND2_X1 U12414 ( .A1(n17582), .A2(n9821), .ZN(n9864) );
  INV_X1 U12415 ( .A(n11592), .ZN(n10147) );
  AND2_X1 U12416 ( .A1(n13934), .A2(n12302), .ZN(n11970) );
  INV_X1 U12417 ( .A(n10168), .ZN(n14818) );
  INV_X1 U12418 ( .A(n10238), .ZN(n15486) );
  AND2_X1 U12419 ( .A1(n9765), .A2(n9819), .ZN(n9753) );
  INV_X1 U12420 ( .A(n10656), .ZN(n13451) );
  INV_X1 U12422 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13043) );
  INV_X2 U12424 ( .A(n12230), .ZN(n12232) );
  INV_X1 U12425 ( .A(n10562), .ZN(n13071) );
  NAND2_X1 U12426 ( .A1(n15460), .A2(n10237), .ZN(n15450) );
  OR2_X1 U12427 ( .A1(n13034), .A2(n10046), .ZN(n9754) );
  AND2_X1 U12428 ( .A1(n13121), .A2(n9807), .ZN(n9755) );
  NAND2_X1 U12429 ( .A1(n12674), .A2(n12673), .ZN(n14880) );
  AND2_X1 U12430 ( .A1(n13029), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13049) );
  NOR2_X1 U12431 ( .A1(n9717), .A2(n14156), .ZN(n11980) );
  NAND2_X1 U12432 ( .A1(n14854), .A2(n14855), .ZN(n14817) );
  OR2_X1 U12433 ( .A1(n12232), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9757) );
  AND2_X1 U12434 ( .A1(n11440), .A2(n9815), .ZN(n9758) );
  NAND2_X1 U12435 ( .A1(n12674), .A2(n10166), .ZN(n14871) );
  NOR2_X1 U12436 ( .A1(n16962), .A2(n9965), .ZN(n16952) );
  NOR2_X1 U12437 ( .A1(n15440), .A2(n13318), .ZN(n15429) );
  AND2_X1 U12438 ( .A1(n10220), .A2(n13402), .ZN(n9759) );
  INV_X1 U12439 ( .A(n9997), .ZN(n9996) );
  NOR2_X1 U12440 ( .A1(n15711), .A2(n9999), .ZN(n9997) );
  NAND2_X1 U12441 ( .A1(n11567), .A2(n11593), .ZN(n9760) );
  NAND2_X1 U12442 ( .A1(n14854), .A2(n10170), .ZN(n10168) );
  OAI21_X1 U12443 ( .B1(n10205), .B2(n10249), .A(n16356), .ZN(n10204) );
  AND2_X1 U12444 ( .A1(n10106), .A2(n9817), .ZN(n9761) );
  INV_X1 U12445 ( .A(n11259), .ZN(n11374) );
  INV_X1 U12446 ( .A(n13461), .ZN(n15499) );
  AND2_X1 U12447 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9762) );
  AND2_X1 U12448 ( .A1(n9959), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9763) );
  AND2_X1 U12449 ( .A1(n10034), .A2(n10033), .ZN(n9764) );
  AND2_X1 U12450 ( .A1(n10108), .A2(n16645), .ZN(n9765) );
  AND2_X1 U12451 ( .A1(n9762), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9766) );
  AND2_X1 U12452 ( .A1(n9753), .A2(n9845), .ZN(n9767) );
  AND2_X1 U12453 ( .A1(n13120), .A2(n10239), .ZN(n9768) );
  AND2_X1 U12454 ( .A1(n10124), .A2(n10123), .ZN(n9769) );
  AND2_X1 U12455 ( .A1(n9764), .A2(n11555), .ZN(n9770) );
  AND2_X1 U12456 ( .A1(n9766), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9771) );
  INV_X1 U12457 ( .A(n15401), .ZN(n10226) );
  AND2_X1 U12458 ( .A1(n9836), .A2(n15354), .ZN(n9772) );
  AND2_X1 U12459 ( .A1(n10110), .A2(n10109), .ZN(n9773) );
  AND2_X1 U12460 ( .A1(n9773), .A2(n15326), .ZN(n9774) );
  OR3_X1 U12461 ( .A1(n14885), .A2(n10018), .A3(n14822), .ZN(n9775) );
  NOR2_X1 U12462 ( .A1(n15679), .A2(n15881), .ZN(n15657) );
  NAND2_X1 U12463 ( .A1(n11441), .A2(n9758), .ZN(n10163) );
  NAND2_X1 U12464 ( .A1(n11441), .A2(n11440), .ZN(n15753) );
  NAND2_X1 U12465 ( .A1(n11376), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10590) );
  AND2_X1 U12466 ( .A1(n11477), .A2(n10028), .ZN(n9776) );
  AND2_X1 U12467 ( .A1(n15523), .A2(n9773), .ZN(n9777) );
  NOR2_X1 U12468 ( .A1(n13038), .A2(n13040), .ZN(n13039) );
  AND2_X1 U12469 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13044) );
  INV_X2 U12470 ( .A(n12332), .ZN(n12328) );
  NAND2_X2 U12471 ( .A1(n13934), .A2(n14157), .ZN(n12345) );
  INV_X1 U12472 ( .A(n10004), .ZN(n10003) );
  NAND2_X1 U12473 ( .A1(n11474), .A2(n10005), .ZN(n10004) );
  AND4_X1 U12474 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n9778) );
  AND2_X1 U12475 ( .A1(n14605), .A2(n10174), .ZN(n9779) );
  NAND2_X1 U12476 ( .A1(n14605), .A2(n14604), .ZN(n14603) );
  OR2_X1 U12477 ( .A1(n10555), .A2(n13059), .ZN(n9780) );
  AND2_X1 U12478 ( .A1(n10635), .A2(n10634), .ZN(n9781) );
  OR2_X1 U12480 ( .A1(n15447), .A2(n15352), .ZN(n9782) );
  AND2_X1 U12481 ( .A1(n10161), .A2(n15734), .ZN(n9783) );
  NOR2_X1 U12482 ( .A1(n9908), .A2(n16579), .ZN(n9784) );
  NAND2_X1 U12483 ( .A1(n10006), .A2(n11474), .ZN(n15930) );
  NOR2_X2 U12484 ( .A1(n11815), .A2(n17691), .ZN(n18109) );
  AND2_X1 U12485 ( .A1(n12350), .A2(n10010), .ZN(n9785) );
  INV_X1 U12486 ( .A(n13059), .ZN(n10027) );
  NAND2_X1 U12487 ( .A1(n15692), .A2(n10099), .ZN(n15659) );
  OAI21_X1 U12488 ( .B1(n15440), .B2(n10234), .A(n10233), .ZN(n13360) );
  AND4_X1 U12489 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n9786) );
  NAND2_X1 U12490 ( .A1(n10216), .A2(n10215), .ZN(n13407) );
  NAND2_X1 U12491 ( .A1(n9895), .A2(n12229), .ZN(n14991) );
  AND2_X1 U12492 ( .A1(n10087), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10637) );
  NOR3_X1 U12493 ( .A1(n14749), .A2(n14720), .A3(n14736), .ZN(n14721) );
  AND3_X1 U12494 ( .A1(n16149), .A2(n16148), .A3(n16147), .ZN(n9787) );
  INV_X1 U12495 ( .A(n10219), .ZN(n15417) );
  OR2_X1 U12496 ( .A1(n10071), .A2(n11727), .ZN(n9788) );
  OR2_X1 U12497 ( .A1(n13360), .A2(n13361), .ZN(n9789) );
  INV_X1 U12498 ( .A(n10128), .ZN(n15425) );
  NOR3_X1 U12499 ( .A1(n15447), .A2(n10132), .A3(n15352), .ZN(n10128) );
  INV_X1 U12500 ( .A(n14661), .ZN(n11962) );
  OR2_X1 U12501 ( .A1(n15586), .A2(n15585), .ZN(n9790) );
  AND2_X1 U12502 ( .A1(n13406), .A2(n13405), .ZN(n9791) );
  AND3_X1 U12503 ( .A1(n10102), .A2(n15775), .A3(n10100), .ZN(n9792) );
  AND2_X1 U12504 ( .A1(n10125), .A2(n14202), .ZN(n9793) );
  AND2_X1 U12505 ( .A1(n10197), .A2(n12211), .ZN(n9794) );
  AND2_X1 U12506 ( .A1(n10873), .A2(n10872), .ZN(n10878) );
  AND2_X1 U12507 ( .A1(n21407), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9795) );
  AND2_X1 U12508 ( .A1(n15044), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9796) );
  INV_X1 U12509 ( .A(n15722), .ZN(n9999) );
  NOR2_X1 U12510 ( .A1(n10631), .A2(n9985), .ZN(n9797) );
  NAND2_X1 U12511 ( .A1(n15609), .A2(n10095), .ZN(n11597) );
  OAI21_X1 U12512 ( .B1(n9998), .B2(n9997), .A(n15699), .ZN(n9995) );
  NAND2_X1 U12513 ( .A1(n13066), .A2(n13067), .ZN(n15777) );
  NAND2_X1 U12514 ( .A1(n15612), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15613) );
  OR3_X1 U12515 ( .A1(n11623), .A2(n11622), .A3(n11621), .ZN(P3_U2640) );
  NAND2_X1 U12516 ( .A1(n14854), .A2(n10169), .ZN(n14840) );
  OR2_X1 U12517 ( .A1(n15151), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9799) );
  AND2_X1 U12518 ( .A1(n11680), .A2(n11679), .ZN(n9800) );
  AND2_X1 U12519 ( .A1(n10084), .A2(n18359), .ZN(n9801) );
  INV_X1 U12520 ( .A(n9750), .ZN(n19629) );
  AND2_X1 U12522 ( .A1(n9947), .A2(n9945), .ZN(n9802) );
  AND2_X1 U12523 ( .A1(n15012), .A2(n15035), .ZN(n9803) );
  AND2_X1 U12524 ( .A1(n10050), .A2(n10049), .ZN(n9804) );
  NAND2_X1 U12525 ( .A1(n11426), .A2(n9936), .ZN(n9805) );
  INV_X1 U12526 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10087) );
  BUF_X1 U12527 ( .A(n9737), .Z(n12742) );
  NOR2_X1 U12528 ( .A1(n10244), .A2(n10243), .ZN(n14114) );
  NAND2_X1 U12529 ( .A1(n15460), .A2(n15462), .ZN(n15455) );
  NOR2_X1 U12530 ( .A1(n13032), .A2(n19318), .ZN(n13028) );
  INV_X1 U12531 ( .A(n14284), .ZN(n9897) );
  NOR2_X1 U12532 ( .A1(n13034), .A2(n15737), .ZN(n13035) );
  AND2_X1 U12533 ( .A1(n13028), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13029) );
  NOR2_X1 U12534 ( .A1(n13036), .A2(n16637), .ZN(n13037) );
  NOR2_X1 U12535 ( .A1(n13034), .A2(n10048), .ZN(n13033) );
  AND2_X1 U12536 ( .A1(n15485), .A2(n9769), .ZN(n9806) );
  AND2_X1 U12537 ( .A1(n9768), .A2(n13163), .ZN(n9807) );
  AND2_X1 U12538 ( .A1(n13029), .A2(n9766), .ZN(n9808) );
  AND2_X1 U12539 ( .A1(n14255), .A2(n14256), .ZN(n14254) );
  NAND2_X1 U12540 ( .A1(n13029), .A2(n9762), .ZN(n13025) );
  XNOR2_X1 U12541 ( .A(n14034), .B(n14286), .ZN(n13630) );
  INV_X1 U12542 ( .A(n11447), .ZN(n10037) );
  AND2_X1 U12543 ( .A1(n11961), .A2(n12306), .ZN(n9809) );
  AND2_X1 U12544 ( .A1(n9976), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9810) );
  AND2_X1 U12545 ( .A1(n10031), .A2(n11333), .ZN(n9811) );
  AND2_X1 U12546 ( .A1(n16659), .A2(n9765), .ZN(n9812) );
  XNOR2_X1 U12547 ( .A(n16010), .B(n13102), .ZN(n13627) );
  OR2_X1 U12548 ( .A1(n12204), .A2(n16458), .ZN(n9813) );
  NOR2_X1 U12549 ( .A1(n17994), .A2(n17995), .ZN(n10281) );
  OAI21_X1 U12550 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n16971) );
  INV_X1 U12551 ( .A(n15640), .ZN(n10158) );
  NOR2_X1 U12552 ( .A1(n16693), .A2(n10114), .ZN(n9814) );
  NOR2_X1 U12553 ( .A1(n16629), .A2(n16625), .ZN(n9815) );
  NAND2_X1 U12554 ( .A1(n13121), .A2(n9768), .ZN(n10238) );
  AND2_X1 U12555 ( .A1(n13118), .A2(n13991), .ZN(n9816) );
  AOI21_X1 U12556 ( .B1(n17990), .B2(n18251), .A(n11741), .ZN(n11742) );
  INV_X1 U12557 ( .A(n11742), .ZN(n10062) );
  AND2_X1 U12558 ( .A1(n10105), .A2(n15979), .ZN(n9817) );
  AND2_X1 U12559 ( .A1(n11455), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11517) );
  NAND2_X1 U12560 ( .A1(n14242), .A2(n14239), .ZN(n9818) );
  AND2_X1 U12561 ( .A1(n15572), .A2(n15561), .ZN(n9819) );
  OR2_X1 U12562 ( .A1(n12223), .A2(n16329), .ZN(n9820) );
  INV_X1 U12563 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15737) );
  OR2_X1 U12564 ( .A1(n17583), .A2(n17711), .ZN(n9821) );
  NOR2_X1 U12565 ( .A1(n16936), .A2(n9980), .ZN(n9822) );
  AND2_X1 U12566 ( .A1(n10028), .A2(n11481), .ZN(n9823) );
  NOR2_X1 U12567 ( .A1(n15429), .A2(n15430), .ZN(n9824) );
  OR2_X1 U12568 ( .A1(n14885), .A2(n10018), .ZN(n9825) );
  AND2_X1 U12569 ( .A1(n10169), .A2(n10167), .ZN(n9826) );
  AND2_X1 U12570 ( .A1(n10113), .A2(n10112), .ZN(n9827) );
  AND2_X1 U12571 ( .A1(n9807), .A2(n15473), .ZN(n9828) );
  AND2_X1 U12572 ( .A1(n9763), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9829) );
  AND2_X1 U12573 ( .A1(n9811), .A2(n11494), .ZN(n9830) );
  INV_X1 U12574 ( .A(n12169), .ZN(n10190) );
  NAND2_X1 U12575 ( .A1(n12105), .A2(n12104), .ZN(n12169) );
  AND2_X1 U12576 ( .A1(n10185), .A2(n10186), .ZN(n9831) );
  AOI21_X1 U12577 ( .B1(n16963), .B2(n9958), .A(n9954), .ZN(n9951) );
  AND2_X1 U12578 ( .A1(n10783), .A2(n10782), .ZN(n11422) );
  INV_X1 U12579 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n9961) );
  NOR2_X1 U12580 ( .A1(n11011), .A2(n10107), .ZN(n10106) );
  INV_X1 U12581 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U12582 ( .A1(n10243), .A2(n10241), .ZN(n14201) );
  OR3_X1 U12583 ( .A1(n13340), .A2(n13339), .A3(n15432), .ZN(n9832) );
  NOR3_X1 U12584 ( .A1(n13017), .A2(n12999), .A3(n13018), .ZN(n13013) );
  AND2_X1 U12585 ( .A1(n10011), .A2(n9785), .ZN(n9833) );
  NAND2_X1 U12586 ( .A1(n10103), .A2(n10106), .ZN(n14329) );
  NAND2_X1 U12587 ( .A1(n10053), .A2(n10052), .ZN(n9834) );
  NOR2_X1 U12588 ( .A1(n13024), .A2(n13494), .ZN(n13022) );
  NOR2_X1 U12589 ( .A1(n13023), .A2(n13055), .ZN(n13054) );
  NAND2_X1 U12590 ( .A1(n14120), .A2(n10125), .ZN(n9835) );
  INV_X1 U12591 ( .A(n15415), .ZN(n10130) );
  NAND2_X1 U12592 ( .A1(n13969), .A2(n12505), .ZN(n13971) );
  AND2_X1 U12593 ( .A1(n10116), .A2(n13497), .ZN(n9836) );
  AND2_X1 U12594 ( .A1(n13069), .A2(n10951), .ZN(n9837) );
  OR2_X1 U12595 ( .A1(n16514), .A2(n16522), .ZN(n9838) );
  AND2_X1 U12596 ( .A1(n10073), .A2(n10071), .ZN(n9839) );
  INV_X1 U12597 ( .A(n10022), .ZN(n14902) );
  AND2_X1 U12598 ( .A1(n9772), .A2(n10115), .ZN(n9840) );
  INV_X1 U12599 ( .A(n9914), .ZN(n13920) );
  INV_X1 U12600 ( .A(n20507), .ZN(n16424) );
  AND2_X1 U12601 ( .A1(n12461), .A2(n12325), .ZN(n20507) );
  INV_X1 U12602 ( .A(n9971), .ZN(n9970) );
  OAI21_X1 U12603 ( .B1(n9965), .B2(n9972), .A(n17895), .ZN(n9971) );
  OR2_X1 U12604 ( .A1(n13017), .A2(n13018), .ZN(n9841) );
  NOR2_X1 U12605 ( .A1(n17054), .A2(n9965), .ZN(n9842) );
  XOR2_X2 U12606 ( .A(n10288), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n9968) );
  INV_X1 U12607 ( .A(n9965), .ZN(n9958) );
  AND2_X2 U12608 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13638) );
  AND2_X1 U12609 ( .A1(n17866), .A2(n9959), .ZN(n9844) );
  INV_X1 U12610 ( .A(n17970), .ZN(n9966) );
  NAND2_X1 U12611 ( .A1(n11203), .A2(n11202), .ZN(n9845) );
  XNOR2_X1 U12612 ( .A(n13000), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13011) );
  NAND2_X1 U12613 ( .A1(n11732), .A2(n11731), .ZN(n9846) );
  NAND2_X1 U12614 ( .A1(n11455), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n9847) );
  INV_X1 U12615 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12616 ( .A1(n10281), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17955) );
  AND2_X1 U12617 ( .A1(n9802), .A2(n9943), .ZN(n17112) );
  AND2_X1 U12618 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17185) );
  NOR2_X1 U12619 ( .A1(n18118), .A2(n17166), .ZN(n18065) );
  NOR2_X1 U12620 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9848) );
  INV_X1 U12621 ( .A(n9934), .ZN(n9930) );
  NOR2_X1 U12622 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n9934) );
  AND2_X1 U12623 ( .A1(n9942), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9849) );
  INV_X1 U12624 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10033) );
  INV_X1 U12625 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9946) );
  INV_X1 U12626 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17222) );
  INV_X1 U12627 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9985) );
  INV_X1 U12628 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9933) );
  OAI22_X1 U12629 ( .A1(n19702), .A2(n14021), .B1(n13916), .B2(n14022), .ZN(
        n9850) );
  NOR2_X2 U12630 ( .A1(n18578), .A2(n18557), .ZN(n18982) );
  OR2_X1 U12631 ( .A1(n18657), .A2(n18798), .ZN(n18557) );
  NOR2_X2 U12632 ( .A1(n18572), .A2(n18557), .ZN(n18976) );
  NOR3_X2 U12633 ( .A1(n19072), .A2(n18848), .A3(n18800), .ZN(n18818) );
  NOR3_X2 U12634 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19072), .A3(
        n18594), .ZN(n18610) );
  NOR3_X2 U12635 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19072), .A3(
        n18800), .ZN(n18791) );
  OAI22_X2 U12636 ( .A1(n16818), .A2(n14021), .B1(n13932), .B2(n14022), .ZN(
        n20940) );
  INV_X1 U12637 ( .A(n20920), .ZN(n9851) );
  INV_X1 U12638 ( .A(n9851), .ZN(n9852) );
  INV_X1 U12639 ( .A(n20933), .ZN(n9853) );
  INV_X1 U12640 ( .A(n9853), .ZN(n9854) );
  INV_X1 U12641 ( .A(n20971), .ZN(n9855) );
  INV_X1 U12642 ( .A(n9855), .ZN(n9856) );
  INV_X1 U12643 ( .A(n20926), .ZN(n9857) );
  INV_X1 U12644 ( .A(n9857), .ZN(n9858) );
  INV_X1 U12645 ( .A(n20961), .ZN(n9859) );
  INV_X1 U12646 ( .A(n9859), .ZN(n9860) );
  NOR3_X2 U12647 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19072), .A3(
        n18703), .ZN(n18698) );
  OAI22_X2 U12648 ( .A1(n16814), .A2(n14021), .B1(n14015), .B2(n14022), .ZN(
        n20954) );
  OAI22_X2 U12649 ( .A1(n16816), .A2(n14021), .B1(n13927), .B2(n14022), .ZN(
        n20947) );
  NOR2_X2 U12650 ( .A1(n19682), .A2(n19695), .ZN(n20136) );
  INV_X1 U12651 ( .A(n9863), .ZN(n17588) );
  INV_X1 U12652 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n9862) );
  INV_X2 U12653 ( .A(n14469), .ZN(n10308) );
  INV_X1 U12654 ( .A(n17781), .ZN(n9868) );
  NAND3_X1 U12655 ( .A1(n9869), .A2(n10748), .A3(n9909), .ZN(n10833) );
  NAND2_X2 U12656 ( .A1(n9781), .A2(n10636), .ZN(n9869) );
  AND2_X4 U12657 ( .A1(n13821), .A2(n13848), .ZN(n10661) );
  AND2_X2 U12658 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13821) );
  NAND2_X1 U12659 ( .A1(n9874), .A2(n9873), .ZN(n15766) );
  NAND3_X1 U12660 ( .A1(n14321), .A2(n14322), .A3(n19615), .ZN(n9873) );
  NAND2_X1 U12661 ( .A1(n9876), .A2(n11419), .ZN(n19614) );
  INV_X1 U12662 ( .A(n19615), .ZN(n9877) );
  OAI21_X2 U12663 ( .B1(n11441), .B2(n9880), .A(n9878), .ZN(n15664) );
  NAND2_X1 U12664 ( .A1(n9883), .A2(n16314), .ZN(n12219) );
  XNOR2_X1 U12665 ( .A(n16315), .B(n9883), .ZN(n16371) );
  OAI21_X1 U12666 ( .B1(n12063), .B2(n9884), .A(n14034), .ZN(n13678) );
  NAND2_X1 U12667 ( .A1(n15080), .A2(n9932), .ZN(n9928) );
  NAND2_X1 U12668 ( .A1(n15080), .A2(n12225), .ZN(n9931) );
  OAI21_X1 U12669 ( .B1(n15080), .B2(n12232), .A(n9932), .ZN(n12227) );
  NOR2_X4 U12670 ( .A1(n15096), .A2(n21077), .ZN(n15080) );
  NAND3_X1 U12671 ( .A1(n9897), .A2(n10189), .A3(n9896), .ZN(n12186) );
  AND2_X2 U12672 ( .A1(n10566), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10587) );
  AND3_X4 U12673 ( .A1(n9900), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10656) );
  NAND3_X1 U12674 ( .A1(n9903), .A2(n9901), .A3(n9805), .ZN(n15965) );
  NAND3_X1 U12675 ( .A1(n9902), .A2(n15762), .A3(n15760), .ZN(n9901) );
  NAND3_X1 U12676 ( .A1(n9750), .A2(n9904), .A3(n9988), .ZN(n9991) );
  NAND2_X1 U12677 ( .A1(n12480), .A2(n20507), .ZN(n10196) );
  XNOR2_X2 U12678 ( .A(n9910), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12480) );
  OAI211_X2 U12679 ( .C1(n15004), .C2(n12234), .A(n9911), .B(n12233), .ZN(
        n9910) );
  NAND2_X1 U12680 ( .A1(n12435), .A2(n12337), .ZN(n9912) );
  AND2_X2 U12681 ( .A1(n11967), .A2(n14661), .ZN(n12435) );
  NAND2_X1 U12682 ( .A1(n12056), .A2(n20548), .ZN(n14172) );
  NAND2_X2 U12683 ( .A1(n9928), .A2(n9924), .ZN(n15033) );
  AND3_X2 U12684 ( .A1(n11961), .A2(n12306), .A3(n14157), .ZN(n12318) );
  NOR2_X2 U12685 ( .A1(n16347), .A2(n12212), .ZN(n15112) );
  NOR2_X1 U12686 ( .A1(n16963), .A2(n9954), .ZN(n9950) );
  INV_X1 U12687 ( .A(n16992), .ZN(n9969) );
  NAND3_X1 U12688 ( .A1(n10530), .A2(n10551), .A3(n9728), .ZN(n10537) );
  OAI211_X1 U12689 ( .C1(n20010), .C2(n13142), .A(n9990), .B(n9989), .ZN(
        n10632) );
  NAND2_X1 U12690 ( .A1(n15667), .A2(n10000), .ZN(n16124) );
  AND2_X2 U12691 ( .A1(n13644), .A2(n13638), .ZN(n11934) );
  AND2_X2 U12692 ( .A1(n12237), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13644) );
  NAND3_X1 U12693 ( .A1(n12337), .A2(n14055), .A3(n14155), .ZN(n10016) );
  NOR2_X2 U12694 ( .A1(n11411), .A2(n11412), .ZN(n11410) );
  NAND2_X1 U12695 ( .A1(n11477), .A2(n9823), .ZN(n11510) );
  NAND2_X1 U12696 ( .A1(n11518), .A2(n9830), .ZN(n11539) );
  AND2_X1 U12697 ( .A1(n11518), .A2(n11483), .ZN(n11491) );
  AND2_X1 U12698 ( .A1(n11538), .A2(n9764), .ZN(n11556) );
  NAND2_X1 U12699 ( .A1(n11538), .A2(n9770), .ZN(n11558) );
  NAND2_X1 U12700 ( .A1(n11538), .A2(n10034), .ZN(n11548) );
  NAND2_X1 U12701 ( .A1(n11538), .A2(n11537), .ZN(n11547) );
  XNOR2_X1 U12702 ( .A(n11574), .B(n9847), .ZN(n11577) );
  NAND3_X1 U12703 ( .A1(n10038), .A2(n14124), .A3(n10037), .ZN(n10036) );
  NAND2_X1 U12704 ( .A1(n13029), .A2(n9771), .ZN(n13024) );
  AOI21_X1 U12705 ( .B1(n13492), .B2(n15654), .A(n19410), .ZN(n10044) );
  INV_X1 U12706 ( .A(n10050), .ZN(n16520) );
  INV_X1 U12707 ( .A(n19410), .ZN(n10049) );
  NAND3_X1 U12708 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U12709 ( .A1(n15347), .A2(n19410), .ZN(n16500) );
  AOI21_X1 U12710 ( .B1(n15347), .B2(n15604), .A(n19410), .ZN(n10061) );
  NAND2_X1 U12711 ( .A1(n19410), .A2(n10059), .ZN(n10057) );
  INV_X1 U12712 ( .A(n15347), .ZN(n10060) );
  INV_X1 U12713 ( .A(n10063), .ZN(n17889) );
  NAND3_X1 U12714 ( .A1(n17944), .A2(n10062), .A3(n18250), .ZN(n10063) );
  NAND2_X2 U12715 ( .A1(n17985), .A2(n18107), .ZN(n17944) );
  NAND2_X1 U12716 ( .A1(n17944), .A2(n10062), .ZN(n17890) );
  NAND2_X1 U12717 ( .A1(n10063), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10066) );
  NAND2_X1 U12718 ( .A1(n17944), .A2(n17937), .ZN(n10065) );
  OAI21_X2 U12719 ( .B1(n18007), .B2(n9846), .A(n18107), .ZN(n11739) );
  NOR2_X1 U12720 ( .A1(n16101), .A2(n16190), .ZN(n17856) );
  NAND2_X1 U12721 ( .A1(n18138), .A2(n10069), .ZN(n10068) );
  NAND2_X1 U12722 ( .A1(n10073), .A2(n10074), .ZN(n18128) );
  NOR2_X1 U12723 ( .A1(n18127), .A2(n10072), .ZN(n10071) );
  NAND2_X1 U12724 ( .A1(n18138), .A2(n18139), .ZN(n18137) );
  INV_X1 U12725 ( .A(n18139), .ZN(n10076) );
  INV_X1 U12726 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10077) );
  XNOR2_X1 U12727 ( .A(n17715), .B(n17709), .ZN(n11715) );
  NAND2_X1 U12728 ( .A1(n15965), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10877) );
  NAND2_X2 U12729 ( .A1(n10750), .A2(n10749), .ZN(n10092) );
  NAND2_X1 U12730 ( .A1(n10092), .A2(n10784), .ZN(n14325) );
  AND2_X1 U12731 ( .A1(n10101), .A2(n15776), .ZN(n10100) );
  INV_X1 U12732 ( .A(n14558), .ZN(n10103) );
  NAND2_X1 U12733 ( .A1(n10103), .A2(n9761), .ZN(n15978) );
  NAND2_X1 U12734 ( .A1(n15523), .A2(n15522), .ZN(n15340) );
  NAND3_X1 U12735 ( .A1(n10140), .A2(n10951), .A3(n13069), .ZN(n10567) );
  NAND2_X1 U12736 ( .A1(n10567), .A2(n9736), .ZN(n10117) );
  NAND4_X1 U12737 ( .A1(n10120), .A2(n10519), .A3(n10521), .A4(n10520), .ZN(
        n10118) );
  NAND4_X1 U12738 ( .A1(n10121), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10119) );
  NAND2_X1 U12739 ( .A1(n15485), .A2(n10122), .ZN(n15445) );
  NOR3_X2 U12740 ( .A1(n15447), .A2(n10132), .A3(n10129), .ZN(n10134) );
  INV_X1 U12741 ( .A(n10134), .ZN(n15416) );
  NAND2_X1 U12742 ( .A1(n15336), .A2(n10137), .ZN(n15325) );
  NAND2_X1 U12743 ( .A1(n15336), .A2(n10135), .ZN(n10139) );
  AND2_X2 U12744 ( .A1(n15336), .A2(n11599), .ZN(n15320) );
  INV_X1 U12745 ( .A(n11375), .ZN(n10138) );
  NAND4_X1 U12746 ( .A1(n10554), .A2(n11247), .A3(n11241), .A4(n9756), .ZN(
        n10140) );
  NAND2_X1 U12747 ( .A1(n15595), .A2(n10141), .ZN(n10145) );
  INV_X1 U12748 ( .A(n15593), .ZN(n10142) );
  NAND2_X1 U12749 ( .A1(n11590), .A2(n11572), .ZN(n10143) );
  NAND2_X1 U12750 ( .A1(n10145), .A2(n10149), .ZN(n11586) );
  NAND2_X1 U12751 ( .A1(n11572), .A2(n11573), .ZN(n10148) );
  NAND2_X1 U12752 ( .A1(n10152), .A2(n11536), .ZN(n15652) );
  NAND2_X1 U12753 ( .A1(n15664), .A2(n11524), .ZN(n10152) );
  OAI21_X1 U12754 ( .B1(n15664), .B2(n10155), .A(n10153), .ZN(n11542) );
  INV_X1 U12756 ( .A(n11536), .ZN(n10155) );
  NAND2_X1 U12757 ( .A1(n15847), .A2(n11545), .ZN(n15643) );
  INV_X1 U12758 ( .A(n11545), .ZN(n10160) );
  AND2_X2 U12759 ( .A1(n14854), .A2(n9826), .ZN(n14797) );
  NAND2_X1 U12760 ( .A1(n14605), .A2(n10172), .ZN(n14887) );
  NAND2_X1 U12761 ( .A1(n10179), .A2(n12490), .ZN(n10177) );
  NAND2_X1 U12762 ( .A1(n10179), .A2(n10178), .ZN(n12489) );
  INV_X1 U12763 ( .A(n12076), .ZN(n12153) );
  AND3_X2 U12764 ( .A1(n14255), .A2(n10180), .A3(n14256), .ZN(n12596) );
  NAND3_X1 U12765 ( .A1(n14255), .A2(n14256), .A3(n10182), .ZN(n10184) );
  NAND3_X1 U12766 ( .A1(n14255), .A2(n14256), .A3(n14393), .ZN(n14392) );
  INV_X1 U12767 ( .A(n10184), .ZN(n14420) );
  NAND2_X1 U12768 ( .A1(n14756), .A2(n10186), .ZN(n14723) );
  AND2_X1 U12769 ( .A1(n14756), .A2(n10187), .ZN(n14732) );
  NAND2_X1 U12770 ( .A1(n14756), .A2(n14757), .ZN(n14745) );
  INV_X1 U12771 ( .A(n12160), .ZN(n10189) );
  NAND2_X1 U12772 ( .A1(n13999), .A2(n14001), .ZN(n14000) );
  XNOR2_X1 U12773 ( .A(n12157), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13999) );
  NAND2_X1 U12774 ( .A1(n9803), .A2(n12229), .ZN(n15024) );
  NAND2_X1 U12775 ( .A1(n10193), .A2(n14016), .ZN(n13632) );
  INV_X1 U12776 ( .A(n13645), .ZN(n10193) );
  NAND2_X1 U12777 ( .A1(n10195), .A2(n10194), .ZN(n13645) );
  NAND2_X1 U12778 ( .A1(n10196), .A2(n12478), .ZN(P1_U3000) );
  INV_X1 U12779 ( .A(n9729), .ZN(n13917) );
  NAND2_X2 U12780 ( .A1(n13611), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12149) );
  NAND2_X1 U12781 ( .A1(n14584), .A2(n10199), .ZN(n10198) );
  OAI21_X2 U12782 ( .B1(n15112), .B2(n10210), .A(n10207), .ZN(n15096) );
  NAND2_X1 U12783 ( .A1(n10220), .A2(n15419), .ZN(n10215) );
  INV_X1 U12784 ( .A(n13383), .ZN(n10220) );
  NAND2_X1 U12785 ( .A1(n13406), .A2(n10223), .ZN(n10222) );
  NAND3_X1 U12786 ( .A1(n10228), .A2(n13441), .A3(n10222), .ZN(n13460) );
  INV_X1 U12787 ( .A(n13407), .ZN(n10227) );
  NAND2_X1 U12788 ( .A1(n15402), .A2(n15401), .ZN(n15403) );
  NAND2_X1 U12789 ( .A1(n10230), .A2(n10229), .ZN(n15402) );
  INV_X1 U12790 ( .A(n13318), .ZN(n10232) );
  NAND2_X1 U12791 ( .A1(n10232), .A2(n9832), .ZN(n10234) );
  AND2_X2 U12792 ( .A1(n15460), .A2(n10235), .ZN(n13317) );
  NAND2_X1 U12793 ( .A1(n10266), .A2(n13987), .ZN(n13986) );
  INV_X1 U12794 ( .A(n12186), .ZN(n12133) );
  OAI211_X1 U12795 ( .C1(n21059), .C2(n12156), .A(n12155), .B(n12154), .ZN(
        n14001) );
  OAI21_X1 U12796 ( .B1(n21059), .B2(n12142), .A(n12154), .ZN(n12139) );
  NAND2_X1 U12797 ( .A1(n10835), .A2(n10834), .ZN(n10879) );
  AND2_X2 U12798 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11846) );
  INV_X1 U12799 ( .A(n12306), .ZN(n11984) );
  NAND2_X1 U12800 ( .A1(n11983), .A2(n14661), .ZN(n11966) );
  INV_X1 U12801 ( .A(n11966), .ZN(n11897) );
  OR3_X2 U12802 ( .A1(n10631), .A2(n10630), .A3(n15396), .ZN(n19842) );
  NAND2_X1 U12803 ( .A1(n11897), .A2(n11896), .ZN(n11969) );
  NAND2_X1 U12804 ( .A1(n12523), .A2(n12522), .ZN(n14006) );
  OR2_X1 U12805 ( .A1(n13692), .A2(n13691), .ZN(n13694) );
  AND2_X1 U12806 ( .A1(n20516), .A2(n20515), .ZN(n20623) );
  OAI21_X2 U12807 ( .B1(n20515), .B2(n12671), .A(n12514), .ZN(n13972) );
  INV_X1 U12808 ( .A(n11957), .ZN(n11983) );
  INV_X1 U12809 ( .A(n14008), .ZN(n12523) );
  XNOR2_X1 U12810 ( .A(n12198), .B(n12197), .ZN(n12541) );
  CLKBUF_X1 U12811 ( .A(n14595), .Z(n14598) );
  AND2_X2 U12812 ( .A1(n13894), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10266) );
  NAND3_X1 U12813 ( .A1(n10488), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10562), 
        .ZN(n13376) );
  NAND2_X1 U12814 ( .A1(n14710), .A2(n14636), .ZN(n14639) );
  AOI22_X1 U12815 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10431) );
  INV_X1 U12816 ( .A(n11426), .ZN(n10832) );
  NAND2_X1 U12817 ( .A1(n10597), .A2(n10598), .ZN(n10601) );
  INV_X1 U12818 ( .A(n14156), .ZN(n11972) );
  AND2_X1 U12819 ( .A1(n14661), .A2(n14156), .ZN(n12256) );
  NOR2_X1 U12820 ( .A1(n10301), .A2(n10300), .ZN(n11624) );
  NOR2_X1 U12821 ( .A1(n10296), .A2(n10301), .ZN(n11661) );
  BUF_X4 U12822 ( .A(n10342), .Z(n17505) );
  AND2_X1 U12823 ( .A1(n13086), .A2(n13085), .ZN(n10246) );
  AND2_X1 U12824 ( .A1(n11587), .A2(n20308), .ZN(n19663) );
  INV_X1 U12825 ( .A(n20465), .ZN(n13796) );
  OR2_X2 U12826 ( .A1(n16166), .A2(n13953), .ZN(n20321) );
  INV_X1 U12827 ( .A(n20321), .ZN(n12479) );
  NAND2_X1 U12828 ( .A1(n13977), .A2(n13976), .ZN(n14905) );
  INV_X1 U12829 ( .A(n14905), .ZN(n13978) );
  OR2_X1 U12830 ( .A1(n16489), .A2(n16143), .ZN(n10247) );
  INV_X1 U12831 ( .A(n15467), .ZN(n15472) );
  INV_X1 U12832 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n13514) );
  INV_X1 U12833 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11569) );
  INV_X1 U12834 ( .A(n19450), .ZN(n19416) );
  INV_X1 U12835 ( .A(n15812), .ZN(n10908) );
  INV_X1 U12836 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12159) );
  AND2_X1 U12837 ( .A1(n12230), .A2(n15172), .ZN(n10248) );
  OR2_X1 U12838 ( .A1(n14582), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10249) );
  AND2_X1 U12839 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10250) );
  AND2_X1 U12840 ( .A1(n11047), .A2(n11046), .ZN(n13985) );
  AND3_X1 U12841 ( .A1(n10456), .A2(n10455), .A3(n10429), .ZN(n10251) );
  INV_X1 U12842 ( .A(n10661), .ZN(n10662) );
  NOR2_X1 U12843 ( .A1(n13012), .A2(n13014), .ZN(n10253) );
  AND3_X1 U12844 ( .A1(n10467), .A2(n10466), .A3(n10429), .ZN(n10254) );
  NAND2_X2 U12845 ( .A1(n17659), .A2(n16207), .ZN(n17719) );
  AND3_X1 U12846 ( .A1(n10444), .A2(n10443), .A3(n10429), .ZN(n10255) );
  OR2_X1 U12847 ( .A1(n17881), .A2(n18107), .ZN(n10256) );
  OR2_X1 U12848 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n11614), .ZN(n10257) );
  CLKBUF_X1 U12849 ( .A(n16903), .Z(n16904) );
  INV_X1 U12850 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12168) );
  INV_X1 U12851 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n21240) );
  INV_X1 U12852 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16622) );
  XOR2_X1 U12853 ( .A(n11585), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n10258) );
  AND4_X1 U12854 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(
        n10259) );
  NOR2_X1 U12855 ( .A1(n16749), .A2(n16744), .ZN(n10260) );
  AND2_X1 U12856 ( .A1(n18030), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10261) );
  INV_X1 U12857 ( .A(n10878), .ZN(n10874) );
  NOR2_X1 U12858 ( .A1(n20741), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10262) );
  NAND2_X1 U12859 ( .A1(n13966), .A2(n13965), .ZN(n13968) );
  INV_X1 U12860 ( .A(n13968), .ZN(n12504) );
  INV_X1 U12861 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21171) );
  INV_X1 U12862 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20582) );
  NOR2_X1 U12863 ( .A1(n19080), .A2(n18183), .ZN(n17980) );
  AND2_X1 U12864 ( .A1(n13380), .A2(n13399), .ZN(n10265) );
  INV_X1 U12865 ( .A(n10570), .ZN(n10571) );
  INV_X1 U12866 ( .A(n11889), .ZN(n13648) );
  AND3_X1 U12867 ( .A1(n11853), .A2(n11852), .A3(n11851), .ZN(n10267) );
  AND4_X1 U12868 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n10268) );
  AND4_X1 U12869 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n10269) );
  AND4_X1 U12870 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n10270) );
  INV_X1 U12871 ( .A(n11939), .ZN(n12870) );
  NAND2_X1 U12872 ( .A1(n11909), .A2(n14637), .ZN(n10271) );
  AND2_X1 U12873 ( .A1(n12271), .A2(n12258), .ZN(n12278) );
  OR2_X1 U12874 ( .A1(n12271), .A2(n12270), .ZN(n12289) );
  NAND2_X1 U12875 ( .A1(n11957), .A2(n14661), .ZN(n11882) );
  NAND2_X1 U12876 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10474) );
  INV_X1 U12877 ( .A(n12952), .ZN(n12868) );
  NAND2_X1 U12878 ( .A1(n12302), .A2(n11882), .ZN(n11883) );
  NOR2_X2 U12879 ( .A1(n13069), .A2(n13376), .ZN(n10570) );
  AOI22_X1 U12880 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10656), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U12881 ( .A1(n10536), .A2(n10535), .ZN(n11244) );
  AND2_X1 U12882 ( .A1(n20905), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12262) );
  INV_X1 U12883 ( .A(n14978), .ZN(n12673) );
  OR2_X1 U12884 ( .A1(n12283), .A2(n12106), .ZN(n12119) );
  NAND2_X1 U12885 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12224) );
  INV_X1 U12886 ( .A(n12187), .ZN(n12132) );
  NAND2_X1 U12887 ( .A1(n11969), .A2(n12138), .ZN(n11910) );
  NAND2_X1 U12888 ( .A1(n13954), .A2(n14157), .ZN(n12064) );
  INV_X1 U12889 ( .A(n10965), .ZN(n10658) );
  AND2_X1 U12890 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  OR3_X1 U12891 ( .A1(n10857), .A2(n10856), .A3(n10855), .ZN(n10864) );
  NAND2_X1 U12892 ( .A1(n11259), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10594) );
  NAND2_X1 U12893 ( .A1(n10991), .A2(n10544), .ZN(n10545) );
  OR2_X1 U12894 ( .A1(n11762), .A2(n11757), .ZN(n10396) );
  NOR2_X1 U12895 ( .A1(n12245), .A2(n12244), .ZN(n12290) );
  INV_X1 U12896 ( .A(n12826), .ZN(n12825) );
  NOR2_X1 U12897 ( .A1(n12706), .A2(n16253), .ZN(n12707) );
  NAND2_X1 U12898 ( .A1(n12119), .A2(n12118), .ZN(n12177) );
  OR2_X1 U12899 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20514), .ZN(
        n12244) );
  AND2_X1 U12900 ( .A1(n12150), .A2(n13612), .ZN(n12151) );
  AND2_X1 U12901 ( .A1(n12131), .A2(n12130), .ZN(n12187) );
  NAND2_X1 U12902 ( .A1(n12302), .A2(n12138), .ZN(n11965) );
  OR2_X1 U12904 ( .A1(n10933), .A2(n10931), .ZN(n10929) );
  NAND2_X1 U12905 ( .A1(n13088), .A2(n13103), .ZN(n13092) );
  AND2_X1 U12906 ( .A1(n13382), .A2(n10265), .ZN(n13383) );
  AND2_X1 U12907 ( .A1(n13315), .A2(n13314), .ZN(n13333) );
  INV_X1 U12908 ( .A(n13267), .ZN(n13818) );
  NAND2_X1 U12909 ( .A1(n13113), .A2(n10490), .ZN(n10491) );
  INV_X1 U12910 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11568) );
  AND2_X1 U12911 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  AND3_X1 U12912 ( .A1(n11241), .A2(n10533), .A3(n11245), .ZN(n10534) );
  NAND2_X1 U12913 ( .A1(n12825), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12845) );
  AND2_X1 U12914 ( .A1(n12372), .A2(n12371), .ZN(n14901) );
  OR2_X1 U12915 ( .A1(n12210), .A2(n12358), .ZN(n12211) );
  INV_X1 U12916 ( .A(n12150), .ZN(n12148) );
  NAND2_X1 U12917 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11946) );
  NAND2_X1 U12918 ( .A1(n12024), .A2(n12023), .ZN(n12136) );
  INV_X1 U12919 ( .A(n15469), .ZN(n13200) );
  INV_X1 U12920 ( .A(n15411), .ZN(n13405) );
  INV_X1 U12921 ( .A(n11595), .ZN(n11572) );
  INV_X1 U12922 ( .A(n11006), .ZN(n11218) );
  INV_X1 U12923 ( .A(n19539), .ZN(n10941) );
  NOR2_X1 U12924 ( .A1(n10543), .A2(n10493), .ZN(n10529) );
  NAND2_X1 U12925 ( .A1(n18109), .A2(n18341), .ZN(n11734) );
  INV_X1 U12926 ( .A(n18563), .ZN(n10391) );
  AOI211_X1 U12927 ( .C1(n9718), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n10317), .B(n10316), .ZN(n10318) );
  INV_X1 U12928 ( .A(n14165), .ZN(n14175) );
  AND2_X1 U12929 ( .A1(n12362), .A2(n12361), .ZN(n14409) );
  OR2_X1 U12930 ( .A1(n12985), .A2(n21215), .ZN(n12987) );
  OR2_X1 U12931 ( .A1(n12887), .A2(n12886), .ZN(n12921) );
  NAND2_X1 U12932 ( .A1(n12562), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12577) );
  NAND2_X1 U12933 ( .A1(n12287), .A2(n12257), .ZN(n12300) );
  AND2_X1 U12934 ( .A1(n12381), .A2(n12380), .ZN(n16270) );
  OR2_X1 U12936 ( .A1(n12103), .A2(n12102), .ZN(n12179) );
  INV_X1 U12937 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20653) );
  INV_X1 U12938 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20740) );
  XNOR2_X1 U12939 ( .A(n12490), .B(n12489), .ZN(n13915) );
  INV_X1 U12940 ( .A(n20304), .ZN(n10964) );
  AND2_X1 U12941 ( .A1(n11459), .A2(n11458), .ZN(n11470) );
  OR2_X1 U12942 ( .A1(n13399), .A2(n13398), .ZN(n15406) );
  INV_X1 U12943 ( .A(n14324), .ZN(n10758) );
  INV_X1 U12944 ( .A(n11590), .ZN(n11591) );
  INV_X1 U12945 ( .A(n11663), .ZN(n11668) );
  AND2_X1 U12946 ( .A1(n18109), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16100) );
  NAND2_X1 U12947 ( .A1(n11735), .A2(n11734), .ZN(n11736) );
  NOR2_X1 U12948 ( .A1(n18121), .A2(n11730), .ZN(n11733) );
  AND2_X1 U12949 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11722), .ZN(
        n11723) );
  INV_X1 U12950 ( .A(n18178), .ZN(n18179) );
  NOR2_X1 U12951 ( .A1(n11801), .A2(n16914), .ZN(n14607) );
  AOI21_X1 U12952 ( .B1(n10406), .B2(n11766), .A(n10405), .ZN(n11763) );
  NAND2_X1 U12953 ( .A1(n12758), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12791) );
  INV_X1 U12954 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16253) );
  INV_X1 U12955 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20344) );
  AND2_X1 U12956 ( .A1(n14167), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14168) );
  NAND2_X1 U12957 ( .A1(n20376), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14165) );
  AND2_X1 U12958 ( .A1(n12413), .A2(n12412), .ZN(n14787) );
  NOR2_X1 U12959 ( .A1(n13667), .A2(n13666), .ZN(n13974) );
  XNOR2_X1 U12960 ( .A(n12987), .B(n12986), .ZN(n14167) );
  INV_X1 U12962 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12506) );
  NOR2_X1 U12963 ( .A1(n10248), .A2(n12231), .ZN(n12233) );
  AND2_X1 U12964 ( .A1(n12401), .A2(n12400), .ZN(n14822) );
  OR2_X1 U12965 ( .A1(n15243), .A2(n16399), .ZN(n12454) );
  NAND2_X1 U12966 ( .A1(n12184), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12185) );
  AND2_X1 U12967 ( .A1(n12078), .A2(n14027), .ZN(n20742) );
  AND2_X1 U12968 ( .A1(n20620), .A2(n20624), .ZN(n20625) );
  AND2_X1 U12969 ( .A1(n20652), .A2(n14285), .ZN(n15315) );
  OR2_X1 U12970 ( .A1(n20784), .A2(n20783), .ZN(n20853) );
  OR2_X1 U12971 ( .A1(n20784), .A2(n14072), .ZN(n20860) );
  INV_X1 U12972 ( .A(n20910), .ZN(n20781) );
  NOR2_X1 U12973 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16184) );
  OR3_X1 U12974 ( .A1(n11233), .A2(n11232), .A3(n11231), .ZN(n13867) );
  NOR2_X1 U12975 ( .A1(n15616), .A2(n15348), .ZN(n15347) );
  NOR2_X1 U12976 ( .A1(n16534), .A2(n16535), .ZN(n16533) );
  NAND2_X1 U12977 ( .A1(n13491), .A2(n13052), .ZN(n13053) );
  AND2_X1 U12978 ( .A1(n19287), .A2(n11530), .ZN(n15721) );
  INV_X1 U12979 ( .A(n19669), .ZN(n16143) );
  INV_X1 U12980 ( .A(n13867), .ZN(n13541) );
  AND3_X1 U12981 ( .A1(n13546), .A2(n13573), .A3(n13545), .ZN(n13875) );
  NAND2_X1 U12982 ( .A1(n10943), .A2(n10942), .ZN(n13868) );
  INV_X1 U12983 ( .A(n19745), .ZN(n19835) );
  INV_X1 U12984 ( .A(n19744), .ZN(n20260) );
  OR2_X1 U12985 ( .A1(n20271), .A2(n20284), .ZN(n20046) );
  INV_X1 U12986 ( .A(n19693), .ZN(n19699) );
  NOR2_X1 U12987 ( .A1(n11763), .A2(n11758), .ZN(n16913) );
  OR2_X1 U12988 ( .A1(n16937), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U12989 ( .A1(n19130), .A2(n17053), .ZN(n17043) );
  INV_X1 U12990 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17166) );
  NAND2_X1 U12991 ( .A1(n19231), .A2(n17206), .ZN(n10414) );
  INV_X1 U12992 ( .A(n17402), .ZN(n17400) );
  INV_X1 U12993 ( .A(n18208), .ZN(n17840) );
  NOR2_X1 U12994 ( .A1(n9961), .A2(n17924), .ZN(n10283) );
  AOI21_X1 U12995 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17980), .A(
        n18585), .ZN(n18028) );
  NAND2_X1 U12996 ( .A1(n11799), .A2(n18099), .ZN(n18396) );
  INV_X1 U12997 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18144) );
  INV_X1 U12998 ( .A(n18552), .ZN(n19215) );
  NAND2_X1 U12999 ( .A1(n16101), .A2(n16100), .ZN(n16188) );
  NOR2_X1 U13000 ( .A1(n11731), .A2(n18020), .ZN(n18263) );
  INV_X1 U13001 ( .A(n18396), .ZN(n18021) );
  OR2_X1 U13002 ( .A1(n18312), .A2(n18488), .ZN(n18447) );
  NOR2_X1 U13003 ( .A1(n19230), .A2(n14438), .ZN(n19010) );
  NOR2_X1 U13004 ( .A1(n10307), .A2(n10306), .ZN(n18563) );
  INV_X1 U13005 ( .A(n19003), .ZN(n16741) );
  INV_X1 U13006 ( .A(n13953), .ZN(n14709) );
  INV_X1 U13007 ( .A(n21391), .ZN(n20378) );
  NOR2_X1 U13008 ( .A1(n14647), .A2(n20373), .ZN(n16304) );
  INV_X1 U13009 ( .A(n20379), .ZN(n21393) );
  NOR2_X1 U13010 ( .A1(n14165), .A2(n14159), .ZN(n20353) );
  INV_X1 U13011 ( .A(n14906), .ZN(n20404) );
  AND2_X1 U13012 ( .A1(n14985), .A2(n14662), .ZN(n14636) );
  AOI21_X1 U13013 ( .B1(n13959), .B2(n13958), .A(n13957), .ZN(n13960) );
  NAND2_X1 U13014 ( .A1(n12676), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12706) );
  NOR2_X1 U13015 ( .A1(n12507), .A2(n12506), .ZN(n12524) );
  AND2_X1 U13016 ( .A1(n12395), .A2(n12394), .ZN(n14857) );
  OR2_X1 U13017 ( .A1(n14430), .A2(n15300), .ZN(n16436) );
  INV_X1 U13018 ( .A(n12460), .ZN(n20473) );
  AND2_X1 U13019 ( .A1(n12461), .A2(n14696), .ZN(n14433) );
  INV_X1 U13020 ( .A(n20526), .ZN(n20543) );
  INV_X1 U13021 ( .A(n20783), .ZN(n20547) );
  OAI211_X1 U13022 ( .C1(n20817), .C2(n20585), .A(n20584), .B(n20583), .ZN(
        n20609) );
  AND2_X1 U13023 ( .A1(n20623), .A2(n20574), .ZN(n20645) );
  OAI21_X1 U13024 ( .B1(n20660), .B2(n20676), .A(n20874), .ZN(n20678) );
  OAI211_X1 U13025 ( .C1(n20911), .C2(n14293), .A(n14292), .B(n20781), .ZN(
        n14317) );
  INV_X1 U13026 ( .A(n20853), .ZN(n20805) );
  OAI21_X1 U13027 ( .B1(n20821), .B2(n20820), .A(n20819), .ZN(n20856) );
  NOR2_X2 U13028 ( .A1(n20784), .A2(n14071), .ZN(n20855) );
  INV_X1 U13029 ( .A(n20860), .ZN(n20899) );
  INV_X1 U13030 ( .A(n14342), .ZN(n20522) );
  INV_X1 U13031 ( .A(n20517), .ZN(n20542) );
  INV_X1 U13032 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20992) );
  INV_X1 U13033 ( .A(n21034), .ZN(n21038) );
  AND2_X1 U13034 ( .A1(n13862), .A2(n13899), .ZN(n13503) );
  INV_X1 U13035 ( .A(n19414), .ZN(n19449) );
  AND2_X1 U13036 ( .A1(n11194), .A2(n11193), .ZN(n14249) );
  AND2_X1 U13037 ( .A1(n14686), .A2(n14688), .ZN(n19460) );
  AND3_X1 U13038 ( .A1(n11137), .A2(n11136), .A3(n11135), .ZN(n15935) );
  INV_X1 U13039 ( .A(n20292), .ZN(n19453) );
  INV_X1 U13040 ( .A(n13702), .ZN(n19604) );
  INV_X1 U13041 ( .A(n19642), .ZN(n16638) );
  NAND2_X1 U13042 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  INV_X1 U13043 ( .A(n19650), .ZN(n19660) );
  OAI21_X1 U13044 ( .B1(n16034), .B2(n16033), .A(n16032), .ZN(n19703) );
  INV_X1 U13045 ( .A(n19739), .ZN(n19731) );
  AND2_X1 U13046 ( .A1(n20264), .A2(n20292), .ZN(n19745) );
  AND2_X1 U13047 ( .A1(n19745), .A2(n19744), .ZN(n19792) );
  NAND2_X1 U13048 ( .A1(n16059), .A2(n16058), .ZN(n19814) );
  NOR2_X2 U13049 ( .A1(n19835), .A2(n20046), .ZN(n19830) );
  NOR2_X2 U13050 ( .A1(n19866), .A2(n20046), .ZN(n19857) );
  NOR2_X1 U13051 ( .A1(n20257), .A2(n19835), .ZN(n19892) );
  INV_X1 U13052 ( .A(n19962), .ZN(n19954) );
  AND2_X1 U13053 ( .A1(n20048), .A2(n19931), .ZN(n19974) );
  AND2_X1 U13054 ( .A1(n14189), .A2(n14188), .ZN(n19997) );
  INV_X1 U13055 ( .A(n20038), .ZN(n20030) );
  NOR2_X1 U13056 ( .A1(n20002), .A2(n20046), .ZN(n20062) );
  OAI21_X1 U13057 ( .B1(n20085), .B2(n20084), .A(n20083), .ZN(n20111) );
  INV_X1 U13058 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20200) );
  NAND2_X1 U13059 ( .A1(n19213), .A2(n19001), .ZN(n17784) );
  NAND2_X1 U13060 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  INV_X1 U13061 ( .A(n17265), .ZN(n17258) );
  NOR2_X1 U13062 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17039), .ZN(n17024) );
  NOR2_X1 U13063 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17056), .ZN(n17047) );
  NOR2_X1 U13064 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17107), .ZN(n17088) );
  NOR2_X1 U13065 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17198), .ZN(n17184) );
  NOR2_X2 U13066 ( .A1(n19169), .A2(n17246), .ZN(n17244) );
  NAND2_X1 U13067 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17349), .ZN(n17332) );
  AND2_X1 U13068 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17362), .ZN(n17349) );
  INV_X1 U13069 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17542) );
  OAI21_X1 U13070 ( .B1(n14610), .B2(n14441), .A(n19213), .ZN(n16204) );
  INV_X1 U13071 ( .A(n17642), .ZN(n17638) );
  NAND4_X1 U13072 ( .A1(n17686), .A2(P3_EAX_REG_10__SCAN_IN), .A3(
        P3_EAX_REG_9__SCAN_IN), .A4(n17573), .ZN(n17661) );
  NOR2_X1 U13073 ( .A1(n17659), .A2(n17658), .ZN(n17708) );
  CLKBUF_X1 U13074 ( .A(n17824), .Z(n17821) );
  NOR2_X1 U13075 ( .A1(n17897), .A2(n17898), .ZN(n17876) );
  INV_X1 U13076 ( .A(n18001), .ZN(n17976) );
  NAND2_X1 U13077 ( .A1(n16773), .A2(n18396), .ZN(n18348) );
  NOR2_X2 U13078 ( .A1(n18201), .A2(n17691), .ZN(n18110) );
  INV_X1 U13079 ( .A(n18194), .ZN(n18169) );
  INV_X1 U13080 ( .A(n18197), .ZN(n18183) );
  NAND2_X1 U13081 ( .A1(n16745), .A2(n10260), .ZN(n16751) );
  AND2_X1 U13082 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18406) );
  INV_X1 U13083 ( .A(n18325), .ZN(n18441) );
  NOR2_X1 U13084 ( .A1(n11770), .A2(n11755), .ZN(n18452) );
  NAND2_X1 U13085 ( .A1(n19022), .A2(n11803), .ZN(n19020) );
  NOR2_X1 U13086 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19169), .ZN(
        n19193) );
  INV_X1 U13087 ( .A(n18913), .ZN(n18798) );
  INV_X1 U13088 ( .A(n18650), .ZN(n18652) );
  INV_X1 U13089 ( .A(n18668), .ZN(n18699) );
  INV_X1 U13090 ( .A(n18557), .ZN(n18585) );
  INV_X1 U13091 ( .A(n18996), .ZN(n18969) );
  NOR2_X1 U13092 ( .A1(n19218), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18198) );
  INV_X1 U13093 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19218) );
  INV_X1 U13094 ( .A(n14685), .ZN(n14688) );
  NOR2_X1 U13095 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13490), .ZN(n16890)
         );
  NAND2_X1 U13096 ( .A1(n13555), .A2(n13554), .ZN(n21064) );
  INV_X1 U13097 ( .A(n20377), .ZN(n21390) );
  NAND2_X1 U13098 ( .A1(n20376), .A2(n14153), .ZN(n21403) );
  INV_X1 U13099 ( .A(n13978), .ZN(n20408) );
  NAND2_X1 U13100 ( .A1(n20408), .A2(n11958), .ZN(n14899) );
  OR2_X1 U13101 ( .A1(n20414), .A2(n21067), .ZN(n20412) );
  INV_X1 U13102 ( .A(n20414), .ZN(n20440) );
  AND2_X1 U13103 ( .A1(n13959), .A2(n13759), .ZN(n13768) );
  INV_X1 U13104 ( .A(n20486), .ZN(n20504) );
  INV_X1 U13105 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20514) );
  AOI22_X1 U13106 ( .A1(n20525), .A2(n20521), .B1(n20808), .B2(n20654), .ZN(
        n20546) );
  NAND2_X1 U13107 ( .A1(n20623), .A2(n20547), .ZN(n20607) );
  AOI22_X1 U13108 ( .A1(n20581), .A2(n20578), .B1(n10262), .B2(n20808), .ZN(
        n20612) );
  INV_X1 U13109 ( .A(n20621), .ZN(n20649) );
  NAND2_X1 U13110 ( .A1(n20687), .A2(n9729), .ZN(n20707) );
  AOI22_X1 U13111 ( .A1(n20710), .A2(n20715), .B1(n20868), .B2(n10262), .ZN(
        n20737) );
  INV_X1 U13112 ( .A(n20772), .ZN(n14320) );
  NAND2_X1 U13113 ( .A1(n20739), .A2(n20861), .ZN(n20804) );
  AOI22_X1 U13114 ( .A1(n20810), .A2(n20820), .B1(n20809), .B2(n20808), .ZN(
        n20859) );
  AOI211_X2 U13115 ( .C1(n14070), .C2(n14073), .A(n14069), .B(n20910), .ZN(
        n14108) );
  AOI22_X1 U13116 ( .A1(n20869), .A2(n20875), .B1(n20868), .B2(n20867), .ZN(
        n20904) );
  NAND2_X1 U13117 ( .A1(n20862), .A2(n20574), .ZN(n14381) );
  INV_X1 U13118 ( .A(n21048), .ZN(n20980) );
  INV_X1 U13119 ( .A(n21056), .ZN(n21058) );
  NAND2_X1 U13120 ( .A1(n13864), .A2(n13503), .ZN(n13510) );
  OR2_X1 U13121 ( .A1(n12994), .A2(n12993), .ZN(n13524) );
  NAND2_X1 U13122 ( .A1(n13080), .A2(n13060), .ZN(n19414) );
  NAND2_X1 U13123 ( .A1(n13080), .A2(n13079), .ZN(n19447) );
  INV_X1 U13124 ( .A(n19379), .ZN(n19442) );
  INV_X1 U13125 ( .A(n13463), .ZN(n13464) );
  NAND2_X1 U13126 ( .A1(n13694), .A2(n13693), .ZN(n20264) );
  INV_X1 U13127 ( .A(n19505), .ZN(n19527) );
  AOI21_X2 U13128 ( .B1(n13573), .B2(n13572), .A(n19533), .ZN(n19489) );
  NOR2_X1 U13129 ( .A1(n19523), .A2(n19505), .ZN(n19501) );
  INV_X1 U13130 ( .A(n19491), .ZN(n19531) );
  NAND2_X1 U13131 ( .A1(n19602), .A2(n19540), .ZN(n19558) );
  INV_X1 U13132 ( .A(n19556), .ZN(n19569) );
  NAND2_X1 U13133 ( .A1(n19537), .A2(n20188), .ZN(n19602) );
  INV_X1 U13134 ( .A(n13007), .ZN(n13008) );
  NAND2_X1 U13135 ( .A1(n12996), .A2(n14195), .ZN(n19619) );
  NOR2_X1 U13136 ( .A1(n11610), .A2(n11609), .ZN(n11611) );
  INV_X1 U13137 ( .A(n19663), .ZN(n16702) );
  NAND2_X1 U13138 ( .A1(n11587), .A2(n10983), .ZN(n19650) );
  AND2_X1 U13139 ( .A1(n16112), .A2(n16117), .ZN(n16726) );
  INV_X1 U13140 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20278) );
  INV_X1 U13141 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13552) );
  AOI211_X2 U13142 ( .C1(n16030), .C2(n16033), .A(n16029), .B(n19874), .ZN(
        n19707) );
  INV_X1 U13143 ( .A(n19762), .ZN(n19770) );
  INV_X1 U13144 ( .A(n19792), .ZN(n19800) );
  INV_X1 U13145 ( .A(n19814), .ZN(n19805) );
  AND2_X1 U13146 ( .A1(n14134), .A2(n14133), .ZN(n19834) );
  INV_X1 U13147 ( .A(n19892), .ZN(n19899) );
  INV_X1 U13148 ( .A(n19922), .ZN(n19930) );
  NAND2_X1 U13149 ( .A1(n20072), .A2(n19931), .ZN(n19962) );
  INV_X1 U13150 ( .A(n19974), .ZN(n19982) );
  INV_X1 U13151 ( .A(n19998), .ZN(n19995) );
  INV_X1 U13152 ( .A(n20109), .ZN(n20073) );
  INV_X1 U13153 ( .A(n20062), .ZN(n20070) );
  AOI21_X1 U13154 ( .B1(n20081), .B2(n20084), .A(n20079), .ZN(n20115) );
  INV_X1 U13155 ( .A(n20105), .ZN(n20167) );
  INV_X1 U13156 ( .A(n20256), .ZN(n20179) );
  NOR2_X1 U13157 ( .A1(n19000), .A2(n17784), .ZN(n19231) );
  INV_X1 U13158 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16911) );
  NOR2_X1 U13159 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17148), .ZN(n17146) );
  NAND4_X1 U13160 ( .A1(n18418), .A2(n17205), .A3(n19076), .A4(n19066), .ZN(
        n17268) );
  NOR2_X1 U13161 ( .A1(n16980), .A2(n14532), .ZN(n17310) );
  NOR2_X2 U13162 ( .A1(n17560), .A2(n18589), .ZN(n17569) );
  INV_X1 U13163 ( .A(n17719), .ZN(n17654) );
  INV_X1 U13164 ( .A(n11810), .ZN(n17691) );
  NOR2_X1 U13165 ( .A1(n11655), .A2(n11654), .ZN(n17705) );
  INV_X1 U13166 ( .A(n17729), .ZN(n17748) );
  INV_X1 U13167 ( .A(n17770), .ZN(n17780) );
  INV_X1 U13168 ( .A(n17831), .ZN(n17826) );
  NAND2_X1 U13169 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18193), .ZN(n18035) );
  INV_X1 U13170 ( .A(n18110), .ZN(n17979) );
  NOR2_X1 U13171 ( .A1(n18183), .A2(n18031), .ZN(n18193) );
  NAND2_X1 U13172 ( .A1(n16751), .A2(n16750), .ZN(n16806) );
  NAND2_X1 U13173 ( .A1(n11817), .A2(n18512), .ZN(n18325) );
  INV_X1 U13174 ( .A(n18458), .ZN(n18513) );
  INV_X1 U13175 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18577) );
  INV_X1 U13176 ( .A(n18934), .ZN(n18910) );
  INV_X1 U13177 ( .A(n18878), .ZN(n18948) );
  INV_X1 U13178 ( .A(n18864), .ZN(n18980) );
  INV_X1 U13179 ( .A(n19166), .ZN(n19081) );
  INV_X1 U13180 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19096) );
  OAI21_X1 U13181 ( .B1(n15608), .B2(n16702), .A(n11611), .ZN(P2_U3018) );
  INV_X1 U13182 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16768) );
  INV_X1 U13183 ( .A(n18065), .ZN(n18101) );
  NAND2_X1 U13184 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18066) );
  NAND2_X1 U13185 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17995) );
  NAND2_X1 U13186 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17963) );
  NAND2_X1 U13187 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17925) );
  NAND2_X1 U13188 ( .A1(n17902), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17875) );
  NAND2_X1 U13189 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17884) );
  NAND2_X1 U13190 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17843) );
  INV_X1 U13191 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16934) );
  XNOR2_X1 U13192 ( .A(n16768), .B(n10287), .ZN(n16772) );
  AOI21_X1 U13193 ( .B1(n16934), .B2(n16752), .A(n10287), .ZN(n16933) );
  INV_X1 U13194 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17857) );
  INV_X1 U13195 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17897) );
  INV_X1 U13196 ( .A(n10283), .ZN(n10280) );
  NOR2_X1 U13197 ( .A1(n17925), .A2(n10280), .ZN(n10278) );
  INV_X1 U13198 ( .A(n10278), .ZN(n17898) );
  INV_X1 U13199 ( .A(n17876), .ZN(n10277) );
  NAND2_X1 U13200 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17838), .ZN(
        n10274) );
  NOR2_X1 U13201 ( .A1(n17857), .A2(n10274), .ZN(n10273) );
  OAI21_X1 U13202 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n10273), .A(
        n16752), .ZN(n17846) );
  INV_X1 U13203 ( .A(n17846), .ZN(n16945) );
  AOI21_X1 U13204 ( .B1(n17857), .B2(n10274), .A(n10273), .ZN(n17853) );
  OAI21_X1 U13205 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17838), .A(
        n10274), .ZN(n10275) );
  INV_X1 U13206 ( .A(n10275), .ZN(n17867) );
  INV_X1 U13207 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16973) );
  NAND2_X1 U13208 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17876), .ZN(
        n10276) );
  AOI21_X1 U13209 ( .B1(n16973), .B2(n10276), .A(n17838), .ZN(n17877) );
  INV_X1 U13210 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21279) );
  OAI22_X1 U13211 ( .A1(n21279), .A2(n10277), .B1(n17876), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17895) );
  INV_X1 U13212 ( .A(n17895), .ZN(n16986) );
  AOI21_X1 U13213 ( .B1(n17897), .B2(n17898), .A(n17876), .ZN(n17903) );
  INV_X1 U13214 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17927) );
  NAND2_X1 U13215 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10283), .ZN(
        n10279) );
  AOI21_X1 U13216 ( .B1(n17927), .B2(n10279), .A(n10278), .ZN(n17929) );
  INV_X1 U13217 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17933) );
  AOI22_X1 U13218 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10283), .B1(
        n10280), .B2(n17933), .ZN(n17936) );
  INV_X1 U13219 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17923) );
  NAND2_X1 U13220 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10281), .ZN(
        n10286) );
  NOR2_X1 U13221 ( .A1(n9977), .A2(n10286), .ZN(n17956) );
  INV_X1 U13222 ( .A(n17956), .ZN(n10282) );
  NOR2_X1 U13223 ( .A1(n17963), .A2(n10282), .ZN(n10284) );
  INV_X1 U13224 ( .A(n10284), .ZN(n17920) );
  AOI21_X1 U13225 ( .B1(n17923), .B2(n17920), .A(n10283), .ZN(n17951) );
  INV_X1 U13226 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17035) );
  NAND2_X1 U13227 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17956), .ZN(
        n10285) );
  AOI21_X1 U13228 ( .B1(n17035), .B2(n10285), .A(n10284), .ZN(n17957) );
  INV_X1 U13229 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17973) );
  XNOR2_X1 U13230 ( .A(n17973), .B(n17956), .ZN(n17970) );
  AOI21_X1 U13231 ( .B1(n9977), .B2(n10286), .A(n17956), .ZN(n17984) );
  NOR2_X1 U13232 ( .A1(n9961), .A2(n17994), .ZN(n17992) );
  NAND2_X1 U13233 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17992), .ZN(
        n17075) );
  INV_X1 U13234 ( .A(n17075), .ZN(n10289) );
  INV_X1 U13235 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17256) );
  NAND2_X1 U13236 ( .A1(n10287), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10288) );
  INV_X1 U13237 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16755) );
  INV_X1 U13238 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13239 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10281), .B1(
        n10290), .B2(n17075), .ZN(n17993) );
  NOR2_X1 U13240 ( .A1(n17066), .A2(n17993), .ZN(n17065) );
  NOR2_X1 U13241 ( .A1(n17046), .A2(n9965), .ZN(n17032) );
  NOR2_X1 U13242 ( .A1(n17957), .A2(n17032), .ZN(n17033) );
  NOR2_X1 U13243 ( .A1(n17033), .A2(n9968), .ZN(n17023) );
  NOR2_X1 U13244 ( .A1(n17951), .A2(n17023), .ZN(n17022) );
  NOR2_X1 U13245 ( .A1(n17022), .A2(n9968), .ZN(n17011) );
  NOR2_X1 U13246 ( .A1(n17936), .A2(n17011), .ZN(n17012) );
  NOR2_X1 U13247 ( .A1(n17012), .A2(n9968), .ZN(n17003) );
  NOR2_X1 U13248 ( .A1(n17929), .A2(n17003), .ZN(n17004) );
  NOR2_X1 U13249 ( .A1(n17004), .A2(n9968), .ZN(n16992) );
  NOR2_X1 U13250 ( .A1(n16972), .A2(n9968), .ZN(n16963) );
  NOR2_X1 U13251 ( .A1(n16945), .A2(n16944), .ZN(n16943) );
  NOR2_X1 U13252 ( .A1(n16943), .A2(n9968), .ZN(n16931) );
  NOR2_X1 U13253 ( .A1(n16932), .A2(n9968), .ZN(n11612) );
  XOR2_X1 U13254 ( .A(n16772), .B(n11612), .Z(n10291) );
  INV_X1 U13255 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19228) );
  AND4_X1 U13256 ( .A1(n19218), .A2(n19228), .A3(n16911), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17229) );
  NAND2_X1 U13257 ( .A1(n10291), .A2(n17229), .ZN(n10422) );
  NOR2_X1 U13258 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19229) );
  NAND3_X1 U13259 ( .A1(n19218), .A2(n19228), .A3(n19229), .ZN(n18418) );
  NOR2_X2 U13260 ( .A1(n10296), .A2(n10297), .ZN(n11656) );
  AOI22_X1 U13261 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13262 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13263 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10293) );
  BUF_X2 U13264 ( .A(n11661), .Z(n14519) );
  AOI22_X1 U13265 ( .A1(n11673), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10292) );
  NAND4_X1 U13266 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10307) );
  NOR2_X2 U13267 ( .A1(n10299), .A2(n10296), .ZN(n11704) );
  INV_X4 U13268 ( .A(n10374), .ZN(n14520) );
  AOI22_X1 U13269 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10305) );
  INV_X2 U13270 ( .A(n10245), .ZN(n17423) );
  AOI22_X1 U13271 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13272 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10303) );
  NOR2_X2 U13273 ( .A1(n10299), .A2(n19033), .ZN(n11671) );
  AOI22_X1 U13274 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10302) );
  NAND4_X1 U13275 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10306) );
  AOI22_X1 U13276 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10320) );
  BUF_X2 U13277 ( .A(n11624), .Z(n17523) );
  AOI22_X1 U13278 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10319) );
  INV_X4 U13279 ( .A(n10309), .ZN(n17503) );
  INV_X4 U13280 ( .A(n10310), .ZN(n17526) );
  AOI22_X1 U13281 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10311) );
  OAI21_X1 U13282 ( .B1(n14469), .B2(n21223), .A(n10311), .ZN(n10317) );
  AOI22_X1 U13283 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13284 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13285 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13286 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10312) );
  NAND4_X1 U13287 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10316) );
  AOI22_X1 U13288 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13289 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10329) );
  INV_X1 U13290 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18550) );
  AOI22_X1 U13291 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10321) );
  OAI21_X1 U13292 ( .B1(n17525), .B2(n18550), .A(n10321), .ZN(n10327) );
  INV_X2 U13293 ( .A(n14458), .ZN(n17504) );
  AOI22_X1 U13294 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13295 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13296 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13297 ( .A1(n11673), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13298 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  AOI22_X1 U13299 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13300 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13301 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13302 ( .A1(n17533), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10332) );
  NAND4_X1 U13303 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(
        n10341) );
  AOI22_X1 U13304 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13305 ( .A1(n11704), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13306 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13307 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10336) );
  NAND4_X1 U13308 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10340) );
  NOR2_X1 U13309 ( .A1(n17206), .A2(n18589), .ZN(n10388) );
  INV_X1 U13310 ( .A(n10388), .ZN(n10392) );
  AOI22_X1 U13311 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9731), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13312 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10351) );
  INV_X1 U13313 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18584) );
  AOI22_X1 U13314 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17504), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10343) );
  OAI21_X1 U13315 ( .B1(n17525), .B2(n18584), .A(n10343), .ZN(n10349) );
  AOI22_X1 U13316 ( .A1(n17526), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13317 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13318 ( .A1(n10308), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13319 ( .A1(n11673), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13320 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  AOI22_X1 U13321 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13322 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13323 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10353) );
  OAI21_X1 U13324 ( .B1(n17525), .B2(n18577), .A(n10353), .ZN(n10359) );
  AOI22_X1 U13325 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13326 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13327 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13328 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10354) );
  NAND4_X1 U13329 ( .A1(n10357), .A2(n10356), .A3(n10355), .A4(n10354), .ZN(
        n10358) );
  AOI211_X1 U13330 ( .C1(n17423), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n10359), .B(n10358), .ZN(n10360) );
  NAND3_X1 U13331 ( .A1(n10362), .A2(n10361), .A3(n10360), .ZN(n17578) );
  NOR4_X2 U13332 ( .A1(n10391), .A2(n14440), .A3(n10392), .A4(n10390), .ZN(
        n10394) );
  AOI22_X1 U13333 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13334 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13335 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13336 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13337 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10372) );
  AOI22_X1 U13338 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13339 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13340 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13341 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10367) );
  NAND4_X1 U13342 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10371) );
  AOI22_X1 U13343 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13344 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13345 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10373) );
  OAI21_X1 U13346 ( .B1(n10374), .B2(n21174), .A(n10373), .ZN(n10380) );
  AOI22_X1 U13347 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13348 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13349 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13350 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13351 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  AOI211_X1 U13352 ( .C1(n17504), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n10380), .B(n10379), .ZN(n10381) );
  NAND3_X1 U13353 ( .A1(n10383), .A2(n10382), .A3(n10381), .ZN(n11746) );
  INV_X1 U13354 ( .A(n11746), .ZN(n18558) );
  NAND2_X1 U13355 ( .A1(n11801), .A2(n18558), .ZN(n11748) );
  NAND2_X1 U13356 ( .A1(n17578), .A2(n18558), .ZN(n11760) );
  INV_X1 U13357 ( .A(n11760), .ZN(n11802) );
  NAND2_X1 U13358 ( .A1(n18552), .A2(n17206), .ZN(n11800) );
  AOI21_X1 U13359 ( .B1(n17659), .B2(n16209), .A(n11800), .ZN(n11752) );
  INV_X1 U13360 ( .A(n11752), .ZN(n10384) );
  AOI221_X1 U13361 ( .B1(n11802), .B2(n10384), .C1(n10393), .C2(n10384), .A(
        n18563), .ZN(n10389) );
  NAND2_X1 U13362 ( .A1(n10390), .A2(n14440), .ZN(n10385) );
  OAI22_X1 U13363 ( .A1(n18589), .A2(n10385), .B1(n19037), .B2(n14440), .ZN(
        n10387) );
  INV_X1 U13364 ( .A(n17575), .ZN(n18580) );
  NOR2_X1 U13365 ( .A1(n18580), .A2(n11760), .ZN(n11767) );
  OAI21_X1 U13366 ( .B1(n10393), .B2(n11767), .A(n18547), .ZN(n10386) );
  OAI211_X1 U13367 ( .C1(n10388), .C2(n10391), .A(n10387), .B(n10386), .ZN(
        n11753) );
  NAND2_X1 U13368 ( .A1(n10394), .A2(n11809), .ZN(n11803) );
  NOR2_X1 U13369 ( .A1(n18580), .A2(n17578), .ZN(n11749) );
  NAND2_X1 U13370 ( .A1(n11749), .A2(n19015), .ZN(n14439) );
  NOR2_X1 U13371 ( .A1(n10392), .A2(n14439), .ZN(n10395) );
  NAND2_X1 U13372 ( .A1(n10394), .A2(n11746), .ZN(n11754) );
  NAND2_X1 U13373 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18198), .ZN(n19068) );
  AOI22_X1 U13374 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19049), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19186), .ZN(n10398) );
  INV_X1 U13375 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19044) );
  OAI22_X1 U13376 ( .A1(n19192), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n19044), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11762) );
  XOR2_X1 U13377 ( .A(n10398), .B(n10397), .Z(n10406) );
  NAND2_X1 U13378 ( .A1(n10398), .A2(n10397), .ZN(n10399) );
  OAI21_X1 U13379 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19186), .A(
        n10399), .ZN(n10400) );
  OAI22_X1 U13380 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19053), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10400), .ZN(n10402) );
  NOR2_X1 U13381 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19053), .ZN(
        n10401) );
  NAND2_X1 U13382 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10400), .ZN(
        n10403) );
  AOI22_X1 U13383 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10402), .B1(
        n10401), .B2(n10403), .ZN(n11766) );
  AOI21_X1 U13384 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10403), .A(
        n10402), .ZN(n10404) );
  AOI21_X1 U13385 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19053), .A(
        n10404), .ZN(n10407) );
  INV_X1 U13386 ( .A(n10407), .ZN(n10405) );
  INV_X1 U13387 ( .A(n11762), .ZN(n10409) );
  OAI21_X1 U13388 ( .B1(n10409), .B2(n11757), .A(n10407), .ZN(n10408) );
  NOR2_X2 U13389 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19169), .ZN(n19072) );
  NAND2_X1 U13390 ( .A1(n18198), .A2(n19072), .ZN(n19066) );
  INV_X2 U13391 ( .A(n19226), .ZN(n19225) );
  NAND2_X2 U13392 ( .A1(n19225), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19156) );
  OAI211_X1 U13393 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19096), .B(n19156), .ZN(n19088) );
  NAND2_X1 U13394 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19210) );
  INV_X1 U13395 ( .A(n19210), .ZN(n19216) );
  AOI211_X1 U13396 ( .C1(n19088), .C2(n18552), .A(n19216), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n10412) );
  INV_X1 U13397 ( .A(n10412), .ZN(n19061) );
  NOR2_X1 U13398 ( .A1(n17246), .A2(n17247), .ZN(n17070) );
  INV_X1 U13399 ( .A(n17070), .ZN(n17267) );
  NAND3_X1 U13400 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n10411) );
  INV_X1 U13401 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19144) );
  NAND2_X1 U13402 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n10415) );
  INV_X1 U13403 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19142) );
  INV_X1 U13404 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19136) );
  INV_X1 U13405 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19130) );
  INV_X1 U13406 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19127) );
  INV_X1 U13407 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19122) );
  INV_X1 U13408 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19118) );
  INV_X1 U13409 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19113) );
  INV_X1 U13410 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19110) );
  INV_X1 U13411 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19106) );
  INV_X1 U13412 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n21303) );
  INV_X1 U13413 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19102) );
  INV_X1 U13414 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19099) );
  NOR3_X1 U13415 ( .A1(n21303), .A2(n19102), .A3(n19099), .ZN(n17217) );
  NAND2_X1 U13416 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17217), .ZN(n17197) );
  NOR2_X1 U13417 ( .A1(n19106), .A2(n17197), .ZN(n17172) );
  NAND2_X1 U13418 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17172), .ZN(n17176) );
  NOR3_X1 U13419 ( .A1(n19113), .A2(n19110), .A3(n17176), .ZN(n17141) );
  NAND3_X1 U13420 ( .A1(n17141), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n17124) );
  NOR2_X1 U13421 ( .A1(n19118), .A2(n17124), .ZN(n17117) );
  NAND2_X1 U13422 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17117), .ZN(n17098) );
  NOR2_X1 U13423 ( .A1(n19122), .A2(n17098), .ZN(n17090) );
  NAND2_X1 U13424 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17090), .ZN(n17071) );
  NOR2_X1 U13425 ( .A1(n19127), .A2(n17071), .ZN(n17064) );
  NAND2_X1 U13426 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17064), .ZN(n17053) );
  NAND3_X1 U13427 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n17043), .ZN(n17021) );
  NAND3_X1 U13428 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n17020), .ZN(n16995) );
  NOR2_X1 U13429 ( .A1(n19142), .A2(n16995), .ZN(n16982) );
  OAI21_X1 U13430 ( .B1(n17245), .B2(n16982), .A(n17268), .ZN(n16989) );
  AOI221_X1 U13431 ( .B1(n17267), .B2(n19144), .C1(n17267), .C2(n10415), .A(
        n16989), .ZN(n16969) );
  INV_X1 U13432 ( .A(n16969), .ZN(n10410) );
  AOI21_X1 U13433 ( .B1(n17267), .B2(n10411), .A(n10410), .ZN(n16940) );
  INV_X1 U13434 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19157) );
  OAI22_X1 U13435 ( .A1(n16940), .A2(n19157), .B1(n16768), .B2(n17254), .ZN(
        n10420) );
  AOI211_X4 U13436 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19215), .A(n10412), .B(
        n10414), .ZN(n17266) );
  NAND2_X1 U13437 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19215), .ZN(n10413) );
  AOI211_X4 U13438 ( .C1(n19210), .C2(n16911), .A(n10414), .B(n10413), .ZN(
        n17265) );
  NOR3_X1 U13439 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17238) );
  INV_X1 U13440 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17552) );
  NAND2_X1 U13441 ( .A1(n17238), .A2(n17552), .ZN(n17230) );
  NOR2_X1 U13442 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17230), .ZN(n17207) );
  INV_X1 U13443 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17204) );
  NAND2_X1 U13444 ( .A1(n17207), .A2(n17204), .ZN(n17198) );
  NAND2_X1 U13445 ( .A1(n17184), .A2(n17542), .ZN(n17181) );
  INV_X1 U13446 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17430) );
  NAND2_X1 U13447 ( .A1(n17162), .A2(n17430), .ZN(n17148) );
  INV_X1 U13448 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17135) );
  NAND2_X1 U13449 ( .A1(n17146), .A2(n17135), .ZN(n17128) );
  INV_X1 U13450 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17110) );
  NAND2_X1 U13451 ( .A1(n17111), .A2(n17110), .ZN(n17107) );
  INV_X1 U13452 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17085) );
  NAND2_X1 U13453 ( .A1(n17088), .A2(n17085), .ZN(n17082) );
  INV_X1 U13454 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17401) );
  NAND2_X1 U13455 ( .A1(n17067), .A2(n17401), .ZN(n17056) );
  INV_X1 U13456 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17042) );
  NAND2_X1 U13457 ( .A1(n17047), .A2(n17042), .ZN(n17039) );
  INV_X1 U13458 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17348) );
  NAND2_X1 U13459 ( .A1(n17024), .A2(n17348), .ZN(n17014) );
  INV_X1 U13460 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17274) );
  NAND2_X1 U13461 ( .A1(n17002), .A2(n17274), .ZN(n16998) );
  NOR2_X1 U13462 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16998), .ZN(n16970) );
  INV_X1 U13463 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16980) );
  NAND2_X1 U13464 ( .A1(n16970), .A2(n16980), .ZN(n16961) );
  NOR2_X1 U13465 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16961), .ZN(n16960) );
  INV_X1 U13466 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17300) );
  NAND2_X1 U13467 ( .A1(n16960), .A2(n17300), .ZN(n16956) );
  NOR2_X1 U13468 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16956), .ZN(n16942) );
  INV_X1 U13469 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17275) );
  NAND2_X1 U13470 ( .A1(n16942), .A2(n17275), .ZN(n10416) );
  NOR2_X1 U13471 ( .A1(n17258), .A2(n10416), .ZN(n11613) );
  OAI21_X1 U13472 ( .B1(n17266), .B2(n11613), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n10418) );
  NAND3_X1 U13473 ( .A1(n17247), .A2(n16982), .A3(P3_REIP_REG_24__SCAN_IN), 
        .ZN(n16974) );
  NOR2_X1 U13474 ( .A1(n10415), .A2(n16974), .ZN(n16941) );
  NAND4_X1 U13475 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16941), .ZN(n11614) );
  NAND2_X1 U13476 ( .A1(n17265), .A2(n10416), .ZN(n16937) );
  NAND3_X1 U13477 ( .A1(n10418), .A2(n10257), .A3(n10417), .ZN(n10419) );
  NOR2_X1 U13478 ( .A1(n10420), .A2(n10419), .ZN(n10421) );
  NAND2_X1 U13479 ( .A1(n10422), .A2(n10421), .ZN(P3_U2641) );
  AOI22_X1 U13480 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10428) );
  AND2_X4 U13481 ( .A1(n10645), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10644) );
  AOI22_X1 U13482 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10423) );
  AND2_X4 U13483 ( .A1(n10655), .A2(n9716), .ZN(n10639) );
  AOI22_X1 U13484 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13485 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10424) );
  AND2_X1 U13486 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NAND3_X1 U13487 ( .A1(n10428), .A2(n10427), .A3(n10426), .ZN(n10437) );
  AOI22_X1 U13488 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13489 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13490 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13491 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13492 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13493 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13494 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10440) );
  NAND3_X1 U13495 ( .A1(n10442), .A2(n10441), .A3(n10440), .ZN(n10448) );
  AOI22_X1 U13496 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13497 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13498 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__5__SCAN_IN), .B2(n10656), .ZN(n10444) );
  AOI22_X1 U13499 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10443) );
  NAND3_X1 U13500 ( .A1(n10446), .A2(n10445), .A3(n10255), .ZN(n10447) );
  INV_X1 U13501 ( .A(n10490), .ZN(n10449) );
  AOI22_X1 U13502 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n10656), .ZN(n10450) );
  AOI22_X1 U13503 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13504 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13505 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10451) );
  NAND4_X1 U13506 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10461) );
  AOI22_X1 U13507 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13508 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13509 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U13510 ( .A1(n16038), .A2(n10991), .ZN(n10952) );
  AOI22_X1 U13511 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13512 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13513 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13514 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13515 ( .A1(n9786), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10472) );
  AOI22_X1 U13516 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13517 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13518 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13519 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10468) );
  NAND2_X1 U13520 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10473) );
  AOI22_X1 U13521 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13522 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10477) );
  NAND4_X1 U13523 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10480) );
  AOI22_X1 U13524 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U13525 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10482) );
  NAND4_X1 U13526 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .ZN(
        n10485) );
  NAND2_X1 U13527 ( .A1(n10485), .A2(n10429), .ZN(n10486) );
  NAND2_X1 U13528 ( .A1(n10488), .A2(n10494), .ZN(n10492) );
  NAND2_X1 U13529 ( .A1(n10493), .A2(n10494), .ZN(n10495) );
  INV_X1 U13530 ( .A(n11249), .ZN(n10496) );
  AOI22_X1 U13531 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13532 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13533 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10498) );
  NAND4_X1 U13534 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10506) );
  AOI22_X1 U13535 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13536 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10656), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13537 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10502) );
  NAND4_X1 U13538 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10505) );
  AOI22_X1 U13539 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13540 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13541 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13542 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13543 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13544 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13545 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13546 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10512) );
  AND2_X1 U13547 ( .A1(n10991), .A2(n9736), .ZN(n11236) );
  NAND2_X1 U13548 ( .A1(n11238), .A2(n11236), .ZN(n10556) );
  NAND2_X1 U13549 ( .A1(n10556), .A2(n13873), .ZN(n10538) );
  AOI22_X1 U13550 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13551 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13552 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13553 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n10656), .ZN(n10522) );
  AOI22_X1 U13554 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13555 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13556 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10524) );
  NAND3_X1 U13557 ( .A1(n13872), .A2(n19682), .A3(n14195), .ZN(n10530) );
  AOI21_X1 U13558 ( .B1(n10544), .B2(n10991), .A(n10533), .ZN(n10531) );
  NAND2_X1 U13559 ( .A1(n10532), .A2(n10531), .ZN(n10536) );
  NOR2_X1 U13560 ( .A1(n10553), .A2(n9728), .ZN(n10535) );
  NOR2_X1 U13561 ( .A1(n13059), .A2(n10544), .ZN(n10541) );
  NOR2_X1 U13562 ( .A1(n13059), .A2(n10533), .ZN(n10539) );
  AND2_X1 U13563 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10540) );
  NOR2_X1 U13564 ( .A1(n10544), .A2(n10533), .ZN(n10547) );
  OAI22_X1 U13565 ( .A1(n9725), .A2(n21192), .B1(n13511), .B2(n20298), .ZN(
        n10548) );
  INV_X1 U13566 ( .A(n10548), .ZN(n10549) );
  NAND2_X1 U13567 ( .A1(n10550), .A2(n10549), .ZN(n10597) );
  NOR2_X1 U13568 ( .A1(n10562), .A2(n10533), .ZN(n11247) );
  NOR2_X1 U13569 ( .A1(n9728), .A2(n10449), .ZN(n10554) );
  NAND2_X1 U13570 ( .A1(n9751), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10560) );
  INV_X1 U13571 ( .A(n10555), .ZN(n10557) );
  NAND2_X1 U13572 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  NAND3_X1 U13573 ( .A1(n10560), .A2(n10559), .A3(n10558), .ZN(n10561) );
  NAND2_X1 U13574 ( .A1(n10561), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10565) );
  MUX2_X1 U13575 ( .A(n21192), .B(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .S(
        P2_STATE2_REG_1__SCAN_IN), .Z(n10563) );
  AOI21_X1 U13576 ( .B1(n10570), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10563), .ZN(
        n10564) );
  NAND2_X1 U13577 ( .A1(n13841), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10568) );
  OAI21_X1 U13578 ( .B1(n20288), .B2(n13511), .A(n10568), .ZN(n10569) );
  INV_X1 U13579 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U13580 ( .A1(n10570), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10573) );
  NAND2_X1 U13581 ( .A1(n11330), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10572) );
  NAND2_X1 U13582 ( .A1(n10601), .A2(n10604), .ZN(n10575) );
  INV_X1 U13583 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13584 ( .A1(n10570), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10579) );
  NAND2_X1 U13585 ( .A1(n11330), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10578) );
  AND3_X2 U13586 ( .A1(n10580), .A2(n10579), .A3(n10578), .ZN(n10582) );
  AOI21_X1 U13587 ( .B1(n21192), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10581) );
  XNOR2_X2 U13588 ( .A(n10582), .B(n10583), .ZN(n10595) );
  NAND2_X1 U13589 ( .A1(n10596), .A2(n10595), .ZN(n10586) );
  INV_X1 U13590 ( .A(n10582), .ZN(n10584) );
  NAND2_X1 U13591 ( .A1(n10587), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10589) );
  INV_X1 U13592 ( .A(n13511), .ZN(n11229) );
  NAND2_X1 U13593 ( .A1(n11229), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10588) );
  INV_X2 U13594 ( .A(n10590), .ZN(n11259) );
  INV_X1 U13595 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13596 ( .A1(n10570), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10593) );
  NAND2_X1 U13597 ( .A1(n11330), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10592) );
  XNOR2_X2 U13598 ( .A(n11288), .B(n11287), .ZN(n13088) );
  BUF_X4 U13599 ( .A(n13088), .Z(n10631) );
  INV_X1 U13600 ( .A(n10597), .ZN(n10600) );
  INV_X1 U13601 ( .A(n10598), .ZN(n10599) );
  NAND2_X1 U13602 ( .A1(n10600), .A2(n10599), .ZN(n10602) );
  AND2_X2 U13603 ( .A1(n10602), .A2(n10603), .ZN(n13096) );
  INV_X1 U13604 ( .A(n10604), .ZN(n10606) );
  NOR2_X1 U13605 ( .A1(n10618), .A2(n16001), .ZN(n10607) );
  INV_X1 U13606 ( .A(n10845), .ZN(n16028) );
  INV_X1 U13607 ( .A(n13096), .ZN(n13625) );
  INV_X1 U13608 ( .A(n19842), .ZN(n19836) );
  AOI22_X1 U13609 ( .A1(n16028), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n19836), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10617) );
  NOR2_X1 U13610 ( .A1(n10618), .A2(n15396), .ZN(n10608) );
  INV_X1 U13611 ( .A(n10801), .ZN(n19740) );
  AND2_X1 U13612 ( .A1(n10609), .A2(n13096), .ZN(n10623) );
  INV_X1 U13613 ( .A(n10623), .ZN(n10629) );
  INV_X1 U13614 ( .A(n19773), .ZN(n19776) );
  INV_X1 U13615 ( .A(n10609), .ZN(n10610) );
  INV_X1 U13616 ( .A(n10622), .ZN(n10611) );
  INV_X1 U13617 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10676) );
  OR3_X1 U13618 ( .A1(n10631), .A2(n9750), .A3(n10611), .ZN(n10797) );
  INV_X1 U13619 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10677) );
  INV_X1 U13620 ( .A(n10612), .ZN(n10615) );
  NAND2_X1 U13621 ( .A1(n10631), .A2(n10613), .ZN(n10628) );
  INV_X1 U13622 ( .A(n20076), .ZN(n20082) );
  NAND2_X1 U13623 ( .A1(n20082), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10614) );
  AND4_X2 U13624 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10636) );
  INV_X1 U13625 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13143) );
  INV_X1 U13626 ( .A(n10618), .ZN(n10619) );
  NAND2_X1 U13627 ( .A1(n10619), .A2(n10631), .ZN(n10620) );
  OR2_X2 U13628 ( .A1(n10620), .A2(n16001), .ZN(n19905) );
  OR2_X2 U13629 ( .A1(n10620), .A2(n15396), .ZN(n16078) );
  INV_X1 U13630 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10621) );
  INV_X1 U13631 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13632 ( .A1(n10631), .A2(n10622), .ZN(n10627) );
  OR2_X2 U13633 ( .A1(n10627), .A2(n19629), .ZN(n20042) );
  NAND2_X1 U13634 ( .A1(n10631), .A2(n10623), .ZN(n10626) );
  OR2_X2 U13635 ( .A1(n10626), .A2(n9750), .ZN(n14183) );
  INV_X1 U13636 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14200) );
  OAI22_X1 U13637 ( .A1(n10674), .A2(n20042), .B1(n14183), .B2(n14200), .ZN(
        n10624) );
  NOR2_X1 U13638 ( .A1(n10625), .A2(n10624), .ZN(n10635) );
  INV_X1 U13639 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13154) );
  OR2_X2 U13640 ( .A1(n10626), .A2(n19629), .ZN(n20123) );
  OR2_X2 U13641 ( .A1(n10627), .A2(n9750), .ZN(n19933) );
  INV_X1 U13642 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13146) );
  OAI22_X1 U13643 ( .A1(n13154), .A2(n20123), .B1(n19933), .B2(n13146), .ZN(
        n10633) );
  INV_X1 U13644 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13142) );
  INV_X1 U13645 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13153) );
  NOR2_X1 U13646 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  INV_X1 U13647 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16086) );
  OR2_X1 U13648 ( .A1(n13287), .A2(n16086), .ZN(n10643) );
  NAND2_X1 U13649 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13269) );
  INV_X1 U13650 ( .A(n13269), .ZN(n10657) );
  NAND2_X1 U13651 ( .A1(n10637), .A2(n10657), .ZN(n11036) );
  AND2_X1 U13652 ( .A1(n10638), .A2(n13268), .ZN(n10668) );
  AOI22_X1 U13653 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10642) );
  AND2_X2 U13654 ( .A1(n9715), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13295) );
  NAND2_X1 U13655 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10641) );
  AND2_X2 U13656 ( .A1(n10639), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U13657 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10640) );
  NAND4_X1 U13658 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10654) );
  INV_X1 U13659 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10649) );
  NAND2_X1 U13660 ( .A1(n13268), .A2(n10645), .ZN(n11054) );
  INV_X1 U13661 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10646) );
  OR2_X1 U13662 ( .A1(n11054), .A2(n10646), .ZN(n10648) );
  AND2_X1 U13663 ( .A1(n10637), .A2(n13268), .ZN(n10682) );
  NAND2_X1 U13664 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10647) );
  OAI211_X1 U13665 ( .C1(n11121), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        n10652) );
  NAND2_X1 U13666 ( .A1(n10644), .A2(n10429), .ZN(n10729) );
  INV_X1 U13667 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14148) );
  INV_X1 U13668 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13125) );
  OAI22_X1 U13669 ( .A1(n10729), .A2(n14148), .B1(n11074), .B2(n13125), .ZN(
        n10651) );
  OR2_X1 U13670 ( .A1(n10652), .A2(n10651), .ZN(n10653) );
  NOR2_X1 U13671 ( .A1(n10654), .A2(n10653), .ZN(n10667) );
  INV_X1 U13672 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16066) );
  INV_X1 U13673 ( .A(n10655), .ZN(n13820) );
  NAND2_X1 U13674 ( .A1(n13268), .A2(n10655), .ZN(n10669) );
  NAND2_X1 U13675 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10660) );
  NAND2_X1 U13676 ( .A1(n10965), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10774) );
  AOI22_X1 U13678 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10659) );
  OAI211_X1 U13679 ( .C1(n16066), .C2(n10669), .A(n10660), .B(n10659), .ZN(
        n10665) );
  INV_X1 U13680 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13132) );
  INV_X1 U13681 ( .A(n10663), .ZN(n13267) );
  INV_X1 U13682 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13122) );
  OAI22_X1 U13683 ( .A1(n13292), .A2(n13132), .B1(n13826), .B2(n13122), .ZN(
        n10664) );
  NOR2_X1 U13684 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  INV_X1 U13685 ( .A(n10990), .ZN(n10752) );
  NOR2_X1 U13686 ( .A1(n10752), .A2(n14195), .ZN(n13525) );
  AOI22_X1 U13687 ( .A1(n13201), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13202), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U13688 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10673) );
  INV_X2 U13689 ( .A(n10778), .ZN(n13297) );
  AOI22_X1 U13690 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10672) );
  NAND2_X1 U13691 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U13692 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10670) );
  AND4_X1 U13693 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10688) );
  OR2_X1 U13694 ( .A1(n11121), .A2(n10674), .ZN(n10675) );
  OAI21_X1 U13695 ( .B1(n10729), .B2(n10676), .A(n10675), .ZN(n10681) );
  INV_X1 U13696 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11056) );
  OR2_X1 U13697 ( .A1(n11036), .A2(n11056), .ZN(n10679) );
  OR2_X1 U13698 ( .A1(n11054), .A2(n10677), .ZN(n10678) );
  OAI211_X1 U13699 ( .C1(n11074), .C2(n13146), .A(n10679), .B(n10678), .ZN(
        n10680) );
  NOR2_X1 U13700 ( .A1(n10681), .A2(n10680), .ZN(n10687) );
  INV_X2 U13701 ( .A(n10774), .ZN(n13213) );
  AOI22_X1 U13702 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U13703 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10683) );
  OAI211_X1 U13704 ( .C1(n13292), .C2(n13153), .A(n10684), .B(n10683), .ZN(
        n10685) );
  INV_X1 U13705 ( .A(n10685), .ZN(n10686) );
  NAND2_X1 U13706 ( .A1(n13525), .A2(n11395), .ZN(n10751) );
  INV_X1 U13707 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11073) );
  OR2_X1 U13708 ( .A1(n13287), .A2(n11073), .ZN(n10693) );
  AOI22_X1 U13709 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10682), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U13710 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10691) );
  NAND2_X1 U13711 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10690) );
  NAND4_X1 U13712 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10690), .ZN(
        n10701) );
  INV_X1 U13713 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10694) );
  INV_X1 U13714 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13176) );
  OAI22_X1 U13715 ( .A1(n11121), .A2(n10694), .B1(n11074), .B2(n13176), .ZN(
        n10699) );
  INV_X1 U13716 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11072) );
  INV_X1 U13717 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10695) );
  OAI22_X1 U13718 ( .A1(n11072), .A2(n11036), .B1(n11054), .B2(n10695), .ZN(
        n10698) );
  INV_X1 U13719 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10696) );
  NOR2_X1 U13720 ( .A1(n10729), .A2(n10696), .ZN(n10697) );
  OR3_X1 U13721 ( .A1(n10699), .A2(n10698), .A3(n10697), .ZN(n10700) );
  NOR2_X1 U13722 ( .A1(n10701), .A2(n10700), .ZN(n10708) );
  INV_X1 U13723 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U13724 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10702) );
  OAI21_X1 U13725 ( .B1(n13826), .B2(n11084), .A(n10702), .ZN(n10706) );
  INV_X1 U13726 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U13727 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U13728 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10703) );
  OAI211_X1 U13729 ( .C1(n13292), .C2(n13168), .A(n10704), .B(n10703), .ZN(
        n10705) );
  NOR2_X1 U13730 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  NAND2_X1 U13731 ( .A1(n10751), .A2(n11004), .ZN(n10709) );
  INV_X1 U13732 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11106) );
  INV_X1 U13733 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13194) );
  OAI22_X1 U13734 ( .A1(n11106), .A2(n20076), .B1(n19933), .B2(n13194), .ZN(
        n10712) );
  INV_X1 U13735 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13187) );
  INV_X1 U13736 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10710) );
  OAI22_X1 U13737 ( .A1(n13187), .A2(n20123), .B1(n20042), .B2(n10710), .ZN(
        n10711) );
  NOR2_X1 U13738 ( .A1(n10712), .A2(n10711), .ZN(n10726) );
  INV_X1 U13739 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10727) );
  INV_X1 U13740 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11093) );
  OAI22_X1 U13741 ( .A1(n10727), .A2(n16078), .B1(n20010), .B2(n11093), .ZN(
        n10715) );
  INV_X1 U13742 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11103) );
  INV_X1 U13743 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10713) );
  OAI22_X1 U13744 ( .A1(n11103), .A2(n19905), .B1(n14183), .B2(n10713), .ZN(
        n10714) );
  NOR2_X1 U13745 ( .A1(n10715), .A2(n10714), .ZN(n10725) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10730) );
  INV_X1 U13747 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10716) );
  OAI22_X1 U13748 ( .A1(n10730), .A2(n14139), .B1(n19773), .B2(n10716), .ZN(
        n10718) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13186) );
  INV_X1 U13750 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10737) );
  OAI22_X1 U13751 ( .A1(n13186), .A2(n19868), .B1(n10797), .B2(n10737), .ZN(
        n10717) );
  NOR2_X1 U13752 ( .A1(n10718), .A2(n10717), .ZN(n10724) );
  INV_X1 U13753 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13093) );
  INV_X1 U13754 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11105) );
  OAI22_X1 U13755 ( .A1(n10845), .A2(n13093), .B1(n11105), .B2(n19842), .ZN(
        n10722) );
  INV_X1 U13756 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10720) );
  INV_X1 U13757 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10719) );
  OAI22_X1 U13758 ( .A1(n10801), .A2(n10720), .B1(n10719), .B2(n16055), .ZN(
        n10721) );
  NOR2_X1 U13759 ( .A1(n10722), .A2(n10721), .ZN(n10723) );
  NAND4_X1 U13760 ( .A1(n10726), .A2(n10725), .A3(n10724), .A4(n10723), .ZN(
        n10748) );
  INV_X1 U13761 ( .A(n13292), .ZN(n10767) );
  AOI22_X1 U13762 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10767), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10735) );
  OAI22_X1 U13763 ( .A1(n13287), .A2(n10727), .B1(n13826), .B2(n11103), .ZN(
        n10728) );
  INV_X1 U13764 ( .A(n10728), .ZN(n10734) );
  OAI22_X1 U13765 ( .A1(n10729), .A2(n10730), .B1(n10774), .B2(n13093), .ZN(
        n10731) );
  INV_X1 U13766 ( .A(n10731), .ZN(n10733) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n13307), .B1(
        n11095), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10732) );
  NAND4_X1 U13768 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(
        n10745) );
  NAND2_X1 U13769 ( .A1(n13288), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10736) );
  OAI21_X1 U13770 ( .B1(n11054), .B2(n10737), .A(n10736), .ZN(n10738) );
  AOI21_X1 U13771 ( .B1(n10739), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n10738), .ZN(n10743) );
  AOI22_X1 U13772 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10682), .B1(
        n13297), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13773 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10741) );
  NAND2_X1 U13774 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10740) );
  NAND4_X1 U13775 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10744) );
  INV_X1 U13776 ( .A(n11402), .ZN(n10746) );
  NAND2_X1 U13777 ( .A1(n9736), .A2(n10746), .ZN(n10747) );
  XOR2_X1 U13778 ( .A(n11004), .B(n10751), .Z(n19632) );
  INV_X1 U13779 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13532) );
  OR2_X1 U13780 ( .A1(n13525), .A2(n13532), .ZN(n13527) );
  XOR2_X1 U13781 ( .A(n10752), .B(n11395), .Z(n10753) );
  NOR2_X1 U13782 ( .A1(n13527), .A2(n10753), .ZN(n10755) );
  INV_X1 U13783 ( .A(n13527), .ZN(n10754) );
  XOR2_X1 U13784 ( .A(n10754), .B(n10753), .Z(n13562) );
  NOR2_X1 U13785 ( .A1(n16014), .A2(n13562), .ZN(n13561) );
  NOR2_X1 U13786 ( .A1(n10755), .A2(n13561), .ZN(n10756) );
  XOR2_X1 U13787 ( .A(n10756), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(
        n19631) );
  NOR2_X1 U13788 ( .A1(n19632), .A2(n19631), .ZN(n19630) );
  NOR2_X1 U13789 ( .A1(n10756), .A2(n10577), .ZN(n10757) );
  OR2_X1 U13790 ( .A1(n19630), .A2(n10757), .ZN(n10759) );
  XNOR2_X1 U13791 ( .A(n10759), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14324) );
  NAND2_X1 U13792 ( .A1(n10759), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10760) );
  NAND2_X1 U13793 ( .A1(n19618), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10786) );
  INV_X1 U13794 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10762) );
  INV_X1 U13795 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10761) );
  OAI22_X1 U13796 ( .A1(n10762), .A2(n10729), .B1(n11121), .B2(n10761), .ZN(
        n10766) );
  INV_X1 U13797 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13216) );
  NOR2_X1 U13798 ( .A1(n11074), .A2(n13216), .ZN(n10765) );
  INV_X1 U13799 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10763) );
  OAI22_X1 U13800 ( .A1(n20101), .A2(n11036), .B1(n11054), .B2(n10763), .ZN(
        n10764) );
  OR3_X1 U13801 ( .A1(n10766), .A2(n10765), .A3(n10764), .ZN(n10773) );
  NAND2_X1 U13802 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10771) );
  AOI22_X1 U13803 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10682), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U13804 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10769) );
  NAND2_X1 U13805 ( .A1(n10767), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10768) );
  NAND4_X1 U13806 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n10772) );
  NOR2_X1 U13807 ( .A1(n10773), .A2(n10772), .ZN(n10783) );
  INV_X1 U13808 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U13809 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10776) );
  AOI22_X1 U13810 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U13811 ( .C1(n10778), .C2(n10777), .A(n10776), .B(n10775), .ZN(
        n10781) );
  INV_X1 U13812 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10779) );
  INV_X1 U13813 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11129) );
  OAI22_X1 U13814 ( .A1(n13287), .A2(n10779), .B1(n13826), .B2(n11129), .ZN(
        n10780) );
  NOR2_X1 U13815 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  INV_X1 U13816 ( .A(n11422), .ZN(n11016) );
  NAND2_X1 U13817 ( .A1(n10784), .A2(n11422), .ZN(n10785) );
  NAND2_X1 U13818 ( .A1(n10833), .A2(n10785), .ZN(n19616) );
  NAND2_X1 U13819 ( .A1(n10786), .A2(n19616), .ZN(n10790) );
  INV_X1 U13820 ( .A(n19618), .ZN(n10788) );
  INV_X1 U13821 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13822 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  INV_X1 U13823 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13222) );
  INV_X1 U13824 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10791) );
  OAI22_X1 U13825 ( .A1(n13222), .A2(n19905), .B1(n16078), .B2(n10791), .ZN(
        n10794) );
  INV_X1 U13826 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10792) );
  INV_X1 U13827 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13226) );
  OAI22_X1 U13828 ( .A1(n10792), .A2(n14183), .B1(n19933), .B2(n13226), .ZN(
        n10793) );
  NOR2_X1 U13829 ( .A1(n10794), .A2(n10793), .ZN(n10809) );
  INV_X1 U13830 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11143) );
  INV_X1 U13831 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10814) );
  OAI22_X1 U13832 ( .A1(n11143), .A2(n20076), .B1(n20042), .B2(n10814), .ZN(
        n10796) );
  INV_X1 U13833 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13234) );
  INV_X1 U13834 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13223) );
  OAI22_X1 U13835 ( .A1(n13234), .A2(n20123), .B1(n20010), .B2(n13223), .ZN(
        n10795) );
  NOR2_X1 U13836 ( .A1(n10796), .A2(n10795), .ZN(n10808) );
  INV_X1 U13837 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13233) );
  INV_X1 U13838 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10817) );
  OAI22_X1 U13839 ( .A1(n13233), .A2(n19868), .B1(n10797), .B2(n10817), .ZN(
        n10800) );
  INV_X1 U13840 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10816) );
  INV_X1 U13841 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10798) );
  OAI22_X1 U13842 ( .A1(n10816), .A2(n14139), .B1(n19773), .B2(n10798), .ZN(
        n10799) );
  NOR2_X1 U13843 ( .A1(n10800), .A2(n10799), .ZN(n10807) );
  INV_X1 U13844 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13908) );
  INV_X1 U13845 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11142) );
  OAI22_X1 U13846 ( .A1(n10845), .A2(n13908), .B1(n11142), .B2(n19842), .ZN(
        n10805) );
  INV_X1 U13847 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10803) );
  INV_X1 U13848 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10802) );
  OAI22_X1 U13849 ( .A1(n10801), .A2(n10803), .B1(n10802), .B2(n16055), .ZN(
        n10804) );
  NOR2_X1 U13850 ( .A1(n10805), .A2(n10804), .ZN(n10806) );
  NAND4_X1 U13851 ( .A1(n10809), .A2(n10808), .A3(n10807), .A4(n10806), .ZN(
        n10831) );
  AOI22_X1 U13852 ( .A1(n13201), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13202), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13853 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10813) );
  AOI22_X1 U13854 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13855 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10811) );
  NAND2_X1 U13856 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10810) );
  AND4_X1 U13857 ( .A1(n10813), .A2(n10812), .A3(n10811), .A4(n10810), .ZN(
        n10827) );
  OR2_X1 U13858 ( .A1(n11121), .A2(n10814), .ZN(n10815) );
  OAI21_X1 U13859 ( .B1(n10729), .B2(n10816), .A(n10815), .ZN(n10821) );
  OR2_X1 U13860 ( .A1(n11036), .A2(n11143), .ZN(n10819) );
  OR2_X1 U13861 ( .A1(n11054), .A2(n10817), .ZN(n10818) );
  OAI211_X1 U13862 ( .C1(n11074), .C2(n13226), .A(n10819), .B(n10818), .ZN(
        n10820) );
  NOR2_X1 U13863 ( .A1(n10821), .A2(n10820), .ZN(n10826) );
  AOI22_X1 U13864 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13865 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10822) );
  OAI211_X1 U13866 ( .C1(n13233), .C2(n13292), .A(n10823), .B(n10822), .ZN(
        n10824) );
  INV_X1 U13867 ( .A(n10824), .ZN(n10825) );
  NAND4_X1 U13868 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n11429) );
  INV_X1 U13869 ( .A(n11429), .ZN(n10829) );
  NAND2_X1 U13870 ( .A1(n9736), .A2(n10829), .ZN(n10830) );
  INV_X1 U13871 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10858) );
  INV_X1 U13872 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13257) );
  OAI22_X1 U13873 ( .A1(n10858), .A2(n16078), .B1(n20123), .B2(n13257), .ZN(
        n10838) );
  INV_X1 U13874 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13245) );
  INV_X1 U13875 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10836) );
  OAI22_X1 U13876 ( .A1(n13245), .A2(n20010), .B1(n14183), .B2(n10836), .ZN(
        n10837) );
  NOR2_X1 U13877 ( .A1(n10838), .A2(n10837), .ZN(n10851) );
  INV_X1 U13878 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13244) );
  INV_X1 U13879 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13249) );
  OAI22_X1 U13880 ( .A1(n13244), .A2(n19905), .B1(n19933), .B2(n13249), .ZN(
        n10840) );
  INV_X1 U13881 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11161) );
  INV_X1 U13882 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10852) );
  OAI22_X1 U13883 ( .A1(n11161), .A2(n20076), .B1(n20042), .B2(n10852), .ZN(
        n10839) );
  NOR2_X1 U13884 ( .A1(n10840), .A2(n10839), .ZN(n10850) );
  INV_X1 U13885 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13256) );
  INV_X1 U13886 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10854) );
  OAI22_X1 U13887 ( .A1(n13256), .A2(n19868), .B1(n10797), .B2(n10854), .ZN(
        n10843) );
  INV_X1 U13888 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10841) );
  INV_X1 U13889 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10853) );
  OAI22_X1 U13890 ( .A1(n10841), .A2(n19773), .B1(n14139), .B2(n10853), .ZN(
        n10842) );
  NOR2_X1 U13891 ( .A1(n10843), .A2(n10842), .ZN(n10849) );
  INV_X1 U13892 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16045) );
  INV_X1 U13893 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10844) );
  OAI22_X1 U13894 ( .A1(n16045), .A2(n10845), .B1(n10801), .B2(n10844), .ZN(
        n10847) );
  INV_X1 U13895 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11162) );
  INV_X1 U13896 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16074) );
  OAI22_X1 U13897 ( .A1(n11162), .A2(n19842), .B1(n16055), .B2(n16074), .ZN(
        n10846) );
  NOR2_X1 U13898 ( .A1(n10847), .A2(n10846), .ZN(n10848) );
  NAND4_X1 U13899 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n10873) );
  OAI22_X1 U13900 ( .A1(n10853), .A2(n10729), .B1(n11121), .B2(n10852), .ZN(
        n10857) );
  NOR2_X1 U13901 ( .A1(n11074), .A2(n13249), .ZN(n10856) );
  OAI22_X1 U13902 ( .A1(n11161), .A2(n11036), .B1(n11054), .B2(n10854), .ZN(
        n10855) );
  OR2_X1 U13903 ( .A1(n13287), .A2(n10858), .ZN(n10862) );
  AOI22_X1 U13904 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10682), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U13905 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10860) );
  NAND2_X1 U13906 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10859) );
  NAND4_X1 U13907 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(
        n10863) );
  NOR2_X1 U13908 ( .A1(n10864), .A2(n10863), .ZN(n10871) );
  NAND2_X1 U13909 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10865) );
  OAI21_X1 U13910 ( .B1(n13826), .B2(n13244), .A(n10865), .ZN(n10869) );
  AOI22_X1 U13911 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10867) );
  NAND2_X1 U13912 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10866) );
  OAI211_X1 U13913 ( .C1(n13292), .C2(n13256), .A(n10867), .B(n10866), .ZN(
        n10868) );
  NOR2_X1 U13914 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  NAND2_X1 U13915 ( .A1(n11437), .A2(n9736), .ZN(n10872) );
  NAND2_X1 U13916 ( .A1(n10875), .A2(n11434), .ZN(n10876) );
  NAND2_X1 U13917 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10883) );
  AOI22_X1 U13918 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10682), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U13919 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10881) );
  NAND2_X1 U13920 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10880) );
  INV_X1 U13921 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10886) );
  INV_X1 U13922 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10884) );
  OR2_X1 U13923 ( .A1(n11121), .A2(n10884), .ZN(n10885) );
  OAI21_X1 U13924 ( .B1(n10729), .B2(n10886), .A(n10885), .ZN(n10890) );
  INV_X1 U13925 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13291) );
  INV_X1 U13926 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20114) );
  OR2_X1 U13927 ( .A1(n11036), .A2(n20114), .ZN(n10888) );
  INV_X1 U13928 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13452) );
  OR2_X1 U13929 ( .A1(n11054), .A2(n13452), .ZN(n10887) );
  OAI211_X1 U13930 ( .C1(n11074), .C2(n13291), .A(n10888), .B(n10887), .ZN(
        n10889) );
  NOR2_X1 U13931 ( .A1(n10890), .A2(n10889), .ZN(n10898) );
  NAND2_X1 U13932 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10892) );
  INV_X1 U13933 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13445) );
  OR2_X1 U13934 ( .A1(n13287), .A2(n13445), .ZN(n10891) );
  AND2_X1 U13935 ( .A1(n10892), .A2(n10891), .ZN(n10897) );
  INV_X1 U13936 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U13937 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U13938 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10893) );
  OAI211_X1 U13939 ( .C1(n13292), .C2(n13305), .A(n10894), .B(n10893), .ZN(
        n10895) );
  INV_X1 U13940 ( .A(n10895), .ZN(n10896) );
  XNOR2_X1 U13941 ( .A(n10905), .B(n11444), .ZN(n10899) );
  NAND2_X1 U13942 ( .A1(n15752), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10903) );
  INV_X1 U13943 ( .A(n10899), .ZN(n10900) );
  NAND2_X1 U13944 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  NOR2_X1 U13945 ( .A1(n10905), .A2(n11444), .ZN(n10904) );
  INV_X1 U13946 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11449) );
  XNOR2_X1 U13947 ( .A(n10904), .B(n11449), .ZN(n16624) );
  INV_X1 U13948 ( .A(n10905), .ZN(n10906) );
  NAND3_X1 U13949 ( .A1(n10906), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11584), .ZN(n10907) );
  NAND2_X1 U13950 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16684) );
  NOR2_X1 U13951 ( .A1(n11274), .A2(n16684), .ZN(n15937) );
  INV_X1 U13952 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11266) );
  NAND2_X1 U13953 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16656) );
  NOR2_X1 U13954 ( .A1(n11266), .A2(n16656), .ZN(n15886) );
  NAND2_X1 U13955 ( .A1(n15937), .A2(n15886), .ZN(n16114) );
  NAND3_X1 U13956 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15917) );
  NOR2_X1 U13957 ( .A1(n16114), .A2(n15917), .ZN(n15885) );
  AND2_X1 U13958 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15885), .ZN(
        n15887) );
  INV_X1 U13959 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15881) );
  INV_X1 U13960 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15853) );
  INV_X1 U13961 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15644) );
  NAND2_X1 U13962 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15812) );
  INV_X1 U13963 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15589) );
  XNOR2_X2 U13964 ( .A(n10909), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12995) );
  NAND2_X1 U13965 ( .A1(n19539), .A2(n14195), .ZN(n10912) );
  XNOR2_X1 U13966 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U13967 ( .A1(n10915), .A2(n10913), .ZN(n10917) );
  NAND2_X1 U13968 ( .A1(n20288), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10910) );
  NAND2_X1 U13969 ( .A1(n10917), .A2(n10910), .ZN(n10927) );
  XNOR2_X1 U13970 ( .A(n13819), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10911) );
  XNOR2_X1 U13971 ( .A(n10927), .B(n10911), .ZN(n10946) );
  MUX2_X1 U13972 ( .A(n10912), .B(n13059), .S(n10946), .Z(n10925) );
  INV_X1 U13973 ( .A(n10946), .ZN(n10960) );
  INV_X1 U13974 ( .A(n10913), .ZN(n10916) );
  NAND2_X1 U13975 ( .A1(n13848), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10914) );
  NAND2_X1 U13976 ( .A1(n10916), .A2(n10914), .ZN(n10969) );
  INV_X1 U13977 ( .A(n10969), .ZN(n10958) );
  INV_X1 U13978 ( .A(n10915), .ZN(n10921) );
  NAND2_X1 U13979 ( .A1(n10921), .A2(n10916), .ZN(n10959) );
  NAND2_X1 U13980 ( .A1(n10959), .A2(n10917), .ZN(n10947) );
  INV_X1 U13981 ( .A(n10947), .ZN(n10918) );
  OAI21_X1 U13982 ( .B1(n14195), .B2(n10958), .A(n10918), .ZN(n10919) );
  OAI21_X1 U13983 ( .B1(n14195), .B2(n10960), .A(n10919), .ZN(n10920) );
  NAND2_X1 U13984 ( .A1(n10920), .A2(n13873), .ZN(n10923) );
  OAI21_X1 U13985 ( .B1(n10921), .B2(n10969), .A(n10027), .ZN(n10922) );
  NAND2_X1 U13986 ( .A1(n10923), .A2(n10922), .ZN(n10924) );
  NAND2_X1 U13987 ( .A1(n10925), .A2(n10924), .ZN(n10934) );
  MUX2_X1 U13988 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n21171), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10931) );
  NAND2_X1 U13989 ( .A1(n21171), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10928) );
  NOR2_X1 U13990 ( .A1(n16203), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10930) );
  NAND2_X1 U13991 ( .A1(n10936), .A2(n10930), .ZN(n11420) );
  INV_X1 U13992 ( .A(n10931), .ZN(n10932) );
  XNOR2_X1 U13993 ( .A(n10933), .B(n10932), .ZN(n11399) );
  MUX2_X1 U13994 ( .A(n13059), .B(n10934), .S(n10962), .Z(n10939) );
  NAND2_X1 U13995 ( .A1(n16203), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U13996 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13552), .ZN(
        n10937) );
  NAND2_X1 U13997 ( .A1(n10939), .A2(n20304), .ZN(n10940) );
  MUX2_X1 U13998 ( .A(n10940), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21192), .Z(n10943) );
  NAND2_X1 U13999 ( .A1(n13868), .A2(n14195), .ZN(n19536) );
  INV_X1 U14000 ( .A(n10943), .ZN(n10945) );
  INV_X1 U14001 ( .A(n13868), .ZN(n10944) );
  AOI22_X1 U14002 ( .A1(n19536), .A2(n10945), .B1(n10944), .B2(n9728), .ZN(
        n10980) );
  INV_X1 U14003 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20189) );
  INV_X1 U14004 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20182) );
  NAND2_X2 U14005 ( .A1(n20314), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20247) );
  NAND2_X1 U14006 ( .A1(n20182), .A2(n20200), .ZN(n20194) );
  NAND2_X1 U14007 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20183) );
  NAND2_X1 U14008 ( .A1(n20188), .A2(n20183), .ZN(n13538) );
  OR3_X1 U14009 ( .A1(n19536), .A2(n19682), .A3(n13538), .ZN(n10979) );
  NAND2_X1 U14010 ( .A1(n9728), .A2(n9736), .ZN(n13062) );
  AOI21_X1 U14011 ( .B1(n10950), .B2(n10527), .A(n13062), .ZN(n11232) );
  INV_X1 U14012 ( .A(n11232), .ZN(n11235) );
  NAND2_X1 U14013 ( .A1(n10946), .A2(n10962), .ZN(n10968) );
  OR2_X1 U14014 ( .A1(n10947), .A2(n10968), .ZN(n10948) );
  INV_X1 U14015 ( .A(n13538), .ZN(n13061) );
  NAND3_X1 U14016 ( .A1(n10552), .A2(n13862), .A3(n13061), .ZN(n10949) );
  OAI211_X1 U14017 ( .C1(n10950), .C2(n16038), .A(n11235), .B(n10949), .ZN(
        n10957) );
  NAND2_X1 U14018 ( .A1(n10952), .A2(n19682), .ZN(n10953) );
  NAND2_X1 U14019 ( .A1(n10951), .A2(n10953), .ZN(n10956) );
  NOR2_X1 U14020 ( .A1(n11245), .A2(n14195), .ZN(n11230) );
  OAI211_X1 U14021 ( .C1(n11230), .C2(n9728), .A(n10544), .B(n10527), .ZN(
        n10954) );
  NAND2_X1 U14022 ( .A1(n10954), .A2(n19682), .ZN(n10955) );
  NAND2_X1 U14023 ( .A1(n10956), .A2(n10955), .ZN(n11233) );
  NOR2_X1 U14024 ( .A1(n10957), .A2(n11233), .ZN(n13542) );
  MUX2_X1 U14025 ( .A(n10990), .B(n10958), .S(n13059), .Z(n11407) );
  NAND2_X1 U14026 ( .A1(n11407), .A2(n10959), .ZN(n10961) );
  NAND2_X1 U14027 ( .A1(n10961), .A2(n11394), .ZN(n10963) );
  NAND2_X1 U14028 ( .A1(n10963), .A2(n10962), .ZN(n20305) );
  NOR2_X1 U14029 ( .A1(n20303), .A2(n10964), .ZN(n10974) );
  NOR2_X1 U14030 ( .A1(n10965), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13548) );
  NAND2_X1 U14031 ( .A1(n13548), .A2(n11036), .ZN(n10967) );
  INV_X1 U14032 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n16202) );
  AND2_X1 U14033 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16202), .ZN(n10966) );
  NAND2_X1 U14034 ( .A1(n10967), .A2(n10966), .ZN(n20294) );
  OAI21_X1 U14035 ( .B1(n10969), .B2(n10968), .A(n13862), .ZN(n10970) );
  NAND2_X1 U14036 ( .A1(n10591), .A2(n10970), .ZN(n10971) );
  NAND2_X1 U14037 ( .A1(n14195), .A2(n20302), .ZN(n10972) );
  NOR2_X1 U14038 ( .A1(n13872), .A2(n10972), .ZN(n10973) );
  AOI21_X1 U14039 ( .B1(n20305), .B2(n10974), .A(n10973), .ZN(n12994) );
  NAND2_X1 U14040 ( .A1(n10551), .A2(n14195), .ZN(n10976) );
  INV_X1 U14041 ( .A(n11247), .ZN(n10975) );
  NAND4_X1 U14042 ( .A1(n10976), .A2(n13862), .A3(n20183), .A4(n10975), .ZN(
        n10977) );
  AND3_X1 U14043 ( .A1(n13542), .A2(n12994), .A3(n10977), .ZN(n10978) );
  OAI211_X1 U14044 ( .C1(n10980), .C2(n11245), .A(n10979), .B(n10978), .ZN(
        n10982) );
  INV_X1 U14045 ( .A(n20303), .ZN(n10983) );
  NAND2_X1 U14046 ( .A1(n12995), .A2(n19660), .ZN(n11393) );
  AND2_X2 U14047 ( .A1(n10996), .A2(n10984), .ZN(n11005) );
  NAND2_X1 U14048 ( .A1(n11005), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10988) );
  AOI21_X1 U14049 ( .B1(n14195), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U14050 ( .A1(n19696), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10985) );
  AND2_X1 U14051 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  NAND2_X1 U14052 ( .A1(n10988), .A2(n10987), .ZN(n13580) );
  AND2_X1 U14053 ( .A1(n20298), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20289) );
  NAND2_X1 U14054 ( .A1(n11195), .A2(n10990), .ZN(n10993) );
  INV_X1 U14055 ( .A(n10991), .ZN(n10992) );
  AND2_X2 U14056 ( .A1(n14195), .A2(n19936), .ZN(n11006) );
  NAND2_X1 U14057 ( .A1(n10992), .A2(n11006), .ZN(n11002) );
  OAI211_X1 U14058 ( .C1(n10996), .C2(n20289), .A(n10993), .B(n11002), .ZN(
        n13579) );
  INV_X1 U14059 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20202) );
  NAND2_X1 U14060 ( .A1(n11005), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10995) );
  AND2_X2 U14061 ( .A1(n19696), .A2(n19936), .ZN(n11210) );
  AOI22_X1 U14062 ( .A1(n11210), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U14063 ( .A1(n10995), .A2(n10994), .ZN(n10999) );
  XNOR2_X1 U14064 ( .A(n13582), .B(n10999), .ZN(n15389) );
  NAND2_X1 U14065 ( .A1(n11195), .A2(n11395), .ZN(n10998) );
  NAND2_X1 U14066 ( .A1(n10996), .A2(n10991), .ZN(n10997) );
  OAI211_X1 U14067 ( .C1(n19936), .C2(n20288), .A(n10998), .B(n10997), .ZN(
        n15388) );
  NOR2_X1 U14068 ( .A1(n15389), .A2(n15388), .ZN(n11001) );
  NOR2_X1 U14069 ( .A1(n13582), .A2(n10999), .ZN(n11000) );
  INV_X1 U14070 ( .A(n11195), .ZN(n11091) );
  NAND2_X1 U14071 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11003) );
  OAI211_X1 U14072 ( .C1(n11091), .C2(n11004), .A(n11003), .B(n11002), .ZN(
        n11009) );
  XNOR2_X1 U14073 ( .A(n11010), .B(n11009), .ZN(n14560) );
  NAND2_X1 U14074 ( .A1(n11005), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14075 ( .A1(n11210), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U14076 ( .A1(n11008), .A2(n11007), .ZN(n14559) );
  NOR2_X1 U14077 ( .A1(n14560), .A2(n14559), .ZN(n14558) );
  NOR2_X1 U14078 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  NAND2_X1 U14079 ( .A1(n11005), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14080 ( .A1(n11006), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11014) );
  NAND2_X1 U14081 ( .A1(n11195), .A2(n11402), .ZN(n11013) );
  NAND2_X1 U14082 ( .A1(n11210), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11012) );
  NAND4_X1 U14083 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n14327) );
  NAND2_X1 U14084 ( .A1(n11005), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14085 ( .A1(n11210), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U14086 ( .A1(n11195), .A2(n11016), .ZN(n11017) );
  AOI22_X1 U14087 ( .A1(n11005), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11195), 
        .B2(n11429), .ZN(n11021) );
  AOI22_X1 U14088 ( .A1(n11210), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11020) );
  NAND2_X1 U14089 ( .A1(n11021), .A2(n11020), .ZN(n15979) );
  INV_X1 U14090 ( .A(n11437), .ZN(n11022) );
  NAND2_X1 U14091 ( .A1(n11195), .A2(n11022), .ZN(n11023) );
  NAND2_X1 U14092 ( .A1(n15978), .A2(n11023), .ZN(n15969) );
  NAND2_X1 U14093 ( .A1(n11005), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U14094 ( .A1(n11210), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U14095 ( .A1(n11025), .A2(n11024), .ZN(n15968) );
  NAND2_X1 U14096 ( .A1(n15969), .A2(n15968), .ZN(n11027) );
  INV_X2 U14097 ( .A(n11444), .ZN(n11584) );
  NAND2_X1 U14098 ( .A1(n11195), .A2(n11584), .ZN(n11026) );
  NAND2_X1 U14099 ( .A1(n11027), .A2(n11026), .ZN(n15958) );
  NAND2_X1 U14100 ( .A1(n11005), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14101 ( .A1(n11210), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U14102 ( .A1(n11029), .A2(n11028), .ZN(n15957) );
  NAND2_X1 U14103 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11033) );
  NAND2_X1 U14104 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11032) );
  AOI22_X1 U14105 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11031) );
  NAND2_X1 U14106 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11030) );
  NAND4_X1 U14107 ( .A1(n11033), .A2(n11032), .A3(n11031), .A4(n11030), .ZN(
        n11041) );
  INV_X1 U14108 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11034) );
  OAI22_X1 U14109 ( .A1(n10729), .A2(n11034), .B1(n11074), .B2(n16086), .ZN(
        n11039) );
  INV_X1 U14110 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13133) );
  INV_X1 U14111 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11035) );
  OAI22_X1 U14112 ( .A1(n11036), .A2(n13133), .B1(n11054), .B2(n11035), .ZN(
        n11038) );
  INV_X1 U14113 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20088) );
  NOR2_X1 U14114 ( .A1(n11121), .A2(n20088), .ZN(n11037) );
  OR3_X1 U14115 ( .A1(n11039), .A2(n11038), .A3(n11037), .ZN(n11040) );
  NOR2_X1 U14116 ( .A1(n11041), .A2(n11040), .ZN(n11047) );
  INV_X1 U14117 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14193) );
  OAI22_X1 U14118 ( .A1(n13287), .A2(n14193), .B1(n13826), .B2(n13125), .ZN(
        n11045) );
  AOI22_X1 U14119 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14120 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11042) );
  OAI211_X1 U14121 ( .C1(n13122), .C2(n13292), .A(n11043), .B(n11042), .ZN(
        n11044) );
  NOR2_X1 U14122 ( .A1(n11045), .A2(n11044), .ZN(n11046) );
  AOI22_X1 U14123 ( .A1(n11210), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11048) );
  OAI21_X1 U14124 ( .B1(n11091), .B2(n13985), .A(n11048), .ZN(n11049) );
  AOI21_X1 U14125 ( .B1(n11005), .B2(P2_REIP_REG_8__SCAN_IN), .A(n11049), .ZN(
        n16706) );
  AOI22_X1 U14126 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U14127 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11053) );
  AOI22_X1 U14128 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U14129 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11051) );
  NAND2_X1 U14130 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11050) );
  AND4_X1 U14131 ( .A1(n11053), .A2(n11052), .A3(n11051), .A4(n11050), .ZN(
        n11066) );
  AOI22_X1 U14132 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11060) );
  INV_X1 U14133 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11055) );
  OR2_X1 U14134 ( .A1(n10729), .A2(n11055), .ZN(n11059) );
  OR2_X1 U14135 ( .A1(n11121), .A2(n11056), .ZN(n11058) );
  NAND2_X1 U14136 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11057) );
  AND4_X1 U14137 ( .A1(n11060), .A2(n11059), .A3(n11058), .A4(n11057), .ZN(
        n11065) );
  AOI22_X1 U14138 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14139 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11061) );
  OAI211_X1 U14140 ( .C1(n13292), .C2(n13143), .A(n11062), .B(n11061), .ZN(
        n11063) );
  INV_X1 U14141 ( .A(n11063), .ZN(n11064) );
  NAND4_X1 U14142 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n13991) );
  AOI22_X1 U14143 ( .A1(n11005), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11195), 
        .B2(n13991), .ZN(n11069) );
  AOI22_X1 U14144 ( .A1(n11210), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11006), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11068) );
  NAND2_X1 U14145 ( .A1(n11069), .A2(n11068), .ZN(n15948) );
  AOI22_X1 U14146 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11089) );
  NAND2_X1 U14147 ( .A1(n13303), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U14148 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11070) );
  OAI211_X1 U14149 ( .C1(n11121), .C2(n11072), .A(n11071), .B(n11070), .ZN(
        n11077) );
  INV_X1 U14150 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11075) );
  OAI22_X1 U14151 ( .A1(n10729), .A2(n11075), .B1(n11074), .B2(n11073), .ZN(
        n11076) );
  NOR2_X1 U14152 ( .A1(n11077), .A2(n11076), .ZN(n11088) );
  NAND2_X1 U14153 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11081) );
  AOI22_X1 U14154 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11080) );
  NAND2_X1 U14155 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11079) );
  NAND2_X1 U14156 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11078) );
  AND4_X1 U14157 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11087) );
  AOI22_X1 U14158 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14159 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11082) );
  OAI211_X1 U14160 ( .C1(n13292), .C2(n11084), .A(n11083), .B(n11082), .ZN(
        n11085) );
  INV_X1 U14161 ( .A(n11085), .ZN(n11086) );
  NAND4_X1 U14162 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n13118) );
  INV_X1 U14163 ( .A(n13118), .ZN(n14115) );
  AOI22_X1 U14164 ( .A1(n11210), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11090) );
  OAI21_X1 U14165 ( .B1(n11091), .B2(n14115), .A(n11090), .ZN(n11092) );
  AOI21_X1 U14166 ( .B1(n11005), .B2(P2_REIP_REG_10__SCAN_IN), .A(n11092), 
        .ZN(n16693) );
  AOI22_X1 U14167 ( .A1(n11005), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14168 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11114) );
  INV_X1 U14169 ( .A(n13295), .ZN(n11094) );
  OAI22_X1 U14170 ( .A1(n11094), .A2(n11093), .B1(n13826), .B2(n13194), .ZN(
        n11100) );
  INV_X1 U14171 ( .A(n11095), .ZN(n11098) );
  NAND2_X1 U14172 ( .A1(n13296), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14173 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11096) );
  OAI211_X1 U14174 ( .C1(n11098), .C2(n10710), .A(n11097), .B(n11096), .ZN(
        n11099) );
  NOR2_X1 U14175 ( .A1(n11100), .A2(n11099), .ZN(n11113) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U14177 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11101) );
  OAI211_X1 U14178 ( .C1(n13292), .C2(n11103), .A(n11102), .B(n11101), .ZN(
        n11104) );
  INV_X1 U14179 ( .A(n11104), .ZN(n11112) );
  AOI22_X1 U14180 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11110) );
  OR2_X1 U14181 ( .A1(n10729), .A2(n11105), .ZN(n11109) );
  OR2_X1 U14182 ( .A1(n11121), .A2(n11106), .ZN(n11108) );
  NAND2_X1 U14183 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11107) );
  AND4_X1 U14184 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n11111) );
  NAND4_X1 U14185 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n14226) );
  AOI22_X1 U14186 ( .A1(n11195), .A2(n14226), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n11210), .ZN(n11115) );
  NAND2_X1 U14187 ( .A1(n11116), .A2(n11115), .ZN(n15378) );
  NAND2_X1 U14188 ( .A1(n11005), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U14189 ( .A1(n11210), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14190 ( .A1(n13201), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U14191 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11119) );
  AOI22_X1 U14192 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10682), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U14193 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11117) );
  AND4_X1 U14194 ( .A1(n11120), .A2(n11119), .A3(n11118), .A4(n11117), .ZN(
        n11134) );
  AOI22_X1 U14195 ( .A1(n13202), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13298), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14196 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11126) );
  OR2_X1 U14197 ( .A1(n11121), .A2(n20101), .ZN(n11125) );
  INV_X1 U14198 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11122) );
  OR2_X1 U14199 ( .A1(n10729), .A2(n11122), .ZN(n11124) );
  NAND2_X1 U14200 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11123) );
  AND4_X1 U14201 ( .A1(n11126), .A2(n11125), .A3(n11124), .A4(n11123), .ZN(
        n11132) );
  AOI22_X1 U14202 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U14203 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11127) );
  OAI211_X1 U14204 ( .C1(n13292), .C2(n11129), .A(n11128), .B(n11127), .ZN(
        n11130) );
  INV_X1 U14205 ( .A(n11130), .ZN(n11131) );
  NAND4_X1 U14206 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n14225) );
  NAND2_X1 U14207 ( .A1(n11195), .A2(n14225), .ZN(n11135) );
  AOI22_X1 U14208 ( .A1(n11005), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11156) );
  AOI22_X1 U14209 ( .A1(n13201), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13202), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U14210 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11141) );
  AOI22_X1 U14211 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U14212 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14213 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11138) );
  AND4_X1 U14214 ( .A1(n11141), .A2(n11140), .A3(n11139), .A4(n11138), .ZN(
        n11153) );
  AOI22_X1 U14215 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11147) );
  OR2_X1 U14216 ( .A1(n10729), .A2(n11142), .ZN(n11146) );
  OR2_X1 U14217 ( .A1(n11121), .A2(n11143), .ZN(n11145) );
  NAND2_X1 U14218 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11144) );
  AND4_X1 U14219 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11152) );
  AOI22_X1 U14220 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U14221 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11148) );
  OAI211_X1 U14222 ( .C1(n13222), .C2(n13292), .A(n11149), .B(n11148), .ZN(
        n11150) );
  INV_X1 U14223 ( .A(n11150), .ZN(n11151) );
  NAND4_X1 U14224 ( .A1(n11154), .A2(n11153), .A3(n11152), .A4(n11151), .ZN(
        n14239) );
  AOI22_X1 U14225 ( .A1(n11195), .A2(n14239), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n11210), .ZN(n11155) );
  NAND2_X1 U14226 ( .A1(n11156), .A2(n11155), .ZN(n16671) );
  NAND2_X1 U14227 ( .A1(n11005), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14228 ( .A1(n11210), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11175) );
  AOI22_X1 U14229 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U14230 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11160) );
  AOI22_X1 U14231 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10682), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14232 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11158) );
  NAND2_X1 U14233 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11157) );
  AND4_X1 U14234 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n11157), .ZN(
        n11172) );
  AOI22_X1 U14235 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11166) );
  OR2_X1 U14236 ( .A1(n11121), .A2(n11161), .ZN(n11165) );
  OR2_X1 U14237 ( .A1(n10729), .A2(n11162), .ZN(n11164) );
  NAND2_X1 U14238 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11163) );
  AND4_X1 U14239 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n11171) );
  AOI22_X1 U14240 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11168) );
  NAND2_X1 U14241 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11167) );
  OAI211_X1 U14242 ( .C1(n13292), .C2(n13244), .A(n11168), .B(n11167), .ZN(
        n11169) );
  INV_X1 U14243 ( .A(n11169), .ZN(n11170) );
  NAND4_X1 U14244 ( .A1(n11173), .A2(n11172), .A3(n11171), .A4(n11170), .ZN(
        n14242) );
  NAND2_X1 U14245 ( .A1(n11195), .A2(n14242), .ZN(n11174) );
  AOI22_X1 U14246 ( .A1(n11005), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11197) );
  INV_X1 U14247 ( .A(n13202), .ZN(n13286) );
  INV_X1 U14248 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11177) );
  OAI22_X1 U14249 ( .A1(n13305), .A2(n13286), .B1(n13287), .B2(n11177), .ZN(
        n11181) );
  INV_X1 U14250 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13285) );
  INV_X1 U14251 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19706) );
  AOI22_X1 U14252 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11179) );
  NAND2_X1 U14253 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11178) );
  OAI211_X1 U14254 ( .C1(n13292), .C2(n13285), .A(n11179), .B(n11178), .ZN(
        n11180) );
  NOR2_X1 U14255 ( .A1(n11181), .A2(n11180), .ZN(n11194) );
  NAND2_X1 U14256 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11185) );
  AOI22_X1 U14257 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U14258 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U14259 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11182) );
  NAND4_X1 U14260 ( .A1(n11185), .A2(n11184), .A3(n11183), .A4(n11182), .ZN(
        n11192) );
  AOI22_X1 U14261 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11190) );
  INV_X1 U14262 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11186) );
  OR2_X1 U14263 ( .A1(n10729), .A2(n11186), .ZN(n11189) );
  OR2_X1 U14264 ( .A1(n11121), .A2(n20114), .ZN(n11188) );
  NAND2_X1 U14265 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11187) );
  NAND4_X1 U14266 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11191) );
  NOR2_X1 U14267 ( .A1(n11192), .A2(n11191), .ZN(n11193) );
  AOI22_X1 U14268 ( .A1(n11195), .A2(n13120), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n11210), .ZN(n11196) );
  NAND2_X1 U14269 ( .A1(n11197), .A2(n11196), .ZN(n16645) );
  AOI222_X1 U14270 ( .A1(n11005), .A2(P2_REIP_REG_16__SCAN_IN), .B1(n11210), 
        .B2(P2_EAX_REG_16__SCAN_IN), .C1(n11006), .C2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16111) );
  NAND2_X1 U14271 ( .A1(n11005), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14272 ( .A1(n11210), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U14273 ( .A1(n11199), .A2(n11198), .ZN(n15572) );
  NAND2_X1 U14274 ( .A1(n11005), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14275 ( .A1(n11210), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U14276 ( .A1(n11201), .A2(n11200), .ZN(n15561) );
  NAND2_X1 U14277 ( .A1(n11005), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14278 ( .A1(n11210), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U14279 ( .A1(n11005), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14280 ( .A1(n11210), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11204) );
  NAND2_X1 U14281 ( .A1(n11005), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14282 ( .A1(n11210), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14283 ( .A1(n11207), .A2(n11206), .ZN(n13497) );
  AOI222_X1 U14284 ( .A1(n11005), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n11210), 
        .B2(P2_EAX_REG_22__SCAN_IN), .C1(n11006), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15861) );
  NAND2_X1 U14285 ( .A1(n11005), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14286 ( .A1(n11210), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14287 ( .A1(n11209), .A2(n11208), .ZN(n15354) );
  INV_X1 U14288 ( .A(n11210), .ZN(n11219) );
  INV_X1 U14289 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19553) );
  NAND2_X1 U14290 ( .A1(n11006), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11211) );
  OAI21_X1 U14291 ( .B1(n11219), .B2(n19553), .A(n11211), .ZN(n11212) );
  AOI21_X1 U14292 ( .B1(n11005), .B2(P2_REIP_REG_24__SCAN_IN), .A(n11212), 
        .ZN(n15535) );
  INV_X1 U14293 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19551) );
  INV_X1 U14294 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15813) );
  OAI22_X1 U14295 ( .A1(n11219), .A2(n19551), .B1(n11218), .B2(n15813), .ZN(
        n11213) );
  AOI21_X1 U14296 ( .B1(n11005), .B2(P2_REIP_REG_25__SCAN_IN), .A(n11213), 
        .ZN(n15529) );
  NAND2_X1 U14297 ( .A1(n11005), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14298 ( .A1(n11210), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U14299 ( .A1(n11215), .A2(n11214), .ZN(n15522) );
  INV_X1 U14300 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19548) );
  NAND2_X1 U14301 ( .A1(n11006), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11216) );
  OAI21_X1 U14302 ( .B1(n11219), .B2(n19548), .A(n11216), .ZN(n11217) );
  AOI21_X1 U14303 ( .B1(n11005), .B2(P2_REIP_REG_27__SCAN_IN), .A(n11217), 
        .ZN(n15341) );
  INV_X1 U14304 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19546) );
  OAI22_X1 U14305 ( .A1(n11219), .A2(n19546), .B1(n11218), .B2(n11568), .ZN(
        n11220) );
  AOI21_X1 U14306 ( .B1(n11005), .B2(P2_REIP_REG_28__SCAN_IN), .A(n11220), 
        .ZN(n11603) );
  NAND2_X1 U14307 ( .A1(n11005), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14308 ( .A1(n11210), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11221) );
  NAND2_X1 U14309 ( .A1(n11222), .A2(n11221), .ZN(n15326) );
  NAND2_X1 U14310 ( .A1(n11005), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14311 ( .A1(n11210), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11006), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U14312 ( .A1(n11224), .A2(n11223), .ZN(n13063) );
  NAND2_X1 U14313 ( .A1(n15328), .A2(n13063), .ZN(n13067) );
  AOI222_X1 U14314 ( .A1(n11005), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11210), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11006), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11225) );
  XNOR2_X1 U14315 ( .A(n13067), .B(n11225), .ZN(n15500) );
  NAND2_X1 U14316 ( .A1(n11227), .A2(n11226), .ZN(n13861) );
  OAI21_X1 U14317 ( .B1(n9736), .B2(n9837), .A(n13861), .ZN(n11228) );
  NAND2_X1 U14318 ( .A1(n11587), .A2(n11228), .ZN(n19667) );
  NAND2_X1 U14319 ( .A1(n11229), .A2(n20259), .ZN(n19388) );
  INV_X2 U14320 ( .A(n19388), .ZN(n19643) );
  INV_X2 U14321 ( .A(n19643), .ZN(n19272) );
  INV_X1 U14322 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n21234) );
  NOR2_X1 U14323 ( .A1(n19272), .A2(n21234), .ZN(n13004) );
  INV_X1 U14324 ( .A(n13004), .ZN(n11258) );
  NAND2_X1 U14325 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11384) );
  NAND2_X1 U14326 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16710) );
  INV_X1 U14327 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15987) );
  NOR2_X1 U14328 ( .A1(n10787), .A2(n15987), .ZN(n15986) );
  INV_X1 U14329 ( .A(n15986), .ZN(n11380) );
  INV_X1 U14330 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U14331 ( .A1(n11587), .A2(n13541), .ZN(n16112) );
  NOR2_X1 U14332 ( .A1(n16014), .A2(n13532), .ZN(n11377) );
  INV_X1 U14333 ( .A(n11377), .ZN(n19670) );
  NOR2_X1 U14334 ( .A1(n10577), .A2(n19670), .ZN(n19657) );
  INV_X1 U14335 ( .A(n19657), .ZN(n11256) );
  NOR2_X1 U14336 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11377), .ZN(
        n11255) );
  NAND2_X1 U14337 ( .A1(n11234), .A2(n14195), .ZN(n13842) );
  NAND2_X1 U14338 ( .A1(n13842), .A2(n11235), .ZN(n11243) );
  INV_X1 U14339 ( .A(n11236), .ZN(n11237) );
  NAND2_X1 U14340 ( .A1(n11238), .A2(n11237), .ZN(n11240) );
  AOI21_X1 U14341 ( .B1(n11240), .B2(n11239), .A(n10533), .ZN(n11242) );
  MUX2_X1 U14342 ( .A(n11243), .B(n11242), .S(n11241), .Z(n11252) );
  OAI22_X1 U14343 ( .A1(n11239), .A2(n11245), .B1(n13873), .B2(n19682), .ZN(
        n11246) );
  INV_X1 U14344 ( .A(n11246), .ZN(n11250) );
  AND2_X1 U14345 ( .A1(n11247), .A2(n13873), .ZN(n11248) );
  NAND2_X1 U14346 ( .A1(n11249), .A2(n11248), .ZN(n13572) );
  NAND3_X1 U14347 ( .A1(n11244), .A2(n11250), .A3(n13572), .ZN(n11251) );
  NOR2_X1 U14348 ( .A1(n11252), .A2(n11251), .ZN(n13815) );
  INV_X1 U14349 ( .A(n11253), .ZN(n13817) );
  NAND2_X1 U14350 ( .A1(n13815), .A2(n13817), .ZN(n11254) );
  NAND2_X1 U14351 ( .A1(n11587), .A2(n11254), .ZN(n16117) );
  AOI211_X1 U14352 ( .C1(n16112), .C2(n11256), .A(n11255), .B(n16726), .ZN(
        n14326) );
  NAND2_X1 U14353 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14326), .ZN(
        n19656) );
  NOR2_X1 U14354 ( .A1(n11380), .A2(n19656), .ZN(n15972) );
  NAND2_X1 U14355 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15972), .ZN(
        n15954) );
  NAND2_X1 U14356 ( .A1(n15887), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15889) );
  INV_X1 U14357 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15890) );
  NOR2_X1 U14358 ( .A1(n15889), .A2(n15890), .ZN(n11382) );
  AND2_X1 U14359 ( .A1(n16683), .A2(n11382), .ZN(n15882) );
  NAND2_X1 U14360 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15882), .ZN(
        n15865) );
  NOR2_X1 U14361 ( .A1(n11384), .A2(n15865), .ZN(n15836) );
  NAND2_X1 U14362 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15836), .ZN(
        n15824) );
  NOR2_X1 U14363 ( .A1(n15812), .A2(n15824), .ZN(n15799) );
  NAND2_X1 U14364 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11560) );
  NOR2_X1 U14365 ( .A1(n15589), .A2(n11560), .ZN(n15774) );
  INV_X1 U14366 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14367 ( .A1(n15799), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15774), .A4(n11373), .ZN(n11257) );
  OAI211_X1 U14368 ( .C1(n15500), .C2(n19667), .A(n11258), .B(n11257), .ZN(
        n11391) );
  INV_X1 U14369 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16148) );
  OR2_X1 U14370 ( .A1(n11374), .A2(n16148), .ZN(n11263) );
  AOI22_X1 U14371 ( .A1(n11367), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11261) );
  NAND2_X1 U14372 ( .A1(n9752), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11260) );
  AND2_X1 U14373 ( .A1(n11261), .A2(n11260), .ZN(n11262) );
  NAND2_X1 U14374 ( .A1(n11263), .A2(n11262), .ZN(n15483) );
  INV_X1 U14375 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11265) );
  INV_X1 U14376 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11264) );
  OAI22_X1 U14377 ( .A1(n10571), .A2(n11265), .B1(n10591), .B2(n11264), .ZN(
        n11268) );
  NOR2_X1 U14378 ( .A1(n11374), .A2(n11266), .ZN(n11267) );
  AOI211_X1 U14379 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n9752), .A(n11268), .B(
        n11267), .ZN(n14245) );
  INV_X1 U14380 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11269) );
  OR2_X1 U14381 ( .A1(n11374), .A2(n11269), .ZN(n11273) );
  AOI22_X1 U14382 ( .A1(n11367), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11271) );
  NAND2_X1 U14383 ( .A1(n9752), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11270) );
  AND2_X1 U14384 ( .A1(n11271), .A2(n11270), .ZN(n11272) );
  NAND2_X1 U14385 ( .A1(n11273), .A2(n11272), .ZN(n14202) );
  INV_X1 U14386 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11274) );
  OR2_X1 U14387 ( .A1(n11374), .A2(n11274), .ZN(n11278) );
  AOI22_X1 U14388 ( .A1(n11367), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14389 ( .A1(n11330), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11275) );
  AND2_X1 U14390 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  NAND2_X1 U14391 ( .A1(n11278), .A2(n11277), .ZN(n13992) );
  OR2_X1 U14392 ( .A1(n11374), .A2(n15987), .ZN(n11282) );
  AOI22_X1 U14393 ( .A1(n11367), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14394 ( .A1(n11330), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11279) );
  AND2_X1 U14395 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  NAND2_X1 U14396 ( .A1(n11282), .A2(n11281), .ZN(n13887) );
  OR2_X1 U14397 ( .A1(n11374), .A2(n10787), .ZN(n11286) );
  AOI22_X1 U14398 ( .A1(n11367), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11284) );
  NAND2_X1 U14399 ( .A1(n11330), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11283) );
  AND2_X1 U14400 ( .A1(n11284), .A2(n11283), .ZN(n11285) );
  NAND2_X1 U14401 ( .A1(n11288), .A2(n11287), .ZN(n11293) );
  INV_X1 U14402 ( .A(n11289), .ZN(n11291) );
  NAND2_X1 U14403 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  NAND2_X1 U14404 ( .A1(n11293), .A2(n11292), .ZN(n13780) );
  INV_X1 U14405 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15971) );
  OR2_X1 U14406 ( .A1(n11374), .A2(n15971), .ZN(n11297) );
  AOI22_X1 U14407 ( .A1(n11367), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11295) );
  NAND2_X1 U14408 ( .A1(n11330), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11294) );
  AND2_X1 U14409 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  NAND2_X1 U14410 ( .A1(n11297), .A2(n11296), .ZN(n13904) );
  INV_X1 U14411 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11451) );
  OR2_X1 U14412 ( .A1(n11374), .A2(n11451), .ZN(n11301) );
  AOI22_X1 U14413 ( .A1(n11367), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U14414 ( .A1(n11330), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11298) );
  AND2_X1 U14415 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  NAND2_X1 U14416 ( .A1(n11301), .A2(n11300), .ZN(n13895) );
  OR2_X1 U14417 ( .A1(n11374), .A2(n11449), .ZN(n11305) );
  AOI22_X1 U14418 ( .A1(n11367), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11303) );
  NAND2_X1 U14419 ( .A1(n11330), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11302) );
  AND2_X1 U14420 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  INV_X1 U14421 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15730) );
  OR2_X1 U14422 ( .A1(n11374), .A2(n15730), .ZN(n11309) );
  AOI22_X1 U14423 ( .A1(n11367), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11307) );
  NAND2_X1 U14424 ( .A1(n11330), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11306) );
  AND2_X1 U14425 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  NAND2_X1 U14426 ( .A1(n11309), .A2(n11308), .ZN(n14119) );
  INV_X1 U14427 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16615) );
  OR2_X1 U14428 ( .A1(n11374), .A2(n16615), .ZN(n11313) );
  AOI22_X1 U14429 ( .A1(n11367), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11311) );
  NAND2_X1 U14430 ( .A1(n11330), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11310) );
  AND2_X1 U14431 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  NAND2_X1 U14432 ( .A1(n11313), .A2(n11312), .ZN(n14125) );
  INV_X1 U14433 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15939) );
  OR2_X1 U14434 ( .A1(n11374), .A2(n15939), .ZN(n11317) );
  AOI22_X1 U14435 ( .A1(n11367), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11315) );
  NAND2_X1 U14436 ( .A1(n9752), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11314) );
  AND2_X1 U14437 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  INV_X1 U14438 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14439 ( .A1(n11367), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11319) );
  NAND2_X1 U14440 ( .A1(n9752), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11318) );
  OAI211_X1 U14441 ( .C1(n11374), .C2(n11507), .A(n11319), .B(n11318), .ZN(
        n14250) );
  INV_X1 U14442 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16125) );
  OR2_X1 U14443 ( .A1(n11374), .A2(n16125), .ZN(n11323) );
  AOI22_X1 U14444 ( .A1(n11367), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11321) );
  NAND2_X1 U14445 ( .A1(n11330), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11320) );
  AND2_X1 U14446 ( .A1(n11321), .A2(n11320), .ZN(n11322) );
  NOR2_X2 U14447 ( .A1(n15494), .A2(n15495), .ZN(n15493) );
  AND2_X2 U14448 ( .A1(n15483), .A2(n15493), .ZN(n15485) );
  INV_X1 U14449 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15718) );
  OR2_X1 U14450 ( .A1(n11374), .A2(n15718), .ZN(n11327) );
  AOI22_X1 U14451 ( .A1(n11367), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11325) );
  NAND2_X1 U14452 ( .A1(n9752), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11324) );
  AND2_X1 U14453 ( .A1(n11325), .A2(n11324), .ZN(n11326) );
  NAND2_X1 U14454 ( .A1(n11327), .A2(n11326), .ZN(n15475) );
  INV_X1 U14455 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15910) );
  AOI22_X1 U14456 ( .A1(n11367), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11329) );
  NAND2_X1 U14457 ( .A1(n11330), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11328) );
  OAI211_X1 U14458 ( .C1(n11374), .C2(n15910), .A(n11329), .B(n11328), .ZN(
        n15367) );
  INV_X1 U14459 ( .A(n11330), .ZN(n11357) );
  INV_X1 U14460 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U14461 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14462 ( .A1(n11367), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11331) );
  OAI211_X1 U14463 ( .C1(n11357), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        n11334) );
  AOI21_X1 U14464 ( .B1(n11259), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11334), .ZN(n15464) );
  AOI22_X1 U14465 ( .A1(n11367), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11336) );
  NAND2_X1 U14466 ( .A1(n11330), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11335) );
  OAI211_X1 U14467 ( .C1(n11374), .C2(n15881), .A(n11336), .B(n11335), .ZN(
        n13496) );
  INV_X1 U14468 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U14469 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U14470 ( .A1(n11367), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11337) );
  OAI211_X1 U14471 ( .C1(n11357), .C2(n11339), .A(n11338), .B(n11337), .ZN(
        n11340) );
  AOI21_X1 U14472 ( .B1(n11259), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11340), .ZN(n15446) );
  OR2_X2 U14473 ( .A1(n15445), .A2(n15446), .ZN(n15447) );
  INV_X1 U14474 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11343) );
  NAND2_X1 U14475 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14476 ( .A1(n11367), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11341) );
  OAI211_X1 U14477 ( .C1(n11357), .C2(n11343), .A(n11342), .B(n11341), .ZN(
        n11344) );
  AOI21_X1 U14478 ( .B1(n11259), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11344), .ZN(n15352) );
  NAND2_X1 U14479 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11346) );
  NAND2_X1 U14480 ( .A1(n11367), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11345) );
  OAI211_X1 U14481 ( .C1(n11357), .C2(n10033), .A(n11346), .B(n11345), .ZN(
        n11347) );
  AOI21_X1 U14482 ( .B1(n11259), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11347), .ZN(n15434) );
  AOI22_X1 U14483 ( .A1(n11367), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11349) );
  NAND2_X1 U14484 ( .A1(n9752), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11348) );
  OAI211_X1 U14485 ( .C1(n11374), .C2(n15813), .A(n11349), .B(n11348), .ZN(
        n15426) );
  INV_X1 U14486 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U14487 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U14488 ( .A1(n11367), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11350) );
  OAI211_X1 U14489 ( .C1(n11357), .C2(n11352), .A(n11351), .B(n11350), .ZN(
        n11353) );
  AOI21_X1 U14490 ( .B1(n11259), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11353), .ZN(n15415) );
  INV_X1 U14491 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U14492 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14493 ( .A1(n11367), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11354) );
  OAI211_X1 U14494 ( .C1(n11357), .C2(n11356), .A(n11355), .B(n11354), .ZN(
        n11358) );
  AOI21_X1 U14495 ( .B1(n11259), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11358), .ZN(n15337) );
  NOR2_X2 U14496 ( .A1(n15416), .A2(n15337), .ZN(n15336) );
  OR2_X1 U14497 ( .A1(n11374), .A2(n11568), .ZN(n11362) );
  AOI22_X1 U14498 ( .A1(n11367), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11360) );
  NAND2_X1 U14499 ( .A1(n11330), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11359) );
  AND2_X1 U14500 ( .A1(n11360), .A2(n11359), .ZN(n11361) );
  NAND2_X1 U14501 ( .A1(n11362), .A2(n11361), .ZN(n11599) );
  OR2_X1 U14502 ( .A1(n11374), .A2(n15589), .ZN(n11366) );
  AOI22_X1 U14503 ( .A1(n11367), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11364) );
  NAND2_X1 U14504 ( .A1(n9752), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11363) );
  AND2_X1 U14505 ( .A1(n11364), .A2(n11363), .ZN(n11365) );
  NAND2_X1 U14506 ( .A1(n11366), .A2(n11365), .ZN(n15321) );
  INV_X1 U14507 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15779) );
  OR2_X1 U14508 ( .A1(n11374), .A2(n15779), .ZN(n11370) );
  AOI22_X1 U14509 ( .A1(n11367), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11369) );
  NAND2_X1 U14510 ( .A1(n11330), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11368) );
  AND3_X1 U14511 ( .A1(n11370), .A2(n11369), .A3(n11368), .ZN(n13058) );
  AOI22_X1 U14512 ( .A1(n11367), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11372) );
  NAND2_X1 U14513 ( .A1(n9752), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11371) );
  OAI211_X1 U14514 ( .C1(n11374), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        n11375) );
  AND2_X1 U14515 ( .A1(n9723), .A2(n11587), .ZN(n19669) );
  INV_X1 U14516 ( .A(n16726), .ZN(n15995) );
  INV_X1 U14517 ( .A(n15774), .ZN(n15787) );
  NOR2_X1 U14518 ( .A1(n16117), .A2(n11377), .ZN(n11378) );
  NOR2_X1 U14519 ( .A1(n11587), .A2(n19643), .ZN(n16717) );
  NOR2_X1 U14520 ( .A1(n11378), .A2(n16717), .ZN(n19677) );
  NAND2_X1 U14521 ( .A1(n19677), .A2(n16726), .ZN(n16115) );
  INV_X1 U14522 ( .A(n16112), .ZN(n19658) );
  NAND3_X1 U14523 ( .A1(n19658), .A2(n10577), .A3(n19670), .ZN(n19662) );
  INV_X1 U14524 ( .A(n16117), .ZN(n11379) );
  NAND2_X1 U14525 ( .A1(n11379), .A2(n10577), .ZN(n19671) );
  NAND4_X1 U14526 ( .A1(n19677), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19662), .A4(n19671), .ZN(n15980) );
  NOR3_X1 U14527 ( .A1(n11380), .A2(n15971), .A3(n15980), .ZN(n11381) );
  INV_X1 U14528 ( .A(n16115), .ZN(n16681) );
  NOR2_X1 U14529 ( .A1(n11381), .A2(n16681), .ZN(n16707) );
  AOI21_X1 U14530 ( .B1(n16115), .B2(n16710), .A(n16707), .ZN(n16682) );
  NAND2_X1 U14531 ( .A1(n16682), .A2(n11382), .ZN(n15872) );
  OR2_X1 U14532 ( .A1(n15872), .A2(n15881), .ZN(n11383) );
  NAND2_X1 U14533 ( .A1(n11383), .A2(n16115), .ZN(n15863) );
  INV_X1 U14534 ( .A(n11384), .ZN(n15848) );
  OAI21_X1 U14535 ( .B1(n16726), .B2(n15848), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11385) );
  INV_X1 U14536 ( .A(n11385), .ZN(n11386) );
  NAND2_X1 U14537 ( .A1(n15863), .A2(n11386), .ZN(n15835) );
  NAND2_X1 U14538 ( .A1(n15835), .A2(n16115), .ZN(n15823) );
  NAND2_X1 U14539 ( .A1(n16115), .A2(n15812), .ZN(n11387) );
  NAND2_X1 U14540 ( .A1(n15823), .A2(n11387), .ZN(n15807) );
  AOI21_X1 U14541 ( .B1(n15995), .B2(n15787), .A(n15807), .ZN(n15780) );
  OAI21_X1 U14542 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16726), .A(
        n15780), .ZN(n11388) );
  NAND2_X1 U14543 ( .A1(n11388), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11389) );
  NAND2_X1 U14544 ( .A1(n10247), .A2(n11389), .ZN(n11390) );
  INV_X1 U14545 ( .A(n11395), .ZN(n11398) );
  INV_X1 U14546 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11396) );
  INV_X1 U14547 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13624) );
  NAND2_X1 U14548 ( .A1(n11396), .A2(n13624), .ZN(n11397) );
  MUX2_X1 U14549 ( .A(n11398), .B(n11397), .S(n11455), .Z(n11411) );
  INV_X1 U14550 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14574) );
  INV_X1 U14551 ( .A(n11399), .ZN(n11400) );
  NAND2_X1 U14552 ( .A1(n13059), .A2(n11400), .ZN(n11401) );
  OAI21_X1 U14553 ( .B1(n13059), .B2(n11402), .A(n11401), .ZN(n11403) );
  INV_X1 U14554 ( .A(n11403), .ZN(n11404) );
  MUX2_X1 U14555 ( .A(n14574), .B(n11404), .S(n10449), .Z(n11405) );
  OAI21_X1 U14556 ( .B1(n11410), .B2(n11405), .A(n11428), .ZN(n14573) );
  OAI21_X2 U14557 ( .B1(n14325), .B2(n11584), .A(n14573), .ZN(n11418) );
  INV_X1 U14558 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11406) );
  MUX2_X1 U14559 ( .A(n11407), .B(P2_EBX_REG_0__SCAN_IN), .S(n11455), .Z(
        n13533) );
  INV_X1 U14560 ( .A(n13533), .ZN(n19446) );
  NOR2_X1 U14561 ( .A1(n19446), .A2(n13532), .ZN(n13559) );
  NAND3_X1 U14562 ( .A1(n11455), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11408) );
  AND2_X1 U14563 ( .A1(n11411), .A2(n11408), .ZN(n15390) );
  NAND2_X1 U14564 ( .A1(n13559), .A2(n15390), .ZN(n11409) );
  NOR2_X1 U14565 ( .A1(n13559), .A2(n15390), .ZN(n13558) );
  AOI21_X1 U14566 ( .B1(n16014), .B2(n11409), .A(n13558), .ZN(n19628) );
  INV_X1 U14567 ( .A(n11410), .ZN(n11414) );
  NAND2_X1 U14568 ( .A1(n11412), .A2(n11411), .ZN(n11413) );
  NAND2_X1 U14569 ( .A1(n11414), .A2(n11413), .ZN(n14561) );
  XNOR2_X1 U14570 ( .A(n14561), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19626) );
  NAND2_X1 U14571 ( .A1(n19628), .A2(n19626), .ZN(n11417) );
  INV_X1 U14572 ( .A(n14561), .ZN(n11415) );
  NAND2_X1 U14573 ( .A1(n11415), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11416) );
  NAND2_X1 U14574 ( .A1(n11417), .A2(n11416), .ZN(n14322) );
  NAND2_X1 U14575 ( .A1(n11418), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11419) );
  INV_X1 U14576 ( .A(n11420), .ZN(n11421) );
  MUX2_X1 U14577 ( .A(n11422), .B(n11421), .S(n13059), .Z(n11423) );
  MUX2_X1 U14578 ( .A(n11423), .B(P2_EBX_REG_4__SCAN_IN), .S(n11455), .Z(
        n11427) );
  XNOR2_X1 U14579 ( .A(n11428), .B(n11427), .ZN(n11424) );
  XNOR2_X1 U14580 ( .A(n11424), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19615) );
  INV_X1 U14581 ( .A(n11424), .ZN(n19423) );
  NAND2_X1 U14582 ( .A1(n19423), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11425) );
  NAND2_X1 U14583 ( .A1(n11426), .A2(n11444), .ZN(n11430) );
  NOR2_X2 U14584 ( .A1(n11428), .A2(n11427), .ZN(n11436) );
  INV_X1 U14585 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19406) );
  MUX2_X1 U14586 ( .A(n11429), .B(n19406), .S(n11455), .Z(n11435) );
  XNOR2_X1 U14587 ( .A(n11436), .B(n11435), .ZN(n19407) );
  NAND2_X1 U14588 ( .A1(n11430), .A2(n19407), .ZN(n11431) );
  XNOR2_X1 U14589 ( .A(n11431), .B(n15987), .ZN(n15767) );
  NAND2_X1 U14590 ( .A1(n15766), .A2(n15767), .ZN(n11433) );
  NAND2_X1 U14591 ( .A1(n11431), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11432) );
  NAND2_X1 U14592 ( .A1(n11433), .A2(n11432), .ZN(n15967) );
  NAND2_X1 U14593 ( .A1(n11434), .A2(n11444), .ZN(n11438) );
  NAND2_X1 U14594 ( .A1(n11436), .A2(n11435), .ZN(n11443) );
  MUX2_X1 U14595 ( .A(n11437), .B(P2_EBX_REG_6__SCAN_IN), .S(n11455), .Z(
        n11442) );
  XNOR2_X1 U14596 ( .A(n11443), .B(n11442), .ZN(n19396) );
  NAND2_X1 U14597 ( .A1(n11438), .A2(n19396), .ZN(n11439) );
  XNOR2_X1 U14598 ( .A(n11439), .B(n15971), .ZN(n15966) );
  NAND2_X1 U14599 ( .A1(n15967), .A2(n15966), .ZN(n11441) );
  NAND2_X1 U14600 ( .A1(n11439), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11440) );
  OR2_X2 U14601 ( .A1(n11443), .A2(n11442), .ZN(n11448) );
  MUX2_X1 U14602 ( .A(n11444), .B(P2_EBX_REG_7__SCAN_IN), .S(n11455), .Z(
        n11447) );
  NAND2_X1 U14603 ( .A1(n11455), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11445) );
  NOR2_X1 U14604 ( .A1(n11460), .A2(n11445), .ZN(n11446) );
  OR2_X1 U14605 ( .A1(n11456), .A2(n11446), .ZN(n19377) );
  OR2_X1 U14606 ( .A1(n19377), .A2(n11444), .ZN(n11450) );
  NOR2_X1 U14607 ( .A1(n11450), .A2(n11449), .ZN(n16629) );
  XNOR2_X1 U14608 ( .A(n11448), .B(n10037), .ZN(n19387) );
  NAND2_X1 U14609 ( .A1(n11450), .A2(n11449), .ZN(n16627) );
  INV_X1 U14610 ( .A(n19387), .ZN(n11452) );
  NAND2_X1 U14611 ( .A1(n11452), .A2(n11451), .ZN(n16626) );
  AND2_X1 U14612 ( .A1(n16627), .A2(n16626), .ZN(n11453) );
  INV_X1 U14613 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11454) );
  INV_X1 U14614 ( .A(n11467), .ZN(n11459) );
  NAND2_X1 U14615 ( .A1(n11455), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11457) );
  MUX2_X1 U14616 ( .A(n11457), .B(n11455), .S(n11456), .Z(n11458) );
  AOI21_X1 U14617 ( .B1(n11470), .B2(n11584), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15745) );
  INV_X1 U14618 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U14619 ( .A1(n11467), .A2(n14124), .ZN(n11465) );
  INV_X1 U14620 ( .A(n11460), .ZN(n11461) );
  NOR2_X1 U14621 ( .A1(n11467), .A2(n14124), .ZN(n11462) );
  NAND2_X1 U14622 ( .A1(n11455), .A2(n11462), .ZN(n11463) );
  AND2_X1 U14623 ( .A1(n11557), .A2(n11463), .ZN(n11464) );
  NAND2_X1 U14624 ( .A1(n11465), .A2(n11464), .ZN(n19351) );
  OR2_X1 U14625 ( .A1(n19351), .A2(n11444), .ZN(n11466) );
  NAND2_X1 U14626 ( .A1(n11466), .A2(n15730), .ZN(n15734) );
  INV_X1 U14627 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n14127) );
  NAND2_X1 U14628 ( .A1(n14127), .A2(n11468), .ZN(n11478) );
  NAND3_X1 U14629 ( .A1(n11455), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n11465), 
        .ZN(n11469) );
  AND2_X1 U14630 ( .A1(n11475), .A2(n11469), .ZN(n15383) );
  AOI21_X1 U14631 ( .B1(n15383), .B2(n11584), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16611) );
  INV_X1 U14632 ( .A(n11470), .ZN(n19362) );
  NAND2_X1 U14633 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11471) );
  OR2_X1 U14634 ( .A1(n19362), .A2(n11471), .ZN(n15731) );
  OR3_X1 U14635 ( .A1(n19351), .A2(n11444), .A3(n15730), .ZN(n15733) );
  NAND2_X1 U14636 ( .A1(n15731), .A2(n15733), .ZN(n16607) );
  INV_X1 U14637 ( .A(n15383), .ZN(n11473) );
  NAND2_X1 U14638 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11472) );
  NOR2_X1 U14639 ( .A1(n11473), .A2(n11472), .ZN(n16610) );
  NOR2_X1 U14640 ( .A1(n16607), .A2(n16610), .ZN(n11474) );
  NAND2_X1 U14641 ( .A1(n11455), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11476) );
  NAND3_X1 U14642 ( .A1(n11455), .A2(n11478), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n11479) );
  NAND2_X1 U14643 ( .A1(n11503), .A2(n11479), .ZN(n19341) );
  NAND2_X1 U14644 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11480) );
  NOR2_X1 U14645 ( .A1(n19341), .A2(n11480), .ZN(n15932) );
  NAND2_X1 U14646 ( .A1(n11455), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11484) );
  NAND2_X1 U14647 ( .A1(n11455), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11502) );
  OAI21_X1 U14648 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n11455), .ZN(n11481) );
  OR2_X2 U14649 ( .A1(n11510), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11482) );
  INV_X1 U14650 ( .A(n11517), .ZN(n11483) );
  MUX2_X1 U14651 ( .A(n11484), .B(n11455), .S(n11491), .Z(n11486) );
  INV_X1 U14652 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11485) );
  NAND2_X1 U14653 ( .A1(n11491), .A2(n11485), .ZN(n11489) );
  NAND2_X1 U14654 ( .A1(n11486), .A2(n11489), .ZN(n19278) );
  INV_X1 U14655 ( .A(n19278), .ZN(n11487) );
  NAND2_X1 U14656 ( .A1(n11487), .A2(n11584), .ZN(n11533) );
  NAND2_X1 U14657 ( .A1(n11533), .A2(n15718), .ZN(n15701) );
  AND2_X1 U14658 ( .A1(n11455), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U14659 ( .A1(n11489), .A2(n11488), .ZN(n11492) );
  OAI21_X1 U14660 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n11455), .ZN(n11490) );
  NAND2_X1 U14661 ( .A1(n11492), .A2(n11521), .ZN(n15372) );
  OR2_X1 U14662 ( .A1(n15372), .A2(n11444), .ZN(n11493) );
  NAND2_X1 U14663 ( .A1(n11493), .A2(n15910), .ZN(n15700) );
  AND2_X1 U14664 ( .A1(n15701), .A2(n15700), .ZN(n15673) );
  INV_X1 U14665 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U14666 ( .A1(n11539), .A2(n11557), .ZN(n11538) );
  NAND2_X1 U14667 ( .A1(n11455), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11495) );
  NOR2_X1 U14668 ( .A1(n11496), .A2(n11495), .ZN(n11497) );
  OR2_X1 U14669 ( .A1(n11538), .A2(n11497), .ZN(n13495) );
  OR2_X1 U14670 ( .A1(n13495), .A2(n11444), .ZN(n11498) );
  NAND2_X1 U14671 ( .A1(n11498), .A2(n15881), .ZN(n15663) );
  NAND2_X1 U14672 ( .A1(n11455), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11499) );
  MUX2_X1 U14673 ( .A(n11499), .B(n11455), .S(n9776), .Z(n11500) );
  INV_X1 U14674 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U14675 ( .A1(n9776), .A2(n14248), .ZN(n11505) );
  NAND2_X1 U14676 ( .A1(n19322), .A2(n11584), .ZN(n11501) );
  NAND2_X1 U14677 ( .A1(n11501), .A2(n11266), .ZN(n16585) );
  XNOR2_X1 U14678 ( .A(n11503), .B(n11502), .ZN(n19330) );
  AOI21_X1 U14679 ( .B1(n19330), .B2(n11584), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15665) );
  INV_X1 U14680 ( .A(n15665), .ZN(n16595) );
  AND2_X1 U14681 ( .A1(n11455), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14682 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  NAND2_X1 U14683 ( .A1(n11506), .A2(n11510), .ZN(n19308) );
  OR2_X1 U14684 ( .A1(n19308), .A2(n11444), .ZN(n11508) );
  NAND2_X1 U14685 ( .A1(n11508), .A2(n11507), .ZN(n16575) );
  OR2_X1 U14686 ( .A1(n19341), .A2(n11444), .ZN(n11509) );
  NAND2_X1 U14687 ( .A1(n11509), .A2(n15939), .ZN(n15931) );
  NAND4_X1 U14688 ( .A1(n16585), .A2(n16595), .A3(n16575), .A4(n15931), .ZN(
        n11516) );
  NAND2_X1 U14689 ( .A1(n11455), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11511) );
  MUX2_X1 U14690 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n11511), .S(n11510), .Z(
        n11512) );
  NAND2_X1 U14691 ( .A1(n11512), .A2(n11557), .ZN(n11513) );
  OAI21_X1 U14692 ( .B1(n11513), .B2(n11444), .A(n16125), .ZN(n11515) );
  INV_X1 U14693 ( .A(n11513), .ZN(n19300) );
  AND2_X1 U14694 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11514) );
  NAND2_X1 U14695 ( .A1(n19300), .A2(n11514), .ZN(n15669) );
  NAND2_X1 U14696 ( .A1(n11515), .A2(n15669), .ZN(n16121) );
  OR2_X1 U14697 ( .A1(n11516), .A2(n16121), .ZN(n11519) );
  XNOR2_X1 U14698 ( .A(n11518), .B(n11517), .ZN(n19287) );
  AOI21_X1 U14699 ( .B1(n19287), .B2(n11584), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15722) );
  NOR2_X1 U14700 ( .A1(n11519), .A2(n15722), .ZN(n11523) );
  NAND2_X1 U14701 ( .A1(n11455), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11520) );
  XNOR2_X1 U14702 ( .A(n11521), .B(n11520), .ZN(n19258) );
  NAND2_X1 U14703 ( .A1(n19258), .A2(n11584), .ZN(n11522) );
  NAND2_X1 U14704 ( .A1(n11522), .A2(n15890), .ZN(n15685) );
  AND4_X1 U14705 ( .A1(n15673), .A2(n15663), .A3(n11523), .A4(n15685), .ZN(
        n11524) );
  NAND2_X1 U14706 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11525) );
  OR2_X1 U14707 ( .A1(n13495), .A2(n11525), .ZN(n15662) );
  NAND2_X1 U14708 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11526) );
  OR2_X1 U14709 ( .A1(n15372), .A2(n11526), .ZN(n15699) );
  AND2_X1 U14710 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U14711 ( .A1(n19322), .A2(n11527), .ZN(n16584) );
  NAND2_X1 U14712 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11528) );
  OR2_X1 U14713 ( .A1(n19308), .A2(n11528), .ZN(n16574) );
  AND2_X1 U14714 ( .A1(n16584), .A2(n16574), .ZN(n15666) );
  AND2_X1 U14715 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14716 ( .A1(n19330), .A2(n11529), .ZN(n16594) );
  AND3_X1 U14717 ( .A1(n15666), .A2(n15669), .A3(n16594), .ZN(n11531) );
  AND2_X1 U14718 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11530) );
  INV_X1 U14719 ( .A(n15721), .ZN(n15670) );
  AND3_X1 U14720 ( .A1(n15699), .A2(n11531), .A3(n15670), .ZN(n11535) );
  AND2_X1 U14721 ( .A1(n11584), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U14722 ( .A1(n19258), .A2(n11532), .ZN(n15684) );
  INV_X1 U14723 ( .A(n11533), .ZN(n11534) );
  NAND2_X1 U14724 ( .A1(n11534), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15672) );
  AND4_X1 U14725 ( .A1(n15662), .A2(n11535), .A3(n15684), .A4(n15672), .ZN(
        n11536) );
  NAND2_X1 U14726 ( .A1(n11455), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11537) );
  NAND3_X1 U14727 ( .A1(n11539), .A2(n11455), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n11540) );
  NAND2_X1 U14728 ( .A1(n11547), .A2(n11540), .ZN(n16129) );
  OR2_X1 U14729 ( .A1(n16129), .A2(n11444), .ZN(n11541) );
  INV_X1 U14730 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U14731 ( .A1(n11541), .A2(n15864), .ZN(n15650) );
  OR2_X1 U14732 ( .A1(n11541), .A2(n15864), .ZN(n15651) );
  NAND2_X1 U14733 ( .A1(n11542), .A2(n15651), .ZN(n15846) );
  AND2_X1 U14734 ( .A1(n11455), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11546) );
  INV_X1 U14735 ( .A(n11546), .ZN(n11543) );
  XNOR2_X1 U14736 ( .A(n11547), .B(n11543), .ZN(n15355) );
  NAND2_X1 U14737 ( .A1(n15355), .A2(n11584), .ZN(n11544) );
  XNOR2_X1 U14738 ( .A(n11544), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15845) );
  NAND2_X1 U14739 ( .A1(n15846), .A2(n15845), .ZN(n15847) );
  OR2_X1 U14740 ( .A1(n11544), .A2(n15853), .ZN(n11545) );
  NAND3_X1 U14741 ( .A1(n11548), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n11455), 
        .ZN(n11549) );
  NAND2_X1 U14742 ( .A1(n11549), .A2(n11557), .ZN(n11550) );
  OR2_X1 U14743 ( .A1(n11556), .A2(n11550), .ZN(n16537) );
  NOR2_X1 U14744 ( .A1(n11551), .A2(n15644), .ZN(n15641) );
  NAND2_X1 U14745 ( .A1(n11551), .A2(n15644), .ZN(n15640) );
  INV_X1 U14746 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11555) );
  NOR2_X1 U14747 ( .A1(n11556), .A2(n11555), .ZN(n11552) );
  NAND2_X1 U14748 ( .A1(n11455), .A2(n11552), .ZN(n11553) );
  NAND2_X1 U14749 ( .A1(n11557), .A2(n11553), .ZN(n11554) );
  AOI21_X1 U14750 ( .B1(n11556), .B2(n11555), .A(n11554), .ZN(n11561) );
  AOI21_X1 U14751 ( .B1(n11561), .B2(n11584), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15632) );
  NAND2_X1 U14752 ( .A1(n11557), .A2(n11564), .ZN(n11580) );
  AND3_X1 U14753 ( .A1(n11455), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n11558), .ZN(
        n11559) );
  NOR2_X1 U14754 ( .A1(n11580), .A2(n11559), .ZN(n16509) );
  NAND2_X1 U14755 ( .A1(n16509), .A2(n11584), .ZN(n11562) );
  XNOR2_X1 U14756 ( .A(n11562), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15621) );
  INV_X1 U14757 ( .A(n11560), .ZN(n15788) );
  INV_X1 U14758 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15814) );
  INV_X1 U14759 ( .A(n11561), .ZN(n16528) );
  OAI21_X1 U14760 ( .B1(n11562), .B2(n15814), .A(n15630), .ZN(n11592) );
  NAND2_X1 U14761 ( .A1(n11455), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14762 ( .A1(n11580), .A2(n11563), .ZN(n11570) );
  INV_X1 U14763 ( .A(n11563), .ZN(n11565) );
  NAND2_X1 U14764 ( .A1(n11565), .A2(n11564), .ZN(n11566) );
  AND2_X1 U14765 ( .A1(n11570), .A2(n11566), .ZN(n15344) );
  NAND2_X1 U14766 ( .A1(n15344), .A2(n11584), .ZN(n11593) );
  NAND2_X1 U14767 ( .A1(n11569), .A2(n11568), .ZN(n11573) );
  AND2_X1 U14768 ( .A1(n11455), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11571) );
  AOI21_X1 U14769 ( .B1(n11571), .B2(n11570), .A(n11574), .ZN(n16502) );
  NAND2_X1 U14770 ( .A1(n16502), .A2(n11584), .ZN(n11595) );
  NAND2_X1 U14771 ( .A1(n11574), .A2(n9847), .ZN(n11581) );
  NAND2_X1 U14772 ( .A1(n11455), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11575) );
  XNOR2_X1 U14773 ( .A(n11581), .B(n11575), .ZN(n11576) );
  AOI21_X1 U14774 ( .B1(n11576), .B2(n11584), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15581) );
  INV_X1 U14775 ( .A(n11576), .ZN(n13082) );
  INV_X1 U14776 ( .A(n11577), .ZN(n15329) );
  NAND3_X1 U14777 ( .A1(n15329), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11584), .ZN(n15592) );
  INV_X1 U14778 ( .A(n11580), .ZN(n11583) );
  NOR2_X1 U14779 ( .A1(n11581), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11582) );
  MUX2_X1 U14780 ( .A(n11583), .B(n11582), .S(n11455), .Z(n16491) );
  NAND2_X1 U14781 ( .A1(n16491), .A2(n11584), .ZN(n11585) );
  XNOR2_X1 U14782 ( .A(n11586), .B(n10258), .ZN(n12998) );
  NOR2_X1 U14783 ( .A1(n13872), .A2(n13059), .ZN(n20308) );
  NAND2_X1 U14784 ( .A1(n12998), .A2(n19663), .ZN(n11588) );
  NAND2_X1 U14785 ( .A1(n11589), .A2(n11588), .ZN(P2_U3015) );
  NOR2_X1 U14786 ( .A1(n15622), .A2(n11592), .ZN(n11594) );
  XNOR2_X1 U14787 ( .A(n11595), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11596) );
  INV_X1 U14788 ( .A(n15611), .ZN(n11598) );
  OAI21_X1 U14789 ( .B1(n11598), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11597), .ZN(n15600) );
  NOR2_X1 U14790 ( .A1(n15600), .A2(n19650), .ZN(n11610) );
  NOR2_X1 U14791 ( .A1(n15336), .A2(n11599), .ZN(n11600) );
  OR2_X2 U14792 ( .A1(n15320), .A2(n11600), .ZN(n16496) );
  XOR2_X1 U14793 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n11602) );
  INV_X1 U14794 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n11601) );
  NOR2_X1 U14795 ( .A1(n19272), .A2(n11601), .ZN(n15602) );
  AOI21_X1 U14796 ( .B1(n15799), .B2(n11602), .A(n15602), .ZN(n11605) );
  AOI21_X1 U14797 ( .B1(n11603), .B2(n15343), .A(n9777), .ZN(n16497) );
  NAND2_X1 U14798 ( .A1(n19645), .A2(n16497), .ZN(n11604) );
  OAI211_X1 U14799 ( .C1(n16496), .C2(n16143), .A(n11605), .B(n11604), .ZN(
        n11606) );
  INV_X1 U14800 ( .A(n11606), .ZN(n11608) );
  NAND2_X1 U14801 ( .A1(n15807), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11607) );
  NOR2_X1 U14802 ( .A1(n9968), .A2(n19076), .ZN(n17099) );
  INV_X1 U14803 ( .A(n17099), .ZN(n17255) );
  NOR3_X1 U14804 ( .A1(n16772), .A2(n11612), .A3(n17255), .ZN(n11623) );
  INV_X1 U14805 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21249) );
  AOI21_X1 U14806 ( .B1(n16940), .B2(n10257), .A(n21249), .ZN(n11622) );
  INV_X1 U14807 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17280) );
  NAND2_X1 U14808 ( .A1(n11613), .A2(n17280), .ZN(n11620) );
  NOR2_X1 U14809 ( .A1(n17254), .A2(n16755), .ZN(n11618) );
  NOR3_X1 U14810 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19157), .A3(n11614), 
        .ZN(n11615) );
  AOI21_X1 U14811 ( .B1(n17266), .B2(P3_EBX_REG_31__SCAN_IN), .A(n11615), .ZN(
        n11616) );
  INV_X1 U14812 ( .A(n11616), .ZN(n11617) );
  NOR2_X1 U14813 ( .A1(n11618), .A2(n11617), .ZN(n11619) );
  AOI22_X1 U14814 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n17504), .B1(
        P3_INSTQUEUE_REG_10__6__SCAN_IN), .B2(n14519), .ZN(n11628) );
  AOI22_X1 U14815 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17503), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14816 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14817 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n17523), .B1(
        P3_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n10308), .ZN(n11625) );
  NAND4_X1 U14818 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n11634) );
  AOI22_X1 U14819 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14820 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n17533), .ZN(n11631) );
  AOI22_X1 U14821 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14822 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14517), .ZN(n11629) );
  NAND4_X1 U14823 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11633) );
  AOI22_X1 U14824 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9732), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14825 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14826 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14827 ( .A1(n17533), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U14828 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11644) );
  AOI22_X1 U14829 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14830 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14831 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14832 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11639) );
  NAND4_X1 U14833 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11643) );
  AOI22_X1 U14834 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14835 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14836 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14837 ( .A1(n17533), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11646) );
  NAND4_X1 U14838 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11655) );
  AOI22_X1 U14839 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14840 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14841 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14842 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11650) );
  NAND4_X1 U14843 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11654) );
  AOI22_X1 U14844 ( .A1(n10342), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11656), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14845 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14846 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14847 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9719), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14848 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11670) );
  INV_X1 U14849 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n21310) );
  AOI22_X1 U14850 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11662) );
  OAI21_X1 U14851 ( .B1(n14469), .B2(n21310), .A(n11662), .ZN(n11663) );
  AOI22_X1 U14852 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14853 ( .A1(n11624), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11664) );
  AOI21_X1 U14854 ( .B1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11704), .A(
        n11665), .ZN(n11666) );
  NAND3_X1 U14855 ( .A1(n11668), .A2(n11667), .A3(n11666), .ZN(n11669) );
  OR2_X2 U14856 ( .A1(n11670), .A2(n11669), .ZN(n17715) );
  AOI22_X1 U14857 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14858 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14859 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11672) );
  OAI21_X1 U14860 ( .B1(n14458), .B2(n21174), .A(n11672), .ZN(n11678) );
  AOI22_X1 U14861 ( .A1(n9719), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14862 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14863 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14864 ( .A1(n17715), .A2(n17709), .ZN(n11702) );
  AOI22_X1 U14865 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14866 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14867 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11681) );
  OAI21_X1 U14868 ( .B1(n17476), .B2(n21223), .A(n11681), .ZN(n11687) );
  AOI22_X1 U14869 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14870 ( .A1(n11704), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14871 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14872 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U14873 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11686) );
  AOI211_X1 U14874 ( .C1(n17423), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n11687), .B(n11686), .ZN(n11688) );
  NAND3_X1 U14875 ( .A1(n11690), .A2(n11689), .A3(n11688), .ZN(n17701) );
  NAND2_X1 U14876 ( .A1(n11721), .A2(n17701), .ZN(n11724) );
  AOI22_X1 U14877 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14878 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11700) );
  INV_X1 U14879 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21314) );
  AOI22_X1 U14880 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9731), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11691) );
  OAI21_X1 U14881 ( .B1(n10310), .B2(n21314), .A(n11691), .ZN(n11698) );
  AOI22_X1 U14882 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14883 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14884 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14885 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14886 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11697) );
  AOI211_X1 U14887 ( .C1(n17325), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n11698), .B(n11697), .ZN(n11699) );
  NAND3_X1 U14888 ( .A1(n11701), .A2(n11700), .A3(n11699), .ZN(n11810) );
  NOR2_X1 U14889 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18109), .ZN(
        n16189) );
  AOI21_X1 U14890 ( .B1(n18109), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16189), .ZN(n17837) );
  INV_X1 U14891 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21104) );
  INV_X1 U14892 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18489) );
  XNOR2_X1 U14893 ( .A(n11702), .B(n17705), .ZN(n11718) );
  XOR2_X1 U14894 ( .A(n17715), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n18188) );
  AOI22_X1 U14895 ( .A1(n10342), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14896 ( .A1(n17526), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11712) );
  INV_X1 U14897 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n21295) );
  AOI22_X1 U14898 ( .A1(n9731), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11703) );
  OAI21_X1 U14899 ( .B1(n10245), .B2(n21295), .A(n11703), .ZN(n11710) );
  AOI22_X1 U14900 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11692), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14901 ( .A1(n11704), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14902 ( .A1(n9719), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14903 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U14904 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n11709) );
  AOI211_X1 U14905 ( .C1(n17504), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n11710), .B(n11709), .ZN(n11711) );
  NAND3_X1 U14906 ( .A1(n11713), .A2(n11712), .A3(n11711), .ZN(n18196) );
  NAND2_X1 U14907 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18196), .ZN(
        n18195) );
  NOR2_X1 U14908 ( .A1(n18188), .A2(n18195), .ZN(n18186) );
  INV_X1 U14909 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19181) );
  NOR2_X1 U14910 ( .A1(n17715), .A2(n19181), .ZN(n11714) );
  INV_X1 U14911 ( .A(n18180), .ZN(n11717) );
  INV_X1 U14912 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18510) );
  NOR2_X1 U14913 ( .A1(n18510), .A2(n11715), .ZN(n11716) );
  XNOR2_X1 U14914 ( .A(n11718), .B(n11719), .ZN(n18168) );
  NOR2_X1 U14915 ( .A1(n18489), .A2(n18168), .ZN(n18167) );
  NOR2_X1 U14916 ( .A1(n11719), .A2(n11718), .ZN(n11720) );
  NOR2_X1 U14917 ( .A1(n18167), .A2(n11720), .ZN(n18159) );
  INV_X1 U14918 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18480) );
  XOR2_X1 U14919 ( .A(n11721), .B(n17701), .Z(n11722) );
  XOR2_X1 U14920 ( .A(n18480), .B(n11722), .Z(n18158) );
  NOR2_X1 U14921 ( .A1(n18159), .A2(n18158), .ZN(n18157) );
  XNOR2_X1 U14922 ( .A(n11724), .B(n17697), .ZN(n18139) );
  INV_X1 U14923 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18460) );
  XNOR2_X1 U14924 ( .A(n11725), .B(n17694), .ZN(n11726) );
  XOR2_X1 U14925 ( .A(n18460), .B(n11726), .Z(n18127) );
  INV_X1 U14926 ( .A(n11815), .ZN(n11772) );
  XNOR2_X1 U14927 ( .A(n11729), .B(n11728), .ZN(n18123) );
  INV_X1 U14928 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18122) );
  NOR2_X1 U14929 ( .A1(n18123), .A2(n18122), .ZN(n18121) );
  NOR2_X1 U14930 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  INV_X1 U14931 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18438) );
  AND2_X2 U14932 ( .A1(n11733), .A2(n18438), .ZN(n18106) );
  INV_X1 U14933 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18063) );
  INV_X1 U14934 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18363) );
  NAND2_X1 U14935 ( .A1(n18016), .A2(n18363), .ZN(n18007) );
  INV_X1 U14936 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11732) );
  INV_X1 U14937 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11731) );
  INV_X1 U14938 ( .A(n11739), .ZN(n11737) );
  NAND2_X1 U14939 ( .A1(n18406), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18383) );
  INV_X1 U14940 ( .A(n18383), .ZN(n18408) );
  NAND2_X1 U14941 ( .A1(n18408), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18360) );
  INV_X1 U14942 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18359) );
  NOR2_X1 U14943 ( .A1(n18360), .A2(n18359), .ZN(n18368) );
  INV_X1 U14944 ( .A(n18368), .ZN(n18364) );
  NOR2_X1 U14945 ( .A1(n18363), .A2(n18364), .ZN(n18346) );
  NAND2_X1 U14946 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18346), .ZN(
        n18314) );
  INV_X1 U14947 ( .A(n18314), .ZN(n16773) );
  NOR2_X2 U14948 ( .A1(n11733), .A2(n18438), .ZN(n18399) );
  NAND2_X1 U14949 ( .A1(n16773), .A2(n18399), .ZN(n11738) );
  NAND2_X1 U14950 ( .A1(n11738), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11735) );
  INV_X1 U14951 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18341) );
  NOR2_X2 U14952 ( .A1(n11737), .A2(n11736), .ZN(n17986) );
  INV_X1 U14953 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18327) );
  NAND2_X1 U14954 ( .A1(n17986), .A2(n18327), .ZN(n17985) );
  INV_X1 U14955 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17908) );
  NOR2_X1 U14956 ( .A1(n18341), .A2(n18327), .ZN(n18317) );
  INV_X1 U14957 ( .A(n18317), .ZN(n17975) );
  INV_X1 U14958 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18320) );
  INV_X1 U14959 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18307) );
  INV_X1 U14960 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17946) );
  NOR2_X1 U14961 ( .A1(n18307), .A2(n17946), .ZN(n18287) );
  NAND2_X1 U14962 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18287), .ZN(
        n18272) );
  NOR2_X1 U14963 ( .A1(n18320), .A2(n18272), .ZN(n17917) );
  NAND2_X1 U14964 ( .A1(n17917), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11823) );
  NOR2_X1 U14965 ( .A1(n17975), .A2(n11823), .ZN(n11827) );
  INV_X1 U14966 ( .A(n11827), .ZN(n11821) );
  NOR2_X1 U14967 ( .A1(n17908), .A2(n11821), .ZN(n18251) );
  NOR2_X1 U14968 ( .A1(n18109), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17967) );
  NAND2_X1 U14969 ( .A1(n17967), .A2(n18307), .ZN(n11740) );
  NOR2_X1 U14970 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11740), .ZN(
        n17938) );
  INV_X1 U14971 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18280) );
  NAND2_X1 U14972 ( .A1(n17938), .A2(n18280), .ZN(n17916) );
  NOR3_X1 U14973 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17916), .ZN(n11741) );
  NAND2_X1 U14974 ( .A1(n18317), .A2(n17990), .ZN(n17937) );
  OR2_X1 U14975 ( .A1(n18109), .A2(n17889), .ZN(n17880) );
  OAI221_X1 U14976 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18107), 
        .C1(n21104), .C2(n17881), .A(n17880), .ZN(n17864) );
  NOR2_X1 U14977 ( .A1(n17864), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17863) );
  NAND2_X1 U14978 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18204) );
  NOR2_X2 U14979 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11745), .ZN(
        n16190) );
  INV_X1 U14980 ( .A(n16190), .ZN(n11834) );
  NAND2_X1 U14981 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11745), .ZN(
        n11816) );
  INV_X1 U14982 ( .A(n11816), .ZN(n16101) );
  NOR2_X1 U14983 ( .A1(n18552), .A2(n11746), .ZN(n11747) );
  NAND2_X1 U14984 ( .A1(n11747), .A2(n17575), .ZN(n11770) );
  INV_X1 U14985 ( .A(n11748), .ZN(n11751) );
  OAI21_X1 U14986 ( .B1(n11749), .B2(n14440), .A(n16209), .ZN(n11750) );
  NAND3_X1 U14987 ( .A1(n11751), .A2(n11804), .A3(n11750), .ZN(n11755) );
  NOR2_X1 U14988 ( .A1(n17691), .A2(n19004), .ZN(n11817) );
  AOI211_X1 U14989 ( .C1(n11755), .C2(n11754), .A(n11753), .B(n11752), .ZN(
        n11756) );
  INV_X1 U14990 ( .A(n11756), .ZN(n14609) );
  OAI21_X1 U14991 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19042), .A(
        n11757), .ZN(n11761) );
  AOI21_X1 U14992 ( .B1(n11758), .B2(n11761), .A(n11763), .ZN(n18998) );
  XOR2_X1 U14993 ( .A(n19215), .B(n18558), .Z(n11759) );
  AOI21_X1 U14994 ( .B1(n11759), .B2(n19088), .A(n19216), .ZN(n16912) );
  NAND3_X1 U14995 ( .A1(n16912), .A2(n11760), .A3(n19001), .ZN(n11769) );
  NOR2_X1 U14996 ( .A1(n11762), .A2(n11761), .ZN(n11765) );
  INV_X1 U14997 ( .A(n11763), .ZN(n11764) );
  OAI21_X1 U14998 ( .B1(n11767), .B2(n14440), .A(n19003), .ZN(n11768) );
  OAI211_X1 U14999 ( .C1(n18998), .C2(n11770), .A(n11769), .B(n11768), .ZN(
        n11771) );
  AND3_X1 U15000 ( .A1(n17835), .A2(n11772), .A3(n18441), .ZN(n11814) );
  INV_X1 U15001 ( .A(n17715), .ZN(n11773) );
  NOR2_X1 U15002 ( .A1(n11773), .A2(n18187), .ZN(n11782) );
  NOR2_X1 U15003 ( .A1(n11782), .A2(n17709), .ZN(n11780) );
  NOR2_X1 U15004 ( .A1(n17705), .A2(n11780), .ZN(n11779) );
  NAND2_X1 U15005 ( .A1(n11779), .A2(n17701), .ZN(n11777) );
  NOR2_X1 U15006 ( .A1(n17697), .A2(n11777), .ZN(n11775) );
  NAND2_X1 U15007 ( .A1(n11775), .A2(n11776), .ZN(n11774) );
  NOR2_X1 U15008 ( .A1(n17691), .A2(n11774), .ZN(n11798) );
  XOR2_X1 U15009 ( .A(n17691), .B(n11774), .Z(n18115) );
  XOR2_X1 U15010 ( .A(n11776), .B(n11775), .Z(n11791) );
  XOR2_X1 U15011 ( .A(n17697), .B(n11777), .Z(n11778) );
  NAND2_X1 U15012 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11778), .ZN(
        n11790) );
  XOR2_X1 U15013 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11778), .Z(
        n18142) );
  XOR2_X1 U15014 ( .A(n17701), .B(n11779), .Z(n18152) );
  XOR2_X1 U15015 ( .A(n17705), .B(n11780), .Z(n11781) );
  NAND2_X1 U15016 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11781), .ZN(
        n11787) );
  XOR2_X1 U15017 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11781), .Z(
        n18166) );
  XOR2_X1 U15018 ( .A(n17709), .B(n11782), .Z(n11783) );
  OR2_X1 U15019 ( .A1(n18510), .A2(n11783), .ZN(n11786) );
  XOR2_X1 U15020 ( .A(n18510), .B(n11783), .Z(n18177) );
  AOI21_X1 U15021 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17715), .A(
        n18196), .ZN(n11785) );
  INV_X1 U15022 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19195) );
  NOR2_X1 U15023 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17715), .ZN(
        n11784) );
  AOI221_X1 U15024 ( .B1(n18196), .B2(n17715), .C1(n11785), .C2(n19195), .A(
        n11784), .ZN(n18176) );
  NAND2_X1 U15025 ( .A1(n18177), .A2(n18176), .ZN(n18175) );
  NAND2_X1 U15026 ( .A1(n11786), .A2(n18175), .ZN(n18165) );
  NAND2_X1 U15027 ( .A1(n18166), .A2(n18165), .ZN(n18164) );
  NAND2_X1 U15028 ( .A1(n11787), .A2(n18164), .ZN(n18153) );
  NAND2_X1 U15029 ( .A1(n18152), .A2(n18153), .ZN(n18151) );
  NOR2_X1 U15030 ( .A1(n18152), .A2(n18153), .ZN(n11788) );
  AOI21_X1 U15031 ( .B1(n18480), .B2(n18151), .A(n11788), .ZN(n18141) );
  NAND2_X1 U15032 ( .A1(n18142), .A2(n18141), .ZN(n11789) );
  NAND2_X1 U15033 ( .A1(n11790), .A2(n11789), .ZN(n11792) );
  NAND2_X1 U15034 ( .A1(n11791), .A2(n11792), .ZN(n11793) );
  XOR2_X1 U15035 ( .A(n11792), .B(n11791), .Z(n18131) );
  NAND2_X1 U15036 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18131), .ZN(
        n18130) );
  NAND2_X1 U15037 ( .A1(n11793), .A2(n18130), .ZN(n18116) );
  NOR2_X1 U15038 ( .A1(n18115), .A2(n18116), .ZN(n11794) );
  NOR2_X1 U15039 ( .A1(n11794), .A2(n18122), .ZN(n11795) );
  NAND2_X1 U15040 ( .A1(n11798), .A2(n11795), .ZN(n11799) );
  INV_X1 U15041 ( .A(n11795), .ZN(n11797) );
  NAND2_X1 U15042 ( .A1(n18115), .A2(n18116), .ZN(n18114) );
  NAND2_X1 U15043 ( .A1(n11798), .A2(n11797), .ZN(n11796) );
  NAND2_X1 U15044 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18100), .ZN(
        n18099) );
  NAND2_X1 U15045 ( .A1(n11801), .A2(n11800), .ZN(n19230) );
  INV_X1 U15046 ( .A(n14440), .ZN(n18568) );
  NOR2_X1 U15047 ( .A1(n18568), .A2(n17575), .ZN(n19016) );
  NAND3_X1 U15048 ( .A1(n11804), .A2(n11802), .A3(n19016), .ZN(n14438) );
  INV_X1 U15049 ( .A(n11804), .ZN(n11807) );
  INV_X1 U15050 ( .A(n11805), .ZN(n11806) );
  NAND3_X1 U15051 ( .A1(n11807), .A2(n19215), .A3(n11806), .ZN(n11808) );
  NAND2_X1 U15052 ( .A1(n11809), .A2(n11808), .ZN(n19014) );
  NOR2_X1 U15053 ( .A1(n19004), .A2(n11810), .ZN(n18267) );
  INV_X1 U15054 ( .A(n18267), .ZN(n18398) );
  INV_X1 U15055 ( .A(n18399), .ZN(n18039) );
  OAI22_X1 U15056 ( .A1(n18021), .A2(n18397), .B1(n18398), .B2(n18039), .ZN(
        n18313) );
  AOI21_X1 U15057 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18495) );
  NAND3_X1 U15058 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18312) );
  NOR2_X1 U15059 ( .A1(n18495), .A2(n18312), .ZN(n18433) );
  NAND2_X1 U15060 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18436) );
  INV_X1 U15061 ( .A(n18436), .ZN(n11811) );
  NAND3_X1 U15062 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18433), .A3(
        n11811), .ZN(n18401) );
  NAND2_X1 U15063 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18478) );
  NOR2_X1 U15064 ( .A1(n18312), .A2(n18478), .ZN(n18432) );
  NAND2_X1 U15065 ( .A1(n11811), .A2(n18432), .ZN(n18423) );
  INV_X1 U15066 ( .A(n18423), .ZN(n18336) );
  NAND2_X1 U15067 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18336), .ZN(
        n11822) );
  NAND2_X1 U15068 ( .A1(n19038), .A2(n19195), .ZN(n18517) );
  NOR2_X1 U15069 ( .A1(n19020), .A2(n19036), .ZN(n18431) );
  INV_X1 U15070 ( .A(n18431), .ZN(n18477) );
  NAND2_X1 U15071 ( .A1(n18517), .A2(n18477), .ZN(n18496) );
  OAI22_X1 U15072 ( .A1(n19031), .A2(n18401), .B1(n11822), .B2(n18496), .ZN(
        n11812) );
  OAI21_X1 U15073 ( .B1(n18313), .B2(n11812), .A(n16773), .ZN(n18262) );
  NOR2_X1 U15074 ( .A1(n18530), .A2(n18262), .ZN(n18279) );
  INV_X1 U15075 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18250) );
  NOR2_X1 U15076 ( .A1(n17908), .A2(n18250), .ZN(n18203) );
  INV_X1 U15077 ( .A(n18203), .ZN(n11828) );
  NOR2_X1 U15078 ( .A1(n11828), .A2(n18204), .ZN(n11826) );
  NAND3_X1 U15079 ( .A1(n11827), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n11826), .ZN(n11824) );
  INV_X1 U15080 ( .A(n11824), .ZN(n11813) );
  INV_X1 U15081 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17849) );
  OAI211_X1 U15082 ( .C1(n11814), .C2(n18279), .A(n11813), .B(n17849), .ZN(
        n11837) );
  NOR2_X1 U15083 ( .A1(n11816), .A2(n11815), .ZN(n11819) );
  INV_X1 U15084 ( .A(n11817), .ZN(n11818) );
  NAND2_X1 U15085 ( .A1(n17835), .A2(n11820), .ZN(n11832) );
  INV_X1 U15086 ( .A(n18397), .ZN(n18999) );
  INV_X1 U15087 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21186) );
  NOR2_X1 U15088 ( .A1(n17849), .A2(n21186), .ZN(n16775) );
  NAND2_X1 U15089 ( .A1(n18203), .A2(n18240), .ZN(n17879) );
  NAND2_X1 U15090 ( .A1(n16775), .A2(n18211), .ZN(n16784) );
  OR2_X1 U15091 ( .A1(n18314), .A2(n11822), .ZN(n18315) );
  NOR2_X1 U15092 ( .A1(n11821), .A2(n18315), .ZN(n18242) );
  NOR2_X1 U15093 ( .A1(n19195), .A2(n11822), .ZN(n18422) );
  INV_X1 U15094 ( .A(n18422), .ZN(n18403) );
  NOR2_X1 U15095 ( .A1(n18314), .A2(n18403), .ZN(n18282) );
  INV_X1 U15096 ( .A(n18282), .ZN(n18337) );
  NOR2_X1 U15097 ( .A1(n18314), .A2(n18401), .ZN(n18266) );
  NAND2_X1 U15098 ( .A1(n18317), .A2(n18266), .ZN(n18319) );
  NOR2_X1 U15099 ( .A1(n11823), .A2(n18319), .ZN(n18245) );
  AOI21_X1 U15100 ( .B1(n18245), .B2(n11826), .A(n19031), .ZN(n18207) );
  AOI221_X1 U15101 ( .B1(n18337), .B2(n19036), .C1(n11824), .C2(n19036), .A(
        n18207), .ZN(n11825) );
  OAI221_X1 U15102 ( .B1(n19038), .B2(n11826), .C1(n19038), .C2(n18242), .A(
        n11825), .ZN(n16192) );
  INV_X1 U15103 ( .A(n18413), .ZN(n18407) );
  OAI21_X1 U15104 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18407), .A(
        n18513), .ZN(n16104) );
  AOI211_X1 U15105 ( .C1(n18999), .C2(n16784), .A(n16192), .B(n16104), .ZN(
        n11830) );
  NAND2_X1 U15106 ( .A1(n18399), .A2(n18346), .ZN(n18020) );
  NAND2_X1 U15107 ( .A1(n18263), .A2(n11827), .ZN(n17907) );
  NOR2_X1 U15108 ( .A1(n11828), .A2(n17907), .ZN(n17878) );
  INV_X1 U15109 ( .A(n18204), .ZN(n18205) );
  NAND2_X1 U15110 ( .A1(n17878), .A2(n18205), .ZN(n18208) );
  NAND2_X1 U15111 ( .A1(n17840), .A2(n16775), .ZN(n16781) );
  INV_X1 U15112 ( .A(n16781), .ZN(n16758) );
  OR2_X1 U15113 ( .A1(n16758), .A2(n18398), .ZN(n11829) );
  AND2_X1 U15114 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  NAND2_X1 U15115 ( .A1(n11832), .A2(n11831), .ZN(n11833) );
  NAND3_X1 U15116 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18418), .A3(
        n11833), .ZN(n11836) );
  OR3_X1 U15117 ( .A1(n11834), .A2(n18325), .A3(n17837), .ZN(n11835) );
  NAND2_X1 U15118 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18523), .ZN(n17845) );
  NAND4_X1 U15119 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n17845), .ZN(
        P3_U2834) );
  INV_X1 U15120 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11838) );
  INV_X1 U15121 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11839) );
  AND2_X2 U15122 ( .A1(n11848), .A2(n11850), .ZN(n12111) );
  NOR2_X4 U15123 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14032) );
  AND2_X2 U15124 ( .A1(n11850), .A2(n14032), .ZN(n12009) );
  AOI22_X1 U15125 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11843) );
  AND2_X2 U15126 ( .A1(n11850), .A2(n13638), .ZN(n11889) );
  AND2_X2 U15127 ( .A1(n11847), .A2(n13638), .ZN(n12798) );
  AOI22_X1 U15128 ( .A1(n11889), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11842) );
  AND2_X2 U15129 ( .A1(n13644), .A2(n14032), .ZN(n11939) );
  AND2_X4 U15130 ( .A1(n14032), .A2(n11846), .ZN(n12952) );
  AOI22_X1 U15131 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15132 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U15133 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11854) );
  AND2_X2 U15134 ( .A1(n11845), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11849) );
  AOI22_X1 U15136 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11853) );
  AND2_X2 U15137 ( .A1(n11847), .A2(n14032), .ZN(n11993) );
  AOI22_X1 U15138 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11852) );
  AND2_X2 U15139 ( .A1(n11850), .A2(n11849), .ZN(n11944) );
  AOI22_X1 U15140 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11851) );
  NAND3_X1 U15141 ( .A1(n10270), .A2(n11854), .A3(n10267), .ZN(n12017) );
  AOI22_X1 U15142 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U15143 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U15144 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U15145 ( .A1(n11889), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11855) );
  NAND4_X1 U15146 ( .A1(n11858), .A2(n11857), .A3(n11856), .A4(n11855), .ZN(
        n11864) );
  AOI22_X1 U15147 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U15148 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U15149 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11860) );
  BUF_X2 U15150 ( .A(n12032), .Z(n12948) );
  AOI22_X1 U15151 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11859) );
  NAND4_X1 U15152 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11863) );
  AOI22_X1 U15153 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U15154 ( .A1(n11889), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U15155 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11866) );
  BUF_X2 U15156 ( .A(n12111), .Z(n12612) );
  AOI22_X1 U15157 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U15158 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12004), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U15159 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U15160 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15161 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11869) );
  NAND2_X2 U15162 ( .A1(n10268), .A2(n10269), .ZN(n13665) );
  NAND2_X1 U15163 ( .A1(n12435), .A2(n13665), .ZN(n11884) );
  AOI22_X1 U15164 ( .A1(n11889), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U15165 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12957), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15166 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11844), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U15167 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11902), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U15168 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U15169 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12004), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15170 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15171 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12009), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U15172 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U15173 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U15174 ( .A1(n12957), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U15175 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U15176 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11895) );
  AOI22_X1 U15177 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11889), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15178 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U15179 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15180 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11890) );
  NAND4_X1 U15181 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11894) );
  NAND2_X1 U15182 ( .A1(n11958), .A2(n12017), .ZN(n11909) );
  INV_X1 U15183 ( .A(n11909), .ZN(n11896) );
  AOI22_X1 U15184 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11889), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U15185 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U15186 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15187 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U15188 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11908) );
  AOI22_X1 U15189 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15190 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15191 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15192 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11903) );
  NAND4_X1 U15193 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11907) );
  OR2_X2 U15194 ( .A1(n11908), .A2(n11907), .ZN(n12138) );
  NAND3_X2 U15195 ( .A1(n11911), .A2(n11910), .A3(n10271), .ZN(n11979) );
  NAND2_X1 U15196 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11915) );
  NAND2_X1 U15197 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U15198 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11913) );
  NAND2_X1 U15199 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11912) );
  BUF_X4 U15200 ( .A(n11934), .Z(n12804) );
  NAND2_X1 U15201 ( .A1(n12804), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U15202 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11918) );
  NAND2_X1 U15203 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U15204 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15205 ( .A1(n11889), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15206 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U15207 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U15208 ( .A1(n9727), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15209 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15210 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U15211 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U15212 ( .A1(n11993), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11925) );
  NAND4_X4 U15213 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n14157) );
  NAND2_X1 U15214 ( .A1(n12435), .A2(n9720), .ZN(n11933) );
  NAND2_X1 U15215 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15216 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15217 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U15218 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15219 ( .A1(n11889), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11943) );
  NAND2_X1 U15220 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11942) );
  NAND2_X1 U15221 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U15222 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11940) );
  AND4_X2 U15223 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11955) );
  NAND2_X1 U15224 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U15225 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U15226 ( .A1(n11993), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11945) );
  NAND2_X1 U15227 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11952) );
  NAND2_X1 U15228 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U15229 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U15230 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11949) );
  NAND4_X4 U15231 ( .A1(n11956), .A2(n11955), .A3(n11954), .A4(n11953), .ZN(
        n14156) );
  NAND2_X1 U15232 ( .A1(n12311), .A2(n11972), .ZN(n12319) );
  INV_X1 U15233 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20982) );
  XNOR2_X1 U15234 ( .A(n20982), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12252) );
  NAND2_X1 U15235 ( .A1(n11962), .A2(n11957), .ZN(n11959) );
  AND2_X2 U15236 ( .A1(n11959), .A2(n11958), .ZN(n12306) );
  NAND2_X1 U15237 ( .A1(n11967), .A2(n11962), .ZN(n11960) );
  OAI21_X1 U15238 ( .B1(n12252), .B2(n14156), .A(n12318), .ZN(n11963) );
  NAND3_X1 U15239 ( .A1(n12319), .A2(n11963), .A3(n12431), .ZN(n11964) );
  NAND2_X1 U15240 ( .A1(n11964), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U15241 ( .A1(n13786), .A2(n11965), .ZN(n12439) );
  NAND2_X1 U15242 ( .A1(n13962), .A2(n11967), .ZN(n11968) );
  OAI21_X1 U15243 ( .B1(n11979), .B2(n11970), .A(n9720), .ZN(n11974) );
  NAND2_X1 U15244 ( .A1(n13665), .A2(n14157), .ZN(n11971) );
  NAND2_X2 U15245 ( .A1(n9743), .A2(n14157), .ZN(n21059) );
  NAND2_X1 U15246 ( .A1(n9720), .A2(n14156), .ZN(n14173) );
  OAI21_X1 U15247 ( .B1(n21059), .B2(n11967), .A(n14173), .ZN(n11973) );
  NOR2_X2 U15248 ( .A1(n13631), .A2(n11973), .ZN(n11982) );
  NAND4_X1 U15249 ( .A1(n12439), .A2(n11988), .A3(n11974), .A4(n11982), .ZN(
        n11975) );
  NAND2_X1 U15250 ( .A1(n11975), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U15251 ( .A1(n12057), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11978) );
  INV_X1 U15252 ( .A(n16179), .ZN(n16173) );
  NAND2_X1 U15253 ( .A1(n16471), .A2(n9919), .ZN(n12983) );
  MUX2_X1 U15254 ( .A(n16173), .B(n12983), .S(n20905), .Z(n11977) );
  INV_X1 U15255 ( .A(n11980), .ZN(n14154) );
  NAND3_X1 U15256 ( .A1(n13962), .A2(n14154), .A3(n12138), .ZN(n11981) );
  NAND2_X1 U15257 ( .A1(n11979), .A2(n11981), .ZN(n11992) );
  INV_X1 U15258 ( .A(n11982), .ZN(n11987) );
  NAND2_X1 U15259 ( .A1(n11970), .A2(n14024), .ZN(n12446) );
  INV_X1 U15260 ( .A(n21059), .ZN(n12207) );
  NAND2_X1 U15261 ( .A1(n11984), .A2(n12207), .ZN(n11985) );
  NAND4_X1 U15262 ( .A1(n12446), .A2(n11985), .A3(n16471), .A4(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11986) );
  NOR2_X1 U15263 ( .A1(n11987), .A2(n11986), .ZN(n11991) );
  INV_X1 U15264 ( .A(n11988), .ZN(n11989) );
  NAND2_X1 U15265 ( .A1(n11989), .A2(n14156), .ZN(n11990) );
  XNOR2_X1 U15266 ( .A(n12049), .B(n12047), .ZN(n12497) );
  NAND2_X1 U15267 ( .A1(n12497), .A2(n9919), .ZN(n12020) );
  AOI22_X1 U15268 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15269 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15270 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11995) );
  INV_X2 U15271 ( .A(n12870), .ZN(n12949) );
  AOI22_X1 U15272 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11994) );
  NAND4_X1 U15273 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n12003) );
  AOI22_X1 U15274 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15275 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15276 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15277 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U15278 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12002) );
  INV_X1 U15279 ( .A(n12142), .ZN(n12016) );
  AOI22_X1 U15280 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15281 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15282 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15283 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U15284 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12015) );
  INV_X1 U15285 ( .A(n12009), .ZN(n12027) );
  AOI22_X1 U15286 ( .A1(n12009), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15287 ( .A1(n12804), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15288 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15289 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12010) );
  NAND4_X1 U15290 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12014) );
  XNOR2_X1 U15291 ( .A(n12016), .B(n12206), .ZN(n12018) );
  NAND2_X1 U15292 ( .A1(n12018), .A2(n12134), .ZN(n12019) );
  NAND2_X1 U15293 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12024) );
  INV_X1 U15294 ( .A(n12206), .ZN(n12040) );
  NAND2_X1 U15295 ( .A1(n9720), .A2(n12142), .ZN(n12021) );
  OAI211_X1 U15296 ( .C1(n12040), .C2(n13954), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n12021), .ZN(n12022) );
  INV_X1 U15297 ( .A(n12022), .ZN(n12023) );
  NAND2_X1 U15298 ( .A1(n12137), .A2(n12136), .ZN(n12026) );
  NAND2_X1 U15299 ( .A1(n12134), .A2(n12206), .ZN(n12025) );
  NAND2_X1 U15300 ( .A1(n12026), .A2(n12025), .ZN(n12044) );
  NOR2_X1 U15301 ( .A1(n9717), .A2(n9919), .ZN(n12039) );
  AOI22_X1 U15302 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15303 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15304 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15305 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U15306 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12038) );
  AOI22_X1 U15307 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15308 ( .A1(n12804), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15309 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15310 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U15311 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12037) );
  AOI22_X1 U15312 ( .A1(n12134), .A2(n12040), .B1(n12039), .B2(n12141), .ZN(
        n12042) );
  NAND2_X1 U15313 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U15314 ( .A1(n12042), .A2(n12041), .ZN(n12043) );
  NAND2_X1 U15315 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12059) );
  OAI21_X1 U15316 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n12059), .ZN(n20741) );
  NAND2_X1 U15317 ( .A1(n16179), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12052) );
  OAI21_X1 U15318 ( .B1(n12983), .B2(n20741), .A(n12052), .ZN(n12045) );
  INV_X1 U15319 ( .A(n12047), .ZN(n12048) );
  NAND2_X1 U15320 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  NAND2_X1 U15321 ( .A1(n13920), .A2(n12050), .ZN(n20548) );
  NAND2_X1 U15322 ( .A1(n12134), .A2(n12141), .ZN(n12051) );
  NAND2_X1 U15323 ( .A1(n12052), .A2(n14633), .ZN(n12053) );
  NAND2_X1 U15324 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  NAND2_X1 U15325 ( .A1(n12077), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12062) );
  INV_X1 U15326 ( .A(n12983), .ZN(n12079) );
  INV_X1 U15327 ( .A(n12059), .ZN(n12058) );
  NAND2_X1 U15328 ( .A1(n12058), .A2(n20653), .ZN(n20618) );
  NAND2_X1 U15329 ( .A1(n12059), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12060) );
  NAND2_X1 U15330 ( .A1(n20618), .A2(n12060), .ZN(n14345) );
  AOI22_X1 U15331 ( .A1(n12079), .A2(n14345), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16179), .ZN(n12061) );
  AOI22_X1 U15332 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12912), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15333 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15334 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15335 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12065) );
  NAND4_X1 U15336 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12074) );
  AOI22_X1 U15337 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12009), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15338 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15339 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15340 ( .A1(n9735), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12069) );
  NAND4_X1 U15341 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12073) );
  AOI22_X1 U15342 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12271), .B2(n12162), .ZN(n12075) );
  NAND2_X1 U15343 ( .A1(n12076), .A2(n12152), .ZN(n12160) );
  NAND2_X1 U15344 ( .A1(n12077), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12081) );
  NAND3_X1 U15345 ( .A1(n20740), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20711) );
  NAND2_X1 U15346 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14293), .ZN(
        n14315) );
  NAND2_X1 U15347 ( .A1(n20740), .A2(n14315), .ZN(n12078) );
  NAND3_X1 U15348 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14338) );
  INV_X1 U15349 ( .A(n14338), .ZN(n13921) );
  NAND2_X1 U15350 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13921), .ZN(
        n14027) );
  AOI22_X1 U15351 ( .A1(n12079), .A2(n20742), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16179), .ZN(n12080) );
  AOI22_X1 U15352 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15353 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15354 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15355 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12082) );
  NAND4_X1 U15356 ( .A1(n12085), .A2(n12084), .A3(n12083), .A4(n12082), .ZN(
        n12091) );
  AOI22_X1 U15357 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15358 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15359 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15360 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12086) );
  NAND4_X1 U15361 ( .A1(n12089), .A2(n12088), .A3(n12087), .A4(n12086), .ZN(
        n12090) );
  AOI22_X1 U15362 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12271), .B2(n12171), .ZN(n12092) );
  NAND2_X1 U15363 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12105) );
  AOI22_X1 U15364 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15365 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15366 ( .A1(n12804), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15367 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12094) );
  NAND4_X1 U15368 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        n12103) );
  AOI22_X1 U15369 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15370 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15371 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15372 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12098) );
  NAND4_X1 U15373 ( .A1(n12101), .A2(n12100), .A3(n12099), .A4(n12098), .ZN(
        n12102) );
  NAND2_X1 U15374 ( .A1(n12271), .A2(n12179), .ZN(n12104) );
  INV_X1 U15375 ( .A(n12292), .ZN(n12283) );
  INV_X1 U15376 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15377 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12110) );
  INV_X1 U15378 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U15379 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15380 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15381 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15382 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12117) );
  AOI22_X1 U15383 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15384 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12114) );
  INV_X1 U15385 ( .A(n12868), .ZN(n12799) );
  AOI22_X1 U15386 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15387 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12112) );
  NAND4_X1 U15388 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12116) );
  NAND2_X1 U15389 ( .A1(n12271), .A2(n12188), .ZN(n12118) );
  NAND2_X1 U15390 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12131) );
  AOI22_X1 U15391 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15392 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15393 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15394 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15395 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12129) );
  AOI22_X1 U15396 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12613), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15397 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15398 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15399 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12124) );
  NAND4_X1 U15400 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12128) );
  NAND2_X1 U15401 ( .A1(n12271), .A2(n12200), .ZN(n12130) );
  AND3_X1 U15402 ( .A1(n12134), .A2(n12256), .A3(n12206), .ZN(n12135) );
  NAND2_X1 U15403 ( .A1(n9720), .A2(n12138), .ZN(n12154) );
  INV_X1 U15404 ( .A(n12139), .ZN(n12140) );
  INV_X1 U15405 ( .A(n12256), .ZN(n12147) );
  NAND2_X1 U15406 ( .A1(n12141), .A2(n12142), .ZN(n12164) );
  OAI21_X1 U15407 ( .B1(n12142), .B2(n12141), .A(n12164), .ZN(n12144) );
  INV_X1 U15408 ( .A(n11965), .ZN(n12143) );
  OAI211_X1 U15409 ( .C1(n12144), .C2(n21059), .A(n12143), .B(n14661), .ZN(
        n12145) );
  INV_X1 U15410 ( .A(n12145), .ZN(n12146) );
  INV_X1 U15411 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20498) );
  INV_X1 U15412 ( .A(n12149), .ZN(n13612) );
  NOR2_X2 U15413 ( .A1(n14667), .A2(n12151), .ZN(n12157) );
  XNOR2_X1 U15414 ( .A(n12164), .B(n12162), .ZN(n12156) );
  XNOR2_X1 U15415 ( .A(n12153), .B(n12152), .ZN(n12481) );
  NAND2_X1 U15416 ( .A1(n12481), .A2(n12256), .ZN(n12155) );
  INV_X1 U15417 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20511) );
  OR2_X1 U15418 ( .A1(n12157), .A2(n20511), .ZN(n12158) );
  NAND2_X1 U15419 ( .A1(n12160), .A2(n14284), .ZN(n12161) );
  INV_X1 U15420 ( .A(n12162), .ZN(n12163) );
  NAND2_X1 U15421 ( .A1(n12164), .A2(n12163), .ZN(n12172) );
  XNOR2_X1 U15422 ( .A(n12172), .B(n12171), .ZN(n12165) );
  OAI22_X1 U15423 ( .A1(n20515), .A2(n12147), .B1(n21059), .B2(n12165), .ZN(
        n14220) );
  NAND2_X1 U15424 ( .A1(n14218), .A2(n14220), .ZN(n14219) );
  NAND2_X2 U15425 ( .A1(n14219), .A2(n12167), .ZN(n12175) );
  XNOR2_X1 U15426 ( .A(n12170), .B(n12169), .ZN(n12515) );
  INV_X1 U15427 ( .A(n12515), .ZN(n12174) );
  NAND2_X1 U15428 ( .A1(n12172), .A2(n12171), .ZN(n12181) );
  XOR2_X1 U15429 ( .A(n12179), .B(n12181), .Z(n12173) );
  OAI22_X1 U15430 ( .A1(n12174), .A2(n12147), .B1(n12173), .B2(n21059), .ZN(
        n14429) );
  INV_X1 U15431 ( .A(n12175), .ZN(n12176) );
  INV_X1 U15432 ( .A(n12179), .ZN(n12180) );
  NOR2_X1 U15433 ( .A1(n12181), .A2(n12180), .ZN(n12189) );
  XOR2_X1 U15434 ( .A(n12188), .B(n12189), .Z(n12182) );
  AOI22_X1 U15435 ( .A1(n12530), .A2(n12256), .B1(n12207), .B2(n12182), .ZN(
        n12183) );
  XNOR2_X1 U15436 ( .A(n12183), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16363) );
  INV_X1 U15437 ( .A(n12183), .ZN(n12184) );
  INV_X1 U15438 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16465) );
  NAND2_X1 U15439 ( .A1(n12186), .A2(n12187), .ZN(n12531) );
  NAND3_X1 U15440 ( .A1(n12198), .A2(n12531), .A3(n12256), .ZN(n12192) );
  NAND2_X1 U15441 ( .A1(n12189), .A2(n12188), .ZN(n12199) );
  XNOR2_X1 U15442 ( .A(n12199), .B(n12200), .ZN(n12190) );
  NAND2_X1 U15443 ( .A1(n12190), .A2(n12207), .ZN(n12191) );
  NAND2_X1 U15444 ( .A1(n12192), .A2(n12191), .ZN(n14582) );
  INV_X1 U15445 ( .A(n14582), .ZN(n12193) );
  INV_X1 U15446 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U15447 ( .A1(n12271), .A2(n12206), .ZN(n12195) );
  OAI21_X1 U15448 ( .B1(n12283), .B2(n12196), .A(n12195), .ZN(n12197) );
  INV_X1 U15449 ( .A(n12199), .ZN(n12201) );
  NAND2_X1 U15450 ( .A1(n12201), .A2(n12200), .ZN(n12205) );
  XNOR2_X1 U15451 ( .A(n12205), .B(n12206), .ZN(n12202) );
  AND2_X1 U15452 ( .A1(n12202), .A2(n12207), .ZN(n12203) );
  AOI21_X1 U15453 ( .B1(n12541), .B2(n12256), .A(n12203), .ZN(n12204) );
  INV_X1 U15454 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16458) );
  NAND2_X1 U15455 ( .A1(n12204), .A2(n16458), .ZN(n16356) );
  INV_X4 U15456 ( .A(n21407), .ZN(n12230) );
  INV_X1 U15457 ( .A(n12205), .ZN(n12208) );
  NAND3_X1 U15458 ( .A1(n12208), .A2(n12207), .A3(n12206), .ZN(n12209) );
  INV_X1 U15459 ( .A(n15151), .ZN(n12210) );
  INV_X1 U15460 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12358) );
  NOR2_X1 U15461 ( .A1(n12232), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12212) );
  NAND2_X1 U15462 ( .A1(n21407), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16330) );
  INV_X1 U15463 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16399) );
  NAND2_X1 U15464 ( .A1(n12230), .A2(n16399), .ZN(n12213) );
  NAND2_X1 U15465 ( .A1(n16330), .A2(n12213), .ZN(n15130) );
  INV_X1 U15466 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16420) );
  NAND2_X1 U15467 ( .A1(n12230), .A2(n16420), .ZN(n15128) );
  NAND2_X1 U15468 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U15469 ( .A1(n12230), .A2(n12214), .ZN(n15126) );
  NAND2_X1 U15470 ( .A1(n15128), .A2(n15126), .ZN(n12215) );
  NOR2_X1 U15471 ( .A1(n15130), .A2(n12215), .ZN(n16328) );
  INV_X1 U15472 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12374) );
  NAND2_X1 U15473 ( .A1(n12230), .A2(n12374), .ZN(n12216) );
  NAND2_X1 U15474 ( .A1(n16328), .A2(n12216), .ZN(n16309) );
  NAND2_X1 U15475 ( .A1(n21407), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12217) );
  NAND2_X1 U15476 ( .A1(n16330), .A2(n12217), .ZN(n16310) );
  INV_X1 U15477 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12218) );
  NOR2_X1 U15478 ( .A1(n12230), .A2(n12218), .ZN(n16313) );
  NOR2_X1 U15479 ( .A1(n16310), .A2(n16313), .ZN(n12221) );
  NAND2_X1 U15480 ( .A1(n12230), .A2(n12218), .ZN(n16314) );
  AOI21_X1 U15481 ( .B1(n16309), .B2(n12221), .A(n12219), .ZN(n15113) );
  INV_X1 U15482 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15114) );
  INV_X1 U15483 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15292) );
  AOI21_X1 U15484 ( .B1(n15114), .B2(n15292), .A(n12230), .ZN(n12220) );
  INV_X1 U15485 ( .A(n12221), .ZN(n12223) );
  OAI21_X1 U15486 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n21407), .ZN(n15124) );
  NAND2_X1 U15487 ( .A1(n21407), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15127) );
  NAND2_X1 U15488 ( .A1(n15124), .A2(n15127), .ZN(n16329) );
  XNOR2_X1 U15489 ( .A(n15063), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15107) );
  INV_X1 U15490 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21077) );
  INV_X1 U15491 ( .A(n12224), .ZN(n12225) );
  INV_X1 U15492 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15244) );
  INV_X1 U15493 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15256) );
  AND2_X1 U15494 ( .A1(n15244), .A2(n15256), .ZN(n12226) );
  AND2_X1 U15495 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U15496 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15198) );
  NAND2_X1 U15497 ( .A1(n15033), .A2(n15198), .ZN(n12228) );
  NAND2_X1 U15498 ( .A1(n12227), .A2(n15063), .ZN(n15044) );
  NOR2_X1 U15499 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15046) );
  INV_X1 U15500 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15209) );
  AND2_X1 U15501 ( .A1(n15046), .A2(n15209), .ZN(n15035) );
  AND2_X1 U15502 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12472) );
  INV_X1 U15503 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12234) );
  INV_X1 U15504 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15172) );
  NOR2_X1 U15505 ( .A1(n15172), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12231) );
  INV_X1 U15506 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13686) );
  XNOR2_X1 U15507 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U15508 ( .A1(n12262), .A2(n12250), .ZN(n12236) );
  INV_X1 U15509 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20870) );
  NAND2_X1 U15510 ( .A1(n20870), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12235) );
  NAND2_X1 U15511 ( .A1(n12236), .A2(n12235), .ZN(n12249) );
  NOR2_X1 U15512 ( .A1(n12237), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12238) );
  OAI22_X1 U15513 ( .A1(n12249), .A2(n12238), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20653), .ZN(n12246) );
  NOR2_X1 U15514 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20740), .ZN(
        n12239) );
  OR2_X1 U15515 ( .A1(n12246), .A2(n12239), .ZN(n12241) );
  NAND2_X1 U15516 ( .A1(n20740), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12240) );
  INV_X1 U15517 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16474) );
  NOR2_X1 U15518 ( .A1(n16474), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12242) );
  XNOR2_X1 U15519 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20740), .ZN(
        n12247) );
  XNOR2_X1 U15520 ( .A(n12247), .B(n12246), .ZN(n12286) );
  XNOR2_X1 U15521 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12248) );
  XNOR2_X1 U15522 ( .A(n12249), .B(n12248), .ZN(n12261) );
  XNOR2_X1 U15523 ( .A(n12262), .B(n12250), .ZN(n12274) );
  NOR4_X1 U15524 ( .A1(n12290), .A2(n12286), .A3(n12261), .A4(n12274), .ZN(
        n12251) );
  NOR2_X1 U15525 ( .A1(n12257), .A2(n12251), .ZN(n14703) );
  NAND2_X1 U15526 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21066) );
  NAND2_X1 U15527 ( .A1(n14703), .A2(n21066), .ZN(n13660) );
  AND2_X1 U15528 ( .A1(n12252), .A2(n20992), .ZN(n16197) );
  INV_X1 U15529 ( .A(n16197), .ZN(n13656) );
  AND2_X1 U15530 ( .A1(n14156), .A2(n13656), .ZN(n12253) );
  OR2_X1 U15531 ( .A1(n13660), .A2(n12253), .ZN(n12304) );
  AOI21_X1 U15532 ( .B1(n9809), .B2(n21066), .A(n9720), .ZN(n12255) );
  NOR2_X1 U15533 ( .A1(n21059), .A2(n16197), .ZN(n12254) );
  OAI21_X1 U15534 ( .B1(n12255), .B2(n12254), .A(n14637), .ZN(n12301) );
  NAND2_X1 U15535 ( .A1(n12257), .A2(n12271), .ZN(n12298) );
  INV_X1 U15536 ( .A(n12261), .ZN(n12258) );
  NAND2_X1 U15537 ( .A1(n14016), .A2(n14157), .ZN(n12259) );
  NAND2_X1 U15538 ( .A1(n12259), .A2(n11972), .ZN(n12279) );
  INV_X1 U15539 ( .A(n12279), .ZN(n12260) );
  AOI211_X1 U15540 ( .C1(n12292), .C2(n12261), .A(n12278), .B(n12260), .ZN(
        n12282) );
  INV_X1 U15541 ( .A(n12271), .ZN(n12267) );
  AOI21_X1 U15542 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n11845), .A(
        n12262), .ZN(n12264) );
  INV_X1 U15543 ( .A(n12264), .ZN(n12263) );
  NOR2_X1 U15544 ( .A1(n12267), .A2(n12263), .ZN(n12266) );
  OAI211_X1 U15545 ( .C1(n9720), .C2(n12316), .A(n12264), .B(n12279), .ZN(
        n12265) );
  OAI21_X1 U15546 ( .B1(n12287), .B2(n12266), .A(n12265), .ZN(n12272) );
  INV_X1 U15547 ( .A(n12272), .ZN(n12277) );
  NAND2_X1 U15548 ( .A1(n14016), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12269) );
  OAI21_X1 U15549 ( .B1(n11972), .B2(n12267), .A(n12269), .ZN(n12268) );
  AOI21_X1 U15550 ( .B1(n12292), .B2(n12274), .A(n12268), .ZN(n12273) );
  INV_X1 U15551 ( .A(n12273), .ZN(n12276) );
  NAND2_X1 U15552 ( .A1(n12269), .A2(n14156), .ZN(n12270) );
  AOI22_X1 U15553 ( .A1(n12274), .A2(n12289), .B1(n12273), .B2(n12272), .ZN(
        n12275) );
  AOI21_X1 U15554 ( .B1(n12277), .B2(n12276), .A(n12275), .ZN(n12281) );
  INV_X1 U15555 ( .A(n12278), .ZN(n12280) );
  OAI22_X1 U15556 ( .A1(n12282), .A2(n12281), .B1(n12280), .B2(n12279), .ZN(
        n12285) );
  NAND2_X1 U15557 ( .A1(n12286), .A2(n12283), .ZN(n12284) );
  AOI22_X1 U15558 ( .A1(n12287), .A2(n12286), .B1(n12285), .B2(n12284), .ZN(
        n12295) );
  INV_X1 U15559 ( .A(n12290), .ZN(n12288) );
  NOR2_X1 U15560 ( .A1(n12292), .A2(n12288), .ZN(n12294) );
  INV_X1 U15561 ( .A(n12289), .ZN(n12291) );
  NAND3_X1 U15562 ( .A1(n12292), .A2(n12291), .A3(n12290), .ZN(n12293) );
  OAI21_X1 U15563 ( .B1(n12295), .B2(n12294), .A(n12293), .ZN(n12296) );
  AOI21_X1 U15564 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n9919), .A(
        n12296), .ZN(n12297) );
  NAND2_X1 U15565 ( .A1(n12298), .A2(n12297), .ZN(n12299) );
  NAND2_X1 U15566 ( .A1(n12301), .A2(n13661), .ZN(n12303) );
  MUX2_X1 U15567 ( .A(n12304), .B(n12303), .S(n12302), .Z(n12314) );
  INV_X1 U15568 ( .A(n14621), .ZN(n14615) );
  NAND2_X1 U15569 ( .A1(n14615), .A2(n14156), .ZN(n12305) );
  NOR2_X1 U15570 ( .A1(n14621), .A2(n11965), .ZN(n13637) );
  NOR2_X1 U15571 ( .A1(n11965), .A2(n9720), .ZN(n12445) );
  OR2_X1 U15572 ( .A1(n13637), .A2(n12445), .ZN(n12308) );
  OR2_X1 U15573 ( .A1(n13962), .A2(n13954), .ZN(n12307) );
  AND2_X1 U15574 ( .A1(n12307), .A2(n12306), .ZN(n12440) );
  NAND2_X1 U15575 ( .A1(n12308), .A2(n12440), .ZN(n12317) );
  AOI21_X1 U15576 ( .B1(n11897), .B2(n14156), .A(n9720), .ZN(n12310) );
  AND2_X1 U15577 ( .A1(n12310), .A2(n12309), .ZN(n12438) );
  NOR2_X1 U15578 ( .A1(n12317), .A2(n12438), .ZN(n12313) );
  OR2_X1 U15579 ( .A1(n12313), .A2(n12312), .ZN(n13664) );
  NAND3_X1 U15580 ( .A1(n12314), .A2(n13667), .A3(n13664), .ZN(n12315) );
  NOR2_X1 U15581 ( .A1(n12317), .A2(n12316), .ZN(n14699) );
  INV_X1 U15582 ( .A(n14699), .ZN(n12324) );
  AND2_X1 U15583 ( .A1(n13637), .A2(n11980), .ZN(n14697) );
  AOI21_X1 U15584 ( .B1(n12318), .B2(n14156), .A(n14697), .ZN(n12323) );
  INV_X1 U15585 ( .A(n12431), .ZN(n12321) );
  NAND2_X1 U15586 ( .A1(n12321), .A2(n13954), .ZN(n12322) );
  NAND4_X1 U15587 ( .A1(n12324), .A2(n12323), .A3(n12320), .A4(n12322), .ZN(
        n12325) );
  AND2_X1 U15588 ( .A1(n14054), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12326) );
  AOI21_X1 U15589 ( .B1(n13786), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12326), .ZN(
        n14644) );
  INV_X1 U15590 ( .A(n12345), .ZN(n12332) );
  NAND2_X1 U15591 ( .A1(n12328), .A2(n20498), .ZN(n12330) );
  INV_X1 U15592 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14055) );
  NAND2_X1 U15593 ( .A1(n14155), .A2(n14055), .ZN(n12329) );
  NAND3_X1 U15594 ( .A1(n12330), .A2(n12398), .A3(n12329), .ZN(n12331) );
  NAND2_X1 U15595 ( .A1(n12328), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12334) );
  INV_X1 U15596 ( .A(n12337), .ZN(n12398) );
  INV_X1 U15597 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13979) );
  NAND2_X1 U15598 ( .A1(n12398), .A2(n13979), .ZN(n12333) );
  NAND2_X1 U15599 ( .A1(n12334), .A2(n12333), .ZN(n13787) );
  INV_X1 U15600 ( .A(n12335), .ZN(n12336) );
  AOI21_X1 U15601 ( .B1(n14166), .B2(n14155), .A(n12336), .ZN(n14059) );
  OR2_X1 U15602 ( .A1(n12422), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U15603 ( .A1(n12328), .A2(n20511), .ZN(n12339) );
  INV_X1 U15604 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14212) );
  NAND2_X1 U15605 ( .A1(n14155), .A2(n14212), .ZN(n12338) );
  NAND3_X1 U15606 ( .A1(n12339), .A2(n12398), .A3(n12338), .ZN(n12340) );
  NAND2_X1 U15607 ( .A1(n12341), .A2(n12340), .ZN(n14058) );
  MUX2_X1 U15608 ( .A(n12419), .B(n12398), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12343) );
  OR2_X1 U15609 ( .A1(n13786), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12342) );
  AND2_X1 U15610 ( .A1(n12343), .A2(n12342), .ZN(n14012) );
  INV_X1 U15611 ( .A(n12422), .ZN(n12344) );
  INV_X1 U15612 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20388) );
  NAND2_X1 U15613 ( .A1(n12344), .A2(n20388), .ZN(n12349) );
  NAND2_X1 U15614 ( .A1(n12328), .A2(n12168), .ZN(n12347) );
  NAND2_X1 U15615 ( .A1(n14155), .A2(n20388), .ZN(n12346) );
  NAND3_X1 U15616 ( .A1(n12347), .A2(n12409), .A3(n12346), .ZN(n12348) );
  AND2_X1 U15617 ( .A1(n12349), .A2(n12348), .ZN(n14109) );
  MUX2_X1 U15618 ( .A(n12419), .B(n12398), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12351) );
  OAI21_X1 U15619 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13786), .A(
        n12351), .ZN(n16460) );
  OR2_X1 U15620 ( .A1(n12422), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15621 ( .A1(n12328), .A2(n15301), .ZN(n12353) );
  INV_X1 U15622 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14269) );
  NAND2_X1 U15623 ( .A1(n14155), .A2(n14269), .ZN(n12352) );
  NAND3_X1 U15624 ( .A1(n12353), .A2(n12409), .A3(n12352), .ZN(n12354) );
  NAND2_X1 U15625 ( .A1(n12355), .A2(n12354), .ZN(n14266) );
  MUX2_X1 U15626 ( .A(n12419), .B(n12409), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12356) );
  OAI21_X1 U15627 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n13786), .A(
        n12356), .ZN(n14261) );
  INV_X1 U15628 ( .A(n14261), .ZN(n12357) );
  NAND2_X1 U15629 ( .A1(n14268), .A2(n12357), .ZN(n14258) );
  OR2_X1 U15630 ( .A1(n12422), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U15631 ( .A1(n12328), .A2(n12358), .ZN(n12360) );
  INV_X1 U15632 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14411) );
  NAND2_X1 U15633 ( .A1(n14155), .A2(n14411), .ZN(n12359) );
  NAND3_X1 U15634 ( .A1(n12360), .A2(n12409), .A3(n12359), .ZN(n12361) );
  MUX2_X1 U15635 ( .A(n12419), .B(n12409), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12363) );
  OAI21_X1 U15636 ( .B1(n13786), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12363), .ZN(n14424) );
  NOR2_X2 U15637 ( .A1(n14423), .A2(n14424), .ZN(n14539) );
  OR2_X1 U15638 ( .A1(n12422), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12367) );
  INV_X1 U15639 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16346) );
  NAND2_X1 U15640 ( .A1(n12328), .A2(n16346), .ZN(n12365) );
  INV_X1 U15641 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U15642 ( .A1(n14155), .A2(n14541), .ZN(n12364) );
  NAND3_X1 U15643 ( .A1(n12365), .A2(n12409), .A3(n12364), .ZN(n12366) );
  NAND2_X1 U15644 ( .A1(n12367), .A2(n12366), .ZN(n14538) );
  NAND2_X1 U15645 ( .A1(n14539), .A2(n14538), .ZN(n14600) );
  MUX2_X1 U15646 ( .A(n12419), .B(n12409), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12368) );
  OAI21_X1 U15647 ( .B1(n13786), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12368), .ZN(n14601) );
  OR2_X1 U15648 ( .A1(n12422), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n12372) );
  NAND2_X1 U15649 ( .A1(n12328), .A2(n16420), .ZN(n12370) );
  INV_X1 U15650 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16292) );
  NAND2_X1 U15651 ( .A1(n14155), .A2(n16292), .ZN(n12369) );
  NAND3_X1 U15652 ( .A1(n12370), .A2(n12398), .A3(n12369), .ZN(n12371) );
  MUX2_X1 U15653 ( .A(n12419), .B(n12409), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12373) );
  OAI21_X1 U15654 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13786), .A(
        n12373), .ZN(n14895) );
  OR2_X1 U15655 ( .A1(n12422), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12378) );
  NAND2_X1 U15656 ( .A1(n12328), .A2(n12374), .ZN(n12376) );
  INV_X1 U15657 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21392) );
  NAND2_X1 U15658 ( .A1(n14155), .A2(n21392), .ZN(n12375) );
  NAND3_X1 U15659 ( .A1(n12376), .A2(n12398), .A3(n12375), .ZN(n12377) );
  NAND2_X1 U15660 ( .A1(n12378), .A2(n12377), .ZN(n14889) );
  INV_X1 U15661 ( .A(n12419), .ZN(n12392) );
  INV_X1 U15662 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n16308) );
  NAND2_X1 U15663 ( .A1(n12392), .A2(n16308), .ZN(n12381) );
  INV_X1 U15664 ( .A(n12337), .ZN(n12409) );
  NAND2_X1 U15665 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12379) );
  OAI211_X1 U15666 ( .C1(n14054), .C2(P1_EBX_REG_15__SCAN_IN), .A(n12328), .B(
        n12379), .ZN(n12380) );
  OR2_X1 U15667 ( .A1(n12422), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U15668 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12382) );
  NAND2_X1 U15669 ( .A1(n12328), .A2(n12382), .ZN(n12383) );
  OAI21_X1 U15670 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(n14054), .A(n12383), .ZN(
        n12384) );
  NAND2_X1 U15671 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12386) );
  OAI211_X1 U15672 ( .C1(n14054), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12328), .B(
        n12386), .ZN(n12387) );
  OAI21_X1 U15673 ( .B1(n12419), .B2(P1_EBX_REG_17__SCAN_IN), .A(n12387), .ZN(
        n14874) );
  OR2_X1 U15674 ( .A1(n12422), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n12391) );
  INV_X1 U15675 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15280) );
  NAND2_X1 U15676 ( .A1(n12328), .A2(n15280), .ZN(n12389) );
  INV_X1 U15677 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U15678 ( .A1(n14155), .A2(n14868), .ZN(n12388) );
  NAND3_X1 U15679 ( .A1(n12389), .A2(n12398), .A3(n12388), .ZN(n12390) );
  NAND2_X1 U15680 ( .A1(n12391), .A2(n12390), .ZN(n14865) );
  INV_X1 U15681 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14858) );
  NAND2_X1 U15682 ( .A1(n12392), .A2(n14858), .ZN(n12395) );
  NAND2_X1 U15683 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12393) );
  OAI211_X1 U15684 ( .C1(n14054), .C2(P1_EBX_REG_19__SCAN_IN), .A(n12345), .B(
        n12393), .ZN(n12394) );
  OR2_X1 U15685 ( .A1(n12422), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U15686 ( .A1(n12345), .A2(n15244), .ZN(n12399) );
  INV_X1 U15687 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U15688 ( .A1(n14155), .A2(n12396), .ZN(n12397) );
  NAND3_X1 U15689 ( .A1(n12399), .A2(n12398), .A3(n12397), .ZN(n12400) );
  MUX2_X1 U15690 ( .A(n12419), .B(n12409), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12402) );
  OAI21_X1 U15691 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13786), .A(
        n12402), .ZN(n14849) );
  NOR2_X2 U15692 ( .A1(n9775), .A2(n14849), .ZN(n14851) );
  OR2_X1 U15693 ( .A1(n12422), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15694 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12403) );
  NAND2_X1 U15695 ( .A1(n12345), .A2(n12403), .ZN(n12404) );
  OAI21_X1 U15696 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(n14054), .A(n12404), .ZN(
        n12405) );
  NAND2_X1 U15697 ( .A1(n12406), .A2(n12405), .ZN(n14843) );
  NAND2_X1 U15698 ( .A1(n14851), .A2(n14843), .ZN(n14845) );
  NAND2_X1 U15699 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12407) );
  OAI211_X1 U15700 ( .C1(n14054), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12345), .B(
        n12407), .ZN(n12408) );
  OAI21_X1 U15701 ( .B1(n12419), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12408), .ZN(
        n14804) );
  OR2_X1 U15702 ( .A1(n12422), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12413) );
  NAND2_X1 U15703 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12410) );
  NAND2_X1 U15704 ( .A1(n12345), .A2(n12410), .ZN(n12411) );
  OAI21_X1 U15705 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n14054), .A(n12411), .ZN(
        n12412) );
  OR2_X2 U15706 ( .A1(n14806), .A2(n14787), .ZN(n14789) );
  MUX2_X1 U15707 ( .A(n12419), .B(n12409), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12414) );
  OAI21_X1 U15708 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13786), .A(
        n12414), .ZN(n14773) );
  NOR2_X2 U15709 ( .A1(n14789), .A2(n14773), .ZN(n14774) );
  OR2_X1 U15710 ( .A1(n12422), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12418) );
  NAND2_X1 U15711 ( .A1(n12409), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U15712 ( .A1(n12345), .A2(n12415), .ZN(n12416) );
  OAI21_X1 U15713 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n14054), .A(n12416), .ZN(
        n12417) );
  NAND2_X1 U15714 ( .A1(n12418), .A2(n12417), .ZN(n14759) );
  MUX2_X1 U15715 ( .A(n12419), .B(n12398), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12421) );
  OR2_X1 U15716 ( .A1(n13786), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12420) );
  AND2_X1 U15717 ( .A1(n12421), .A2(n12420), .ZN(n14750) );
  NAND2_X1 U15718 ( .A1(n14761), .A2(n14750), .ZN(n14749) );
  OR2_X1 U15719 ( .A1(n12422), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12425) );
  INV_X1 U15720 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21118) );
  NAND2_X1 U15721 ( .A1(n12345), .A2(n21118), .ZN(n12423) );
  OAI211_X1 U15722 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n14054), .A(n12423), .B(
        n12409), .ZN(n12424) );
  AND2_X1 U15723 ( .A1(n12425), .A2(n12424), .ZN(n14736) );
  INV_X1 U15724 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U15725 ( .A1(n14155), .A2(n14832), .ZN(n12427) );
  OR2_X1 U15726 ( .A1(n13786), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12426) );
  NAND2_X1 U15727 ( .A1(n12426), .A2(n12427), .ZN(n14643) );
  MUX2_X1 U15728 ( .A(n12427), .B(n14643), .S(n12398), .Z(n14720) );
  AOI22_X1 U15729 ( .A1(n13786), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14054), .ZN(n12428) );
  INV_X1 U15730 ( .A(n12428), .ZN(n12429) );
  NAND2_X1 U15731 ( .A1(n12318), .A2(n11972), .ZN(n12430) );
  OAI21_X1 U15732 ( .B1(n12431), .B2(n13954), .A(n12430), .ZN(n12432) );
  AND2_X1 U15733 ( .A1(n12312), .A2(n14156), .ZN(n16154) );
  NAND2_X1 U15734 ( .A1(n12461), .A2(n16154), .ZN(n16396) );
  INV_X1 U15735 ( .A(n11970), .ZN(n12434) );
  INV_X1 U15736 ( .A(n11958), .ZN(n14662) );
  AOI21_X1 U15737 ( .B1(n14024), .B2(n13665), .A(n14662), .ZN(n12433) );
  OAI211_X1 U15738 ( .C1(n12435), .C2(n9717), .A(n12434), .B(n12433), .ZN(
        n12436) );
  AND2_X1 U15739 ( .A1(n12436), .A2(n14156), .ZN(n12437) );
  NOR2_X1 U15740 ( .A1(n12438), .A2(n12437), .ZN(n12444) );
  OAI21_X1 U15741 ( .B1(n12440), .B2(n12409), .A(n12439), .ZN(n12441) );
  INV_X1 U15742 ( .A(n12441), .ZN(n12443) );
  NAND2_X1 U15743 ( .A1(n11979), .A2(n11980), .ZN(n12442) );
  AND3_X1 U15744 ( .A1(n12444), .A2(n12443), .A3(n12442), .ZN(n13634) );
  INV_X1 U15745 ( .A(n12445), .ZN(n13666) );
  INV_X1 U15746 ( .A(n12446), .ZN(n12447) );
  AOI21_X1 U15747 ( .B1(n13666), .B2(n13631), .A(n12447), .ZN(n12448) );
  NAND2_X1 U15748 ( .A1(n13634), .A2(n12448), .ZN(n12449) );
  NAND2_X1 U15749 ( .A1(n12461), .A2(n12449), .ZN(n16385) );
  INV_X1 U15750 ( .A(n16396), .ZN(n12450) );
  NOR2_X1 U15751 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12450), .ZN(
        n14680) );
  NOR2_X1 U15752 ( .A1(n20511), .A2(n20498), .ZN(n14431) );
  NOR2_X1 U15753 ( .A1(n12168), .A2(n12159), .ZN(n16466) );
  NAND2_X1 U15754 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16466), .ZN(
        n12452) );
  INV_X1 U15755 ( .A(n12452), .ZN(n14585) );
  NAND2_X1 U15756 ( .A1(n14431), .A2(n14585), .ZN(n16433) );
  NOR2_X1 U15757 ( .A1(n16420), .A2(n16433), .ZN(n16413) );
  INV_X1 U15758 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12451) );
  NOR2_X1 U15759 ( .A1(n12358), .A2(n16458), .ZN(n16439) );
  NAND4_X1 U15760 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16439), .ZN(n16414) );
  NOR2_X1 U15761 ( .A1(n12451), .A2(n16414), .ZN(n12453) );
  AND2_X1 U15762 ( .A1(n16413), .A2(n12453), .ZN(n16404) );
  INV_X1 U15763 ( .A(n16404), .ZN(n15241) );
  NOR2_X1 U15764 ( .A1(n16399), .A2(n15241), .ZN(n16397) );
  NAND2_X1 U15765 ( .A1(n20493), .A2(n16397), .ZN(n15217) );
  AND2_X1 U15766 ( .A1(n13637), .A2(n14155), .ZN(n14696) );
  AOI21_X1 U15767 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20499) );
  NOR2_X1 U15768 ( .A1(n20499), .A2(n12452), .ZN(n16434) );
  NAND2_X1 U15769 ( .A1(n12453), .A2(n16434), .ZN(n16409) );
  NOR2_X1 U15770 ( .A1(n16420), .A2(n16409), .ZN(n12463) );
  NAND2_X1 U15771 ( .A1(n14433), .A2(n12463), .ZN(n15243) );
  NAND2_X1 U15772 ( .A1(n15217), .A2(n12454), .ZN(n15291) );
  AND2_X1 U15773 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15281) );
  NAND2_X1 U15774 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16368) );
  INV_X1 U15775 ( .A(n16368), .ZN(n15279) );
  AND2_X1 U15776 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15279), .ZN(
        n12455) );
  NAND2_X1 U15777 ( .A1(n15281), .A2(n12455), .ZN(n15238) );
  AND2_X1 U15778 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12469) );
  NAND3_X1 U15779 ( .A1(n12469), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12456) );
  NOR2_X1 U15780 ( .A1(n15238), .A2(n12456), .ZN(n12457) );
  NAND2_X1 U15781 ( .A1(n15291), .A2(n12457), .ZN(n15221) );
  INV_X1 U15782 ( .A(n15198), .ZN(n12458) );
  NAND2_X1 U15783 ( .A1(n12458), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12459) );
  NOR2_X1 U15784 ( .A1(n15221), .A2(n12459), .ZN(n15191) );
  NAND2_X1 U15785 ( .A1(n15191), .A2(n12472), .ZN(n15160) );
  NAND3_X1 U15786 ( .A1(n13686), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12476) );
  OR2_X1 U15787 ( .A1(n12983), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12460) );
  INV_X1 U15788 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14715) );
  NOR2_X1 U15789 ( .A1(n12460), .A2(n14715), .ZN(n12988) );
  INV_X1 U15790 ( .A(n12988), .ZN(n12475) );
  INV_X1 U15791 ( .A(n15300), .ZN(n14681) );
  NOR2_X1 U15792 ( .A1(n16385), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12462) );
  NOR2_X1 U15793 ( .A1(n12461), .A2(n20473), .ZN(n13789) );
  NAND2_X1 U15794 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12463), .ZN(
        n16390) );
  AND2_X1 U15795 ( .A1(n14433), .A2(n16390), .ZN(n12464) );
  NOR2_X1 U15796 ( .A1(n14430), .A2(n12464), .ZN(n16386) );
  NAND2_X1 U15797 ( .A1(n15300), .A2(n15238), .ZN(n12466) );
  INV_X1 U15798 ( .A(n20495), .ZN(n16410) );
  OAI21_X1 U15799 ( .B1(n16399), .B2(n15241), .A(n16410), .ZN(n12465) );
  NAND3_X1 U15800 ( .A1(n16386), .A2(n12466), .A3(n12465), .ZN(n15271) );
  NAND2_X1 U15801 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12467) );
  OR2_X1 U15802 ( .A1(n15271), .A2(n12467), .ZN(n12468) );
  NAND2_X1 U15803 ( .A1(n12468), .A2(n16436), .ZN(n15255) );
  INV_X1 U15804 ( .A(n12469), .ZN(n15245) );
  NAND2_X1 U15805 ( .A1(n15300), .A2(n15245), .ZN(n12470) );
  NAND2_X1 U15806 ( .A1(n15255), .A2(n12470), .ZN(n15228) );
  AND2_X1 U15807 ( .A1(n15300), .A2(n15198), .ZN(n12471) );
  NOR2_X1 U15808 ( .A1(n15228), .A2(n12471), .ZN(n15206) );
  NAND2_X1 U15809 ( .A1(n15206), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15203) );
  INV_X1 U15810 ( .A(n12472), .ZN(n12473) );
  OAI21_X1 U15811 ( .B1(n15203), .B2(n12473), .A(n16436), .ZN(n15169) );
  OAI211_X1 U15812 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14681), .A(
        n15169), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15161) );
  NAND3_X1 U15813 ( .A1(n15161), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16436), .ZN(n12474) );
  OAI211_X1 U15814 ( .C1(n15160), .C2(n12476), .A(n12475), .B(n12474), .ZN(
        n12477) );
  NAND2_X1 U15815 ( .A1(n14699), .A2(n13661), .ZN(n16166) );
  NAND2_X1 U15816 ( .A1(n12480), .A2(n12479), .ZN(n12992) );
  NAND2_X1 U15817 ( .A1(n12481), .A2(n12654), .ZN(n12487) );
  INV_X1 U15818 ( .A(n14637), .ZN(n12482) );
  INV_X1 U15819 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12484) );
  XNOR2_X1 U15820 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14209) );
  AOI21_X1 U15821 ( .B1(n9710), .B2(n14209), .A(n12978), .ZN(n12483) );
  OAI21_X1 U15822 ( .B1(n12943), .B2(n12484), .A(n12483), .ZN(n12485) );
  AOI21_X1 U15823 ( .B1(n12513), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12485), .ZN(n12486) );
  NAND2_X1 U15824 ( .A1(n12487), .A2(n12486), .ZN(n12488) );
  NAND2_X1 U15825 ( .A1(n12978), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12505) );
  NAND2_X1 U15826 ( .A1(n13915), .A2(n12654), .ZN(n12494) );
  INV_X1 U15827 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12491) );
  INV_X1 U15828 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14171) );
  OAI22_X1 U15829 ( .A1(n12943), .A2(n12491), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14171), .ZN(n12492) );
  AOI21_X1 U15830 ( .B1(n12513), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12492), .ZN(n12493) );
  NAND2_X1 U15831 ( .A1(n12494), .A2(n12493), .ZN(n13966) );
  NAND2_X1 U15832 ( .A1(n9729), .A2(n14024), .ZN(n12496) );
  NAND2_X1 U15833 ( .A1(n12496), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13607) );
  INV_X1 U15835 ( .A(n12513), .ZN(n12518) );
  NAND2_X1 U15836 ( .A1(n20913), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12500) );
  NAND2_X1 U15837 ( .A1(n12979), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12499) );
  OAI211_X1 U15838 ( .C1(n12518), .C2(n11845), .A(n12500), .B(n12499), .ZN(
        n12501) );
  AOI21_X1 U15839 ( .B1(n12498), .B2(n12654), .A(n12501), .ZN(n12502) );
  OR2_X1 U15840 ( .A1(n13607), .A2(n12502), .ZN(n13608) );
  INV_X1 U15841 ( .A(n12502), .ZN(n13609) );
  OR2_X1 U15842 ( .A1(n13609), .A2(n12795), .ZN(n12503) );
  NAND2_X1 U15843 ( .A1(n13608), .A2(n12503), .ZN(n13965) );
  INV_X1 U15844 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U15845 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12507) );
  INV_X1 U15846 ( .A(n12507), .ZN(n12509) );
  INV_X1 U15847 ( .A(n12524), .ZN(n12508) );
  OAI21_X1 U15848 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12509), .A(
        n12508), .ZN(n14401) );
  AOI22_X1 U15849 ( .A1(n9710), .A2(n14401), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12510) );
  OAI21_X1 U15850 ( .B1(n12943), .B2(n12511), .A(n12510), .ZN(n12512) );
  AOI21_X1 U15851 ( .B1(n12513), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12512), .ZN(n12514) );
  NAND2_X1 U15852 ( .A1(n13971), .A2(n13972), .ZN(n14008) );
  NAND2_X1 U15853 ( .A1(n12515), .A2(n12654), .ZN(n12521) );
  XNOR2_X1 U15854 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n12524), .ZN(
        n20481) );
  INV_X1 U15855 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20683) );
  OAI21_X1 U15856 ( .B1(n20683), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20913), .ZN(n12517) );
  NAND2_X1 U15857 ( .A1(n12979), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12516) );
  OAI211_X1 U15858 ( .C1(n12518), .C2(n16474), .A(n12517), .B(n12516), .ZN(
        n12519) );
  OAI21_X1 U15859 ( .B1(n12795), .B2(n20481), .A(n12519), .ZN(n12520) );
  INV_X1 U15860 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14236) );
  INV_X1 U15861 ( .A(n12532), .ZN(n12534) );
  INV_X1 U15862 ( .A(n12525), .ZN(n12526) );
  INV_X1 U15863 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20381) );
  NAND2_X1 U15864 ( .A1(n12526), .A2(n20381), .ZN(n12527) );
  NAND2_X1 U15865 ( .A1(n12534), .A2(n12527), .ZN(n20387) );
  AOI22_X1 U15866 ( .A1(n20387), .A2(n9710), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12528) );
  OAI21_X1 U15867 ( .B1(n12943), .B2(n14236), .A(n12528), .ZN(n12529) );
  NAND2_X1 U15868 ( .A1(n12531), .A2(n12654), .ZN(n12540) );
  INV_X1 U15869 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20430) );
  INV_X1 U15870 ( .A(n12542), .ZN(n12536) );
  INV_X1 U15871 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12533) );
  NAND2_X1 U15872 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  NAND2_X1 U15873 ( .A1(n12536), .A2(n12535), .ZN(n20372) );
  AOI22_X1 U15874 ( .A1(n20372), .A2(n9710), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12537) );
  OAI21_X1 U15875 ( .B1(n12943), .B2(n20430), .A(n12537), .ZN(n12538) );
  INV_X1 U15876 ( .A(n12538), .ZN(n12539) );
  NAND2_X1 U15877 ( .A1(n12540), .A2(n12539), .ZN(n14263) );
  AND2_X2 U15878 ( .A1(n14233), .A2(n14263), .ZN(n14255) );
  NAND2_X1 U15879 ( .A1(n12541), .A2(n12654), .ZN(n12547) );
  INV_X1 U15880 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12544) );
  OAI21_X1 U15881 ( .B1(n12542), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12559), .ZN(n20361) );
  AOI22_X1 U15882 ( .A1(n20361), .A2(n9710), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12543) );
  OAI21_X1 U15883 ( .B1(n12943), .B2(n12544), .A(n12543), .ZN(n12545) );
  INV_X1 U15884 ( .A(n12545), .ZN(n12546) );
  NAND2_X1 U15885 ( .A1(n12547), .A2(n12546), .ZN(n14256) );
  INV_X1 U15886 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14394) );
  AOI22_X1 U15887 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15888 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15889 ( .A1(n12804), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15890 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12548) );
  NAND4_X1 U15891 ( .A1(n12551), .A2(n12550), .A3(n12549), .A4(n12548), .ZN(
        n12557) );
  AOI22_X1 U15892 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15893 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15894 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15895 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12552) );
  NAND4_X1 U15896 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12556) );
  OR2_X1 U15897 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  NAND2_X1 U15898 ( .A1(n12654), .A2(n12558), .ZN(n12561) );
  XNOR2_X1 U15899 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12562), .ZN(
        n15156) );
  AOI22_X1 U15900 ( .A1(n9710), .A2(n15156), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12560) );
  OAI211_X1 U15901 ( .C1(n12943), .C2(n14394), .A(n12561), .B(n12560), .ZN(
        n14393) );
  XOR2_X1 U15902 ( .A(n20344), .B(n12577), .Z(n20342) );
  INV_X1 U15903 ( .A(n20342), .ZN(n15147) );
  AOI22_X1 U15904 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12912), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15905 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15906 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15907 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12563) );
  NAND4_X1 U15908 ( .A1(n12566), .A2(n12565), .A3(n12564), .A4(n12563), .ZN(
        n12572) );
  AOI22_X1 U15909 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15910 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15911 ( .A1(n9735), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15912 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12567) );
  NAND4_X1 U15913 ( .A1(n12570), .A2(n12569), .A3(n12568), .A4(n12567), .ZN(
        n12571) );
  NOR2_X1 U15914 ( .A1(n12572), .A2(n12571), .ZN(n12575) );
  NAND2_X1 U15915 ( .A1(n12979), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15916 ( .A1(n12978), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12573) );
  OAI211_X1 U15917 ( .C1(n12671), .C2(n12575), .A(n12574), .B(n12573), .ZN(
        n12576) );
  AOI21_X1 U15918 ( .B1(n15147), .B2(n9710), .A(n12576), .ZN(n14421) );
  XNOR2_X1 U15919 ( .A(n12592), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15139) );
  AOI22_X1 U15920 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15921 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15922 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15923 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12578) );
  NAND4_X1 U15924 ( .A1(n12581), .A2(n12580), .A3(n12579), .A4(n12578), .ZN(
        n12587) );
  AOI22_X1 U15925 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12613), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15926 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15927 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15928 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12582) );
  NAND4_X1 U15929 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12586) );
  NOR2_X1 U15930 ( .A1(n12587), .A2(n12586), .ZN(n12590) );
  NAND2_X1 U15931 ( .A1(n12979), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12589) );
  NAND2_X1 U15932 ( .A1(n12978), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12588) );
  OAI211_X1 U15933 ( .C1(n12671), .C2(n12590), .A(n12589), .B(n12588), .ZN(
        n12591) );
  AOI21_X1 U15934 ( .B1(n15139), .B2(n9710), .A(n12591), .ZN(n14537) );
  INV_X1 U15935 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14986) );
  OAI21_X1 U15936 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12593), .A(
        n12611), .ZN(n16355) );
  AOI22_X1 U15937 ( .A1(n9710), .A2(n16355), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12594) );
  OAI21_X1 U15938 ( .B1(n12943), .B2(n14986), .A(n12594), .ZN(n12595) );
  OAI21_X1 U15939 ( .B1(n12596), .B2(n12595), .A(n12610), .ZN(n14595) );
  INV_X1 U15940 ( .A(n14595), .ZN(n12609) );
  AOI22_X1 U15941 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15942 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15943 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15944 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12597) );
  NAND4_X1 U15945 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12606) );
  AOI22_X1 U15946 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15947 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15948 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15949 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12601) );
  NAND4_X1 U15950 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12605) );
  OR2_X1 U15951 ( .A1(n12606), .A2(n12605), .ZN(n12607) );
  NAND2_X1 U15952 ( .A1(n12654), .A2(n12607), .ZN(n14599) );
  INV_X1 U15953 ( .A(n14599), .ZN(n12608) );
  NAND2_X1 U15954 ( .A1(n12609), .A2(n12608), .ZN(n14596) );
  XOR2_X1 U15955 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12627), .Z(
        n16341) );
  AOI22_X1 U15956 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12742), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15957 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15958 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15959 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12614) );
  NAND4_X1 U15960 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n12623) );
  AOI22_X1 U15961 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15962 ( .A1(n12804), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15963 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15964 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12618) );
  NAND4_X1 U15965 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12622) );
  OR2_X1 U15966 ( .A1(n12623), .A2(n12622), .ZN(n12624) );
  AOI22_X1 U15967 ( .A1(n12654), .A2(n12624), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12626) );
  NAND2_X1 U15968 ( .A1(n12979), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12625) );
  OAI211_X1 U15969 ( .C1(n16341), .C2(n12795), .A(n12626), .B(n12625), .ZN(
        n14604) );
  XNOR2_X1 U15970 ( .A(n12642), .B(n16285), .ZN(n16287) );
  AOI22_X1 U15971 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15972 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15973 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15974 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15975 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12637) );
  AOI22_X1 U15976 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15977 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15978 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15979 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12632) );
  NAND4_X1 U15980 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12636) );
  NOR2_X1 U15981 ( .A1(n12637), .A2(n12636), .ZN(n12640) );
  NAND2_X1 U15982 ( .A1(n12979), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U15983 ( .A1(n12978), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12638) );
  OAI211_X1 U15984 ( .C1(n12671), .C2(n12640), .A(n12639), .B(n12638), .ZN(
        n12641) );
  AOI21_X1 U15985 ( .B1(n16287), .B2(n9710), .A(n12641), .ZN(n14893) );
  XOR2_X1 U15986 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12657), .Z(
        n21388) );
  AOI22_X1 U15987 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15988 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11844), .B1(
        n12742), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U15989 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U15990 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12643) );
  NAND4_X1 U15991 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12652) );
  AOI22_X1 U15992 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12804), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15993 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12928), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15994 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12811), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15995 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12933), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12647) );
  NAND4_X1 U15996 ( .A1(n12650), .A2(n12649), .A3(n12648), .A4(n12647), .ZN(
        n12651) );
  OR2_X1 U15997 ( .A1(n12652), .A2(n12651), .ZN(n12653) );
  AOI22_X1 U15998 ( .A1(n12654), .A2(n12653), .B1(n12978), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12656) );
  NAND2_X1 U15999 ( .A1(n12979), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12655) );
  OAI211_X1 U16000 ( .C1(n21388), .C2(n12795), .A(n12656), .B(n12655), .ZN(
        n14888) );
  INV_X1 U16001 ( .A(n14887), .ZN(n12674) );
  XNOR2_X1 U16002 ( .A(n12675), .B(n16275), .ZN(n16277) );
  AOI22_X1 U16003 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U16004 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U16005 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U16006 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12658) );
  NAND4_X1 U16007 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n12667) );
  AOI22_X1 U16008 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U16009 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U16010 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U16011 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U16012 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12666) );
  NOR2_X1 U16013 ( .A1(n12667), .A2(n12666), .ZN(n12670) );
  NAND2_X1 U16014 ( .A1(n12979), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12669) );
  NAND2_X1 U16015 ( .A1(n12978), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12668) );
  OAI211_X1 U16016 ( .C1(n12671), .C2(n12670), .A(n12669), .B(n12668), .ZN(
        n12672) );
  AOI21_X1 U16017 ( .B1(n16277), .B2(n9710), .A(n12672), .ZN(n14978) );
  OAI21_X1 U16018 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12676), .A(
        n12706), .ZN(n16319) );
  INV_X1 U16019 ( .A(n16319), .ZN(n16266) );
  AOI22_X1 U16020 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U16021 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12679) );
  AOI22_X1 U16022 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U16023 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12677) );
  NAND4_X1 U16024 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        n12686) );
  AOI22_X1 U16025 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12933), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U16026 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U16027 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U16028 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12681) );
  NAND4_X1 U16029 ( .A1(n12684), .A2(n12683), .A3(n12682), .A4(n12681), .ZN(
        n12685) );
  OR2_X1 U16030 ( .A1(n12686), .A2(n12685), .ZN(n12689) );
  INV_X1 U16031 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14968) );
  INV_X1 U16032 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12687) );
  OAI22_X1 U16033 ( .A1(n12943), .A2(n14968), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12687), .ZN(n12688) );
  AOI21_X1 U16034 ( .B1(n12945), .B2(n12689), .A(n12688), .ZN(n12690) );
  MUX2_X1 U16035 ( .A(n16266), .B(n12690), .S(n12795), .Z(n14881) );
  INV_X1 U16036 ( .A(n14881), .ZN(n12691) );
  AOI22_X1 U16037 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U16038 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U16039 ( .A1(n9735), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U16040 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12692) );
  NAND4_X1 U16041 ( .A1(n12695), .A2(n12694), .A3(n12693), .A4(n12692), .ZN(
        n12701) );
  AOI22_X1 U16042 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12742), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U16043 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U16044 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U16045 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12696) );
  NAND4_X1 U16046 ( .A1(n12699), .A2(n12698), .A3(n12697), .A4(n12696), .ZN(
        n12700) );
  OAI21_X1 U16047 ( .B1(n12701), .B2(n12700), .A(n12945), .ZN(n12705) );
  XNOR2_X1 U16048 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12706), .ZN(
        n16251) );
  INV_X1 U16049 ( .A(n12978), .ZN(n12702) );
  OAI22_X1 U16050 ( .A1(n16251), .A2(n12795), .B1(n12702), .B2(n16253), .ZN(
        n12703) );
  AOI21_X1 U16051 ( .B1(n12979), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12703), .ZN(
        n12704) );
  INV_X1 U16052 ( .A(n12757), .ZN(n12710) );
  INV_X1 U16053 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12721) );
  INV_X1 U16054 ( .A(n12707), .ZN(n12708) );
  NAND2_X1 U16055 ( .A1(n12721), .A2(n12708), .ZN(n12709) );
  NAND2_X1 U16056 ( .A1(n12710), .A2(n12709), .ZN(n16245) );
  AOI22_X1 U16057 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U16058 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U16059 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U16060 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12711) );
  NAND4_X1 U16061 ( .A1(n12714), .A2(n12713), .A3(n12712), .A4(n12711), .ZN(
        n12720) );
  AOI22_X1 U16062 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12613), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U16063 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U16064 ( .A1(n9735), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U16065 ( .A1(n12798), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12715) );
  NAND4_X1 U16066 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12719) );
  NOR2_X1 U16067 ( .A1(n12720), .A2(n12719), .ZN(n12725) );
  INV_X1 U16068 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12722) );
  OAI22_X1 U16069 ( .A1(n12943), .A2(n12722), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12721), .ZN(n12723) );
  INV_X1 U16070 ( .A(n12723), .ZN(n12724) );
  OAI21_X1 U16071 ( .B1(n12972), .B2(n12725), .A(n12724), .ZN(n12726) );
  MUX2_X1 U16072 ( .A(n16245), .B(n12726), .S(n12795), .Z(n14863) );
  AND2_X2 U16073 ( .A1(n14861), .A2(n14863), .ZN(n14854) );
  INV_X1 U16074 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16233) );
  XNOR2_X1 U16075 ( .A(n12757), .B(n16233), .ZN(n16231) );
  INV_X1 U16076 ( .A(n16231), .ZN(n15101) );
  AOI22_X1 U16077 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U16078 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U16079 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U16080 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U16081 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12736) );
  AOI22_X1 U16082 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U16083 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U16084 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U16085 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12731) );
  NAND4_X1 U16086 ( .A1(n12734), .A2(n12733), .A3(n12732), .A4(n12731), .ZN(
        n12735) );
  NOR2_X1 U16087 ( .A1(n12736), .A2(n12735), .ZN(n12740) );
  INV_X1 U16088 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12737) );
  OAI22_X1 U16089 ( .A1(n12943), .A2(n12737), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n16233), .ZN(n12738) );
  INV_X1 U16090 ( .A(n12738), .ZN(n12739) );
  OAI21_X1 U16091 ( .B1(n12972), .B2(n12740), .A(n12739), .ZN(n12741) );
  MUX2_X1 U16092 ( .A(n15101), .B(n12741), .S(n12795), .Z(n14855) );
  AOI22_X1 U16093 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12742), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U16094 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U16095 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U16096 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12743) );
  NAND4_X1 U16097 ( .A1(n12746), .A2(n12745), .A3(n12744), .A4(n12743), .ZN(
        n12752) );
  AOI22_X1 U16098 ( .A1(n11844), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U16099 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U16100 ( .A1(n9735), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U16101 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12747) );
  NAND4_X1 U16102 ( .A1(n12750), .A2(n12749), .A3(n12748), .A4(n12747), .ZN(
        n12751) );
  NOR2_X1 U16103 ( .A1(n12752), .A2(n12751), .ZN(n12756) );
  INV_X1 U16104 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21072) );
  OAI21_X1 U16105 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20683), .A(
        n20582), .ZN(n12753) );
  OAI21_X1 U16106 ( .B1(n12943), .B2(n21072), .A(n12753), .ZN(n12754) );
  INV_X1 U16107 ( .A(n12754), .ZN(n12755) );
  OAI21_X1 U16108 ( .B1(n12972), .B2(n12756), .A(n12755), .ZN(n12760) );
  OAI21_X1 U16109 ( .B1(n12758), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12791), .ZN(n15092) );
  OR2_X1 U16110 ( .A1(n15092), .A2(n12795), .ZN(n12759) );
  NAND2_X1 U16111 ( .A1(n12760), .A2(n12759), .ZN(n14819) );
  XNOR2_X1 U16112 ( .A(n12791), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16221) );
  AOI22_X1 U16113 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U16114 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U16115 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U16116 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12761) );
  NAND4_X1 U16117 ( .A1(n12764), .A2(n12763), .A3(n12762), .A4(n12761), .ZN(
        n12770) );
  AOI22_X1 U16118 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U16119 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U16120 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U16121 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12765) );
  NAND4_X1 U16122 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12769) );
  OR2_X1 U16123 ( .A1(n12770), .A2(n12769), .ZN(n12772) );
  INV_X1 U16124 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14946) );
  INV_X1 U16125 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12790) );
  OAI22_X1 U16126 ( .A1(n12943), .A2(n14946), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12790), .ZN(n12771) );
  AOI21_X1 U16127 ( .B1(n12945), .B2(n12772), .A(n12771), .ZN(n12773) );
  MUX2_X1 U16128 ( .A(n16221), .B(n12773), .S(n12795), .Z(n14847) );
  AOI22_X1 U16129 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12935), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16130 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12004), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U16131 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12928), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U16132 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12775) );
  NAND4_X1 U16133 ( .A1(n12778), .A2(n12777), .A3(n12776), .A4(n12775), .ZN(
        n12785) );
  AOI22_X1 U16134 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12934), .B1(
        n12779), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U16135 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U16136 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12933), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12781) );
  AOI22_X1 U16137 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12780) );
  NAND4_X1 U16138 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        n12784) );
  NOR2_X1 U16139 ( .A1(n12785), .A2(n12784), .ZN(n12788) );
  OAI21_X1 U16140 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20683), .A(
        n20582), .ZN(n12787) );
  NAND2_X1 U16141 ( .A1(n12979), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n12786) );
  OAI211_X1 U16142 ( .C1(n12972), .C2(n12788), .A(n12787), .B(n12786), .ZN(
        n12797) );
  INV_X1 U16143 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12789) );
  OAI21_X1 U16144 ( .B1(n12791), .B2(n12790), .A(n12789), .ZN(n12794) );
  AND2_X1 U16145 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U16146 ( .A1(n12794), .A2(n12826), .ZN(n16211) );
  OR2_X1 U16147 ( .A1(n16211), .A2(n12795), .ZN(n12796) );
  NAND2_X1 U16148 ( .A1(n12797), .A2(n12796), .ZN(n14841) );
  AOI22_X1 U16149 ( .A1(n12935), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16150 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12798), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U16151 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12799), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16152 ( .A1(n12933), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12800) );
  NAND4_X1 U16153 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n12810) );
  AOI22_X1 U16154 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U16155 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U16156 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U16157 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12805) );
  NAND4_X1 U16158 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12809) );
  NOR2_X1 U16159 ( .A1(n12810), .A2(n12809), .ZN(n12831) );
  AOI22_X1 U16160 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16161 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16162 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12811), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16163 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12812) );
  NAND4_X1 U16164 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12821) );
  AOI22_X1 U16165 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16166 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U16167 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16168 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U16169 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12820) );
  NOR2_X1 U16170 ( .A1(n12821), .A2(n12820), .ZN(n12830) );
  XOR2_X1 U16171 ( .A(n12831), .B(n12830), .Z(n12824) );
  INV_X1 U16172 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12822) );
  INV_X1 U16173 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21216) );
  OAI22_X1 U16174 ( .A1(n12943), .A2(n12822), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21216), .ZN(n12823) );
  AOI21_X1 U16175 ( .B1(n12945), .B2(n12824), .A(n12823), .ZN(n12828) );
  NAND2_X1 U16176 ( .A1(n12826), .A2(n21216), .ZN(n12827) );
  AND2_X1 U16177 ( .A1(n12845), .A2(n12827), .ZN(n15066) );
  MUX2_X1 U16178 ( .A(n12828), .B(n15066), .S(n9710), .Z(n14802) );
  INV_X1 U16179 ( .A(n14802), .ZN(n12829) );
  NAND2_X1 U16180 ( .A1(n14797), .A2(n12829), .ZN(n14783) );
  NOR2_X1 U16181 ( .A1(n12831), .A2(n12830), .ZN(n12849) );
  AOI22_X1 U16182 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16183 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16184 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16185 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12832) );
  NAND4_X1 U16186 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12841) );
  INV_X1 U16187 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21287) );
  AOI22_X1 U16188 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U16189 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U16190 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16191 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12836) );
  NAND4_X1 U16192 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        n12840) );
  OR2_X1 U16193 ( .A1(n12841), .A2(n12840), .ZN(n12848) );
  INV_X1 U16194 ( .A(n12848), .ZN(n12842) );
  XNOR2_X1 U16195 ( .A(n12849), .B(n12842), .ZN(n12844) );
  INV_X1 U16196 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14930) );
  INV_X1 U16197 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14791) );
  OAI22_X1 U16198 ( .A1(n12943), .A2(n14930), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14791), .ZN(n12843) );
  AOI21_X1 U16199 ( .B1(n12844), .B2(n12945), .A(n12843), .ZN(n12847) );
  NAND2_X1 U16200 ( .A1(n12845), .A2(n14791), .ZN(n12846) );
  AND2_X1 U16201 ( .A1(n12884), .A2(n12846), .ZN(n14790) );
  MUX2_X1 U16202 ( .A(n12847), .B(n14790), .S(n9710), .Z(n14785) );
  NAND2_X1 U16203 ( .A1(n12849), .A2(n12848), .ZN(n12864) );
  AOI22_X1 U16204 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U16205 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U16206 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U16207 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12850) );
  NAND4_X1 U16208 ( .A1(n12853), .A2(n12852), .A3(n12851), .A4(n12850), .ZN(
        n12859) );
  AOI22_X1 U16209 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U16210 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U16211 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16212 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12854) );
  NAND4_X1 U16213 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n12854), .ZN(
        n12858) );
  NOR2_X1 U16214 ( .A1(n12859), .A2(n12858), .ZN(n12865) );
  XOR2_X1 U16215 ( .A(n12864), .B(n12865), .Z(n12861) );
  INV_X1 U16216 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14925) );
  INV_X1 U16217 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14777) );
  OAI22_X1 U16218 ( .A1(n12943), .A2(n14925), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14777), .ZN(n12860) );
  AOI21_X1 U16219 ( .B1(n12861), .B2(n12945), .A(n12860), .ZN(n12862) );
  XNOR2_X1 U16220 ( .A(n12884), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14776) );
  MUX2_X1 U16221 ( .A(n12862), .B(n14776), .S(n9710), .Z(n14770) );
  INV_X1 U16222 ( .A(n14770), .ZN(n12863) );
  NOR2_X1 U16223 ( .A1(n12865), .A2(n12864), .ZN(n12891) );
  INV_X1 U16224 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12866) );
  NOR2_X1 U16225 ( .A1(n12027), .A2(n12866), .ZN(n12872) );
  INV_X1 U16226 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12869) );
  INV_X1 U16227 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12867) );
  OAI22_X1 U16228 ( .A1(n12870), .A2(n12869), .B1(n12868), .B2(n12867), .ZN(
        n12871) );
  AOI211_X1 U16229 ( .C1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .C2(n12935), .A(
        n12872), .B(n12871), .ZN(n12881) );
  AOI22_X1 U16230 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U16231 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16232 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U16233 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U16234 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U16235 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12874) );
  AND4_X1 U16236 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        n12878) );
  NAND4_X1 U16237 ( .A1(n12881), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n12890) );
  XNOR2_X1 U16238 ( .A(n12891), .B(n12890), .ZN(n12883) );
  INV_X1 U16239 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20913) );
  AOI22_X1 U16240 ( .A1(n12979), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20913), .ZN(n12882) );
  OAI21_X1 U16241 ( .B1(n12883), .B2(n12972), .A(n12882), .ZN(n12889) );
  INV_X1 U16242 ( .A(n12884), .ZN(n12885) );
  NAND2_X1 U16243 ( .A1(n12885), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12887) );
  INV_X1 U16244 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U16245 ( .A1(n12887), .A2(n12886), .ZN(n12888) );
  NAND2_X1 U16246 ( .A1(n12921), .A2(n12888), .ZN(n15039) );
  MUX2_X1 U16247 ( .A(n12889), .B(n15039), .S(n9710), .Z(n14757) );
  NAND2_X1 U16248 ( .A1(n12891), .A2(n12890), .ZN(n12906) );
  AOI22_X1 U16249 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16250 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U16251 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U16252 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12892) );
  NAND4_X1 U16253 ( .A1(n12895), .A2(n12894), .A3(n12893), .A4(n12892), .ZN(
        n12901) );
  AOI22_X1 U16254 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16255 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16256 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U16257 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12896) );
  NAND4_X1 U16258 ( .A1(n12899), .A2(n12898), .A3(n12897), .A4(n12896), .ZN(
        n12900) );
  NOR2_X1 U16259 ( .A1(n12901), .A2(n12900), .ZN(n12907) );
  XOR2_X1 U16260 ( .A(n12906), .B(n12907), .Z(n12904) );
  INV_X1 U16261 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14916) );
  INV_X1 U16262 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12902) );
  OAI22_X1 U16263 ( .A1(n12943), .A2(n14916), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12902), .ZN(n12903) );
  AOI21_X1 U16264 ( .B1(n12904), .B2(n12945), .A(n12903), .ZN(n12905) );
  XNOR2_X1 U16265 ( .A(n12921), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15026) );
  MUX2_X1 U16266 ( .A(n12905), .B(n15026), .S(n9710), .Z(n14746) );
  NOR2_X1 U16267 ( .A1(n12907), .A2(n12906), .ZN(n12927) );
  AOI22_X1 U16268 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U16269 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U16270 ( .A1(n9738), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U16271 ( .A1(n12811), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12908) );
  NAND4_X1 U16272 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n12918) );
  AOI22_X1 U16273 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12960), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16274 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U16275 ( .A1(n12949), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12952), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16276 ( .A1(n12912), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12913) );
  NAND4_X1 U16277 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        n12917) );
  OR2_X1 U16278 ( .A1(n12918), .A2(n12917), .ZN(n12926) );
  XNOR2_X1 U16279 ( .A(n12927), .B(n12926), .ZN(n12920) );
  AOI22_X1 U16280 ( .A1(n12979), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20913), .ZN(n12919) );
  OAI21_X1 U16281 ( .B1(n12920), .B2(n12972), .A(n12919), .ZN(n12925) );
  INV_X1 U16282 ( .A(n12921), .ZN(n12922) );
  NAND2_X1 U16283 ( .A1(n12922), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12923) );
  INV_X1 U16284 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U16285 ( .A1(n12923), .A2(n14737), .ZN(n12924) );
  NAND2_X1 U16286 ( .A1(n12974), .A2(n12924), .ZN(n15020) );
  MUX2_X1 U16287 ( .A(n12925), .B(n15020), .S(n9710), .Z(n14733) );
  NAND2_X1 U16288 ( .A1(n12927), .A2(n12926), .ZN(n12967) );
  AOI22_X1 U16289 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U16290 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12960), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16291 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16292 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9727), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12929) );
  NAND4_X1 U16293 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12941) );
  AOI22_X1 U16294 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12933), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16295 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12934), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16296 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12935), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16297 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12936) );
  NAND4_X1 U16298 ( .A1(n12939), .A2(n12938), .A3(n12937), .A4(n12936), .ZN(
        n12940) );
  NOR2_X1 U16299 ( .A1(n12941), .A2(n12940), .ZN(n12968) );
  XOR2_X1 U16300 ( .A(n12967), .B(n12968), .Z(n12946) );
  INV_X1 U16301 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14909) );
  INV_X1 U16302 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12942) );
  OAI22_X1 U16303 ( .A1(n12943), .A2(n14909), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12942), .ZN(n12944) );
  AOI21_X1 U16304 ( .B1(n12946), .B2(n12945), .A(n12944), .ZN(n12947) );
  XNOR2_X1 U16305 ( .A(n12974), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15005) );
  MUX2_X1 U16306 ( .A(n12947), .B(n15005), .S(n9710), .Z(n14724) );
  AOI22_X1 U16307 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U16308 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12949), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16309 ( .A1(n12952), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U16310 ( .A1(n12613), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12873), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12953) );
  NAND4_X1 U16311 ( .A1(n12956), .A2(n12955), .A3(n12954), .A4(n12953), .ZN(
        n12966) );
  AOI22_X1 U16312 ( .A1(n12742), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16313 ( .A1(n12934), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12804), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16314 ( .A1(n12958), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U16315 ( .A1(n12960), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12959), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12961) );
  NAND4_X1 U16316 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n12965) );
  NOR2_X1 U16317 ( .A1(n12966), .A2(n12965), .ZN(n12970) );
  NOR2_X1 U16318 ( .A1(n12968), .A2(n12967), .ZN(n12969) );
  XOR2_X1 U16319 ( .A(n12970), .B(n12969), .Z(n12973) );
  AOI22_X1 U16320 ( .A1(n12979), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20913), .ZN(n12971) );
  OAI21_X1 U16321 ( .B1(n12973), .B2(n12972), .A(n12971), .ZN(n12977) );
  INV_X1 U16322 ( .A(n12974), .ZN(n12975) );
  NAND2_X1 U16323 ( .A1(n12975), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12985) );
  INV_X1 U16324 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21215) );
  XNOR2_X1 U16325 ( .A(n12985), .B(n21215), .ZN(n14999) );
  MUX2_X1 U16326 ( .A(n12977), .B(n14999), .S(n9710), .Z(n14642) );
  AOI22_X1 U16327 ( .A1(n12979), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12978), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12980) );
  INV_X1 U16328 ( .A(n12980), .ZN(n12981) );
  NAND3_X1 U16329 ( .A1(n9919), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16478) );
  INV_X1 U16330 ( .A(n16478), .ZN(n12982) );
  AND2_X2 U16331 ( .A1(n12982), .A2(n20911), .ZN(n20477) );
  NAND2_X1 U16332 ( .A1(n20915), .A2(n12983), .ZN(n21065) );
  NAND2_X1 U16333 ( .A1(n21065), .A2(n9919), .ZN(n12984) );
  NOR2_X1 U16334 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20582), .ZN(n16174) );
  AOI21_X1 U16335 ( .B1(n20683), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n16174), 
        .ZN(n13617) );
  INV_X1 U16336 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12986) );
  AOI21_X1 U16337 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12988), .ZN(n12989) );
  OAI21_X1 U16338 ( .B1(n20482), .B2(n14167), .A(n12989), .ZN(n12990) );
  AOI21_X1 U16339 ( .B1(n14710), .B2(n20477), .A(n12990), .ZN(n12991) );
  NAND2_X1 U16340 ( .A1(n12992), .A2(n12991), .ZN(P1_U2968) );
  NAND2_X1 U16341 ( .A1(n9728), .A2(n13899), .ZN(n12993) );
  NAND2_X1 U16342 ( .A1(n12995), .A2(n16568), .ZN(n13010) );
  INV_X1 U16343 ( .A(n13524), .ZN(n12996) );
  INV_X1 U16344 ( .A(n19619), .ZN(n12997) );
  NAND2_X1 U16345 ( .A1(n12998), .A2(n12997), .ZN(n13009) );
  NOR2_X1 U16346 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16199) );
  INV_X1 U16347 ( .A(n16199), .ZN(n16731) );
  NAND2_X1 U16348 ( .A1(n21192), .A2(n16731), .ZN(n13515) );
  NAND3_X2 U16349 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20259), .A3(n20125), 
        .ZN(n14135) );
  INV_X1 U16350 ( .A(n14135), .ZN(n19622) );
  NAND2_X1 U16351 ( .A1(n13044), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13041) );
  NAND2_X1 U16352 ( .A1(n13042), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13038) );
  NAND2_X1 U16353 ( .A1(n13039), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13036) );
  NAND2_X1 U16354 ( .A1(n13037), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13034) );
  NAND2_X1 U16355 ( .A1(n13031), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13032) );
  INV_X1 U16356 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13026) );
  INV_X1 U16357 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13494) );
  NAND2_X1 U16358 ( .A1(n13022), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13023) );
  INV_X1 U16359 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13055) );
  NAND2_X1 U16360 ( .A1(n13054), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13021) );
  INV_X1 U16361 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16523) );
  NAND2_X1 U16362 ( .A1(n13020), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13017) );
  INV_X1 U16363 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13018) );
  INV_X1 U16364 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16365 ( .A1(n13012), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13000) );
  NAND2_X1 U16366 ( .A1(n10591), .A2(n19936), .ZN(n16023) );
  INV_X1 U16367 ( .A(n16023), .ZN(n20262) );
  OR2_X1 U16368 ( .A1(n20259), .A2(n20262), .ZN(n20279) );
  NAND2_X1 U16369 ( .A1(n20279), .A2(n21192), .ZN(n13001) );
  INV_X1 U16370 ( .A(n13103), .ZN(n13003) );
  INV_X1 U16371 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21288) );
  NAND2_X1 U16372 ( .A1(n21288), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U16373 ( .A1(n13003), .A2(n13002), .ZN(n13528) );
  NAND2_X1 U16374 ( .A1(n13011), .A2(n19613), .ZN(n13006) );
  AOI21_X1 U16375 ( .B1(n16638), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13004), .ZN(n13005) );
  OAI211_X1 U16376 ( .C1(n16489), .C2(n14135), .A(n13006), .B(n13005), .ZN(
        n13007) );
  NAND3_X1 U16377 ( .A1(n13010), .A2(n13009), .A3(n13008), .ZN(P2_U2983) );
  NOR2_X1 U16378 ( .A1(n13013), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13014) );
  INV_X1 U16379 ( .A(n9841), .ZN(n13016) );
  INV_X1 U16380 ( .A(n13013), .ZN(n13015) );
  OAI21_X1 U16381 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n13016), .A(
        n13015), .ZN(n15604) );
  INV_X1 U16382 ( .A(n15604), .ZN(n16501) );
  NAND2_X1 U16383 ( .A1(n13017), .A2(n13018), .ZN(n13019) );
  AND2_X1 U16384 ( .A1(n9841), .A2(n13019), .ZN(n15616) );
  OAI21_X1 U16385 ( .B1(n13020), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n13017), .ZN(n15627) );
  INV_X1 U16386 ( .A(n15627), .ZN(n16514) );
  AOI21_X1 U16387 ( .B1(n13021), .B2(n16523), .A(n13020), .ZN(n16522) );
  OAI21_X1 U16388 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13022), .A(
        n13023), .ZN(n15654) );
  INV_X1 U16389 ( .A(n15654), .ZN(n16135) );
  OAI21_X1 U16390 ( .B1(n9808), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n13024), .ZN(n15696) );
  INV_X1 U16391 ( .A(n15696), .ZN(n19263) );
  AND2_X1 U16392 ( .A1(n13025), .A2(n13026), .ZN(n13027) );
  OR2_X1 U16393 ( .A1(n9808), .A2(n13027), .ZN(n15707) );
  INV_X1 U16394 ( .A(n15707), .ZN(n15364) );
  INV_X1 U16395 ( .A(n13028), .ZN(n13030) );
  AOI21_X1 U16396 ( .B1(n21240), .B2(n13030), .A(n13029), .ZN(n19299) );
  OAI21_X1 U16397 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13031), .A(
        n13032), .ZN(n16591) );
  INV_X1 U16398 ( .A(n16591), .ZN(n19321) );
  OAI21_X1 U16399 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13033), .A(
        n9754), .ZN(n19346) );
  INV_X1 U16400 ( .A(n19346), .ZN(n13046) );
  AOI21_X1 U16401 ( .B1(n15737), .B2(n13034), .A(n13035), .ZN(n19357) );
  AOI21_X1 U16402 ( .B1(n16637), .B2(n13036), .A(n13037), .ZN(n19375) );
  AOI21_X1 U16403 ( .B1(n13040), .B2(n13038), .A(n13039), .ZN(n19401) );
  AOI21_X1 U16404 ( .B1(n19625), .B2(n13041), .A(n13042), .ZN(n19612) );
  AOI21_X1 U16405 ( .B1(n19641), .B2(n13043), .A(n13044), .ZN(n19633) );
  AOI22_X1 U16406 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21192), .ZN(n16006) );
  AOI22_X1 U16407 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13043), .B2(n21192), .ZN(
        n15387) );
  NAND2_X1 U16408 ( .A1(n16006), .A2(n15387), .ZN(n15386) );
  NOR2_X1 U16409 ( .A1(n19633), .A2(n15386), .ZN(n14568) );
  OAI21_X1 U16410 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13044), .A(
        n13041), .ZN(n14569) );
  NAND2_X1 U16411 ( .A1(n14568), .A2(n14569), .ZN(n19432) );
  NOR2_X1 U16412 ( .A1(n19612), .A2(n19432), .ZN(n19409) );
  OAI21_X1 U16413 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13042), .A(
        n13038), .ZN(n19412) );
  NAND2_X1 U16414 ( .A1(n19409), .A2(n19412), .ZN(n19399) );
  NOR2_X1 U16415 ( .A1(n19401), .A2(n19399), .ZN(n19384) );
  OAI21_X1 U16416 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13039), .A(
        n13036), .ZN(n19386) );
  NAND2_X1 U16417 ( .A1(n19384), .A2(n19386), .ZN(n19373) );
  NOR2_X1 U16418 ( .A1(n19375), .A2(n19373), .ZN(n19364) );
  OAI21_X1 U16419 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n13037), .A(
        n13034), .ZN(n19366) );
  NAND2_X1 U16420 ( .A1(n19364), .A2(n19366), .ZN(n19355) );
  NOR2_X1 U16421 ( .A1(n19357), .A2(n19355), .ZN(n15376) );
  INV_X1 U16422 ( .A(n13035), .ZN(n13045) );
  AOI21_X1 U16423 ( .B1(n16622), .B2(n13045), .A(n13033), .ZN(n16606) );
  INV_X1 U16424 ( .A(n16606), .ZN(n15375) );
  NAND2_X1 U16425 ( .A1(n15376), .A2(n15375), .ZN(n15373) );
  NOR2_X1 U16426 ( .A1(n13046), .A2(n15373), .ZN(n19333) );
  AOI21_X1 U16427 ( .B1(n21272), .B2(n9754), .A(n13031), .ZN(n19335) );
  INV_X1 U16428 ( .A(n19335), .ZN(n13047) );
  NAND2_X1 U16429 ( .A1(n19333), .A2(n13047), .ZN(n19319) );
  NOR2_X1 U16430 ( .A1(n19321), .A2(n19319), .ZN(n19310) );
  AOI21_X1 U16431 ( .B1(n19318), .B2(n13032), .A(n13028), .ZN(n19312) );
  INV_X1 U16432 ( .A(n19312), .ZN(n13048) );
  NAND2_X1 U16433 ( .A1(n19310), .A2(n13048), .ZN(n19297) );
  NOR2_X1 U16434 ( .A1(n19299), .A2(n19297), .ZN(n19292) );
  INV_X1 U16435 ( .A(n13049), .ZN(n13050) );
  OAI21_X1 U16436 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13029), .A(
        n13050), .ZN(n19291) );
  AND2_X1 U16437 ( .A1(n19292), .A2(n19291), .ZN(n13051) );
  OAI21_X1 U16438 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13049), .A(
        n13025), .ZN(n15714) );
  INV_X1 U16439 ( .A(n15714), .ZN(n19270) );
  AOI21_X1 U16440 ( .B1(n13024), .B2(n13494), .A(n13022), .ZN(n15682) );
  INV_X1 U16441 ( .A(n15682), .ZN(n13052) );
  INV_X1 U16442 ( .A(n13053), .ZN(n13492) );
  AOI21_X1 U16443 ( .B1(n13055), .B2(n13023), .A(n13054), .ZN(n16558) );
  OAI21_X1 U16444 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n13054), .A(
        n13021), .ZN(n15645) );
  INV_X1 U16445 ( .A(n15645), .ZN(n16535) );
  NOR2_X2 U16446 ( .A1(n16533), .A2(n19410), .ZN(n16521) );
  NOR2_X1 U16447 ( .A1(n19410), .A2(n16493), .ZN(n13057) );
  XNOR2_X1 U16448 ( .A(n13012), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16492) );
  INV_X1 U16449 ( .A(n16492), .ZN(n13056) );
  XNOR2_X1 U16450 ( .A(n13057), .B(n13056), .ZN(n13087) );
  NOR3_X1 U16451 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16200) );
  NAND2_X1 U16452 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16200), .ZN(n19450) );
  INV_X1 U16453 ( .A(n9837), .ZN(n13864) );
  NOR2_X1 U16454 ( .A1(n13510), .A2(n13059), .ZN(n13080) );
  NAND2_X1 U16455 ( .A1(n21288), .A2(n20183), .ZN(n13078) );
  INV_X1 U16456 ( .A(n13078), .ZN(n13060) );
  NAND2_X1 U16457 ( .A1(n21288), .A2(n13061), .ZN(n13072) );
  OR2_X1 U16458 ( .A1(n13062), .A2(n13072), .ZN(n13883) );
  INV_X1 U16459 ( .A(n15328), .ZN(n13065) );
  INV_X1 U16460 ( .A(n13063), .ZN(n13064) );
  NAND2_X1 U16461 ( .A1(n13065), .A2(n13064), .ZN(n13066) );
  OAI22_X1 U16462 ( .A1(n15773), .A2(n19414), .B1(n19442), .B2(n15777), .ZN(
        n13068) );
  INV_X1 U16463 ( .A(n13068), .ZN(n13086) );
  INV_X1 U16464 ( .A(n13503), .ZN(n13070) );
  NOR2_X1 U16465 ( .A1(n13070), .A2(n13069), .ZN(n13697) );
  NAND2_X1 U16466 ( .A1(n13697), .A2(n9736), .ZN(n19534) );
  INV_X1 U16467 ( .A(n13072), .ZN(n13073) );
  OR2_X1 U16468 ( .A1(n19534), .A2(n13073), .ZN(n16486) );
  INV_X1 U16469 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13074) );
  NAND3_X1 U16470 ( .A1(n13697), .A2(n13078), .A3(n13074), .ZN(n13075) );
  INV_X1 U16471 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19936) );
  NOR3_X1 U16472 ( .A1(n21192), .A2(n19936), .A3(n16731), .ZN(n16727) );
  NAND2_X1 U16473 ( .A1(n19272), .A2(n19450), .ZN(n13076) );
  NOR2_X1 U16474 ( .A1(n16727), .A2(n13076), .ZN(n13077) );
  INV_X1 U16475 ( .A(n19431), .ZN(n19440) );
  INV_X1 U16476 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13083) );
  AND2_X1 U16477 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13078), .ZN(n13079) );
  INV_X1 U16478 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13081) );
  OAI222_X1 U16479 ( .A1(n19440), .A2(n13083), .B1(n19447), .B2(n13082), .C1(
        n13081), .C2(n19420), .ZN(n13084) );
  AOI21_X1 U16480 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19444), .A(n13084), .ZN(
        n13085) );
  OAI21_X1 U16481 ( .B1(n13087), .B2(n19450), .A(n10246), .ZN(P2_U2825) );
  NAND2_X1 U16482 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U16483 ( .B1(n19870), .B2(n20278), .A(n21171), .ZN(n13090) );
  INV_X1 U16484 ( .A(n19870), .ZN(n14181) );
  NAND2_X1 U16485 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20120) );
  INV_X1 U16486 ( .A(n20120), .ZN(n13089) );
  NAND2_X1 U16487 ( .A1(n14181), .A2(n13089), .ZN(n20122) );
  AND3_X1 U16488 ( .A1(n13090), .A2(n20122), .A3(n20259), .ZN(n20008) );
  AOI21_X1 U16489 ( .B1(n13105), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20008), .ZN(n13091) );
  NOR2_X1 U16490 ( .A1(n13376), .A2(n13093), .ZN(n13094) );
  NAND2_X1 U16491 ( .A1(n13115), .A2(n13094), .ZN(n13775) );
  NAND2_X1 U16492 ( .A1(n13096), .A2(n13103), .ZN(n13098) );
  AOI22_X1 U16493 ( .A1(n13105), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20259), .B2(n20298), .ZN(n13097) );
  INV_X1 U16494 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16037) );
  NAND2_X1 U16495 ( .A1(n13099), .A2(n13103), .ZN(n13101) );
  NAND2_X1 U16496 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20288), .ZN(
        n20039) );
  NAND2_X1 U16497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20298), .ZN(
        n20077) );
  NAND2_X1 U16498 ( .A1(n20039), .A2(n20077), .ZN(n20075) );
  AND2_X1 U16499 ( .A1(n20259), .A2(n20075), .ZN(n19742) );
  AOI21_X1 U16500 ( .B1(n13105), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19742), .ZN(n13100) );
  NAND2_X1 U16501 ( .A1(n9750), .A2(n13103), .ZN(n13107) );
  XNOR2_X1 U16502 ( .A(n19870), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16051) );
  AOI22_X1 U16503 ( .A1(n13105), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20259), .B2(n16051), .ZN(n13106) );
  NAND2_X1 U16504 ( .A1(n13107), .A2(n13106), .ZN(n13110) );
  INV_X1 U16505 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13108) );
  NOR2_X1 U16506 ( .A1(n13376), .A2(n13108), .ZN(n13109) );
  OR2_X1 U16507 ( .A1(n13110), .A2(n13109), .ZN(n13111) );
  NAND2_X1 U16508 ( .A1(n13110), .A2(n13109), .ZN(n13112) );
  NAND2_X1 U16509 ( .A1(n13111), .A2(n13112), .ZN(n13621) );
  NAND2_X1 U16510 ( .A1(n13691), .A2(n13692), .ZN(n13693) );
  NAND2_X1 U16511 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13113), .ZN(
        n13114) );
  AND2_X1 U16512 ( .A1(n13115), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13116) );
  INV_X1 U16513 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16042) );
  NOR2_X1 U16514 ( .A1(n13376), .A2(n16042), .ZN(n13773) );
  NAND2_X1 U16515 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13117) );
  AND2_X1 U16516 ( .A1(n14226), .A2(n14225), .ZN(n13119) );
  INV_X1 U16517 ( .A(n14249), .ZN(n13120) );
  INV_X1 U16518 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n20017) );
  OAI22_X1 U16519 ( .A1(n13287), .A2(n20017), .B1(n13286), .B2(n13122), .ZN(
        n13127) );
  AOI22_X1 U16520 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U16521 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13123) );
  OAI211_X1 U16522 ( .C1(n13125), .C2(n13292), .A(n13124), .B(n13123), .ZN(
        n13126) );
  NOR2_X1 U16523 ( .A1(n13127), .A2(n13126), .ZN(n13141) );
  NAND2_X1 U16524 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13131) );
  AOI22_X1 U16525 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16526 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13129) );
  NAND2_X1 U16527 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13128) );
  NAND4_X1 U16528 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13139) );
  AOI22_X1 U16529 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13137) );
  OR2_X1 U16530 ( .A1(n10729), .A2(n13132), .ZN(n13136) );
  OR2_X1 U16531 ( .A1(n11121), .A2(n13133), .ZN(n13135) );
  NAND2_X1 U16532 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13134) );
  NAND4_X1 U16533 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13138) );
  NOR2_X1 U16534 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  AND2_X1 U16535 ( .A1(n13141), .A2(n13140), .ZN(n15491) );
  OAI22_X1 U16536 ( .A1(n13143), .A2(n13286), .B1(n13287), .B2(n13142), .ZN(
        n13148) );
  AOI22_X1 U16537 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13145) );
  NAND2_X1 U16538 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13144) );
  OAI211_X1 U16539 ( .C1(n13292), .C2(n13146), .A(n13145), .B(n13144), .ZN(
        n13147) );
  NOR2_X1 U16540 ( .A1(n13148), .A2(n13147), .ZN(n13162) );
  NAND2_X1 U16541 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13152) );
  AOI22_X1 U16542 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U16543 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13150) );
  NAND2_X1 U16544 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13149) );
  NAND4_X1 U16545 ( .A1(n13152), .A2(n13151), .A3(n13150), .A4(n13149), .ZN(
        n13160) );
  AOI22_X1 U16546 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13158) );
  OR2_X1 U16547 ( .A1(n10729), .A2(n13153), .ZN(n13157) );
  OR2_X1 U16548 ( .A1(n11121), .A2(n13154), .ZN(n13156) );
  NAND2_X1 U16549 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13155) );
  NAND4_X1 U16550 ( .A1(n13158), .A2(n13157), .A3(n13156), .A4(n13155), .ZN(
        n13159) );
  NOR2_X1 U16551 ( .A1(n13160), .A2(n13159), .ZN(n13161) );
  AND2_X1 U16552 ( .A1(n13162), .A2(n13161), .ZN(n15487) );
  INV_X1 U16553 ( .A(n15487), .ZN(n13163) );
  AOI22_X1 U16554 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13181) );
  NAND2_X1 U16555 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13167) );
  AOI22_X1 U16556 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U16557 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13165) );
  NAND2_X1 U16558 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13164) );
  AND4_X1 U16559 ( .A1(n13167), .A2(n13166), .A3(n13165), .A4(n13164), .ZN(
        n13180) );
  AOI22_X1 U16560 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13173) );
  OR2_X1 U16561 ( .A1(n10729), .A2(n13168), .ZN(n13172) );
  INV_X1 U16562 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13169) );
  OR2_X1 U16563 ( .A1(n11121), .A2(n13169), .ZN(n13171) );
  NAND2_X1 U16564 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13170) );
  AND4_X1 U16565 ( .A1(n13173), .A2(n13172), .A3(n13171), .A4(n13170), .ZN(
        n13179) );
  AOI22_X1 U16566 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U16567 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13174) );
  OAI211_X1 U16568 ( .C1(n13292), .C2(n13176), .A(n13175), .B(n13174), .ZN(
        n13177) );
  INV_X1 U16569 ( .A(n13177), .ZN(n13178) );
  NAND4_X1 U16570 ( .A1(n13181), .A2(n13180), .A3(n13179), .A4(n13178), .ZN(
        n15473) );
  AOI22_X1 U16571 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U16572 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13185) );
  AOI22_X1 U16573 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U16574 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13183) );
  NAND2_X1 U16575 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13182) );
  AND4_X1 U16576 ( .A1(n13185), .A2(n13184), .A3(n13183), .A4(n13182), .ZN(
        n13198) );
  AOI22_X1 U16577 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13191) );
  OR2_X1 U16578 ( .A1(n10729), .A2(n13186), .ZN(n13190) );
  OR2_X1 U16579 ( .A1(n11121), .A2(n13187), .ZN(n13189) );
  NAND2_X1 U16580 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13188) );
  AND4_X1 U16581 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13197) );
  AOI22_X1 U16582 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13193) );
  NAND2_X1 U16583 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13192) );
  OAI211_X1 U16584 ( .C1(n13292), .C2(n13194), .A(n13193), .B(n13192), .ZN(
        n13195) );
  INV_X1 U16585 ( .A(n13195), .ZN(n13196) );
  NAND4_X1 U16586 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n13196), .ZN(
        n15469) );
  NOR2_X2 U16587 ( .A1(n15466), .A2(n13200), .ZN(n15460) );
  AOI22_X1 U16588 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13202), .B1(
        n13201), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13221) );
  NAND2_X1 U16589 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13206) );
  AOI22_X1 U16590 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U16591 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13204) );
  NAND2_X1 U16592 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13203) );
  AND4_X1 U16593 ( .A1(n13206), .A2(n13205), .A3(n13204), .A4(n13203), .ZN(
        n13220) );
  AOI22_X1 U16594 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13212) );
  INV_X1 U16595 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13207) );
  OR2_X1 U16596 ( .A1(n10729), .A2(n13207), .ZN(n13211) );
  INV_X1 U16597 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13208) );
  OR2_X1 U16598 ( .A1(n11121), .A2(n13208), .ZN(n13210) );
  NAND2_X1 U16599 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13209) );
  AND4_X1 U16600 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n13219) );
  AOI22_X1 U16601 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13215) );
  NAND2_X1 U16602 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13214) );
  OAI211_X1 U16603 ( .C1(n13292), .C2(n13216), .A(n13215), .B(n13214), .ZN(
        n13217) );
  INV_X1 U16604 ( .A(n13217), .ZN(n13218) );
  NAND4_X1 U16605 ( .A1(n13221), .A2(n13220), .A3(n13219), .A4(n13218), .ZN(
        n15462) );
  OAI22_X1 U16606 ( .A1(n13287), .A2(n13223), .B1(n13286), .B2(n13222), .ZN(
        n13228) );
  AOI22_X1 U16607 ( .A1(n13213), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13225) );
  NAND2_X1 U16608 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n13224) );
  OAI211_X1 U16609 ( .C1(n13226), .C2(n13292), .A(n13225), .B(n13224), .ZN(
        n13227) );
  NOR2_X1 U16610 ( .A1(n13228), .A2(n13227), .ZN(n13242) );
  NAND2_X1 U16611 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13232) );
  AOI22_X1 U16612 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13231) );
  NAND2_X1 U16613 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13230) );
  NAND2_X1 U16614 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13229) );
  NAND4_X1 U16615 ( .A1(n13232), .A2(n13231), .A3(n13230), .A4(n13229), .ZN(
        n13240) );
  AOI22_X1 U16616 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13238) );
  OR2_X1 U16617 ( .A1(n10729), .A2(n13233), .ZN(n13237) );
  OR2_X1 U16618 ( .A1(n11121), .A2(n13234), .ZN(n13236) );
  NAND2_X1 U16619 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13235) );
  NAND4_X1 U16620 ( .A1(n13238), .A2(n13237), .A3(n13236), .A4(n13235), .ZN(
        n13239) );
  NOR2_X1 U16621 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  AND2_X1 U16622 ( .A1(n13242), .A2(n13241), .ZN(n15457) );
  INV_X1 U16623 ( .A(n15457), .ZN(n13243) );
  OAI22_X1 U16624 ( .A1(n13245), .A2(n13287), .B1(n13286), .B2(n13244), .ZN(
        n13251) );
  AOI22_X1 U16625 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U16626 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13247) );
  OAI211_X1 U16627 ( .C1(n13292), .C2(n13249), .A(n13248), .B(n13247), .ZN(
        n13250) );
  NOR2_X1 U16628 ( .A1(n13251), .A2(n13250), .ZN(n13265) );
  NAND2_X1 U16629 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13255) );
  AOI22_X1 U16630 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U16631 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n13253) );
  NAND2_X1 U16632 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13252) );
  NAND4_X1 U16633 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13263) );
  AOI22_X1 U16634 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13261) );
  OR2_X1 U16635 ( .A1(n10729), .A2(n13256), .ZN(n13260) );
  OR2_X1 U16636 ( .A1(n11121), .A2(n13257), .ZN(n13259) );
  NAND2_X1 U16637 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13258) );
  NAND4_X1 U16638 ( .A1(n13261), .A2(n13260), .A3(n13259), .A4(n13258), .ZN(
        n13262) );
  NOR2_X1 U16639 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  AOI22_X1 U16640 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10656), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13276) );
  AOI22_X1 U16641 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13275) );
  AOI22_X1 U16642 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U16643 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13272) );
  INV_X1 U16644 ( .A(n13268), .ZN(n13270) );
  AND2_X1 U16645 ( .A1(n13270), .A2(n13269), .ZN(n13448) );
  NAND2_X1 U16646 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13271) );
  AND3_X1 U16647 ( .A1(n13272), .A2(n13448), .A3(n13271), .ZN(n13273) );
  NAND4_X1 U16648 ( .A1(n13276), .A2(n13275), .A3(n13274), .A4(n13273), .ZN(
        n13284) );
  AOI22_X1 U16649 ( .A1(n9715), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16650 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16651 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13280) );
  NAND2_X1 U16652 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13278) );
  INV_X1 U16653 ( .A(n13448), .ZN(n13442) );
  NAND2_X1 U16654 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13277) );
  AND3_X1 U16655 ( .A1(n13278), .A2(n13442), .A3(n13277), .ZN(n13279) );
  NAND4_X1 U16656 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  NAND2_X1 U16657 ( .A1(n13284), .A2(n13283), .ZN(n13339) );
  NOR2_X1 U16658 ( .A1(n9736), .A2(n13339), .ZN(n13316) );
  INV_X1 U16659 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n21206) );
  OAI22_X1 U16660 ( .A1(n21206), .A2(n13287), .B1(n13286), .B2(n13285), .ZN(
        n13294) );
  AOI22_X1 U16661 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13213), .B1(
        n13288), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U16662 ( .A1(n10682), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13289) );
  OAI211_X1 U16663 ( .C1(n13292), .C2(n13291), .A(n13290), .B(n13289), .ZN(
        n13293) );
  NOR2_X1 U16664 ( .A1(n13294), .A2(n13293), .ZN(n13315) );
  NAND2_X1 U16665 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13302) );
  AOI22_X1 U16666 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13297), .B1(
        n13296), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U16667 ( .A1(n11095), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13300) );
  NAND2_X1 U16668 ( .A1(n13298), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13299) );
  NAND4_X1 U16669 ( .A1(n13302), .A2(n13301), .A3(n13300), .A4(n13299), .ZN(
        n13313) );
  AOI22_X1 U16670 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13311) );
  OR2_X1 U16671 ( .A1(n10729), .A2(n13305), .ZN(n13310) );
  INV_X1 U16672 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13306) );
  OR2_X1 U16673 ( .A1(n11121), .A2(n13306), .ZN(n13309) );
  NAND2_X1 U16674 ( .A1(n13307), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13308) );
  NAND4_X1 U16675 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13312) );
  NOR2_X1 U16676 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  XNOR2_X1 U16677 ( .A(n13316), .B(n13333), .ZN(n13337) );
  OR2_X1 U16678 ( .A1(n14195), .A2(n13339), .ZN(n15441) );
  NOR2_X1 U16679 ( .A1(n15439), .A2(n15441), .ZN(n15440) );
  BUF_X1 U16680 ( .A(n13317), .Z(n15451) );
  AOI22_X1 U16681 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16682 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16683 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13322) );
  NAND2_X1 U16684 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13320) );
  NAND2_X1 U16685 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13319) );
  AND3_X1 U16686 ( .A1(n13320), .A2(n13442), .A3(n13319), .ZN(n13321) );
  NAND4_X1 U16687 ( .A1(n13324), .A2(n13323), .A3(n13322), .A4(n13321), .ZN(
        n13332) );
  AOI22_X1 U16688 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13330) );
  AOI22_X1 U16689 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U16690 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13328) );
  NAND2_X1 U16691 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13326) );
  NAND2_X1 U16692 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13325) );
  AND3_X1 U16693 ( .A1(n13326), .A2(n13448), .A3(n13325), .ZN(n13327) );
  NAND4_X1 U16694 ( .A1(n13330), .A2(n13329), .A3(n13328), .A4(n13327), .ZN(
        n13331) );
  AND2_X1 U16695 ( .A1(n13332), .A2(n13331), .ZN(n13338) );
  INV_X1 U16696 ( .A(n13333), .ZN(n13335) );
  INV_X1 U16697 ( .A(n13339), .ZN(n13334) );
  AND2_X1 U16698 ( .A1(n13335), .A2(n13334), .ZN(n13336) );
  INV_X1 U16699 ( .A(n13376), .ZN(n13400) );
  NAND2_X1 U16700 ( .A1(n13336), .A2(n13338), .ZN(n13341) );
  OAI211_X1 U16701 ( .C1(n13338), .C2(n13336), .A(n13400), .B(n13341), .ZN(
        n15430) );
  INV_X1 U16702 ( .A(n13337), .ZN(n13340) );
  NAND2_X1 U16703 ( .A1(n9736), .A2(n13338), .ZN(n15432) );
  INV_X1 U16704 ( .A(n13341), .ZN(n13356) );
  AOI22_X1 U16705 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U16706 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U16707 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13345) );
  NAND2_X1 U16708 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13343) );
  INV_X1 U16709 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19804) );
  NAND2_X1 U16710 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13342) );
  AND3_X1 U16711 ( .A1(n13343), .A2(n13342), .A3(n13442), .ZN(n13344) );
  NAND4_X1 U16712 ( .A1(n13347), .A2(n13346), .A3(n13345), .A4(n13344), .ZN(
        n13355) );
  AOI22_X1 U16713 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U16714 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13352) );
  AOI22_X1 U16715 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U16716 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13349) );
  NAND2_X1 U16717 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13348) );
  AND3_X1 U16718 ( .A1(n13349), .A2(n13448), .A3(n13348), .ZN(n13350) );
  NAND4_X1 U16719 ( .A1(n13353), .A2(n13352), .A3(n13351), .A4(n13350), .ZN(
        n13354) );
  AND2_X1 U16720 ( .A1(n13355), .A2(n13354), .ZN(n13358) );
  NAND2_X1 U16721 ( .A1(n13356), .A2(n13358), .ZN(n13377) );
  OAI211_X1 U16722 ( .C1(n13356), .C2(n13358), .A(n13400), .B(n13377), .ZN(
        n13361) );
  INV_X1 U16723 ( .A(n13361), .ZN(n13357) );
  INV_X1 U16724 ( .A(n13358), .ZN(n13359) );
  NOR2_X1 U16725 ( .A1(n14195), .A2(n13359), .ZN(n15423) );
  NAND2_X1 U16726 ( .A1(n15424), .A2(n15423), .ZN(n15422) );
  AOI22_X1 U16727 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U16728 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U16729 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13365) );
  NAND2_X1 U16730 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13363) );
  NAND2_X1 U16731 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13362) );
  AND3_X1 U16732 ( .A1(n13363), .A2(n13442), .A3(n13362), .ZN(n13364) );
  NAND4_X1 U16733 ( .A1(n13367), .A2(n13366), .A3(n13365), .A4(n13364), .ZN(
        n13375) );
  AOI22_X1 U16734 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U16735 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U16736 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U16737 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13369) );
  NAND2_X1 U16738 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13368) );
  AND3_X1 U16739 ( .A1(n13369), .A2(n13448), .A3(n13368), .ZN(n13370) );
  NAND4_X1 U16740 ( .A1(n13373), .A2(n13372), .A3(n13371), .A4(n13370), .ZN(
        n13374) );
  NAND2_X1 U16741 ( .A1(n13375), .A2(n13374), .ZN(n13378) );
  AOI21_X1 U16742 ( .B1(n13377), .B2(n13378), .A(n13376), .ZN(n13380) );
  INV_X1 U16743 ( .A(n13377), .ZN(n13379) );
  INV_X1 U16744 ( .A(n13378), .ZN(n13381) );
  NAND2_X1 U16745 ( .A1(n13379), .A2(n13381), .ZN(n13399) );
  NAND2_X1 U16746 ( .A1(n9736), .A2(n13381), .ZN(n15418) );
  AOI22_X1 U16747 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U16748 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U16749 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U16750 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13385) );
  NAND2_X1 U16751 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13384) );
  AND3_X1 U16752 ( .A1(n13385), .A2(n13442), .A3(n13384), .ZN(n13386) );
  NAND4_X1 U16753 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13397) );
  AOI22_X1 U16754 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U16755 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U16756 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13393) );
  NAND2_X1 U16757 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13391) );
  NAND2_X1 U16758 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13390) );
  AND3_X1 U16759 ( .A1(n13391), .A2(n13448), .A3(n13390), .ZN(n13392) );
  NAND4_X1 U16760 ( .A1(n13395), .A2(n13394), .A3(n13393), .A4(n13392), .ZN(
        n13396) );
  NAND2_X1 U16761 ( .A1(n13397), .A2(n13396), .ZN(n13398) );
  INV_X1 U16762 ( .A(n13398), .ZN(n13404) );
  INV_X1 U16763 ( .A(n13399), .ZN(n13401) );
  OAI211_X1 U16764 ( .C1(n13404), .C2(n13401), .A(n15406), .B(n13400), .ZN(
        n13402) );
  INV_X1 U16765 ( .A(n13402), .ZN(n13403) );
  INV_X1 U16766 ( .A(n15412), .ZN(n13406) );
  NAND2_X1 U16767 ( .A1(n9736), .A2(n13404), .ZN(n15411) );
  AOI22_X1 U16768 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U16769 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U16770 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U16771 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13409) );
  NAND2_X1 U16772 ( .A1(n9739), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n13408) );
  AND3_X1 U16773 ( .A1(n13409), .A2(n13442), .A3(n13408), .ZN(n13410) );
  NAND4_X1 U16774 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13421) );
  AOI22_X1 U16775 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U16776 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U16777 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U16778 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13415) );
  NAND2_X1 U16779 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13414) );
  AND3_X1 U16780 ( .A1(n13415), .A2(n13448), .A3(n13414), .ZN(n13416) );
  NAND4_X1 U16781 ( .A1(n13419), .A2(n13418), .A3(n13417), .A4(n13416), .ZN(
        n13420) );
  NAND2_X1 U16782 ( .A1(n13421), .A2(n13420), .ZN(n15407) );
  AOI22_X1 U16783 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10656), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U16784 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U16785 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U16786 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13423) );
  NAND2_X1 U16787 ( .A1(n9740), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13422) );
  AND3_X1 U16788 ( .A1(n13423), .A2(n13442), .A3(n13422), .ZN(n13424) );
  NAND4_X1 U16789 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        n13435) );
  NAND2_X1 U16790 ( .A1(n10656), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13429) );
  NAND2_X1 U16791 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13428) );
  AND3_X1 U16792 ( .A1(n13429), .A2(n13448), .A3(n13428), .ZN(n13433) );
  AOI22_X1 U16793 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U16794 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U16795 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13430) );
  NAND4_X1 U16796 ( .A1(n13433), .A2(n13432), .A3(n13431), .A4(n13430), .ZN(
        n13434) );
  NAND2_X1 U16797 ( .A1(n13435), .A2(n13434), .ZN(n13439) );
  INV_X1 U16798 ( .A(n15407), .ZN(n13436) );
  NAND2_X1 U16799 ( .A1(n14195), .A2(n13436), .ZN(n13437) );
  OR2_X1 U16800 ( .A1(n15406), .A2(n13437), .ZN(n13438) );
  NOR2_X1 U16801 ( .A1(n13438), .A2(n13439), .ZN(n13440) );
  AOI21_X1 U16802 ( .B1(n13439), .B2(n13438), .A(n13440), .ZN(n15401) );
  INV_X1 U16803 ( .A(n13440), .ZN(n13441) );
  AOI22_X1 U16804 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10656), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13444) );
  AOI21_X1 U16805 ( .B1(n10644), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13442), .ZN(n13443) );
  OAI211_X1 U16806 ( .C1(n10662), .C2(n13445), .A(n13444), .B(n13443), .ZN(
        n13458) );
  AOI22_X1 U16807 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13818), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13447) );
  AOI22_X1 U16808 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U16809 ( .A1(n13447), .A2(n13446), .ZN(n13457) );
  AOI21_X1 U16810 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n10644), .A(
        n13448), .ZN(n13450) );
  AOI22_X1 U16811 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13449) );
  OAI211_X1 U16812 ( .C1(n13452), .C2(n13451), .A(n13450), .B(n13449), .ZN(
        n13456) );
  AOI22_X1 U16813 ( .A1(n13266), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9740), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U16814 ( .A1(n13818), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13453) );
  NAND2_X1 U16815 ( .A1(n13454), .A2(n13453), .ZN(n13455) );
  OAI22_X1 U16816 ( .A1(n13458), .A2(n13457), .B1(n13456), .B2(n13455), .ZN(
        n13459) );
  XNOR2_X1 U16817 ( .A(n13460), .B(n13459), .ZN(n14694) );
  NOR2_X1 U16818 ( .A1(n13868), .A2(n13861), .ZN(n13544) );
  OAI21_X1 U16819 ( .B1(n13544), .B2(n11253), .A(n13899), .ZN(n13461) );
  INV_X2 U16820 ( .A(n15499), .ZN(n15480) );
  NAND2_X1 U16821 ( .A1(n14694), .A2(n15492), .ZN(n13465) );
  NAND2_X1 U16822 ( .A1(n13461), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U16823 ( .A1(n13465), .A2(n13464), .ZN(P2_U2857) );
  NOR2_X1 U16824 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13467) );
  NOR4_X1 U16825 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13466) );
  NAND4_X1 U16826 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13467), .A4(n13466), .ZN(n13490) );
  NOR4_X1 U16827 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13471) );
  NOR4_X1 U16828 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13470) );
  NOR4_X1 U16829 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13469) );
  NOR4_X1 U16830 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13468) );
  AND4_X1 U16831 ( .A1(n13471), .A2(n13470), .A3(n13469), .A4(n13468), .ZN(
        n13477) );
  NOR4_X1 U16832 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13475) );
  NOR4_X1 U16833 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13474) );
  NOR4_X1 U16834 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13473) );
  INV_X1 U16835 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n13472) );
  AND4_X1 U16836 ( .A1(n13475), .A2(n13474), .A3(n13473), .A4(n13472), .ZN(
        n13476) );
  NAND2_X1 U16837 ( .A1(n13477), .A2(n13476), .ZN(n13478) );
  INV_X1 U16838 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21057) );
  NOR3_X1 U16839 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21057), .ZN(n13480) );
  NOR4_X1 U16840 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13479) );
  NAND4_X1 U16841 ( .A1(n14918), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13480), .A4(
        n13479), .ZN(U214) );
  NOR4_X1 U16842 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n13484) );
  NOR4_X1 U16843 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13483) );
  NOR4_X1 U16844 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13482) );
  NOR4_X1 U16845 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_12__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n13481) );
  NAND4_X1 U16846 ( .A1(n13484), .A2(n13483), .A3(n13482), .A4(n13481), .ZN(
        n13489) );
  NOR4_X1 U16847 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n13487) );
  NOR4_X1 U16848 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13486) );
  NOR4_X1 U16849 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13485) );
  INV_X1 U16850 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20207) );
  NAND4_X1 U16851 ( .A1(n13487), .A2(n13486), .A3(n13485), .A4(n20207), .ZN(
        n13488) );
  NOR2_X1 U16852 ( .A1(n14688), .A2(n13490), .ZN(n16809) );
  NAND2_X1 U16853 ( .A1(n16809), .A2(U214), .ZN(U212) );
  INV_X1 U16854 ( .A(n13491), .ZN(n13493) );
  AOI211_X1 U16855 ( .C1(n15682), .C2(n13493), .A(n13492), .B(n19450), .ZN(
        n13502) );
  INV_X1 U16856 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20232) );
  OAI22_X1 U16857 ( .A1(n20232), .A2(n19440), .B1(n13494), .B2(n19420), .ZN(
        n13501) );
  INV_X1 U16858 ( .A(n19444), .ZN(n19429) );
  OAI22_X1 U16859 ( .A1(n13495), .A2(n19447), .B1(n11494), .B2(n19429), .ZN(
        n13500) );
  OAI21_X1 U16860 ( .B1(n9806), .B2(n13496), .A(n15445), .ZN(n15678) );
  OR2_X1 U16861 ( .A1(n15892), .A2(n13497), .ZN(n13498) );
  NAND2_X1 U16862 ( .A1(n13498), .A2(n15860), .ZN(n15877) );
  OAI22_X1 U16863 ( .A1(n15678), .A2(n19414), .B1(n15877), .B2(n19442), .ZN(
        n13499) );
  OR4_X1 U16864 ( .A1(n13502), .A2(n13501), .A3(n13500), .A4(n13499), .ZN(
        P2_U2834) );
  INV_X1 U16865 ( .A(n10951), .ZN(n13504) );
  AND2_X1 U16866 ( .A1(n13504), .A2(n13503), .ZN(n19452) );
  INV_X1 U16867 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13506) );
  INV_X1 U16868 ( .A(n13697), .ZN(n13698) );
  INV_X1 U16869 ( .A(n20259), .ZN(n20261) );
  NOR2_X1 U16870 ( .A1(n20261), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13507) );
  INV_X1 U16871 ( .A(n13507), .ZN(n13505) );
  OAI211_X1 U16872 ( .C1(n19452), .C2(n13506), .A(n13698), .B(n13505), .ZN(
        P2_U2814) );
  INV_X1 U16873 ( .A(n11239), .ZN(n13517) );
  OAI21_X1 U16874 ( .B1(n13507), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13510), 
        .ZN(n13508) );
  OAI21_X1 U16875 ( .B1(n13517), .B2(n13510), .A(n13508), .ZN(P2_U3612) );
  NOR2_X1 U16876 ( .A1(n21192), .A2(n16023), .ZN(n13900) );
  AOI22_X1 U16877 ( .A1(n13510), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n13900), 
        .B2(n13514), .ZN(n13509) );
  INV_X1 U16878 ( .A(n13509), .ZN(P2_U2816) );
  INV_X1 U16879 ( .A(n13510), .ZN(n13513) );
  NAND2_X1 U16880 ( .A1(n20295), .A2(n21192), .ZN(n19540) );
  INV_X1 U16881 ( .A(n20183), .ZN(n16734) );
  AND2_X1 U16882 ( .A1(n13511), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13882) );
  OAI22_X1 U16883 ( .A1(n19540), .A2(n16734), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n13882), .ZN(n13512) );
  NOR2_X1 U16884 ( .A1(n13513), .A2(n13512), .ZN(n13521) );
  OAI22_X1 U16885 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19539), .B1(n20188), 
        .B2(n21192), .ZN(n13518) );
  NAND2_X1 U16886 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20183), .ZN(n13516) );
  AOI22_X1 U16887 ( .A1(n13518), .A2(n13517), .B1(n13516), .B2(n13515), .ZN(
        n13520) );
  NAND2_X1 U16888 ( .A1(n13521), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n13519) );
  OAI21_X1 U16889 ( .B1(n13521), .B2(n13520), .A(n13519), .ZN(P2_U3610) );
  AND2_X1 U16890 ( .A1(n11239), .A2(n20183), .ZN(n13539) );
  INV_X1 U16891 ( .A(n13539), .ZN(n13522) );
  NAND3_X1 U16892 ( .A1(n13522), .A2(n13862), .A3(n13538), .ZN(n13523) );
  NOR2_X1 U16893 ( .A1(n9837), .A2(n13523), .ZN(n13869) );
  NOR2_X1 U16894 ( .A1(n13869), .A2(n19533), .ZN(n20301) );
  OAI21_X1 U16895 ( .B1(n20301), .B2(n16202), .A(n13524), .ZN(P2_U2819) );
  NAND2_X1 U16896 ( .A1(n13525), .A2(n13532), .ZN(n13526) );
  AND2_X1 U16897 ( .A1(n13527), .A2(n13526), .ZN(n16719) );
  INV_X1 U16898 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19439) );
  NOR2_X1 U16899 ( .A1(n19272), .A2(n19439), .ZN(n16718) );
  INV_X1 U16900 ( .A(n13528), .ZN(n13530) );
  INV_X1 U16901 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13529) );
  AOI21_X1 U16902 ( .B1(n19642), .B2(n13530), .A(n13529), .ZN(n13531) );
  AOI211_X1 U16903 ( .C1(n16568), .C2(n16719), .A(n16718), .B(n13531), .ZN(
        n13535) );
  XNOR2_X1 U16904 ( .A(n13533), .B(n13532), .ZN(n16716) );
  NAND2_X1 U16905 ( .A1(n12997), .A2(n16716), .ZN(n13534) );
  OAI211_X1 U16906 ( .C1(n13625), .C2(n14135), .A(n13535), .B(n13534), .ZN(
        P2_U3014) );
  NAND2_X1 U16907 ( .A1(n12312), .A2(n14703), .ZN(n13568) );
  AND2_X1 U16908 ( .A1(n20911), .A2(n21247), .ZN(n14414) );
  INV_X1 U16909 ( .A(n12318), .ZN(n13567) );
  NOR2_X1 U16910 ( .A1(n13567), .A2(n13953), .ZN(n13536) );
  AOI211_X1 U16911 ( .C1(n13555), .C2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14414), 
        .B(n13959), .ZN(n13537) );
  INV_X1 U16912 ( .A(n13537), .ZN(P1_U2801) );
  OR3_X1 U16913 ( .A1(n19536), .A2(n13538), .A3(n10951), .ZN(n13546) );
  AND2_X1 U16914 ( .A1(n13539), .A2(n13862), .ZN(n13540) );
  INV_X1 U16915 ( .A(n13542), .ZN(n13543) );
  NOR2_X1 U16916 ( .A1(n13544), .A2(n13543), .ZN(n13545) );
  NAND2_X1 U16917 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20295), .ZN(n16201) );
  OAI22_X1 U16918 ( .A1(n13875), .A2(n19533), .B1(n16202), .B2(n16201), .ZN(
        n13547) );
  AOI21_X1 U16919 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21192), .A(n13547), 
        .ZN(n16025) );
  INV_X1 U16920 ( .A(n16025), .ZN(n13553) );
  INV_X1 U16921 ( .A(n13548), .ZN(n13549) );
  NAND2_X1 U16922 ( .A1(n9736), .A2(n13549), .ZN(n13550) );
  OR2_X1 U16923 ( .A1(n10951), .A2(n13550), .ZN(n13870) );
  OR3_X1 U16924 ( .A1(n16025), .A2(n16023), .A3(n13870), .ZN(n13551) );
  OAI21_X1 U16925 ( .B1(n13553), .B2(n13552), .A(n13551), .ZN(P2_U3595) );
  NOR2_X1 U16926 ( .A1(n14414), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13557)
         );
  OAI21_X1 U16927 ( .B1(n12337), .B2(n11980), .A(n21064), .ZN(n13556) );
  OAI21_X1 U16928 ( .B1(n13557), .B2(n21064), .A(n13556), .ZN(P1_U3487) );
  AOI21_X1 U16929 ( .B1(n13559), .B2(n15390), .A(n13558), .ZN(n13560) );
  XOR2_X1 U16930 ( .A(n13560), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n15996) );
  NOR2_X1 U16931 ( .A1(n19272), .A2(n20202), .ZN(n15999) );
  AOI21_X1 U16932 ( .B1(n16638), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15999), .ZN(n13564) );
  AOI21_X1 U16933 ( .B1(n16014), .B2(n13562), .A(n13561), .ZN(n16000) );
  NAND2_X1 U16934 ( .A1(n16000), .A2(n16632), .ZN(n13563) );
  OAI211_X1 U16935 ( .C1(n19634), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13564), .B(n13563), .ZN(n13565) );
  AOI21_X1 U16936 ( .B1(n15996), .B2(n12997), .A(n13565), .ZN(n13566) );
  OAI21_X1 U16937 ( .B1(n15396), .B2(n14135), .A(n13566), .ZN(P2_U3013) );
  INV_X1 U16938 ( .A(n13661), .ZN(n14700) );
  AOI22_X1 U16939 ( .A1(n13568), .A2(n13567), .B1(n14700), .B2(n14154), .ZN(
        n14708) );
  INV_X1 U16940 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n13569) );
  AOI21_X1 U16941 ( .B1(n14708), .B2(n14709), .A(n13569), .ZN(n13571) );
  INV_X1 U16942 ( .A(n16471), .ZN(n14625) );
  NOR3_X1 U16943 ( .A1(n14625), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n9919), 
        .ZN(n13570) );
  OR2_X1 U16944 ( .A1(n13571), .A2(n13570), .ZN(P1_U2803) );
  AND2_X1 U16945 ( .A1(n10527), .A2(n11455), .ZN(n13575) );
  INV_X1 U16946 ( .A(n19459), .ZN(n15543) );
  AND2_X1 U16947 ( .A1(n19489), .A2(n9756), .ZN(n14686) );
  INV_X1 U16948 ( .A(n14686), .ZN(n13576) );
  NAND2_X1 U16949 ( .A1(n15543), .A2(n13576), .ZN(n19491) );
  OAI22_X1 U16950 ( .A1(n14688), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14685), .ZN(n14144) );
  NAND2_X1 U16951 ( .A1(n14195), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13577) );
  AND4_X1 U16952 ( .A1(n13577), .A2(n10489), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19936), .ZN(n13578) );
  NOR2_X1 U16953 ( .A1(n13580), .A2(n13579), .ZN(n13581) );
  OR2_X1 U16954 ( .A1(n13582), .A2(n13581), .ZN(n19441) );
  INV_X1 U16955 ( .A(n19441), .ZN(n16720) );
  NOR2_X1 U16956 ( .A1(n20292), .A2(n19441), .ZN(n19526) );
  INV_X1 U16957 ( .A(n19526), .ZN(n13583) );
  OAI211_X1 U16958 ( .C1(n19453), .C2(n16720), .A(n13583), .B(n19505), .ZN(
        n13585) );
  NAND2_X1 U16959 ( .A1(n19489), .A2(n19696), .ZN(n15576) );
  AOI22_X1 U16960 ( .A1(n19523), .A2(n16720), .B1(n19522), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13584) );
  OAI211_X1 U16961 ( .C1(n19531), .C2(n14144), .A(n13585), .B(n13584), .ZN(
        P2_U2919) );
  NAND2_X1 U16962 ( .A1(n16154), .A2(n16197), .ZN(n13658) );
  NOR2_X1 U16963 ( .A1(n14156), .A2(n13656), .ZN(n13586) );
  AND2_X1 U16964 ( .A1(n12318), .A2(n13586), .ZN(n16176) );
  INV_X1 U16965 ( .A(n16176), .ZN(n13587) );
  NAND2_X1 U16966 ( .A1(n13658), .A2(n13587), .ZN(n13589) );
  AND2_X1 U16967 ( .A1(n13661), .A2(n14709), .ZN(n13588) );
  NAND2_X1 U16968 ( .A1(n20414), .A2(n14157), .ZN(n20409) );
  NOR2_X1 U16969 ( .A1(n21247), .A2(n20582), .ZN(n14048) );
  INV_X1 U16970 ( .A(n14048), .ZN(n16480) );
  NOR2_X1 U16971 ( .A1(n16480), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20432) );
  CLKBUF_X1 U16972 ( .A(n20432), .Z(n21067) );
  INV_X2 U16973 ( .A(n20412), .ZN(n20437) );
  AOI22_X1 U16974 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20437), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n21067), .ZN(n13590) );
  OAI21_X1 U16975 ( .B1(n12722), .B2(n20409), .A(n13590), .ZN(P1_U2918) );
  AOI22_X1 U16976 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U16977 ( .B1(n12822), .B2(n20409), .A(n13591), .ZN(P1_U2913) );
  AOI22_X1 U16978 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13592) );
  OAI21_X1 U16979 ( .B1(n14925), .B2(n20409), .A(n13592), .ZN(P1_U2911) );
  AOI22_X1 U16980 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13593) );
  OAI21_X1 U16981 ( .B1(n14946), .B2(n20409), .A(n13593), .ZN(P1_U2915) );
  INV_X1 U16982 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14940) );
  AOI22_X1 U16983 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13594) );
  OAI21_X1 U16984 ( .B1(n14940), .B2(n20409), .A(n13594), .ZN(P1_U2914) );
  INV_X1 U16985 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U16986 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U16987 ( .B1(n13596), .B2(n20409), .A(n13595), .ZN(P1_U2919) );
  AOI22_X1 U16988 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13597) );
  OAI21_X1 U16989 ( .B1(n14916), .B2(n20409), .A(n13597), .ZN(P1_U2909) );
  AOI22_X1 U16990 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13598) );
  OAI21_X1 U16991 ( .B1(n14968), .B2(n20409), .A(n13598), .ZN(P1_U2920) );
  AOI22_X1 U16992 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13599) );
  OAI21_X1 U16993 ( .B1(n21072), .B2(n20409), .A(n13599), .ZN(P1_U2916) );
  AOI22_X1 U16994 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13600) );
  OAI21_X1 U16995 ( .B1(n12737), .B2(n20409), .A(n13600), .ZN(P1_U2917) );
  AOI22_X1 U16996 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U16997 ( .B1(n14930), .B2(n20409), .A(n13601), .ZN(P1_U2912) );
  INV_X1 U16998 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13603) );
  AOI22_X1 U16999 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13602) );
  OAI21_X1 U17000 ( .B1(n13603), .B2(n20409), .A(n13602), .ZN(P1_U2910) );
  INV_X1 U17001 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U17002 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20432), .B1(n20437), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13604) );
  OAI21_X1 U17003 ( .B1(n13605), .B2(n20409), .A(n13604), .ZN(P1_U2908) );
  AOI22_X1 U17004 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13606) );
  OAI21_X1 U17005 ( .B1(n14909), .B2(n20409), .A(n13606), .ZN(P1_U2907) );
  INV_X1 U17006 ( .A(n20477), .ZN(n15136) );
  INV_X1 U17007 ( .A(n13607), .ZN(n13610) );
  OAI21_X1 U17008 ( .B1(n13610), .B2(n13609), .A(n13608), .ZN(n14277) );
  INV_X1 U17009 ( .A(n13611), .ZN(n13614) );
  INV_X1 U17010 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13613) );
  AOI21_X1 U17011 ( .B1(n13614), .B2(n13613), .A(n13612), .ZN(n13785) );
  INV_X1 U17012 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13615) );
  NOR2_X1 U17013 ( .A1(n12460), .A2(n13615), .ZN(n13793) );
  INV_X1 U17014 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13616) );
  AOI21_X1 U17015 ( .B1(n15131), .B2(n13617), .A(n13616), .ZN(n13618) );
  AOI211_X1 U17016 ( .C1(n13785), .C2(n12479), .A(n13793), .B(n13618), .ZN(
        n13619) );
  OAI21_X1 U17017 ( .B1(n15136), .B2(n14277), .A(n13619), .ZN(P1_U2999) );
  INV_X1 U17018 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13622) );
  MUX2_X1 U17019 ( .A(n13622), .B(n19629), .S(n15499), .Z(n13623) );
  OAI21_X1 U17020 ( .B1(n20271), .B2(n15482), .A(n13623), .ZN(P2_U2885) );
  MUX2_X1 U17021 ( .A(n13625), .B(n13624), .S(n15480), .Z(n13626) );
  OAI21_X1 U17022 ( .B1(n20292), .B2(n15482), .A(n13626), .ZN(P2_U2887) );
  MUX2_X1 U17023 ( .A(n11396), .B(n15396), .S(n15499), .Z(n13629) );
  OAI21_X1 U17024 ( .B1(n20281), .B2(n15482), .A(n13629), .ZN(P2_U2886) );
  NOR2_X1 U17025 ( .A1(n9809), .A2(n13631), .ZN(n13633) );
  NAND4_X1 U17026 ( .A1(n13634), .A2(n12320), .A3(n13633), .A4(n13632), .ZN(
        n14616) );
  NAND2_X1 U17027 ( .A1(n9749), .A2(n14616), .ZN(n13654) );
  AND2_X1 U17028 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13641) );
  INV_X1 U17029 ( .A(n13641), .ZN(n13635) );
  NAND2_X1 U17030 ( .A1(n16154), .A2(n13635), .ZN(n13643) );
  OR2_X1 U17031 ( .A1(n14155), .A2(n11980), .ZN(n13636) );
  NAND2_X1 U17032 ( .A1(n13637), .A2(n13636), .ZN(n13681) );
  NOR2_X1 U17033 ( .A1(n13638), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13639) );
  NOR2_X1 U17034 ( .A1(n13681), .A2(n13639), .ZN(n13640) );
  AOI21_X1 U17035 ( .B1(n16154), .B2(n13641), .A(n13640), .ZN(n13642) );
  MUX2_X1 U17036 ( .A(n13643), .B(n13642), .S(n11839), .Z(n13652) );
  INV_X1 U17037 ( .A(n13681), .ZN(n13650) );
  INV_X1 U17038 ( .A(n13638), .ZN(n14626) );
  AND2_X1 U17039 ( .A1(n14626), .A2(n13644), .ZN(n13649) );
  NOR2_X1 U17040 ( .A1(n13645), .A2(n14621), .ZN(n13679) );
  NAND2_X1 U17041 ( .A1(n13638), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13646) );
  NAND2_X1 U17042 ( .A1(n13646), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13647) );
  NAND2_X1 U17043 ( .A1(n13648), .A2(n13647), .ZN(n13655) );
  AOI22_X1 U17044 ( .A1(n13650), .A2(n13649), .B1(n13679), .B2(n13655), .ZN(
        n13651) );
  AND2_X1 U17045 ( .A1(n13652), .A2(n13651), .ZN(n13653) );
  NAND2_X1 U17046 ( .A1(n13654), .A2(n13653), .ZN(n14039) );
  INV_X1 U17047 ( .A(n13918), .ZN(n16183) );
  AOI22_X1 U17048 ( .A1(n14039), .A2(n16471), .B1(n13655), .B2(n16183), .ZN(
        n13676) );
  NAND2_X1 U17049 ( .A1(n14054), .A2(n13656), .ZN(n14707) );
  NAND2_X1 U17050 ( .A1(n9809), .A2(n14707), .ZN(n13657) );
  NAND2_X1 U17051 ( .A1(n13658), .A2(n13657), .ZN(n13659) );
  NAND3_X1 U17052 ( .A1(n13659), .A2(n21066), .A3(n13661), .ZN(n13671) );
  OR2_X1 U17053 ( .A1(n12320), .A2(n13660), .ZN(n13663) );
  NAND2_X1 U17054 ( .A1(n14697), .A2(n13661), .ZN(n13662) );
  NAND2_X1 U17055 ( .A1(n13663), .A2(n13662), .ZN(n13952) );
  INV_X1 U17056 ( .A(n13952), .ZN(n13670) );
  OAI21_X1 U17057 ( .B1(n14173), .B2(n13665), .A(n13664), .ZN(n13668) );
  NOR2_X1 U17058 ( .A1(n13668), .A2(n13974), .ZN(n13669) );
  NAND3_X1 U17059 ( .A1(n13671), .A2(n13670), .A3(n13669), .ZN(n16155) );
  NAND2_X1 U17060 ( .A1(n16155), .A2(n14709), .ZN(n13674) );
  NAND2_X1 U17061 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14048), .ZN(n16484) );
  INV_X1 U17062 ( .A(n16484), .ZN(n13672) );
  NAND2_X1 U17063 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13672), .ZN(n13673) );
  NAND2_X1 U17064 ( .A1(n13674), .A2(n13673), .ZN(n16470) );
  AND2_X1 U17065 ( .A1(n9919), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13675) );
  OR2_X1 U17066 ( .A1(n16470), .A2(n13675), .ZN(n16475) );
  MUX2_X1 U17067 ( .A(n11839), .B(n13676), .S(n16475), .Z(n13677) );
  INV_X1 U17068 ( .A(n13677), .ZN(P1_U3469) );
  INV_X1 U17069 ( .A(n14616), .ZN(n14622) );
  OR2_X1 U17070 ( .A1(n9748), .A2(n14622), .ZN(n13685) );
  XNOR2_X1 U17071 ( .A(n14633), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13683) );
  XNOR2_X1 U17072 ( .A(n13638), .B(n12237), .ZN(n13687) );
  NAND2_X1 U17073 ( .A1(n13679), .A2(n13687), .ZN(n13680) );
  OAI21_X1 U17074 ( .B1(n13681), .B2(n13687), .A(n13680), .ZN(n13682) );
  AOI21_X1 U17075 ( .B1(n16154), .B2(n13683), .A(n13682), .ZN(n13684) );
  NAND2_X1 U17076 ( .A1(n13685), .A2(n13684), .ZN(n14040) );
  AOI22_X1 U17077 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20498), .B2(n13686), .ZN(
        n14628) );
  NAND2_X1 U17078 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14627) );
  INV_X1 U17079 ( .A(n14627), .ZN(n13688) );
  AOI222_X1 U17080 ( .A1(n14040), .A2(n16471), .B1(n14628), .B2(n13688), .C1(
        n16183), .C2(n13687), .ZN(n13689) );
  MUX2_X1 U17081 ( .A(n12237), .B(n13689), .S(n16475), .Z(n13690) );
  INV_X1 U17082 ( .A(n13690), .ZN(P1_U3472) );
  NOR2_X1 U17083 ( .A1(n9904), .A2(n15480), .ZN(n13695) );
  AOI21_X1 U17084 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n13461), .A(n13695), .ZN(
        n13696) );
  OAI21_X1 U17085 ( .B1(n20264), .B2(n15482), .A(n13696), .ZN(P2_U2884) );
  INV_X1 U17086 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13701) );
  INV_X1 U17087 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13700) );
  OAI21_X1 U17088 ( .B1(n9736), .B2(n20183), .A(n13697), .ZN(n19608) );
  INV_X1 U17089 ( .A(n19608), .ZN(n13702) );
  NOR3_X4 U17090 ( .A1(n13698), .A2(n9736), .A3(n16734), .ZN(n19606) );
  INV_X1 U17091 ( .A(n19606), .ZN(n13699) );
  AOI22_X1 U17092 ( .A1(n14685), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13715), .ZN(n19467) );
  OAI222_X1 U17093 ( .A1(n13701), .A2(n19534), .B1(n13700), .B2(n13702), .C1(
        n13699), .C2(n19467), .ZN(P2_U2982) );
  AOI22_X1 U17094 ( .A1(n14685), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14688), .ZN(n19532) );
  INV_X1 U17095 ( .A(n19532), .ZN(n15573) );
  NAND2_X1 U17096 ( .A1(n19606), .A2(n15573), .ZN(n13719) );
  INV_X2 U17097 ( .A(n19534), .ZN(n19609) );
  AOI22_X1 U17098 ( .A1(n19609), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13703) );
  NAND2_X1 U17099 ( .A1(n13719), .A2(n13703), .ZN(P2_U2953) );
  AOI22_X1 U17100 ( .A1(n14685), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n14688), .ZN(n19474) );
  INV_X1 U17101 ( .A(n19474), .ZN(n13704) );
  NAND2_X1 U17102 ( .A1(n19606), .A2(n13704), .ZN(n13707) );
  AOI22_X1 U17103 ( .A1(n19609), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n19608), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13705) );
  NAND2_X1 U17104 ( .A1(n13707), .A2(n13705), .ZN(P2_U2979) );
  AOI22_X1 U17105 ( .A1(n19609), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U17106 ( .A1(n13707), .A2(n13706), .ZN(P2_U2964) );
  INV_X1 U17107 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13708) );
  OR2_X1 U17108 ( .A1(n14688), .A2(n13708), .ZN(n13710) );
  NAND2_X1 U17109 ( .A1(n14688), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13709) );
  AND2_X1 U17110 ( .A1(n13710), .A2(n13709), .ZN(n19472) );
  INV_X1 U17111 ( .A(n19472), .ZN(n13711) );
  NAND2_X1 U17112 ( .A1(n19606), .A2(n13711), .ZN(n13714) );
  AOI22_X1 U17113 ( .A1(n19609), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n19604), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13712) );
  NAND2_X1 U17114 ( .A1(n13714), .A2(n13712), .ZN(P2_U2980) );
  AOI22_X1 U17115 ( .A1(n19609), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13713) );
  NAND2_X1 U17116 ( .A1(n13714), .A2(n13713), .ZN(P2_U2965) );
  AOI22_X1 U17117 ( .A1(n14685), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13715), .ZN(n19485) );
  INV_X1 U17118 ( .A(n19485), .ZN(n13716) );
  NAND2_X1 U17119 ( .A1(n19606), .A2(n13716), .ZN(n13734) );
  AOI22_X1 U17120 ( .A1(n19609), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n19608), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U17121 ( .A1(n13734), .A2(n13717), .ZN(P2_U2975) );
  AOI22_X1 U17122 ( .A1(n19609), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n19604), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13718) );
  NAND2_X1 U17123 ( .A1(n13719), .A2(n13718), .ZN(P2_U2968) );
  INV_X1 U17124 ( .A(n14144), .ZN(n19458) );
  NAND2_X1 U17125 ( .A1(n19606), .A2(n19458), .ZN(n13729) );
  AOI22_X1 U17126 ( .A1(n19609), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19608), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U17127 ( .A1(n13729), .A2(n13720), .ZN(P2_U2952) );
  OAI22_X1 U17128 ( .A1(n14688), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14685), .ZN(n19488) );
  INV_X1 U17129 ( .A(n19488), .ZN(n16546) );
  NAND2_X1 U17130 ( .A1(n19606), .A2(n16546), .ZN(n13748) );
  AOI22_X1 U17131 ( .A1(n19609), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19608), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13721) );
  NAND2_X1 U17132 ( .A1(n13748), .A2(n13721), .ZN(P2_U2973) );
  AOI22_X1 U17133 ( .A1(n14685), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14688), .ZN(n19690) );
  INV_X1 U17134 ( .A(n19690), .ZN(n19492) );
  NAND2_X1 U17135 ( .A1(n19606), .A2(n19492), .ZN(n13746) );
  AOI22_X1 U17136 ( .A1(n19609), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n19604), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13722) );
  NAND2_X1 U17137 ( .A1(n13746), .A2(n13722), .ZN(P2_U2972) );
  INV_X1 U17138 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16857) );
  INV_X1 U17139 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18567) );
  AOI22_X1 U17140 ( .A1(n14685), .A2(n16857), .B1(n18567), .B2(n14688), .ZN(
        n16552) );
  NAND2_X1 U17141 ( .A1(n19606), .A2(n16552), .ZN(n13727) );
  AOI22_X1 U17142 ( .A1(n19609), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n19608), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13723) );
  NAND2_X1 U17143 ( .A1(n13727), .A2(n13723), .ZN(P2_U2971) );
  AOI22_X1 U17144 ( .A1(n14685), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14688), .ZN(n19687) );
  INV_X1 U17145 ( .A(n19687), .ZN(n15556) );
  NAND2_X1 U17146 ( .A1(n19606), .A2(n15556), .ZN(n13744) );
  AOI22_X1 U17147 ( .A1(n19609), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n19604), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13724) );
  NAND2_X1 U17148 ( .A1(n13744), .A2(n13724), .ZN(P2_U2970) );
  AOI22_X1 U17149 ( .A1(n14685), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14688), .ZN(n19683) );
  INV_X1 U17150 ( .A(n19683), .ZN(n15566) );
  NAND2_X1 U17151 ( .A1(n19606), .A2(n15566), .ZN(n13742) );
  AOI22_X1 U17152 ( .A1(n19609), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n19604), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U17153 ( .A1(n13742), .A2(n13725), .ZN(P2_U2969) );
  AOI22_X1 U17154 ( .A1(n19609), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U17155 ( .A1(n13727), .A2(n13726), .ZN(P2_U2956) );
  AOI22_X1 U17156 ( .A1(n19609), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n19604), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13728) );
  NAND2_X1 U17157 ( .A1(n13729), .A2(n13728), .ZN(P2_U2967) );
  INV_X1 U17158 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16843) );
  OR2_X1 U17159 ( .A1(n14688), .A2(n16843), .ZN(n13731) );
  NAND2_X1 U17160 ( .A1(n14688), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13730) );
  AND2_X1 U17161 ( .A1(n13731), .A2(n13730), .ZN(n19476) );
  INV_X1 U17162 ( .A(n19476), .ZN(n15516) );
  NAND2_X1 U17163 ( .A1(n19606), .A2(n15516), .ZN(n13740) );
  AOI22_X1 U17164 ( .A1(n19609), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n19608), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U17165 ( .A1(n13740), .A2(n13732), .ZN(P2_U2978) );
  AOI22_X1 U17166 ( .A1(n19609), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U17167 ( .A1(n13734), .A2(n13733), .ZN(P2_U2960) );
  AOI22_X1 U17168 ( .A1(n14685), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14688), .ZN(n19698) );
  INV_X1 U17169 ( .A(n19698), .ZN(n13735) );
  NAND2_X1 U17170 ( .A1(n19606), .A2(n13735), .ZN(n13738) );
  AOI22_X1 U17171 ( .A1(n19609), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U17172 ( .A1(n13738), .A2(n13736), .ZN(P2_U2959) );
  AOI22_X1 U17173 ( .A1(n19609), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19608), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13737) );
  NAND2_X1 U17174 ( .A1(n13738), .A2(n13737), .ZN(P2_U2974) );
  AOI22_X1 U17175 ( .A1(n19609), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13739) );
  NAND2_X1 U17176 ( .A1(n13740), .A2(n13739), .ZN(P2_U2963) );
  AOI22_X1 U17177 ( .A1(n19609), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19608), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13741) );
  NAND2_X1 U17178 ( .A1(n13742), .A2(n13741), .ZN(P2_U2954) );
  AOI22_X1 U17179 ( .A1(n19609), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19608), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13743) );
  NAND2_X1 U17180 ( .A1(n13744), .A2(n13743), .ZN(P2_U2955) );
  AOI22_X1 U17181 ( .A1(n19609), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13745) );
  NAND2_X1 U17182 ( .A1(n13746), .A2(n13745), .ZN(P2_U2957) );
  AOI22_X1 U17183 ( .A1(n19609), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13747) );
  NAND2_X1 U17184 ( .A1(n13748), .A2(n13747), .ZN(P2_U2958) );
  NAND2_X1 U17185 ( .A1(n14688), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13750) );
  INV_X1 U17186 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16847) );
  OR2_X1 U17187 ( .A1(n14688), .A2(n16847), .ZN(n13749) );
  NAND2_X1 U17188 ( .A1(n13750), .A2(n13749), .ZN(n19481) );
  NAND2_X1 U17189 ( .A1(n19606), .A2(n19481), .ZN(n13753) );
  AOI22_X1 U17190 ( .A1(n19609), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13751) );
  NAND2_X1 U17191 ( .A1(n13753), .A2(n13751), .ZN(P2_U2961) );
  INV_X1 U17192 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19582) );
  NAND2_X1 U17193 ( .A1(n19604), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13752) );
  OAI211_X1 U17194 ( .C1(n19582), .C2(n19534), .A(n13753), .B(n13752), .ZN(
        P2_U2976) );
  INV_X1 U17195 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n21071) );
  NAND2_X1 U17196 ( .A1(n14688), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13755) );
  INV_X1 U17197 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16845) );
  OR2_X1 U17198 ( .A1(n14688), .A2(n16845), .ZN(n13754) );
  NAND2_X1 U17199 ( .A1(n13755), .A2(n13754), .ZN(n19478) );
  NAND2_X1 U17200 ( .A1(n19606), .A2(n19478), .ZN(n13758) );
  NAND2_X1 U17201 ( .A1(n19604), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13756) );
  OAI211_X1 U17202 ( .C1(n21071), .C2(n19534), .A(n13758), .B(n13756), .ZN(
        P2_U2962) );
  INV_X1 U17203 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19580) );
  NAND2_X1 U17204 ( .A1(n19604), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13757) );
  OAI211_X1 U17205 ( .C1(n19580), .C2(n19534), .A(n13758), .B(n13757), .ZN(
        P2_U2977) );
  INV_X1 U17206 ( .A(n21066), .ZN(n20985) );
  NAND2_X1 U17207 ( .A1(n21059), .A2(n20985), .ZN(n13759) );
  NOR2_X2 U17208 ( .A1(n20470), .A2(n11972), .ZN(n20455) );
  MUX2_X1 U17209 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n14918), .Z(
        n14957) );
  NAND2_X1 U17210 ( .A1(n20455), .A2(n14957), .ZN(n13805) );
  AND2_X2 U17211 ( .A1(n13768), .A2(n11972), .ZN(n20465) );
  AOI22_X1 U17212 ( .A1(n20465), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13760) );
  NAND2_X1 U17213 ( .A1(n13805), .A2(n13760), .ZN(P1_U2955) );
  MUX2_X1 U17214 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n14918), .Z(
        n14961) );
  NAND2_X1 U17215 ( .A1(n20455), .A2(n14961), .ZN(n13801) );
  AOI22_X1 U17216 ( .A1(n20465), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13761) );
  NAND2_X1 U17217 ( .A1(n13801), .A2(n13761), .ZN(P1_U2954) );
  MUX2_X1 U17218 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n14918), .Z(
        n14942) );
  NAND2_X1 U17219 ( .A1(n20455), .A2(n14942), .ZN(n13809) );
  AOI22_X1 U17220 ( .A1(n20465), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U17221 ( .A1(n13809), .A2(n13762), .ZN(P1_U2958) );
  MUX2_X1 U17222 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n14918), .Z(
        n14953) );
  NAND2_X1 U17223 ( .A1(n20455), .A2(n14953), .ZN(n13807) );
  AOI22_X1 U17224 ( .A1(n20465), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13763) );
  NAND2_X1 U17225 ( .A1(n13807), .A2(n13763), .ZN(P1_U2956) );
  MUX2_X1 U17226 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n14918), .Z(
        n14936) );
  NAND2_X1 U17227 ( .A1(n20455), .A2(n14936), .ZN(n13814) );
  AOI22_X1 U17228 ( .A1(n20465), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U17229 ( .A1(n13814), .A2(n13764), .ZN(P1_U2959) );
  MUX2_X1 U17230 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n14918), .Z(
        n14948) );
  NAND2_X1 U17231 ( .A1(n20455), .A2(n14948), .ZN(n13799) );
  AOI22_X1 U17232 ( .A1(n20465), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13765) );
  NAND2_X1 U17233 ( .A1(n13799), .A2(n13765), .ZN(P1_U2957) );
  INV_X1 U17234 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13771) );
  INV_X1 U17235 ( .A(n20455), .ZN(n13770) );
  INV_X1 U17236 ( .A(n14918), .ZN(n14634) );
  INV_X1 U17237 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13766) );
  NOR2_X1 U17238 ( .A1(n14634), .A2(n13766), .ZN(n13767) );
  AOI21_X1 U17239 ( .B1(DATAI_15_), .B2(n14634), .A(n13767), .ZN(n14979) );
  INV_X1 U17240 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13769) );
  OAI222_X1 U17241 ( .A1(n13796), .A2(n13771), .B1(n13770), .B2(n14979), .C1(
        n13769), .C2(n13768), .ZN(P1_U2967) );
  INV_X1 U17242 ( .A(n13773), .ZN(n13774) );
  NAND2_X1 U17243 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  OR2_X1 U17244 ( .A1(n13777), .A2(n13776), .ZN(n13778) );
  NAND2_X1 U17245 ( .A1(n13772), .A2(n13778), .ZN(n19503) );
  NAND2_X1 U17246 ( .A1(n13780), .A2(n13779), .ZN(n13782) );
  INV_X1 U17247 ( .A(n13781), .ZN(n13888) );
  AND2_X1 U17248 ( .A1(n13782), .A2(n13888), .ZN(n19648) );
  INV_X1 U17249 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19428) );
  NOR2_X1 U17250 ( .A1(n15499), .A2(n19428), .ZN(n13783) );
  AOI21_X1 U17251 ( .B1(n19648), .B2(n15499), .A(n13783), .ZN(n13784) );
  OAI21_X1 U17252 ( .B1(n19503), .B2(n15482), .A(n13784), .ZN(P2_U2883) );
  INV_X1 U17253 ( .A(n13785), .ZN(n13795) );
  OR2_X1 U17254 ( .A1(n13786), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13788) );
  NAND2_X1 U17255 ( .A1(n13788), .A2(n13787), .ZN(n13980) );
  INV_X1 U17256 ( .A(n13980), .ZN(n14272) );
  NAND2_X1 U17257 ( .A1(n20502), .A2(n16385), .ZN(n13790) );
  INV_X1 U17258 ( .A(n13790), .ZN(n13791) );
  AOI21_X1 U17259 ( .B1(n13613), .B2(n13790), .A(n13789), .ZN(n14676) );
  AOI22_X1 U17260 ( .A1(n13791), .A2(n13613), .B1(n14676), .B2(n16396), .ZN(
        n13792) );
  AOI211_X1 U17261 ( .C1(n20486), .C2(n14272), .A(n13793), .B(n13792), .ZN(
        n13794) );
  OAI21_X1 U17262 ( .B1(n13795), .B2(n16424), .A(n13794), .ZN(P1_U3031) );
  MUX2_X1 U17263 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n14918), .Z(
        n14972) );
  NAND2_X1 U17264 ( .A1(n20455), .A2(n14972), .ZN(n13803) );
  AOI22_X1 U17265 ( .A1(n20465), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U17266 ( .A1(n13803), .A2(n13797), .ZN(P1_U2937) );
  AOI22_X1 U17267 ( .A1(n20465), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13798) );
  NAND2_X1 U17268 ( .A1(n13799), .A2(n13798), .ZN(P1_U2942) );
  AOI22_X1 U17269 ( .A1(n20465), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U17270 ( .A1(n13801), .A2(n13800), .ZN(P1_U2939) );
  AOI22_X1 U17271 ( .A1(n20465), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13802) );
  NAND2_X1 U17272 ( .A1(n13803), .A2(n13802), .ZN(P1_U2952) );
  AOI22_X1 U17273 ( .A1(n20465), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13804) );
  NAND2_X1 U17274 ( .A1(n13805), .A2(n13804), .ZN(P1_U2940) );
  AOI22_X1 U17275 ( .A1(n20465), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U17276 ( .A1(n13807), .A2(n13806), .ZN(P1_U2941) );
  AOI22_X1 U17277 ( .A1(n20465), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13808) );
  NAND2_X1 U17278 ( .A1(n13809), .A2(n13808), .ZN(P1_U2943) );
  MUX2_X1 U17279 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n14918), .Z(
        n14965) );
  NAND2_X1 U17280 ( .A1(n20455), .A2(n14965), .ZN(n13812) );
  AOI22_X1 U17281 ( .A1(n20465), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U17282 ( .A1(n13812), .A2(n13810), .ZN(P1_U2953) );
  AOI22_X1 U17283 ( .A1(n20465), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13811) );
  NAND2_X1 U17284 ( .A1(n13812), .A2(n13811), .ZN(P1_U2938) );
  AOI22_X1 U17285 ( .A1(n20465), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13813) );
  NAND2_X1 U17286 ( .A1(n13814), .A2(n13813), .ZN(P1_U2944) );
  INV_X1 U17287 ( .A(n13815), .ZN(n13846) );
  NAND2_X1 U17288 ( .A1(n13817), .A2(n9725), .ZN(n13833) );
  NAND2_X1 U17289 ( .A1(n13833), .A2(n13267), .ZN(n13823) );
  NAND2_X1 U17290 ( .A1(n13820), .A2(n13819), .ZN(n13829) );
  INV_X1 U17291 ( .A(n13821), .ZN(n13822) );
  NAND2_X1 U17292 ( .A1(n13841), .A2(n13822), .ZN(n13837) );
  AND3_X1 U17293 ( .A1(n13823), .A2(n13829), .A3(n13837), .ZN(n13825) );
  NAND2_X1 U17294 ( .A1(n13861), .A2(n13867), .ZN(n13830) );
  AOI22_X1 U17295 ( .A1(n13830), .A2(n13829), .B1(n13821), .B2(n13841), .ZN(
        n13824) );
  MUX2_X1 U17296 ( .A(n13825), .B(n13824), .S(n10429), .Z(n13827) );
  NAND2_X1 U17297 ( .A1(n13827), .A2(n13826), .ZN(n13828) );
  AOI21_X1 U17298 ( .B1(n10631), .B2(n13846), .A(n13828), .ZN(n16024) );
  INV_X1 U17299 ( .A(n13875), .ZN(n13856) );
  MUX2_X1 U17300 ( .A(n10429), .B(n16024), .S(n13856), .Z(n13879) );
  NAND2_X1 U17301 ( .A1(n9750), .A2(n13846), .ZN(n13840) );
  NOR2_X1 U17302 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U17303 ( .A1(n13267), .A2(n13829), .ZN(n13831) );
  NAND2_X1 U17304 ( .A1(n13830), .A2(n13831), .ZN(n13835) );
  INV_X1 U17305 ( .A(n13831), .ZN(n13832) );
  NAND2_X1 U17306 ( .A1(n13833), .A2(n13832), .ZN(n13834) );
  OAI211_X1 U17307 ( .C1(n13837), .C2(n13836), .A(n13835), .B(n13834), .ZN(
        n13838) );
  INV_X1 U17308 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U17309 ( .A1(n13840), .A2(n13839), .ZN(n16020) );
  OAI22_X1 U17310 ( .A1(n13856), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16020), .B2(n13875), .ZN(n13878) );
  OR2_X1 U17311 ( .A1(n13878), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13858) );
  INV_X1 U17312 ( .A(n13841), .ZN(n13850) );
  INV_X1 U17313 ( .A(n11226), .ZN(n13843) );
  NAND2_X1 U17314 ( .A1(n13843), .A2(n13842), .ZN(n13847) );
  OAI21_X1 U17315 ( .B1(n10638), .B2(n10637), .A(n13847), .ZN(n13844) );
  OAI21_X1 U17316 ( .B1(n13850), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13844), .ZN(n13845) );
  AOI21_X1 U17317 ( .B1(n16001), .B2(n13846), .A(n13845), .ZN(n16015) );
  INV_X1 U17318 ( .A(n16015), .ZN(n13853) );
  NAND2_X1 U17319 ( .A1(n13853), .A2(n20288), .ZN(n13855) );
  NAND2_X1 U17320 ( .A1(n13096), .A2(n13846), .ZN(n13852) );
  INV_X1 U17321 ( .A(n13847), .ZN(n13849) );
  MUX2_X1 U17322 ( .A(n13850), .B(n13849), .S(n13848), .Z(n13851) );
  NAND2_X1 U17323 ( .A1(n13852), .A2(n13851), .ZN(n16007) );
  OAI22_X1 U17324 ( .A1(n13853), .A2(n20288), .B1(n20298), .B2(n16007), .ZN(
        n13854) );
  NAND2_X1 U17325 ( .A1(n13855), .A2(n13854), .ZN(n13857) );
  OAI211_X1 U17326 ( .C1(n20278), .C2(n16020), .A(n13857), .B(n13856), .ZN(
        n13859) );
  AND3_X1 U17327 ( .A1(n13879), .A2(n13858), .A3(n13859), .ZN(n13860) );
  OAI22_X1 U17328 ( .A1(n13860), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n13859), .B2(n13879), .ZN(n13881) );
  INV_X1 U17329 ( .A(n13861), .ZN(n13865) );
  INV_X1 U17330 ( .A(n13862), .ZN(n13863) );
  AOI22_X1 U17331 ( .A1(n13868), .A2(n13865), .B1(n13864), .B2(n13863), .ZN(
        n13866) );
  OAI21_X1 U17332 ( .B1(n13868), .B2(n13867), .A(n13866), .ZN(n20309) );
  OAI21_X1 U17333 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n13869), .ZN(n13871) );
  OAI211_X1 U17334 ( .C1(n13873), .C2(n13872), .A(n13871), .B(n13870), .ZN(
        n13874) );
  NOR2_X1 U17335 ( .A1(n20309), .A2(n13874), .ZN(n13877) );
  NAND2_X1 U17336 ( .A1(n13875), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13876) );
  OAI211_X1 U17337 ( .C1(n13879), .C2(n13878), .A(n13877), .B(n13876), .ZN(
        n13880) );
  AOI21_X1 U17338 ( .B1(n13881), .B2(n16203), .A(n13880), .ZN(n16740) );
  NAND2_X1 U17339 ( .A1(n16740), .A2(n10591), .ZN(n13885) );
  OAI21_X1 U17340 ( .B1(n10551), .B2(n13883), .A(n13882), .ZN(n13884) );
  AOI21_X1 U17341 ( .B1(n13885), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13884), 
        .ZN(n16735) );
  OAI21_X1 U17342 ( .B1(n16735), .B2(n21192), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13886) );
  NAND2_X1 U17343 ( .A1(n13886), .A2(n16201), .ZN(P2_U3593) );
  XOR2_X1 U17344 ( .A(n13772), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13893)
         );
  INV_X1 U17345 ( .A(n13905), .ZN(n13891) );
  INV_X1 U17346 ( .A(n13887), .ZN(n13889) );
  NAND2_X1 U17347 ( .A1(n13889), .A2(n13888), .ZN(n13890) );
  NAND2_X1 U17348 ( .A1(n13891), .A2(n13890), .ZN(n19413) );
  MUX2_X1 U17349 ( .A(n19413), .B(n19406), .S(n15480), .Z(n13892) );
  OAI21_X1 U17350 ( .B1(n13893), .B2(n15482), .A(n13892), .ZN(P2_U2882) );
  XNOR2_X1 U17351 ( .A(n13894), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13898) );
  INV_X1 U17352 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13896) );
  OAI21_X1 U17353 ( .B1(n13907), .B2(n13895), .A(n13981), .ZN(n19390) );
  MUX2_X1 U17354 ( .A(n13896), .B(n19390), .S(n15499), .Z(n13897) );
  OAI21_X1 U17355 ( .B1(n13898), .B2(n15482), .A(n13897), .ZN(P2_U2880) );
  AOI21_X1 U17356 ( .B1(n20183), .B2(n13900), .A(n13899), .ZN(n13903) );
  NOR2_X1 U17357 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n21192), .ZN(n13901) );
  OAI211_X1 U17358 ( .C1(n16735), .C2(n13901), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n16734), .ZN(n13902) );
  OAI211_X1 U17359 ( .C1(n16735), .C2(n13903), .A(n13902), .B(n19450), .ZN(
        P2_U3177) );
  NOR2_X1 U17360 ( .A1(n13905), .A2(n13904), .ZN(n13906) );
  NOR2_X1 U17361 ( .A1(n13907), .A2(n13906), .ZN(n19402) );
  INV_X1 U17362 ( .A(n19402), .ZN(n13913) );
  NOR2_X1 U17363 ( .A1(n13772), .A2(n13908), .ZN(n13910) );
  INV_X1 U17364 ( .A(n13894), .ZN(n13909) );
  OAI211_X1 U17365 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13910), .A(
        n13909), .B(n15492), .ZN(n13912) );
  NAND2_X1 U17366 ( .A1(n15480), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13911) );
  OAI211_X1 U17367 ( .C1(n13913), .C2(n15480), .A(n13912), .B(n13911), .ZN(
        P2_U2881) );
  INV_X1 U17368 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16811) );
  INV_X1 U17369 ( .A(DATAI_31_), .ZN(n13914) );
  OAI22_X1 U17370 ( .A1(n16811), .A2(n14021), .B1(n13914), .B2(n14022), .ZN(
        n20971) );
  INV_X1 U17371 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19702) );
  INV_X1 U17372 ( .A(DATAI_23_), .ZN(n13916) );
  OAI22_X1 U17373 ( .A1(n19702), .A2(n14021), .B1(n13916), .B2(n14022), .ZN(
        n20969) );
  NAND2_X1 U17374 ( .A1(n20862), .A2(n20622), .ZN(n20517) );
  NOR2_X2 U17375 ( .A1(n14025), .A2(n14662), .ZN(n20968) );
  INV_X1 U17376 ( .A(n20968), .ZN(n20852) );
  NAND2_X1 U17377 ( .A1(n20522), .A2(n14936), .ZN(n20903) );
  INV_X1 U17378 ( .A(n14286), .ZN(n14033) );
  OR2_X1 U17379 ( .A1(n9748), .A2(n14033), .ZN(n20866) );
  NAND2_X1 U17380 ( .A1(n9914), .A2(n12498), .ZN(n20616) );
  OAI21_X1 U17381 ( .B1(n20866), .B2(n20616), .A(n14027), .ZN(n13922) );
  AOI22_X1 U17382 ( .A1(n13922), .A2(n20911), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13921), .ZN(n14026) );
  OAI22_X1 U17383 ( .A1(n20852), .A2(n14027), .B1(n20903), .B2(n14026), .ZN(
        n13923) );
  AOI21_X1 U17384 ( .B1(n9850), .B2(n20542), .A(n13923), .ZN(n13926) );
  INV_X1 U17385 ( .A(n20862), .ZN(n15313) );
  NAND2_X1 U17386 ( .A1(n20650), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14066) );
  OR2_X1 U17387 ( .A1(n14066), .A2(n20915), .ZN(n15310) );
  OAI21_X1 U17388 ( .B1(n15313), .B2(n15310), .A(n14338), .ZN(n13924) );
  INV_X1 U17389 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20817) );
  NAND2_X1 U17390 ( .A1(n13924), .A2(n20781), .ZN(n14029) );
  NAND2_X1 U17391 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13925) );
  OAI211_X1 U17392 ( .C1(n9855), .C2(n14381), .A(n13926), .B(n13925), .ZN(
        P1_U3160) );
  INV_X1 U17393 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16816) );
  INV_X1 U17394 ( .A(DATAI_28_), .ZN(n13927) );
  INV_X1 U17395 ( .A(n20947), .ZN(n20838) );
  INV_X1 U17396 ( .A(DATAI_20_), .ZN(n13928) );
  INV_X1 U17397 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21108) );
  OAI22_X1 U17398 ( .A1(n13928), .A2(n14022), .B1(n21108), .B2(n14021), .ZN(
        n20946) );
  NOR2_X2 U17399 ( .A1(n14025), .A2(n11967), .ZN(n20945) );
  INV_X1 U17400 ( .A(n20945), .ZN(n20837) );
  NAND2_X1 U17401 ( .A1(n20522), .A2(n14953), .ZN(n20891) );
  OAI22_X1 U17402 ( .A1(n20837), .A2(n14027), .B1(n20891), .B2(n14026), .ZN(
        n13929) );
  AOI21_X1 U17403 ( .B1(n20946), .B2(n20542), .A(n13929), .ZN(n13931) );
  NAND2_X1 U17404 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13930) );
  OAI211_X1 U17405 ( .C1(n20838), .C2(n14381), .A(n13931), .B(n13930), .ZN(
        P1_U3157) );
  INV_X1 U17406 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16818) );
  INV_X1 U17407 ( .A(DATAI_27_), .ZN(n13932) );
  INV_X1 U17408 ( .A(n20940), .ZN(n20833) );
  INV_X1 U17409 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n21087) );
  INV_X1 U17410 ( .A(DATAI_19_), .ZN(n13933) );
  OAI22_X1 U17411 ( .A1(n21087), .A2(n14021), .B1(n13933), .B2(n14022), .ZN(
        n20939) );
  NOR2_X2 U17412 ( .A1(n14025), .A2(n13934), .ZN(n20938) );
  INV_X1 U17413 ( .A(n20938), .ZN(n20832) );
  NAND2_X1 U17414 ( .A1(n20522), .A2(n14957), .ZN(n20888) );
  OAI22_X1 U17415 ( .A1(n20832), .A2(n14027), .B1(n20888), .B2(n14026), .ZN(
        n13935) );
  AOI21_X1 U17416 ( .B1(n20939), .B2(n20542), .A(n13935), .ZN(n13937) );
  NAND2_X1 U17417 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13936) );
  OAI211_X1 U17418 ( .C1(n20833), .C2(n14381), .A(n13937), .B(n13936), .ZN(
        P1_U3156) );
  INV_X1 U17419 ( .A(DATAI_24_), .ZN(n13938) );
  OAI22_X1 U17420 ( .A1(n14931), .A2(n14021), .B1(n13938), .B2(n14022), .ZN(
        n20920) );
  INV_X1 U17421 ( .A(DATAI_16_), .ZN(n13939) );
  INV_X1 U17422 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16836) );
  OAI22_X1 U17423 ( .A1(n13939), .A2(n14022), .B1(n16836), .B2(n14021), .ZN(
        n20919) );
  NOR2_X2 U17424 ( .A1(n14025), .A2(n9720), .ZN(n20918) );
  INV_X1 U17425 ( .A(n20918), .ZN(n20812) );
  NAND2_X1 U17426 ( .A1(n20522), .A2(n14972), .ZN(n20879) );
  OAI22_X1 U17427 ( .A1(n20812), .A2(n14027), .B1(n20879), .B2(n14026), .ZN(
        n13940) );
  AOI21_X1 U17428 ( .B1(n20919), .B2(n20542), .A(n13940), .ZN(n13942) );
  NAND2_X1 U17429 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13941) );
  OAI211_X1 U17430 ( .C1(n14381), .C2(n9851), .A(n13942), .B(n13941), .ZN(
        P1_U3153) );
  INV_X1 U17431 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16820) );
  INV_X1 U17432 ( .A(DATAI_26_), .ZN(n13943) );
  OAI22_X1 U17433 ( .A1(n16820), .A2(n14021), .B1(n13943), .B2(n14022), .ZN(
        n20933) );
  INV_X1 U17434 ( .A(DATAI_18_), .ZN(n13944) );
  INV_X1 U17435 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16832) );
  NOR2_X2 U17436 ( .A1(n14025), .A2(n12302), .ZN(n20931) );
  INV_X1 U17437 ( .A(n20931), .ZN(n20828) );
  NAND2_X1 U17438 ( .A1(n20522), .A2(n14961), .ZN(n20885) );
  OAI22_X1 U17439 ( .A1(n20828), .A2(n14027), .B1(n20885), .B2(n14026), .ZN(
        n13945) );
  AOI21_X1 U17440 ( .B1(n20932), .B2(n20542), .A(n13945), .ZN(n13947) );
  NAND2_X1 U17441 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13946) );
  OAI211_X1 U17442 ( .C1(n9853), .C2(n14381), .A(n13947), .B(n13946), .ZN(
        P1_U3155) );
  INV_X1 U17443 ( .A(DATAI_25_), .ZN(n21187) );
  INV_X1 U17444 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16822) );
  OAI22_X1 U17445 ( .A1(n21187), .A2(n14022), .B1(n16822), .B2(n14021), .ZN(
        n20926) );
  INV_X1 U17446 ( .A(DATAI_17_), .ZN(n13948) );
  INV_X1 U17447 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16834) );
  OAI22_X1 U17448 ( .A1(n13948), .A2(n14022), .B1(n16834), .B2(n14021), .ZN(
        n20925) );
  NOR2_X2 U17449 ( .A1(n14025), .A2(n11972), .ZN(n20924) );
  INV_X1 U17450 ( .A(n20924), .ZN(n20824) );
  NAND2_X1 U17451 ( .A1(n20522), .A2(n14965), .ZN(n20882) );
  OAI22_X1 U17452 ( .A1(n20824), .A2(n14027), .B1(n20882), .B2(n14026), .ZN(
        n13949) );
  AOI21_X1 U17453 ( .B1(n20925), .B2(n20542), .A(n13949), .ZN(n13951) );
  NAND2_X1 U17454 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13950) );
  OAI211_X1 U17455 ( .C1(n9857), .C2(n14381), .A(n13951), .B(n13950), .ZN(
        P1_U3154) );
  AND2_X1 U17456 ( .A1(n14156), .A2(n21066), .ZN(n13958) );
  NOR2_X1 U17457 ( .A1(n13954), .A2(n13953), .ZN(n13956) );
  NOR2_X1 U17458 ( .A1(n11958), .A2(n14661), .ZN(n13955) );
  NAND4_X1 U17459 ( .A1(n11970), .A2(n13956), .A3(n13955), .A4(n11957), .ZN(
        n13975) );
  NOR2_X1 U17460 ( .A1(n13975), .A2(n14154), .ZN(n13957) );
  NAND2_X1 U17461 ( .A1(n13962), .A2(n11958), .ZN(n13963) );
  INV_X1 U17462 ( .A(n14972), .ZN(n13964) );
  INV_X1 U17463 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20441) );
  OAI222_X1 U17464 ( .A1(n14277), .A2(n14990), .B1(n14988), .B2(n13964), .C1(
        n14985), .C2(n20441), .ZN(P1_U2904) );
  OAI21_X1 U17465 ( .B1(n13966), .B2(n13965), .A(n13968), .ZN(n14180) );
  INV_X1 U17466 ( .A(n14965), .ZN(n13967) );
  OAI222_X1 U17467 ( .A1(n14180), .A2(n14990), .B1(n14988), .B2(n13967), .C1(
        n14985), .C2(n12491), .ZN(P1_U2903) );
  OAI21_X1 U17468 ( .B1(n10264), .B2(n12504), .A(n13969), .ZN(n14217) );
  INV_X1 U17469 ( .A(n14961), .ZN(n13970) );
  OAI222_X1 U17470 ( .A1(n14217), .A2(n14990), .B1(n14988), .B2(n13970), .C1(
        n14985), .C2(n12484), .ZN(P1_U2902) );
  XOR2_X1 U17471 ( .A(n13971), .B(n13972), .Z(n14223) );
  INV_X1 U17472 ( .A(n14223), .ZN(n14407) );
  INV_X1 U17473 ( .A(n14957), .ZN(n13973) );
  OAI222_X1 U17474 ( .A1(n14407), .A2(n14990), .B1(n14988), .B2(n13973), .C1(
        n14985), .C2(n12511), .ZN(P1_U2901) );
  NAND2_X1 U17475 ( .A1(n13974), .A2(n14709), .ZN(n13977) );
  OR2_X1 U17476 ( .A1(n13975), .A2(n14054), .ZN(n13976) );
  NAND2_X2 U17477 ( .A1(n20408), .A2(n14662), .ZN(n14906) );
  OAI222_X1 U17478 ( .A1(n13980), .A2(n14906), .B1(n14905), .B2(n13979), .C1(
        n14277), .C2(n14899), .ZN(P1_U2872) );
  NAND2_X1 U17479 ( .A1(n13982), .A2(n13981), .ZN(n13984) );
  INV_X1 U17480 ( .A(n13983), .ZN(n13993) );
  AND2_X1 U17481 ( .A1(n13984), .A2(n13993), .ZN(n19380) );
  INV_X1 U17482 ( .A(n19380), .ZN(n13990) );
  INV_X1 U17483 ( .A(n13985), .ZN(n13987) );
  OAI211_X1 U17484 ( .C1(n10266), .C2(n13987), .A(n15492), .B(n13986), .ZN(
        n13989) );
  NAND2_X1 U17485 ( .A1(n15480), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13988) );
  OAI211_X1 U17486 ( .C1(n13990), .C2(n15480), .A(n13989), .B(n13988), .ZN(
        P2_U2879) );
  INV_X1 U17487 ( .A(n13991), .ZN(n14116) );
  XNOR2_X1 U17488 ( .A(n13986), .B(n14116), .ZN(n13998) );
  INV_X1 U17489 ( .A(n14120), .ZN(n13996) );
  INV_X1 U17490 ( .A(n13992), .ZN(n13994) );
  NAND2_X1 U17491 ( .A1(n13994), .A2(n13993), .ZN(n13995) );
  NAND2_X1 U17492 ( .A1(n13996), .A2(n13995), .ZN(n19367) );
  MUX2_X1 U17493 ( .A(n19367), .B(n11454), .S(n15480), .Z(n13997) );
  OAI21_X1 U17494 ( .B1(n13998), .B2(n15482), .A(n13997), .ZN(P2_U2878) );
  CLKBUF_X1 U17495 ( .A(n13999), .Z(n14002) );
  OAI21_X1 U17496 ( .B1(n14002), .B2(n14001), .A(n14000), .ZN(n20497) );
  INV_X1 U17497 ( .A(n14217), .ZN(n14063) );
  AOI22_X1 U17498 ( .A1(n20474), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14003) );
  OAI21_X1 U17499 ( .B1(n20482), .B2(n14209), .A(n14003), .ZN(n14004) );
  AOI21_X1 U17500 ( .B1(n14063), .B2(n20477), .A(n14004), .ZN(n14005) );
  OAI21_X1 U17501 ( .B1(n20497), .B2(n20321), .A(n14005), .ZN(P1_U2997) );
  NAND2_X1 U17502 ( .A1(n14008), .A2(n14007), .ZN(n14009) );
  AND2_X1 U17503 ( .A1(n14006), .A2(n14009), .ZN(n20476) );
  INV_X1 U17504 ( .A(n20476), .ZN(n14011) );
  INV_X1 U17505 ( .A(n14953), .ZN(n14010) );
  INV_X1 U17506 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20434) );
  OAI222_X1 U17507 ( .A1(n14011), .A2(n14990), .B1(n14988), .B2(n14010), .C1(
        n20434), .C2(n14985), .ZN(P1_U2900) );
  OR2_X1 U17508 ( .A1(n14061), .A2(n14012), .ZN(n14013) );
  NAND2_X1 U17509 ( .A1(n14110), .A2(n14013), .ZN(n14397) );
  INV_X1 U17510 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14014) );
  OAI222_X1 U17511 ( .A1(n14397), .A2(n14906), .B1(n14905), .B2(n14014), .C1(
        n14899), .C2(n14407), .ZN(P1_U2869) );
  INV_X1 U17512 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16814) );
  INV_X1 U17513 ( .A(DATAI_29_), .ZN(n14015) );
  INV_X1 U17514 ( .A(n20954), .ZN(n20843) );
  INV_X1 U17515 ( .A(DATAI_21_), .ZN(n21284) );
  INV_X1 U17516 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16828) );
  OAI22_X1 U17517 ( .A1(n21284), .A2(n14022), .B1(n16828), .B2(n14021), .ZN(
        n20953) );
  NOR2_X2 U17518 ( .A1(n14025), .A2(n14016), .ZN(n20952) );
  INV_X1 U17519 ( .A(n20952), .ZN(n20842) );
  NAND2_X1 U17520 ( .A1(n20522), .A2(n14948), .ZN(n20894) );
  OAI22_X1 U17521 ( .A1(n20842), .A2(n14027), .B1(n20894), .B2(n14026), .ZN(
        n14017) );
  AOI21_X1 U17522 ( .B1(n20953), .B2(n20542), .A(n14017), .ZN(n14019) );
  NAND2_X1 U17523 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14018) );
  OAI211_X1 U17524 ( .C1(n20843), .C2(n14381), .A(n14019), .B(n14018), .ZN(
        P1_U3158) );
  INV_X1 U17525 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16812) );
  INV_X1 U17526 ( .A(DATAI_30_), .ZN(n14020) );
  OAI22_X1 U17527 ( .A1(n16812), .A2(n14021), .B1(n14020), .B2(n14022), .ZN(
        n20961) );
  INV_X1 U17528 ( .A(DATAI_22_), .ZN(n14023) );
  INV_X1 U17529 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16825) );
  OAI22_X1 U17530 ( .A1(n14023), .A2(n14022), .B1(n16825), .B2(n14021), .ZN(
        n20960) );
  NOR2_X2 U17531 ( .A1(n14025), .A2(n14024), .ZN(n20959) );
  INV_X1 U17532 ( .A(n20959), .ZN(n20847) );
  NAND2_X1 U17533 ( .A1(n20522), .A2(n14942), .ZN(n20897) );
  OAI22_X1 U17534 ( .A1(n20847), .A2(n14027), .B1(n20897), .B2(n14026), .ZN(
        n14028) );
  AOI21_X1 U17535 ( .B1(n20960), .B2(n20542), .A(n14028), .ZN(n14031) );
  NAND2_X1 U17536 ( .A1(n14029), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14030) );
  OAI211_X1 U17537 ( .C1(n9859), .C2(n14381), .A(n14031), .B(n14030), .ZN(
        P1_U3159) );
  NOR2_X1 U17538 ( .A1(n14034), .A2(n14033), .ZN(n14035) );
  XNOR2_X1 U17539 ( .A(n14035), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20395) );
  NOR2_X1 U17540 ( .A1(n20395), .A2(n12320), .ZN(n16472) );
  NAND2_X1 U17541 ( .A1(n16155), .A2(n21247), .ZN(n14038) );
  NAND2_X1 U17542 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), 
        .ZN(n14037) );
  NAND2_X1 U17543 ( .A1(n14038), .A2(n16474), .ZN(n14036) );
  OAI211_X1 U17544 ( .C1(n16472), .C2(n14038), .A(n14037), .B(n14036), .ZN(
        n14045) );
  NOR2_X1 U17545 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21247), .ZN(n14041) );
  MUX2_X1 U17546 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14039), .S(
        n16155), .Z(n16164) );
  AOI22_X1 U17547 ( .A1(n14041), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16164), .B2(n21247), .ZN(n14043) );
  MUX2_X1 U17548 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14040), .S(
        n16155), .Z(n16151) );
  AOI22_X1 U17549 ( .A1(n14041), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21247), .B2(n16151), .ZN(n14042) );
  OAI21_X1 U17550 ( .B1(n14043), .B2(n14042), .A(n14045), .ZN(n16171) );
  INV_X1 U17551 ( .A(n16171), .ZN(n14044) );
  AOI21_X1 U17552 ( .B1(n14032), .B2(n14045), .A(n14044), .ZN(n14047) );
  NOR2_X1 U17553 ( .A1(n14047), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14046) );
  OAI21_X1 U17554 ( .B1(n14046), .B2(n16484), .A(n14342), .ZN(n20513) );
  INV_X1 U17555 ( .A(n14047), .ZN(n14049) );
  NAND2_X1 U17556 ( .A1(n14049), .A2(n14048), .ZN(n16178) );
  INV_X1 U17557 ( .A(n16178), .ZN(n14052) );
  INV_X1 U17558 ( .A(n12498), .ZN(n14050) );
  AND2_X1 U17559 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20817), .ZN(n15316) );
  OAI22_X1 U17560 ( .A1(n9729), .A2(n20915), .B1(n14050), .B2(n15316), .ZN(
        n14051) );
  OAI21_X1 U17561 ( .B1(n14052), .B2(n14051), .A(n20513), .ZN(n14053) );
  OAI21_X1 U17562 ( .B1(n20513), .B2(n20905), .A(n14053), .ZN(P1_U3478) );
  INV_X1 U17563 ( .A(n14180), .ZN(n14671) );
  XNOR2_X1 U17564 ( .A(n14166), .B(n14054), .ZN(n14675) );
  OAI22_X1 U17565 ( .A1(n14906), .A2(n14675), .B1(n14055), .B2(n14905), .ZN(
        n14056) );
  AOI21_X1 U17566 ( .B1(n14671), .B2(n20405), .A(n14056), .ZN(n14057) );
  INV_X1 U17567 ( .A(n14057), .ZN(P1_U2871) );
  NOR2_X1 U17568 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  OR2_X1 U17569 ( .A1(n14061), .A2(n14060), .ZN(n20503) );
  OAI22_X1 U17570 ( .A1(n14906), .A2(n20503), .B1(n14212), .B2(n14905), .ZN(
        n14062) );
  AOI21_X1 U17571 ( .B1(n14063), .B2(n20405), .A(n14062), .ZN(n14064) );
  INV_X1 U17572 ( .A(n14064), .ZN(P1_U2870) );
  INV_X1 U17573 ( .A(n20515), .ZN(n14065) );
  INV_X1 U17574 ( .A(n20784), .ZN(n20739) );
  NAND2_X1 U17575 ( .A1(n14066), .A2(n20911), .ZN(n20613) );
  OAI21_X1 U17576 ( .B1(n20739), .B2(n20915), .A(n20613), .ZN(n14070) );
  AND2_X1 U17577 ( .A1(n9749), .A2(n9748), .ZN(n20807) );
  INV_X1 U17578 ( .A(n20616), .ZN(n14067) );
  NOR2_X1 U17579 ( .A1(n20618), .A2(n20740), .ZN(n14103) );
  AOI21_X1 U17580 ( .B1(n20807), .B2(n14067), .A(n14103), .ZN(n14073) );
  NAND3_X1 U17581 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20653), .ZN(n20811) );
  INV_X1 U17582 ( .A(n20811), .ZN(n14068) );
  NOR2_X1 U17583 ( .A1(n20911), .A2(n14068), .ZN(n14069) );
  INV_X1 U17584 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14077) );
  INV_X1 U17585 ( .A(n20574), .ZN(n14071) );
  INV_X1 U17586 ( .A(n20622), .ZN(n14072) );
  INV_X1 U17587 ( .A(n20919), .ZN(n20751) );
  OAI22_X1 U17588 ( .A1(n14073), .A2(n20915), .B1(n20811), .B2(n20913), .ZN(
        n14102) );
  INV_X1 U17589 ( .A(n20879), .ZN(n20917) );
  AOI22_X1 U17590 ( .A1(n20918), .A2(n14103), .B1(n14102), .B2(n20917), .ZN(
        n14074) );
  OAI21_X1 U17591 ( .B1(n20860), .B2(n20751), .A(n14074), .ZN(n14075) );
  AOI21_X1 U17592 ( .B1(n9852), .B2(n20855), .A(n14075), .ZN(n14076) );
  OAI21_X1 U17593 ( .B1(n14108), .B2(n14077), .A(n14076), .ZN(P1_U3121) );
  INV_X1 U17594 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14081) );
  INV_X1 U17595 ( .A(n20925), .ZN(n20754) );
  INV_X1 U17596 ( .A(n20882), .ZN(n20923) );
  AOI22_X1 U17597 ( .A1(n20924), .A2(n14103), .B1(n14102), .B2(n20923), .ZN(
        n14078) );
  OAI21_X1 U17598 ( .B1(n20860), .B2(n20754), .A(n14078), .ZN(n14079) );
  AOI21_X1 U17599 ( .B1(n9858), .B2(n20855), .A(n14079), .ZN(n14080) );
  OAI21_X1 U17600 ( .B1(n14108), .B2(n14081), .A(n14080), .ZN(P1_U3122) );
  INV_X1 U17601 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14085) );
  INV_X1 U17602 ( .A(n20960), .ZN(n20769) );
  INV_X1 U17603 ( .A(n20897), .ZN(n20958) );
  AOI22_X1 U17604 ( .A1(n20959), .A2(n14103), .B1(n14102), .B2(n20958), .ZN(
        n14082) );
  OAI21_X1 U17605 ( .B1(n20860), .B2(n20769), .A(n14082), .ZN(n14083) );
  AOI21_X1 U17606 ( .B1(n9860), .B2(n20855), .A(n14083), .ZN(n14084) );
  OAI21_X1 U17607 ( .B1(n14108), .B2(n14085), .A(n14084), .ZN(P1_U3127) );
  INV_X1 U17608 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14089) );
  INV_X1 U17609 ( .A(n20932), .ZN(n20757) );
  INV_X1 U17610 ( .A(n20885), .ZN(n20930) );
  AOI22_X1 U17611 ( .A1(n20931), .A2(n14103), .B1(n14102), .B2(n20930), .ZN(
        n14086) );
  OAI21_X1 U17612 ( .B1(n20860), .B2(n20757), .A(n14086), .ZN(n14087) );
  AOI21_X1 U17613 ( .B1(n9854), .B2(n20855), .A(n14087), .ZN(n14088) );
  OAI21_X1 U17614 ( .B1(n14108), .B2(n14089), .A(n14088), .ZN(P1_U3123) );
  INV_X1 U17615 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14093) );
  INV_X1 U17616 ( .A(n20946), .ZN(n20763) );
  INV_X1 U17617 ( .A(n20891), .ZN(n20944) );
  AOI22_X1 U17618 ( .A1(n20945), .A2(n14103), .B1(n14102), .B2(n20944), .ZN(
        n14090) );
  OAI21_X1 U17619 ( .B1(n20860), .B2(n20763), .A(n14090), .ZN(n14091) );
  AOI21_X1 U17620 ( .B1(n20947), .B2(n20855), .A(n14091), .ZN(n14092) );
  OAI21_X1 U17621 ( .B1(n14108), .B2(n14093), .A(n14092), .ZN(P1_U3125) );
  INV_X1 U17622 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14097) );
  INV_X1 U17623 ( .A(n20953), .ZN(n20766) );
  INV_X1 U17624 ( .A(n20894), .ZN(n20951) );
  AOI22_X1 U17625 ( .A1(n20952), .A2(n14103), .B1(n14102), .B2(n20951), .ZN(
        n14094) );
  OAI21_X1 U17626 ( .B1(n20860), .B2(n20766), .A(n14094), .ZN(n14095) );
  AOI21_X1 U17627 ( .B1(n20954), .B2(n20855), .A(n14095), .ZN(n14096) );
  OAI21_X1 U17628 ( .B1(n14108), .B2(n14097), .A(n14096), .ZN(P1_U3126) );
  INV_X1 U17629 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14101) );
  INV_X1 U17630 ( .A(n20969), .ZN(n20776) );
  INV_X1 U17631 ( .A(n20903), .ZN(n20966) );
  AOI22_X1 U17632 ( .A1(n20968), .A2(n14103), .B1(n14102), .B2(n20966), .ZN(
        n14098) );
  OAI21_X1 U17633 ( .B1(n20860), .B2(n20776), .A(n14098), .ZN(n14099) );
  AOI21_X1 U17634 ( .B1(n9856), .B2(n20855), .A(n14099), .ZN(n14100) );
  OAI21_X1 U17635 ( .B1(n14108), .B2(n14101), .A(n14100), .ZN(P1_U3128) );
  INV_X1 U17636 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14107) );
  INV_X1 U17637 ( .A(n20939), .ZN(n20760) );
  INV_X1 U17638 ( .A(n20888), .ZN(n20937) );
  AOI22_X1 U17639 ( .A1(n20938), .A2(n14103), .B1(n14102), .B2(n20937), .ZN(
        n14104) );
  OAI21_X1 U17640 ( .B1(n20860), .B2(n20760), .A(n14104), .ZN(n14105) );
  AOI21_X1 U17641 ( .B1(n20940), .B2(n20855), .A(n14105), .ZN(n14106) );
  OAI21_X1 U17642 ( .B1(n14108), .B2(n14107), .A(n14106), .ZN(P1_U3124) );
  NAND2_X1 U17643 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  NAND2_X1 U17644 ( .A1(n16461), .A2(n14111), .ZN(n20393) );
  OAI22_X1 U17645 ( .A1(n20393), .A2(n14906), .B1(n20388), .B2(n14905), .ZN(
        n14112) );
  AOI21_X1 U17646 ( .B1(n20476), .B2(n20405), .A(n14112), .ZN(n14113) );
  INV_X1 U17647 ( .A(n14113), .ZN(P1_U2868) );
  INV_X1 U17648 ( .A(n14114), .ZN(n14118) );
  OAI21_X1 U17649 ( .B1(n13986), .B2(n14116), .A(n14115), .ZN(n14117) );
  NAND3_X1 U17650 ( .A1(n14118), .A2(n15492), .A3(n14117), .ZN(n14123) );
  NOR2_X1 U17651 ( .A1(n14120), .A2(n14119), .ZN(n14121) );
  NOR2_X1 U17652 ( .A1(n14126), .A2(n14121), .ZN(n19358) );
  NAND2_X1 U17653 ( .A1(n19358), .A2(n15499), .ZN(n14122) );
  OAI211_X1 U17654 ( .C1(n15499), .C2(n14124), .A(n14123), .B(n14122), .ZN(
        P2_U2877) );
  XNOR2_X1 U17655 ( .A(n14114), .B(n14226), .ZN(n14129) );
  OAI21_X1 U17656 ( .B1(n14126), .B2(n14125), .A(n14228), .ZN(n16614) );
  MUX2_X1 U17657 ( .A(n14127), .B(n16614), .S(n15499), .Z(n14128) );
  OAI21_X1 U17658 ( .B1(n14129), .B2(n15482), .A(n14128), .ZN(P2_U2876) );
  NAND2_X1 U17659 ( .A1(n20264), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20258) );
  OAI21_X1 U17660 ( .B1(n20258), .B2(n20046), .A(n20259), .ZN(n14143) );
  NOR2_X1 U17661 ( .A1(n20278), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19867) );
  NAND2_X1 U17662 ( .A1(n19867), .A2(n20288), .ZN(n14142) );
  INV_X1 U17663 ( .A(n14142), .ZN(n14130) );
  OR2_X1 U17664 ( .A1(n14143), .A2(n14130), .ZN(n14134) );
  NAND2_X1 U17665 ( .A1(n14139), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14131) );
  INV_X1 U17666 ( .A(n19867), .ZN(n19869) );
  NOR2_X1 U17667 ( .A1(n20039), .A2(n19869), .ZN(n19839) );
  AOI21_X1 U17668 ( .B1(n14131), .B2(n19936), .A(n19839), .ZN(n14132) );
  NOR2_X1 U17669 ( .A1(n14132), .A2(n19874), .ZN(n14133) );
  AOI22_X1 U17670 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19693), .ZN(n20130) );
  AOI22_X1 U17671 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19693), .ZN(n19881) );
  INV_X1 U17672 ( .A(n19857), .ZN(n19865) );
  NAND2_X1 U17673 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20125), .ZN(n19695) );
  NAND2_X1 U17674 ( .A1(n9728), .A2(n19686), .ZN(n19678) );
  INV_X1 U17675 ( .A(n19839), .ZN(n14137) );
  OAI22_X1 U17676 ( .A1(n19881), .A2(n19865), .B1(n19678), .B2(n14137), .ZN(
        n14138) );
  AOI21_X1 U17677 ( .B1(n19830), .B2(n20080), .A(n14138), .ZN(n14147) );
  INV_X1 U17678 ( .A(n14139), .ZN(n14140) );
  OAI21_X1 U17679 ( .B1(n14140), .B2(n19839), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14141) );
  OAI21_X1 U17680 ( .B1(n14143), .B2(n14142), .A(n14141), .ZN(n19831) );
  NAND2_X1 U17681 ( .A1(n19831), .A2(n14145), .ZN(n14146) );
  OAI211_X1 U17682 ( .C1(n19834), .C2(n14148), .A(n14147), .B(n14146), .ZN(
        P2_U3088) );
  AND2_X1 U17683 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20683), .ZN(n14149) );
  OAI21_X1 U17684 ( .B1(n16471), .B2(n14149), .A(n20913), .ZN(n14151) );
  INV_X1 U17685 ( .A(n16184), .ZN(n21062) );
  OAI21_X1 U17686 ( .B1(n20817), .B2(n21062), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n16182) );
  INV_X1 U17687 ( .A(n16182), .ZN(n14150) );
  AOI21_X1 U17688 ( .B1(n14151), .B2(n9919), .A(n14150), .ZN(n14152) );
  NOR2_X1 U17689 ( .A1(n14167), .A2(n21247), .ZN(n14153) );
  OAI21_X1 U17690 ( .B1(n14165), .B2(n14154), .A(n21403), .ZN(n20400) );
  INV_X1 U17691 ( .A(n20400), .ZN(n14406) );
  AND2_X1 U17692 ( .A1(n14155), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14163) );
  INV_X1 U17693 ( .A(n14163), .ZN(n14158) );
  AND2_X1 U17694 ( .A1(n21066), .A2(n20683), .ZN(n16177) );
  OAI21_X1 U17695 ( .B1(n14156), .B2(n16197), .A(n16177), .ZN(n14160) );
  NAND3_X1 U17696 ( .A1(n14158), .A2(n14157), .A3(n14160), .ZN(n14159) );
  INV_X1 U17697 ( .A(n20376), .ZN(n14547) );
  AOI22_X1 U17698 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20353), .B1(n14547), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14179) );
  NOR2_X1 U17699 ( .A1(n14160), .A2(n9720), .ZN(n14161) );
  INV_X1 U17700 ( .A(n20373), .ZN(n20375) );
  INV_X1 U17701 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20337) );
  INV_X1 U17702 ( .A(n16177), .ZN(n14162) );
  NAND2_X1 U17703 ( .A1(n14163), .A2(n14162), .ZN(n14164) );
  NOR2_X2 U17704 ( .A1(n14165), .A2(n14164), .ZN(n20377) );
  NAND2_X1 U17705 ( .A1(n20377), .A2(n14166), .ZN(n14170) );
  NAND2_X1 U17706 ( .A1(n20341), .A2(n14171), .ZN(n14169) );
  OAI211_X1 U17707 ( .C1(n20389), .C2(n14171), .A(n14170), .B(n14169), .ZN(
        n14177) );
  INV_X1 U17708 ( .A(n14173), .ZN(n14174) );
  NAND2_X1 U17709 ( .A1(n14175), .A2(n14174), .ZN(n20394) );
  NOR2_X1 U17710 ( .A1(n14172), .A2(n20394), .ZN(n14176) );
  AOI211_X1 U17711 ( .C1(n20375), .C2(n20337), .A(n14177), .B(n14176), .ZN(
        n14178) );
  OAI211_X1 U17712 ( .C1(n14406), .C2(n14180), .A(n14179), .B(n14178), .ZN(
        P1_U2839) );
  INV_X1 U17713 ( .A(n20264), .ZN(n19495) );
  NAND2_X1 U17714 ( .A1(n19495), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20121) );
  NAND2_X1 U17715 ( .A1(n20278), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16081) );
  INV_X1 U17716 ( .A(n16081), .ZN(n19900) );
  NAND2_X1 U17717 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19900), .ZN(
        n14187) );
  OAI21_X1 U17718 ( .B1(n20121), .B2(n20260), .A(n14187), .ZN(n14186) );
  NAND2_X1 U17719 ( .A1(n14181), .A2(n19900), .ZN(n14197) );
  INV_X1 U17720 ( .A(n14197), .ZN(n19996) );
  AND2_X1 U17721 ( .A1(n14197), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14182) );
  NAND2_X1 U17722 ( .A1(n14183), .A2(n14182), .ZN(n14189) );
  OAI211_X1 U17723 ( .C1(n19996), .C2(n19936), .A(n14189), .B(n20125), .ZN(
        n14184) );
  INV_X1 U17724 ( .A(n14184), .ZN(n14185) );
  NAND2_X1 U17725 ( .A1(n14186), .A2(n14185), .ZN(n19998) );
  OAI21_X1 U17726 ( .B1(n14187), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13514), 
        .ZN(n14188) );
  NAND2_X1 U17727 ( .A1(n20048), .A2(n19744), .ZN(n20038) );
  INV_X1 U17728 ( .A(n20072), .ZN(n20002) );
  AOI22_X1 U17729 ( .A1(n20030), .A2(n20127), .B1(n19992), .B2(n20080), .ZN(
        n14190) );
  OAI21_X1 U17730 ( .B1(n19678), .B2(n14197), .A(n14190), .ZN(n14191) );
  AOI21_X1 U17731 ( .B1(n19997), .B2(n14145), .A(n14191), .ZN(n14192) );
  OAI21_X1 U17732 ( .B1(n19995), .B2(n14193), .A(n14192), .ZN(P2_U3136) );
  NAND2_X1 U17733 ( .A1(n14195), .A2(n19686), .ZN(n19718) );
  INV_X1 U17734 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18551) );
  OAI22_X2 U17735 ( .A1(n16822), .A2(n19701), .B1(n18551), .B2(n19699), .ZN(
        n20132) );
  AOI22_X2 U17736 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19693), .ZN(n20135) );
  INV_X1 U17737 ( .A(n20135), .ZN(n20089) );
  AOI22_X1 U17738 ( .A1(n19992), .A2(n20132), .B1(n20030), .B2(n20089), .ZN(
        n14196) );
  OAI21_X1 U17739 ( .B1(n19718), .B2(n14197), .A(n14196), .ZN(n14198) );
  AOI21_X1 U17740 ( .B1(n19997), .B2(n14194), .A(n14198), .ZN(n14199) );
  OAI21_X1 U17741 ( .B1(n19995), .B2(n14200), .A(n14199), .ZN(P2_U3137) );
  XNOR2_X1 U17742 ( .A(n14201), .B(n14239), .ZN(n14206) );
  INV_X1 U17743 ( .A(n14202), .ZN(n14203) );
  NAND2_X1 U17744 ( .A1(n14203), .A2(n9835), .ZN(n14204) );
  AND2_X1 U17745 ( .A1(n14204), .A2(n14244), .ZN(n16676) );
  INV_X1 U17746 ( .A(n16676), .ZN(n19336) );
  INV_X1 U17747 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n21151) );
  MUX2_X1 U17748 ( .A(n19336), .B(n21151), .S(n15480), .Z(n14205) );
  OAI21_X1 U17749 ( .B1(n14206), .B2(n15482), .A(n14205), .ZN(P2_U2874) );
  NOR2_X1 U17750 ( .A1(n20337), .A2(n20373), .ZN(n14208) );
  NAND2_X1 U17751 ( .A1(n20373), .A2(n20376), .ZN(n20356) );
  NAND2_X1 U17752 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n14207) );
  OR2_X1 U17753 ( .A1(n20373), .A2(n14207), .ZN(n14396) );
  AND2_X1 U17754 ( .A1(n20356), .A2(n14396), .ZN(n14398) );
  OAI21_X1 U17755 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n14208), .A(n14398), .ZN(
        n14216) );
  INV_X1 U17756 ( .A(n9748), .ZN(n20519) );
  INV_X1 U17757 ( .A(n20394), .ZN(n14404) );
  NOR2_X1 U17758 ( .A1(n21390), .A2(n20503), .ZN(n14214) );
  INV_X1 U17759 ( .A(n14209), .ZN(n14210) );
  AOI22_X1 U17760 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n21395), .B1(
        n20341), .B2(n14210), .ZN(n14211) );
  OAI21_X1 U17761 ( .B1(n21391), .B2(n14212), .A(n14211), .ZN(n14213) );
  AOI211_X1 U17762 ( .C1(n20519), .C2(n14404), .A(n14214), .B(n14213), .ZN(
        n14215) );
  OAI211_X1 U17763 ( .C1(n14406), .C2(n14217), .A(n14216), .B(n14215), .ZN(
        P1_U2838) );
  OAI21_X1 U17764 ( .B1(n14218), .B2(n14220), .A(n14219), .ZN(n20487) );
  NAND2_X1 U17765 ( .A1(n20473), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20483) );
  NAND2_X1 U17766 ( .A1(n20474), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14221) );
  OAI211_X1 U17767 ( .C1(n20482), .C2(n14401), .A(n20483), .B(n14221), .ZN(
        n14222) );
  AOI21_X1 U17768 ( .B1(n14223), .B2(n20477), .A(n14222), .ZN(n14224) );
  OAI21_X1 U17769 ( .B1(n20487), .B2(n20321), .A(n14224), .ZN(P1_U2996) );
  INV_X1 U17770 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n21145) );
  AOI21_X1 U17771 ( .B1(n14114), .B2(n14226), .A(n14225), .ZN(n14227) );
  OR3_X1 U17772 ( .A1(n14201), .A2(n14227), .A3(n15482), .ZN(n14232) );
  NAND2_X1 U17773 ( .A1(n14229), .A2(n14228), .ZN(n14230) );
  AND2_X1 U17774 ( .A1(n14230), .A2(n9835), .ZN(n19347) );
  NAND2_X1 U17775 ( .A1(n15499), .A2(n19347), .ZN(n14231) );
  OAI211_X1 U17776 ( .C1(n15499), .C2(n21145), .A(n14232), .B(n14231), .ZN(
        P2_U2875) );
  AND2_X1 U17777 ( .A1(n14006), .A2(n14234), .ZN(n14235) );
  NOR2_X1 U17778 ( .A1(n14233), .A2(n14235), .ZN(n20406) );
  INV_X1 U17779 ( .A(n20406), .ZN(n14238) );
  INV_X1 U17780 ( .A(n14948), .ZN(n14237) );
  OAI222_X1 U17781 ( .A1(n14238), .A2(n14990), .B1(n14988), .B2(n14237), .C1(
        n14236), .C2(n14985), .ZN(P1_U2899) );
  AND2_X1 U17782 ( .A1(n14201), .A2(n14239), .ZN(n14243) );
  OAI211_X1 U17783 ( .C1(n14243), .C2(n14242), .A(n15492), .B(n14241), .ZN(
        n14247) );
  AOI21_X1 U17784 ( .B1(n14245), .B2(n14244), .A(n14251), .ZN(n19326) );
  NAND2_X1 U17785 ( .A1(n19326), .A2(n15499), .ZN(n14246) );
  OAI211_X1 U17786 ( .C1(n15499), .C2(n14248), .A(n14247), .B(n14246), .ZN(
        P2_U2873) );
  XNOR2_X1 U17787 ( .A(n14241), .B(n14249), .ZN(n14253) );
  INV_X1 U17788 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19307) );
  OAI21_X1 U17789 ( .B1(n14251), .B2(n14250), .A(n15494), .ZN(n19313) );
  MUX2_X1 U17790 ( .A(n19307), .B(n19313), .S(n15499), .Z(n14252) );
  OAI21_X1 U17791 ( .B1(n14253), .B2(n15482), .A(n14252), .ZN(P2_U2872) );
  NOR2_X1 U17792 ( .A1(n14255), .A2(n14256), .ZN(n14257) );
  OR2_X1 U17793 ( .A1(n14254), .A2(n14257), .ZN(n16359) );
  INV_X1 U17794 ( .A(n9722), .ZN(n14260) );
  INV_X1 U17795 ( .A(n14258), .ZN(n14259) );
  AOI21_X1 U17796 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n20352) );
  AOI22_X1 U17797 ( .A1(n20352), .A2(n20404), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n13978), .ZN(n14262) );
  OAI21_X1 U17798 ( .B1(n16359), .B2(n14899), .A(n14262), .ZN(P1_U2865) );
  INV_X1 U17799 ( .A(n14263), .ZN(n14265) );
  INV_X1 U17800 ( .A(n14233), .ZN(n14264) );
  AOI21_X1 U17801 ( .B1(n14265), .B2(n14264), .A(n14255), .ZN(n20369) );
  NOR2_X1 U17802 ( .A1(n9833), .A2(n14266), .ZN(n14267) );
  OR2_X1 U17803 ( .A1(n9722), .A2(n14267), .ZN(n20365) );
  OAI22_X1 U17804 ( .A1(n20365), .A2(n14906), .B1(n14269), .B2(n14905), .ZN(
        n14270) );
  AOI21_X1 U17805 ( .B1(n20369), .B2(n20405), .A(n14270), .ZN(n14271) );
  INV_X1 U17806 ( .A(n14271), .ZN(P1_U2866) );
  NAND2_X1 U17807 ( .A1(n20356), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14276) );
  NAND2_X1 U17808 ( .A1(n20377), .A2(n14272), .ZN(n14275) );
  NAND2_X1 U17809 ( .A1(n20378), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n14274) );
  OAI21_X1 U17810 ( .B1(n21395), .B2(n20341), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14273) );
  NAND4_X1 U17811 ( .A1(n14276), .A2(n14275), .A3(n14274), .A4(n14273), .ZN(
        n14279) );
  NOR2_X1 U17812 ( .A1(n14277), .A2(n14406), .ZN(n14278) );
  AOI211_X1 U17813 ( .C1(n14404), .C2(n12498), .A(n14279), .B(n14278), .ZN(
        n14280) );
  INV_X1 U17814 ( .A(n14280), .ZN(P1_U2840) );
  INV_X1 U17815 ( .A(n20369), .ZN(n14282) );
  INV_X1 U17816 ( .A(n14942), .ZN(n14281) );
  OAI222_X1 U17817 ( .A1(n14282), .A2(n14990), .B1(n14988), .B2(n14281), .C1(
        n20430), .C2(n14985), .ZN(P1_U2898) );
  INV_X1 U17818 ( .A(n14936), .ZN(n14283) );
  OAI222_X1 U17819 ( .A1(n16359), .A2(n14990), .B1(n14988), .B2(n14283), .C1(
        n14985), .C2(n12544), .ZN(P1_U2897) );
  AND2_X1 U17820 ( .A1(n20650), .A2(n14284), .ZN(n14285) );
  INV_X1 U17821 ( .A(n15315), .ZN(n14291) );
  NOR2_X1 U17822 ( .A1(n9748), .A2(n14286), .ZN(n20709) );
  INV_X1 U17823 ( .A(n20709), .ZN(n14287) );
  OAI21_X1 U17824 ( .B1(n14287), .B2(n20616), .A(n14315), .ZN(n14289) );
  AOI22_X1 U17825 ( .A1(n14289), .A2(n20911), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14293), .ZN(n14314) );
  OAI22_X1 U17826 ( .A1(n20837), .A2(n14315), .B1(n20891), .B2(n14314), .ZN(
        n14288) );
  AOI21_X1 U17827 ( .B1(n20947), .B2(n20733), .A(n14288), .ZN(n14295) );
  INV_X1 U17828 ( .A(n14289), .ZN(n14290) );
  OAI211_X1 U17829 ( .C1(n14291), .C2(n20683), .A(n20911), .B(n14290), .ZN(
        n14292) );
  NAND2_X1 U17830 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14294) );
  OAI211_X1 U17831 ( .C1(n14320), .C2(n20763), .A(n14295), .B(n14294), .ZN(
        P1_U3093) );
  OAI22_X1 U17832 ( .A1(n20842), .A2(n14315), .B1(n20894), .B2(n14314), .ZN(
        n14296) );
  AOI21_X1 U17833 ( .B1(n20954), .B2(n20733), .A(n14296), .ZN(n14298) );
  NAND2_X1 U17834 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14297) );
  OAI211_X1 U17835 ( .C1(n14320), .C2(n20766), .A(n14298), .B(n14297), .ZN(
        P1_U3094) );
  OAI22_X1 U17836 ( .A1(n20828), .A2(n14315), .B1(n20885), .B2(n14314), .ZN(
        n14299) );
  AOI21_X1 U17837 ( .B1(n9854), .B2(n20733), .A(n14299), .ZN(n14301) );
  NAND2_X1 U17838 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14300) );
  OAI211_X1 U17839 ( .C1(n14320), .C2(n20757), .A(n14301), .B(n14300), .ZN(
        P1_U3091) );
  OAI22_X1 U17840 ( .A1(n20824), .A2(n14315), .B1(n20882), .B2(n14314), .ZN(
        n14302) );
  AOI21_X1 U17841 ( .B1(n9858), .B2(n20733), .A(n14302), .ZN(n14304) );
  NAND2_X1 U17842 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14303) );
  OAI211_X1 U17843 ( .C1(n14320), .C2(n20754), .A(n14304), .B(n14303), .ZN(
        P1_U3090) );
  OAI22_X1 U17844 ( .A1(n20852), .A2(n14315), .B1(n20903), .B2(n14314), .ZN(
        n14305) );
  AOI21_X1 U17845 ( .B1(n9856), .B2(n20733), .A(n14305), .ZN(n14307) );
  NAND2_X1 U17846 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14306) );
  OAI211_X1 U17847 ( .C1(n14320), .C2(n20776), .A(n14307), .B(n14306), .ZN(
        P1_U3096) );
  OAI22_X1 U17848 ( .A1(n20847), .A2(n14315), .B1(n20897), .B2(n14314), .ZN(
        n14308) );
  AOI21_X1 U17849 ( .B1(n9860), .B2(n20733), .A(n14308), .ZN(n14310) );
  NAND2_X1 U17850 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14309) );
  OAI211_X1 U17851 ( .C1(n14320), .C2(n20769), .A(n14310), .B(n14309), .ZN(
        P1_U3095) );
  OAI22_X1 U17852 ( .A1(n20812), .A2(n14315), .B1(n20879), .B2(n14314), .ZN(
        n14311) );
  AOI21_X1 U17853 ( .B1(n9852), .B2(n20733), .A(n14311), .ZN(n14313) );
  NAND2_X1 U17854 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14312) );
  OAI211_X1 U17855 ( .C1(n14320), .C2(n20751), .A(n14313), .B(n14312), .ZN(
        P1_U3089) );
  OAI22_X1 U17856 ( .A1(n20832), .A2(n14315), .B1(n20888), .B2(n14314), .ZN(
        n14316) );
  AOI21_X1 U17857 ( .B1(n20940), .B2(n20733), .A(n14316), .ZN(n14319) );
  NAND2_X1 U17858 ( .A1(n14317), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14318) );
  OAI211_X1 U17859 ( .C1(n14320), .C2(n20760), .A(n14319), .B(n14318), .ZN(
        P1_U3092) );
  XOR2_X1 U17860 ( .A(n14321), .B(n14322), .Z(n14385) );
  NAND2_X1 U17861 ( .A1(n14325), .A2(n14324), .ZN(n14388) );
  NAND3_X1 U17862 ( .A1(n14323), .A2(n19660), .A3(n14388), .ZN(n14335) );
  OAI21_X1 U17863 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14326), .A(
        n15980), .ZN(n14334) );
  OR2_X1 U17864 ( .A1(n14328), .A2(n14327), .ZN(n14330) );
  NAND2_X1 U17865 ( .A1(n14330), .A2(n14329), .ZN(n19494) );
  INV_X1 U17866 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20205) );
  OAI22_X1 U17867 ( .A1(n19494), .A2(n19667), .B1(n20205), .B2(n19388), .ZN(
        n14331) );
  INV_X1 U17868 ( .A(n14331), .ZN(n14333) );
  NAND2_X1 U17869 ( .A1(n10631), .A2(n19669), .ZN(n14332) );
  NAND4_X1 U17870 ( .A1(n14335), .A2(n14334), .A3(n14333), .A4(n14332), .ZN(
        n14336) );
  AOI21_X1 U17871 ( .B1(n14385), .B2(n19663), .A(n14336), .ZN(n14337) );
  INV_X1 U17872 ( .A(n14337), .ZN(P2_U3043) );
  NOR2_X1 U17873 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14338), .ZN(
        n14378) );
  INV_X1 U17874 ( .A(n20866), .ZN(n20907) );
  INV_X1 U17875 ( .A(n14172), .ZN(n20865) );
  OR2_X1 U17876 ( .A1(n20650), .A2(n9729), .ZN(n20783) );
  INV_X1 U17877 ( .A(n20970), .ZN(n14339) );
  AOI21_X1 U17878 ( .B1(n14339), .B2(n14381), .A(n20683), .ZN(n14340) );
  AOI21_X1 U17879 ( .B1(n20907), .B2(n20865), .A(n14340), .ZN(n14341) );
  NOR2_X1 U17880 ( .A1(n14341), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14343) );
  NOR2_X1 U17881 ( .A1(n14345), .A2(n20913), .ZN(n20808) );
  NOR2_X1 U17882 ( .A1(n20808), .A2(n14342), .ZN(n20874) );
  OR2_X1 U17883 ( .A1(n20741), .A2(n20740), .ZN(n14346) );
  NAND2_X1 U17884 ( .A1(n14346), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20815) );
  OAI211_X1 U17885 ( .C1(n14378), .C2(n14343), .A(n20874), .B(n20815), .ZN(
        n14383) );
  OR2_X1 U17886 ( .A1(n14172), .A2(n20915), .ZN(n14344) );
  OR2_X1 U17887 ( .A1(n20866), .A2(n14344), .ZN(n14348) );
  NAND2_X1 U17888 ( .A1(n14345), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20656) );
  INV_X1 U17889 ( .A(n20656), .ZN(n20868) );
  INV_X1 U17890 ( .A(n14346), .ZN(n20809) );
  NAND2_X1 U17891 ( .A1(n20868), .A2(n20809), .ZN(n14347) );
  NAND2_X1 U17892 ( .A1(n14348), .A2(n14347), .ZN(n14377) );
  AOI22_X1 U17893 ( .A1(n20938), .A2(n14378), .B1(n14377), .B2(n20937), .ZN(
        n14350) );
  NAND2_X1 U17894 ( .A1(n20970), .A2(n20940), .ZN(n14349) );
  OAI211_X1 U17895 ( .C1(n14381), .C2(n20760), .A(n14350), .B(n14349), .ZN(
        n14351) );
  AOI21_X1 U17896 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n14351), .ZN(n14352) );
  INV_X1 U17897 ( .A(n14352), .ZN(P1_U3148) );
  AOI22_X1 U17898 ( .A1(n20931), .A2(n14378), .B1(n14377), .B2(n20930), .ZN(
        n14354) );
  NAND2_X1 U17899 ( .A1(n20970), .A2(n9854), .ZN(n14353) );
  OAI211_X1 U17900 ( .C1(n14381), .C2(n20757), .A(n14354), .B(n14353), .ZN(
        n14355) );
  AOI21_X1 U17901 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n14355), .ZN(n14356) );
  INV_X1 U17902 ( .A(n14356), .ZN(P1_U3147) );
  AOI22_X1 U17903 ( .A1(n20918), .A2(n14378), .B1(n20917), .B2(n14377), .ZN(
        n14358) );
  NAND2_X1 U17904 ( .A1(n20970), .A2(n9852), .ZN(n14357) );
  OAI211_X1 U17905 ( .C1(n20751), .C2(n14381), .A(n14358), .B(n14357), .ZN(
        n14359) );
  AOI21_X1 U17906 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n14359), .ZN(n14360) );
  INV_X1 U17907 ( .A(n14360), .ZN(P1_U3145) );
  AOI22_X1 U17908 ( .A1(n20924), .A2(n14378), .B1(n14377), .B2(n20923), .ZN(
        n14362) );
  NAND2_X1 U17909 ( .A1(n20970), .A2(n9858), .ZN(n14361) );
  OAI211_X1 U17910 ( .C1(n14381), .C2(n20754), .A(n14362), .B(n14361), .ZN(
        n14363) );
  AOI21_X1 U17911 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n14363), .ZN(n14364) );
  INV_X1 U17912 ( .A(n14364), .ZN(P1_U3146) );
  AOI22_X1 U17913 ( .A1(n20945), .A2(n14378), .B1(n14377), .B2(n20944), .ZN(
        n14366) );
  NAND2_X1 U17914 ( .A1(n20970), .A2(n20947), .ZN(n14365) );
  OAI211_X1 U17915 ( .C1(n14381), .C2(n20763), .A(n14366), .B(n14365), .ZN(
        n14367) );
  AOI21_X1 U17916 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n14367), .ZN(n14368) );
  INV_X1 U17917 ( .A(n14368), .ZN(P1_U3149) );
  AOI22_X1 U17918 ( .A1(n20968), .A2(n14378), .B1(n14377), .B2(n20966), .ZN(
        n14370) );
  NAND2_X1 U17919 ( .A1(n20970), .A2(n9856), .ZN(n14369) );
  OAI211_X1 U17920 ( .C1(n14381), .C2(n20776), .A(n14370), .B(n14369), .ZN(
        n14371) );
  AOI21_X1 U17921 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14371), .ZN(n14372) );
  INV_X1 U17922 ( .A(n14372), .ZN(P1_U3152) );
  AOI22_X1 U17923 ( .A1(n20959), .A2(n14378), .B1(n14377), .B2(n20958), .ZN(
        n14374) );
  NAND2_X1 U17924 ( .A1(n20970), .A2(n9860), .ZN(n14373) );
  OAI211_X1 U17925 ( .C1(n14381), .C2(n20769), .A(n14374), .B(n14373), .ZN(
        n14375) );
  AOI21_X1 U17926 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n14375), .ZN(n14376) );
  INV_X1 U17927 ( .A(n14376), .ZN(P1_U3151) );
  AOI22_X1 U17928 ( .A1(n20952), .A2(n14378), .B1(n14377), .B2(n20951), .ZN(
        n14380) );
  NAND2_X1 U17929 ( .A1(n20970), .A2(n20954), .ZN(n14379) );
  OAI211_X1 U17930 ( .C1(n14381), .C2(n20766), .A(n14380), .B(n14379), .ZN(
        n14382) );
  AOI21_X1 U17931 ( .B1(n14383), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14382), .ZN(n14384) );
  INV_X1 U17932 ( .A(n14384), .ZN(P1_U3150) );
  INV_X1 U17933 ( .A(n14385), .ZN(n14391) );
  NOR2_X1 U17934 ( .A1(n9904), .A2(n14135), .ZN(n14387) );
  INV_X1 U17935 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14572) );
  OAI22_X1 U17936 ( .A1(n14572), .A2(n19642), .B1(n19634), .B2(n14569), .ZN(
        n14386) );
  AOI211_X1 U17937 ( .C1(n19643), .C2(P2_REIP_REG_3__SCAN_IN), .A(n14387), .B(
        n14386), .ZN(n14390) );
  NAND3_X1 U17938 ( .A1(n14323), .A2(n14388), .A3(n16632), .ZN(n14389) );
  OAI211_X1 U17939 ( .C1(n14391), .C2(n19619), .A(n14390), .B(n14389), .ZN(
        P2_U3011) );
  OAI21_X1 U17940 ( .B1(n14254), .B2(n14393), .A(n14392), .ZN(n14408) );
  MUX2_X1 U17941 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n14918), .Z(
        n20442) );
  INV_X1 U17942 ( .A(n20442), .ZN(n14395) );
  OAI222_X1 U17943 ( .A1(n14408), .A2(n14990), .B1(n14988), .B2(n14395), .C1(
        n14394), .C2(n14985), .ZN(P1_U2896) );
  NOR2_X1 U17944 ( .A1(n14396), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n14403) );
  INV_X1 U17945 ( .A(n14397), .ZN(n20485) );
  AOI22_X1 U17946 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(n20378), .B1(n20377), .B2(
        n20485), .ZN(n14400) );
  AOI22_X1 U17947 ( .A1(n21395), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n14398), .ZN(n14399) );
  OAI211_X1 U17948 ( .C1(n14401), .C2(n21398), .A(n14400), .B(n14399), .ZN(
        n14402) );
  AOI211_X1 U17949 ( .C1(n9749), .C2(n14404), .A(n14403), .B(n14402), .ZN(
        n14405) );
  OAI21_X1 U17950 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(P1_U2837) );
  INV_X1 U17951 ( .A(n14408), .ZN(n15158) );
  NAND2_X1 U17952 ( .A1(n14258), .A2(n14409), .ZN(n14410) );
  NAND2_X1 U17953 ( .A1(n14423), .A2(n14410), .ZN(n15299) );
  OAI22_X1 U17954 ( .A1(n15299), .A2(n14906), .B1(n14411), .B2(n20408), .ZN(
        n14412) );
  AOI21_X1 U17955 ( .B1(n15158), .B2(n20405), .A(n14412), .ZN(n14413) );
  INV_X1 U17956 ( .A(n14413), .ZN(P1_U2864) );
  AOI22_X1 U17957 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n21395), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n20378), .ZN(n14415) );
  NAND2_X1 U17958 ( .A1(n14414), .A2(n20376), .ZN(n20379) );
  OAI211_X1 U17959 ( .C1(n21390), .C2(n15299), .A(n14415), .B(n20379), .ZN(
        n14418) );
  INV_X1 U17960 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21007) );
  NAND4_X1 U17961 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n20374)
         );
  INV_X1 U17962 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20383) );
  NOR3_X1 U17963 ( .A1(n20374), .A2(n20383), .A3(n20373), .ZN(n20363) );
  NAND2_X1 U17964 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20363), .ZN(n20357) );
  NOR2_X1 U17965 ( .A1(n21007), .A2(n20357), .ZN(n20340) );
  INV_X1 U17966 ( .A(n20356), .ZN(n16281) );
  AOI21_X1 U17967 ( .B1(n20340), .B2(P1_REIP_REG_8__SCAN_IN), .A(n16281), .ZN(
        n20347) );
  OAI21_X1 U17968 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20340), .A(n20347), .ZN(
        n14416) );
  OAI21_X1 U17969 ( .B1(n21398), .B2(n15156), .A(n14416), .ZN(n14417) );
  AOI211_X1 U17970 ( .C1(n15158), .C2(n20368), .A(n14418), .B(n14417), .ZN(
        n14419) );
  INV_X1 U17971 ( .A(n14419), .ZN(P1_U2832) );
  AOI21_X1 U17972 ( .B1(n14421), .B2(n14392), .A(n14420), .ZN(n20348) );
  INV_X1 U17973 ( .A(n20348), .ZN(n14426) );
  MUX2_X1 U17974 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14918), .Z(
        n20444) );
  AOI22_X1 U17975 ( .A1(n14983), .A2(n20444), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14982), .ZN(n14422) );
  OAI21_X1 U17976 ( .B1(n14426), .B2(n14990), .A(n14422), .ZN(P1_U2895) );
  INV_X1 U17977 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14425) );
  AOI21_X1 U17978 ( .B1(n14424), .B2(n14423), .A(n14539), .ZN(n20346) );
  INV_X1 U17979 ( .A(n20346), .ZN(n16447) );
  OAI222_X1 U17980 ( .A1(n14426), .A2(n14899), .B1(n14905), .B2(n14425), .C1(
        n16447), .C2(n14906), .ZN(P1_U2863) );
  OAI21_X1 U17981 ( .B1(n14427), .B2(n14429), .A(n14428), .ZN(n20475) );
  NOR2_X1 U17982 ( .A1(n20504), .A2(n20393), .ZN(n14436) );
  AOI21_X1 U17983 ( .B1(n14431), .B2(n20493), .A(n14433), .ZN(n14586) );
  NOR2_X1 U17984 ( .A1(n20499), .A2(n14586), .ZN(n20488) );
  OAI21_X1 U17985 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20488), .ZN(n14434) );
  INV_X1 U17986 ( .A(n14430), .ZN(n20494) );
  OAI21_X1 U17987 ( .B1(n20495), .B2(n14431), .A(n20494), .ZN(n14432) );
  AOI21_X1 U17988 ( .B1(n14433), .B2(n20499), .A(n14432), .ZN(n20492) );
  OAI22_X1 U17989 ( .A1(n16466), .A2(n14434), .B1(n20492), .B2(n12168), .ZN(
        n14435) );
  AOI211_X1 U17990 ( .C1(n20473), .C2(P1_REIP_REG_4__SCAN_IN), .A(n14436), .B(
        n14435), .ZN(n14437) );
  OAI21_X1 U17991 ( .B1(n20475), .B2(n16424), .A(n14437), .ZN(P1_U3027) );
  AND2_X1 U17992 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n14533) );
  NOR3_X1 U17993 ( .A1(n17659), .A2(n14440), .A3(n14439), .ZN(n14441) );
  NOR2_X1 U17994 ( .A1(n17659), .A2(n17560), .ZN(n17568) );
  INV_X1 U17995 ( .A(n17568), .ZN(n17566) );
  INV_X1 U17996 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17333) );
  INV_X1 U17997 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17559) );
  NAND2_X1 U17998 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17561) );
  NOR2_X1 U17999 ( .A1(n17559), .A2(n17561), .ZN(n17551) );
  NAND3_X1 U18000 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17551), .ZN(n17537) );
  AND2_X1 U18001 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17538) );
  NAND4_X1 U18002 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n17548), .A4(n17538), .ZN(n17539) );
  NAND4_X1 U18003 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n14442)
         );
  NOR2_X1 U18004 ( .A1(n17539), .A2(n14442), .ZN(n14443) );
  NAND4_X1 U18005 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(n14443), .ZN(n17432) );
  NAND3_X1 U18006 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(n17400), .ZN(n17377) );
  NAND2_X1 U18007 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17320), .ZN(n14532) );
  NAND2_X1 U18008 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17310), .ZN(n17301) );
  NAND2_X1 U18009 ( .A1(n17556), .A2(n17301), .ZN(n17299) );
  OAI21_X1 U18010 ( .B1(n14533), .B2(n17566), .A(n17299), .ZN(n16091) );
  AOI22_X1 U18011 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17423), .B1(
        P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n10308), .ZN(n14447) );
  AOI22_X1 U18012 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n9719), .B1(
        P3_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n17325), .ZN(n14446) );
  AOI22_X1 U18013 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n9731), .ZN(n14445) );
  AOI22_X1 U18014 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14444) );
  NAND4_X1 U18015 ( .A1(n14447), .A2(n14446), .A3(n14445), .A4(n14444), .ZN(
        n14453) );
  AOI22_X1 U18016 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n14519), .ZN(n14451) );
  AOI22_X1 U18017 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17503), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U18018 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n17448), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n14517), .ZN(n14449) );
  AOI22_X1 U18019 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n17526), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14448) );
  NAND4_X1 U18020 ( .A1(n14451), .A2(n14450), .A3(n14449), .A4(n14448), .ZN(
        n14452) );
  NOR2_X1 U18021 ( .A1(n14453), .A2(n14452), .ZN(n14531) );
  AOI22_X1 U18022 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14457) );
  AOI22_X1 U18023 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U18024 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U18025 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14454) );
  NAND4_X1 U18026 ( .A1(n14457), .A2(n14456), .A3(n14455), .A4(n14454), .ZN(
        n14464) );
  AOI22_X1 U18027 ( .A1(n14517), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U18028 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14461) );
  AOI22_X1 U18029 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U18030 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14459) );
  NAND4_X1 U18031 ( .A1(n14462), .A2(n14461), .A3(n14460), .A4(n14459), .ZN(
        n14463) );
  NOR2_X1 U18032 ( .A1(n14464), .A2(n14463), .ZN(n17297) );
  AOI22_X1 U18033 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14468) );
  AOI22_X1 U18034 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U18035 ( .A1(n17526), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U18036 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9732), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14465) );
  NAND4_X1 U18037 ( .A1(n14468), .A2(n14467), .A3(n14466), .A4(n14465), .ZN(
        n14475) );
  AOI22_X1 U18038 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U18039 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14472) );
  AOI22_X1 U18040 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U18041 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14470) );
  NAND4_X1 U18042 ( .A1(n14473), .A2(n14472), .A3(n14471), .A4(n14470), .ZN(
        n14474) );
  NOR2_X1 U18043 ( .A1(n14475), .A2(n14474), .ZN(n17307) );
  AOI22_X1 U18044 ( .A1(n10308), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U18045 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U18046 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U18047 ( .A1(n11673), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14476) );
  NAND4_X1 U18048 ( .A1(n14479), .A2(n14478), .A3(n14477), .A4(n14476), .ZN(
        n14486) );
  AOI22_X1 U18049 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U18050 ( .A1(n11704), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U18051 ( .A1(n17533), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U18052 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14481) );
  NAND4_X1 U18053 ( .A1(n14484), .A2(n14483), .A3(n14482), .A4(n14481), .ZN(
        n14485) );
  NOR2_X1 U18054 ( .A1(n14486), .A2(n14485), .ZN(n17316) );
  AOI22_X1 U18055 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14490) );
  AOI22_X1 U18056 ( .A1(n17526), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U18057 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U18058 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14487) );
  NAND4_X1 U18059 ( .A1(n14490), .A2(n14489), .A3(n14488), .A4(n14487), .ZN(
        n14496) );
  AOI22_X1 U18060 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U18061 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17504), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14493) );
  AOI22_X1 U18062 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U18063 ( .A1(n14517), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14491) );
  NAND4_X1 U18064 ( .A1(n14494), .A2(n14493), .A3(n14492), .A4(n14491), .ZN(
        n14495) );
  NOR2_X1 U18065 ( .A1(n14496), .A2(n14495), .ZN(n17317) );
  NOR2_X1 U18066 ( .A1(n17316), .A2(n17317), .ZN(n17315) );
  AOI22_X1 U18067 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U18068 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U18069 ( .A1(n17477), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9731), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14497) );
  OAI21_X1 U18070 ( .B1(n10245), .B2(n21310), .A(n14497), .ZN(n14503) );
  AOI22_X1 U18071 ( .A1(n14517), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14501) );
  AOI22_X1 U18072 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14500) );
  AOI22_X1 U18073 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14499) );
  AOI22_X1 U18074 ( .A1(n17526), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14498) );
  NAND4_X1 U18075 ( .A1(n14501), .A2(n14500), .A3(n14499), .A4(n14498), .ZN(
        n14502) );
  AOI211_X1 U18076 ( .C1(n17325), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n14503), .B(n14502), .ZN(n14504) );
  NAND3_X1 U18077 ( .A1(n14506), .A2(n14505), .A3(n14504), .ZN(n17312) );
  NAND2_X1 U18078 ( .A1(n17315), .A2(n17312), .ZN(n17311) );
  NOR2_X1 U18079 ( .A1(n17307), .A2(n17311), .ZN(n17306) );
  AOI22_X1 U18080 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14516) );
  AOI22_X1 U18081 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14515) );
  INV_X1 U18082 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n21246) );
  AOI22_X1 U18083 ( .A1(n10308), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14507) );
  OAI21_X1 U18084 ( .B1(n10245), .B2(n21246), .A(n14507), .ZN(n14513) );
  AOI22_X1 U18085 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U18086 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U18087 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17448), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U18088 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14508) );
  NAND4_X1 U18089 ( .A1(n14511), .A2(n14510), .A3(n14509), .A4(n14508), .ZN(
        n14512) );
  AOI211_X1 U18090 ( .C1(n11673), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n14513), .B(n14512), .ZN(n14514) );
  NAND3_X1 U18091 ( .A1(n14516), .A2(n14515), .A3(n14514), .ZN(n17303) );
  NAND2_X1 U18092 ( .A1(n17306), .A2(n17303), .ZN(n17302) );
  NOR2_X1 U18093 ( .A1(n17297), .A2(n17302), .ZN(n17296) );
  AOI22_X1 U18094 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U18095 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14529) );
  AOI22_X1 U18096 ( .A1(n17533), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14518) );
  OAI21_X1 U18097 ( .B1(n10245), .B2(n18577), .A(n14518), .ZN(n14527) );
  AOI22_X1 U18098 ( .A1(n11671), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14525) );
  AOI22_X1 U18099 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14524) );
  AOI22_X1 U18100 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14523) );
  AOI22_X1 U18101 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14522) );
  NAND4_X1 U18102 ( .A1(n14525), .A2(n14524), .A3(n14523), .A4(n14522), .ZN(
        n14526) );
  AOI211_X1 U18103 ( .C1(n17505), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n14527), .B(n14526), .ZN(n14528) );
  NAND3_X1 U18104 ( .A1(n14530), .A2(n14529), .A3(n14528), .ZN(n16089) );
  NAND2_X1 U18105 ( .A1(n17296), .A2(n16089), .ZN(n16088) );
  NOR2_X1 U18106 ( .A1(n14531), .A2(n16088), .ZN(n17293) );
  AOI21_X1 U18107 ( .B1(n14531), .B2(n16088), .A(n17293), .ZN(n17584) );
  AOI22_X1 U18108 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16091), .B1(n17584), 
        .B2(n17569), .ZN(n14536) );
  INV_X1 U18109 ( .A(n14532), .ZN(n17314) );
  NAND3_X1 U18110 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(n14533), .ZN(n17273) );
  INV_X1 U18111 ( .A(n17273), .ZN(n14534) );
  NAND3_X1 U18112 ( .A1(n17314), .A2(n17275), .A3(n14534), .ZN(n14535) );
  NAND2_X1 U18113 ( .A1(n14536), .A2(n14535), .ZN(P3_U2674) );
  XOR2_X1 U18114 ( .A(n14537), .B(n10184), .Z(n15141) );
  OR2_X1 U18115 ( .A1(n14539), .A2(n14538), .ZN(n14540) );
  NAND2_X1 U18116 ( .A1(n14600), .A2(n14540), .ZN(n16441) );
  OAI22_X1 U18117 ( .A1(n16441), .A2(n14906), .B1(n14541), .B2(n20408), .ZN(
        n14542) );
  AOI21_X1 U18118 ( .B1(n15141), .B2(n20405), .A(n14542), .ZN(n14543) );
  INV_X1 U18119 ( .A(n14543), .ZN(P1_U2862) );
  INV_X1 U18120 ( .A(n15141), .ZN(n14554) );
  NAND2_X1 U18121 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .ZN(n14545) );
  NOR2_X1 U18122 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14545), .ZN(n14551) );
  AOI21_X1 U18123 ( .B1(n21395), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21393), .ZN(n14544) );
  OAI21_X1 U18124 ( .B1(n21398), .B2(n15139), .A(n14544), .ZN(n14550) );
  INV_X1 U18125 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20362) );
  NOR4_X1 U18126 ( .A1(n20374), .A2(n14545), .A3(n21007), .A4(n20362), .ZN(
        n14546) );
  NAND3_X1 U18127 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(n14546), .ZN(n14647) );
  NOR2_X1 U18128 ( .A1(n14547), .A2(n14647), .ZN(n16282) );
  NOR2_X1 U18129 ( .A1(n16281), .A2(n16282), .ZN(n16302) );
  AOI22_X1 U18130 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n20378), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n16302), .ZN(n14548) );
  OAI21_X1 U18131 ( .B1(n21390), .B2(n16441), .A(n14548), .ZN(n14549) );
  AOI211_X1 U18132 ( .C1(n14551), .C2(n20340), .A(n14550), .B(n14549), .ZN(
        n14552) );
  OAI21_X1 U18133 ( .B1(n14554), .B2(n21403), .A(n14552), .ZN(P1_U2830) );
  MUX2_X1 U18134 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14918), .Z(
        n20446) );
  AOI22_X1 U18135 ( .A1(n14983), .A2(n20446), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14982), .ZN(n14553) );
  OAI21_X1 U18136 ( .B1(n14554), .B2(n14990), .A(n14553), .ZN(P1_U2894) );
  INV_X1 U18137 ( .A(n19452), .ZN(n14581) );
  NAND2_X1 U18138 ( .A1(n10049), .A2(n15386), .ZN(n14556) );
  XNOR2_X1 U18139 ( .A(n19633), .B(n14556), .ZN(n14557) );
  NAND2_X1 U18140 ( .A1(n14557), .A2(n19416), .ZN(n14567) );
  AOI21_X1 U18141 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n19668) );
  NOR2_X1 U18142 ( .A1(n14561), .A2(n19447), .ZN(n14563) );
  INV_X1 U18143 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20204) );
  OAI22_X1 U18144 ( .A1(n20204), .A2(n19440), .B1(n19641), .B2(n19420), .ZN(
        n14562) );
  AOI211_X1 U18145 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n19444), .A(n14563), .B(
        n14562), .ZN(n14564) );
  OAI21_X1 U18146 ( .B1(n19668), .B2(n19442), .A(n14564), .ZN(n14565) );
  AOI21_X1 U18147 ( .B1(n9750), .B2(n19449), .A(n14565), .ZN(n14566) );
  OAI211_X1 U18148 ( .C1(n14581), .C2(n20271), .A(n14567), .B(n14566), .ZN(
        P2_U2853) );
  NOR2_X1 U18149 ( .A1(n19410), .A2(n14568), .ZN(n14570) );
  XNOR2_X1 U18150 ( .A(n14570), .B(n14569), .ZN(n14571) );
  NAND2_X1 U18151 ( .A1(n14571), .A2(n19416), .ZN(n14580) );
  OAI22_X1 U18152 ( .A1(n14572), .A2(n19420), .B1(n20205), .B2(n19440), .ZN(
        n14576) );
  OAI22_X1 U18153 ( .A1(n19429), .A2(n14574), .B1(n14573), .B2(n19447), .ZN(
        n14575) );
  NOR2_X1 U18154 ( .A1(n14576), .A2(n14575), .ZN(n14577) );
  OAI21_X1 U18155 ( .B1(n19494), .B2(n19442), .A(n14577), .ZN(n14578) );
  AOI21_X1 U18156 ( .B1(n13088), .B2(n19449), .A(n14578), .ZN(n14579) );
  OAI211_X1 U18157 ( .C1(n20264), .C2(n14581), .A(n14580), .B(n14579), .ZN(
        P2_U2852) );
  XNOR2_X1 U18158 ( .A(n14582), .B(n15301), .ZN(n14583) );
  XNOR2_X1 U18159 ( .A(n14584), .B(n14583), .ZN(n14594) );
  OAI21_X1 U18160 ( .B1(n14681), .B2(n14585), .A(n20492), .ZN(n16463) );
  NAND2_X1 U18161 ( .A1(n20473), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n14591) );
  OAI21_X1 U18162 ( .B1(n20365), .B2(n20504), .A(n14591), .ZN(n14588) );
  INV_X1 U18163 ( .A(n14586), .ZN(n16419) );
  NAND2_X1 U18164 ( .A1(n16434), .A2(n16419), .ZN(n16432) );
  NOR2_X1 U18165 ( .A1(n16432), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14587) );
  AOI211_X1 U18166 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16463), .A(
        n14588), .B(n14587), .ZN(n14589) );
  OAI21_X1 U18167 ( .B1(n14594), .B2(n16424), .A(n14589), .ZN(P1_U3025) );
  NAND2_X1 U18168 ( .A1(n20474), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14590) );
  OAI211_X1 U18169 ( .C1(n20482), .C2(n20372), .A(n14591), .B(n14590), .ZN(
        n14592) );
  AOI21_X1 U18170 ( .B1(n20369), .B2(n20477), .A(n14592), .ZN(n14593) );
  OAI21_X1 U18171 ( .B1(n14594), .B2(n20321), .A(n14593), .ZN(P1_U2993) );
  INV_X1 U18172 ( .A(n14596), .ZN(n14597) );
  AOI21_X1 U18173 ( .B1(n14599), .B2(n14598), .A(n14597), .ZN(n16352) );
  INV_X1 U18174 ( .A(n16352), .ZN(n14989) );
  AOI21_X1 U18175 ( .B1(n14601), .B2(n14600), .A(n10022), .ZN(n16426) );
  AOI22_X1 U18176 ( .A1(n16426), .A2(n20404), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n13978), .ZN(n14602) );
  OAI21_X1 U18177 ( .B1(n14989), .B2(n14899), .A(n14602), .ZN(P1_U2861) );
  OAI21_X1 U18178 ( .B1(n14605), .B2(n14604), .A(n14603), .ZN(n14900) );
  MUX2_X1 U18179 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14918), .Z(
        n20450) );
  AOI22_X1 U18180 ( .A1(n14983), .A2(n20450), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14982), .ZN(n14606) );
  OAI21_X1 U18181 ( .B1(n14900), .B2(n14990), .A(n14606), .ZN(P1_U2892) );
  INV_X1 U18182 ( .A(n19229), .ZN(n19173) );
  AOI21_X1 U18183 ( .B1(n19012), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16093) );
  OR2_X1 U18184 ( .A1(n14608), .A2(n16093), .ZN(n19007) );
  NOR2_X1 U18185 ( .A1(n19173), .A2(n19007), .ZN(n14614) );
  NAND2_X1 U18186 ( .A1(n19001), .A2(n19210), .ZN(n14612) );
  NOR2_X1 U18187 ( .A1(n19215), .A2(n17781), .ZN(n17783) );
  INV_X1 U18188 ( .A(n19088), .ZN(n19214) );
  OAI21_X1 U18189 ( .B1(n14607), .B2(n17783), .A(n19214), .ZN(n17723) );
  NOR3_X1 U18190 ( .A1(n16206), .A2(n14610), .A3(n14609), .ZN(n14611) );
  OAI21_X1 U18191 ( .B1(n14612), .B2(n17723), .A(n14611), .ZN(n19035) );
  NOR2_X1 U18192 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19169), .ZN(n18546) );
  INV_X1 U18193 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18535) );
  NAND3_X1 U18194 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n19167)
         );
  NOR2_X1 U18195 ( .A1(n18535), .A2(n19167), .ZN(n14613) );
  MUX2_X1 U18196 ( .A(n14614), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19199), .Z(P3_U3284) );
  AOI22_X1 U18197 ( .A1(n12498), .A2(n14616), .B1(n14615), .B2(n11845), .ZN(
        n16152) );
  OAI21_X1 U18198 ( .B1(n16152), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n21247), 
        .ZN(n14617) );
  AOI22_X1 U18199 ( .A1(n14617), .A2(n14627), .B1(n11845), .B2(n16183), .ZN(
        n14620) );
  INV_X1 U18200 ( .A(n16475), .ZN(n14619) );
  AOI21_X1 U18201 ( .B1(n16154), .B2(n16471), .A(n14619), .ZN(n14618) );
  OAI22_X1 U18202 ( .A1(n14620), .A2(n14619), .B1(n14618), .B2(n11845), .ZN(
        P1_U3474) );
  NOR3_X1 U18203 ( .A1(n14621), .A2(n13638), .A3(n14032), .ZN(n14624) );
  NOR2_X1 U18204 ( .A1(n14172), .A2(n14622), .ZN(n14623) );
  AOI211_X1 U18205 ( .C1(n16154), .C2(n14633), .A(n14624), .B(n14623), .ZN(
        n16157) );
  NOR2_X1 U18206 ( .A1(n16157), .A2(n14625), .ZN(n14631) );
  NAND2_X1 U18207 ( .A1(n14626), .A2(n16183), .ZN(n14629) );
  OAI22_X1 U18208 ( .A1(n14629), .A2(n14032), .B1(n14628), .B2(n14627), .ZN(
        n14630) );
  OAI21_X1 U18209 ( .B1(n14631), .B2(n14630), .A(n16475), .ZN(n14632) );
  OAI21_X1 U18210 ( .B1(n16475), .B2(n14633), .A(n14632), .ZN(P1_U3473) );
  NOR2_X1 U18211 ( .A1(n14637), .A2(n14634), .ZN(n14635) );
  NOR3_X4 U18212 ( .A1(n14982), .A2(n14637), .A3(n14918), .ZN(n14971) );
  AOI22_X1 U18213 ( .A1(n14971), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14982), .ZN(n14638) );
  OAI211_X1 U18214 ( .C1(n14969), .C2(n16811), .A(n14639), .B(n14638), .ZN(
        P1_U2873) );
  OAI22_X1 U18215 ( .A1(n9730), .A2(n12409), .B1(n14734), .B2(n14643), .ZN(
        n14646) );
  INV_X1 U18216 ( .A(n14644), .ZN(n14645) );
  XNOR2_X1 U18217 ( .A(n14646), .B(n14645), .ZN(n14665) );
  INV_X1 U18218 ( .A(n14665), .ZN(n15166) );
  INV_X1 U18219 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14666) );
  INV_X1 U18220 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21385) );
  INV_X1 U18221 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21387) );
  INV_X1 U18222 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n16412) );
  INV_X1 U18223 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16303) );
  NOR4_X1 U18224 ( .A1(n21385), .A2(n21387), .A3(n16412), .A4(n16303), .ZN(
        n14649) );
  NAND2_X1 U18225 ( .A1(n16304), .A2(n14649), .ZN(n16273) );
  NAND2_X1 U18226 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16261) );
  NOR2_X1 U18227 ( .A1(n16273), .A2(n16261), .ZN(n16257) );
  NAND2_X1 U18228 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14813) );
  INV_X1 U18229 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21022) );
  NOR2_X1 U18230 ( .A1(n14813), .A2(n21022), .ZN(n14648) );
  NAND2_X1 U18231 ( .A1(n16239), .A2(n14648), .ZN(n16225) );
  NAND3_X1 U18232 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n14650) );
  NOR2_X1 U18233 ( .A1(n16225), .A2(n14650), .ZN(n14758) );
  AND3_X1 U18234 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n14652) );
  NAND2_X1 U18235 ( .A1(n14758), .A2(n14652), .ZN(n14755) );
  NAND2_X1 U18236 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14725) );
  INV_X1 U18237 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n15006) );
  NOR3_X1 U18238 ( .A1(n14755), .A2(n14725), .A3(n15006), .ZN(n14712) );
  AND2_X1 U18239 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14655) );
  INV_X1 U18240 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21018) );
  NAND2_X1 U18241 ( .A1(n14649), .A2(n16282), .ZN(n16262) );
  NOR3_X1 U18242 ( .A1(n21018), .A2(n16261), .A3(n16262), .ZN(n16237) );
  AND2_X1 U18243 ( .A1(n16237), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14815) );
  NOR2_X1 U18244 ( .A1(n14813), .A2(n14650), .ZN(n14651) );
  NAND2_X1 U18245 ( .A1(n14815), .A2(n14651), .ZN(n14771) );
  INV_X1 U18246 ( .A(n14652), .ZN(n14653) );
  OR2_X1 U18247 ( .A1(n14771), .A2(n14653), .ZN(n14747) );
  OR2_X1 U18248 ( .A1(n14725), .A2(n14747), .ZN(n14654) );
  NAND2_X1 U18249 ( .A1(n20356), .A2(n14654), .ZN(n14740) );
  OAI21_X1 U18250 ( .B1(n16281), .B2(n14655), .A(n14740), .ZN(n14711) );
  OAI21_X1 U18251 ( .B1(n14712), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14711), 
        .ZN(n14658) );
  INV_X1 U18252 ( .A(n14999), .ZN(n14656) );
  AOI22_X1 U18253 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21395), .B1(
        n20341), .B2(n14656), .ZN(n14657) );
  OAI211_X1 U18254 ( .C1(n21391), .C2(n14666), .A(n14658), .B(n14657), .ZN(
        n14659) );
  AOI21_X1 U18255 ( .B1(n15166), .B2(n20377), .A(n14659), .ZN(n14660) );
  OAI21_X1 U18256 ( .B1(n14996), .B2(n21403), .A(n14660), .ZN(P1_U2810) );
  AOI22_X1 U18257 ( .A1(n14964), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14982), .ZN(n14664) );
  NOR3_X4 U18258 ( .A1(n14982), .A2(n14662), .A3(n14661), .ZN(n14973) );
  MUX2_X1 U18259 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14918), .Z(
        n20454) );
  AOI22_X1 U18260 ( .A1(n14973), .A2(n20454), .B1(n14971), .B2(DATAI_30_), 
        .ZN(n14663) );
  OAI211_X1 U18261 ( .C1(n14996), .C2(n14990), .A(n14664), .B(n14663), .ZN(
        P1_U2874) );
  OAI222_X1 U18262 ( .A1(n14899), .A2(n14996), .B1(n14905), .B2(n14666), .C1(
        n14665), .C2(n14906), .ZN(P1_U2842) );
  NAND2_X1 U18263 ( .A1(n14668), .A2(n20498), .ZN(n14674) );
  NAND2_X1 U18264 ( .A1(n14674), .A2(n12479), .ZN(n14673) );
  NOR2_X1 U18265 ( .A1(n12460), .A2(n20337), .ZN(n14678) );
  AOI21_X1 U18266 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14678), .ZN(n14669) );
  OAI21_X1 U18267 ( .B1(n20482), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14669), .ZN(n14670) );
  AOI21_X1 U18268 ( .B1(n14671), .B2(n20477), .A(n14670), .ZN(n14672) );
  OAI21_X1 U18269 ( .B1(n14667), .B2(n14673), .A(n14672), .ZN(P1_U2998) );
  NAND2_X1 U18270 ( .A1(n14674), .A2(n20507), .ZN(n14684) );
  INV_X1 U18271 ( .A(n14675), .ZN(n14679) );
  NOR2_X1 U18272 ( .A1(n20498), .A2(n14676), .ZN(n14677) );
  AOI211_X1 U18273 ( .C1(n20486), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        n14683) );
  OR3_X1 U18274 ( .A1(n14681), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14680), .ZN(n14682) );
  OAI211_X1 U18275 ( .C1(n14667), .C2(n14684), .A(n14683), .B(n14682), .ZN(
        P1_U3030) );
  AOI22_X1 U18276 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19461), .B1(n19460), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14692) );
  NAND2_X1 U18277 ( .A1(n14688), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14690) );
  INV_X1 U18278 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14687) );
  OR2_X1 U18279 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  NAND2_X1 U18280 ( .A1(n14690), .A2(n14689), .ZN(n19605) );
  AOI22_X1 U18281 ( .A1(n19459), .A2(n19605), .B1(n19522), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14691) );
  OAI211_X1 U18282 ( .C1(n15777), .C2(n15576), .A(n14692), .B(n14691), .ZN(
        n14693) );
  AOI21_X1 U18283 ( .B1(n14694), .B2(n19505), .A(n14693), .ZN(n14695) );
  INV_X1 U18284 ( .A(n14695), .ZN(P2_U2889) );
  INV_X1 U18285 ( .A(n14696), .ZN(n14702) );
  OR2_X1 U18286 ( .A1(n14697), .A2(n12318), .ZN(n14698) );
  NOR2_X1 U18287 ( .A1(n14699), .A2(n14698), .ZN(n14701) );
  MUX2_X1 U18288 ( .A(n14702), .B(n14701), .S(n14700), .Z(n14706) );
  INV_X1 U18289 ( .A(n14703), .ZN(n14704) );
  NAND2_X1 U18290 ( .A1(n12312), .A2(n14704), .ZN(n14705) );
  NAND2_X1 U18291 ( .A1(n14706), .A2(n14705), .ZN(n16170) );
  NOR2_X1 U18292 ( .A1(n14707), .A2(n11980), .ZN(n21061) );
  OAI21_X1 U18293 ( .B1(n21061), .B2(n20985), .A(n14708), .ZN(n16168) );
  AND2_X1 U18294 ( .A1(n16168), .A2(n14709), .ZN(n20323) );
  MUX2_X1 U18295 ( .A(P1_MORE_REG_SCAN_IN), .B(n16170), .S(n20323), .Z(
        P1_U3484) );
  INV_X1 U18296 ( .A(n14710), .ZN(n14719) );
  INV_X1 U18297 ( .A(n14711), .ZN(n14716) );
  NAND3_X1 U18298 ( .A1(n14712), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n14715), 
        .ZN(n14714) );
  AOI22_X1 U18299 ( .A1(n20378), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21395), .ZN(n14713) );
  OAI211_X1 U18300 ( .C1(n14716), .C2(n14715), .A(n14714), .B(n14713), .ZN(
        n14717) );
  AOI21_X1 U18301 ( .B1(n14829), .B2(n20377), .A(n14717), .ZN(n14718) );
  OAI21_X1 U18302 ( .B1(n14719), .B2(n21403), .A(n14718), .ZN(P1_U2809) );
  AND2_X1 U18303 ( .A1(n14734), .A2(n14720), .ZN(n14722) );
  NAND2_X1 U18304 ( .A1(n15010), .A2(n20368), .ZN(n14731) );
  INV_X1 U18305 ( .A(n14755), .ZN(n14742) );
  NOR2_X1 U18306 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14725), .ZN(n14729) );
  AOI22_X1 U18307 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n21395), .B1(
        n20341), .B2(n15005), .ZN(n14727) );
  NAND2_X1 U18308 ( .A1(n20378), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14726) );
  OAI211_X1 U18309 ( .C1(n14740), .C2(n15006), .A(n14727), .B(n14726), .ZN(
        n14728) );
  AOI21_X1 U18310 ( .B1(n14742), .B2(n14729), .A(n14728), .ZN(n14730) );
  OAI211_X1 U18311 ( .C1(n21390), .C2(n15174), .A(n14731), .B(n14730), .ZN(
        P1_U2811) );
  INV_X1 U18312 ( .A(n14734), .ZN(n14735) );
  AOI21_X1 U18313 ( .B1(n14736), .B2(n14749), .A(n14735), .ZN(n15182) );
  INV_X1 U18314 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21035) );
  OAI22_X1 U18315 ( .A1(n14737), .A2(n20389), .B1(n21398), .B2(n15020), .ZN(
        n14738) );
  AOI21_X1 U18316 ( .B1(n20378), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14738), .ZN(
        n14739) );
  OAI21_X1 U18317 ( .B1(n21035), .B2(n14740), .A(n14739), .ZN(n14741) );
  AOI21_X1 U18318 ( .B1(n15182), .B2(n20377), .A(n14741), .ZN(n14744) );
  NAND3_X1 U18319 ( .A1(n14742), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n21035), 
        .ZN(n14743) );
  OAI211_X1 U18320 ( .C1(n15018), .C2(n21403), .A(n14744), .B(n14743), .ZN(
        P1_U2812) );
  AOI21_X1 U18321 ( .B1(n14746), .B2(n14745), .A(n14732), .ZN(n15031) );
  NAND2_X1 U18322 ( .A1(n15031), .A2(n20368), .ZN(n14754) );
  AND2_X1 U18323 ( .A1(n14747), .A2(n20356), .ZN(n14767) );
  INV_X1 U18324 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14834) );
  AOI22_X1 U18325 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n21395), .B1(
        n20341), .B2(n15026), .ZN(n14748) );
  OAI21_X1 U18326 ( .B1(n21391), .B2(n14834), .A(n14748), .ZN(n14752) );
  OAI21_X1 U18327 ( .B1(n14761), .B2(n14750), .A(n14749), .ZN(n15192) );
  NOR2_X1 U18328 ( .A1(n15192), .A2(n21390), .ZN(n14751) );
  AOI211_X1 U18329 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14767), .A(n14752), 
        .B(n14751), .ZN(n14753) );
  OAI211_X1 U18330 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14755), .A(n14754), 
        .B(n14753), .ZN(P1_U2813) );
  OAI21_X1 U18331 ( .B1(n14756), .B2(n14757), .A(n14745), .ZN(n15037) );
  INV_X1 U18332 ( .A(n14758), .ZN(n14786) );
  INV_X1 U18333 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15049) );
  INV_X1 U18334 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21028) );
  NOR4_X1 U18335 ( .A1(n14786), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n15049), 
        .A4(n21028), .ZN(n14766) );
  NOR2_X1 U18336 ( .A1(n14774), .A2(n14759), .ZN(n14760) );
  OR2_X1 U18337 ( .A1(n14761), .A2(n14760), .ZN(n15199) );
  INV_X1 U18338 ( .A(n15039), .ZN(n14762) );
  AOI22_X1 U18339 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21395), .B1(
        n20341), .B2(n14762), .ZN(n14764) );
  NAND2_X1 U18340 ( .A1(n20378), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14763) );
  OAI211_X1 U18341 ( .C1(n15199), .C2(n21390), .A(n14764), .B(n14763), .ZN(
        n14765) );
  AOI211_X1 U18342 ( .C1(n14767), .C2(P1_REIP_REG_26__SCAN_IN), .A(n14766), 
        .B(n14765), .ZN(n14768) );
  OAI21_X1 U18343 ( .B1(n15037), .B2(n21403), .A(n14768), .ZN(P1_U2814) );
  INV_X1 U18344 ( .A(n14769), .ZN(n14784) );
  AOI21_X1 U18345 ( .B1(n14770), .B2(n14784), .A(n14756), .ZN(n15053) );
  INV_X1 U18346 ( .A(n15053), .ZN(n14929) );
  AND2_X1 U18347 ( .A1(n14771), .A2(n20356), .ZN(n14811) );
  XNOR2_X1 U18348 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14772) );
  NOR2_X1 U18349 ( .A1(n14786), .A2(n14772), .ZN(n14781) );
  AND2_X1 U18350 ( .A1(n14789), .A2(n14773), .ZN(n14775) );
  OR2_X1 U18351 ( .A1(n14775), .A2(n14774), .ZN(n15213) );
  INV_X1 U18352 ( .A(n14776), .ZN(n15051) );
  OAI22_X1 U18353 ( .A1(n14777), .A2(n20389), .B1(n21398), .B2(n15051), .ZN(
        n14778) );
  AOI21_X1 U18354 ( .B1(n20378), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14778), .ZN(
        n14779) );
  OAI21_X1 U18355 ( .B1(n15213), .B2(n21390), .A(n14779), .ZN(n14780) );
  AOI211_X1 U18356 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14811), .A(n14781), 
        .B(n14780), .ZN(n14782) );
  OAI21_X1 U18357 ( .B1(n14929), .B2(n21403), .A(n14782), .ZN(P1_U2815) );
  AOI21_X1 U18358 ( .B1(n14785), .B2(n14799), .A(n14769), .ZN(n15061) );
  INV_X1 U18359 ( .A(n15061), .ZN(n14935) );
  NOR2_X1 U18360 ( .A1(n14786), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14795) );
  NAND2_X1 U18361 ( .A1(n14806), .A2(n14787), .ZN(n14788) );
  NAND2_X1 U18362 ( .A1(n14789), .A2(n14788), .ZN(n15220) );
  INV_X1 U18363 ( .A(n14790), .ZN(n15059) );
  OAI22_X1 U18364 ( .A1(n14791), .A2(n20389), .B1(n21398), .B2(n15059), .ZN(
        n14792) );
  AOI21_X1 U18365 ( .B1(n20378), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14792), .ZN(
        n14793) );
  OAI21_X1 U18366 ( .B1(n15220), .B2(n21390), .A(n14793), .ZN(n14794) );
  AOI211_X1 U18367 ( .C1(n14811), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14795), 
        .B(n14794), .ZN(n14796) );
  OAI21_X1 U18368 ( .B1(n14935), .B2(n21403), .A(n14796), .ZN(P1_U2816) );
  INV_X1 U18369 ( .A(n14798), .ZN(n14801) );
  INV_X1 U18370 ( .A(n14799), .ZN(n14800) );
  AOI21_X1 U18371 ( .B1(n14802), .B2(n14801), .A(n14800), .ZN(n15071) );
  INV_X1 U18372 ( .A(n15071), .ZN(n14939) );
  NAND2_X1 U18373 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14803) );
  INV_X1 U18374 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15067) );
  OAI21_X1 U18375 ( .B1(n16225), .B2(n14803), .A(n15067), .ZN(n14810) );
  NAND2_X1 U18376 ( .A1(n14845), .A2(n14804), .ZN(n14805) );
  NAND2_X1 U18377 ( .A1(n14806), .A2(n14805), .ZN(n15230) );
  AOI22_X1 U18378 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n21395), .B1(
        n20341), .B2(n15066), .ZN(n14808) );
  NAND2_X1 U18379 ( .A1(n20378), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n14807) );
  OAI211_X1 U18380 ( .C1(n15230), .C2(n21390), .A(n14808), .B(n14807), .ZN(
        n14809) );
  AOI21_X1 U18381 ( .B1(n14811), .B2(n14810), .A(n14809), .ZN(n14812) );
  OAI21_X1 U18382 ( .B1(n14939), .B2(n21403), .A(n14812), .ZN(P1_U2817) );
  INV_X1 U18383 ( .A(n14813), .ZN(n14814) );
  AOI21_X1 U18384 ( .B1(n16239), .B2(n14814), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14828) );
  NAND2_X1 U18385 ( .A1(n14815), .A2(n14814), .ZN(n14816) );
  AND2_X1 U18386 ( .A1(n14816), .A2(n20356), .ZN(n16220) );
  INV_X1 U18387 ( .A(n16220), .ZN(n16214) );
  AOI21_X1 U18388 ( .B1(n14819), .B2(n14817), .A(n14818), .ZN(n15094) );
  NAND2_X1 U18389 ( .A1(n15094), .A2(n20368), .ZN(n14827) );
  INV_X1 U18390 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14820) );
  OAI22_X1 U18391 ( .A1(n14820), .A2(n20389), .B1(n21398), .B2(n15092), .ZN(
        n14825) );
  INV_X1 U18392 ( .A(n9775), .ZN(n14821) );
  AOI21_X1 U18393 ( .B1(n14822), .B2(n9825), .A(n14821), .ZN(n15267) );
  INV_X1 U18394 ( .A(n15267), .ZN(n14823) );
  NOR2_X1 U18395 ( .A1(n14823), .A2(n21390), .ZN(n14824) );
  AOI211_X1 U18396 ( .C1(n20378), .C2(P1_EBX_REG_20__SCAN_IN), .A(n14825), .B(
        n14824), .ZN(n14826) );
  OAI211_X1 U18397 ( .C1(n14828), .C2(n16214), .A(n14827), .B(n14826), .ZN(
        P1_U2820) );
  INV_X1 U18398 ( .A(n14829), .ZN(n14831) );
  INV_X1 U18399 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14830) );
  OAI22_X1 U18400 ( .A1(n14831), .A2(n14906), .B1(n14830), .B2(n14905), .ZN(
        P1_U2841) );
  INV_X1 U18401 ( .A(n15010), .ZN(n14913) );
  OAI222_X1 U18402 ( .A1(n14832), .A2(n20408), .B1(n14906), .B2(n15174), .C1(
        n14913), .C2(n14899), .ZN(P1_U2843) );
  AOI22_X1 U18403 ( .A1(n15182), .A2(n20404), .B1(n13978), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n14833) );
  OAI21_X1 U18404 ( .B1(n15018), .B2(n14899), .A(n14833), .ZN(P1_U2844) );
  INV_X1 U18405 ( .A(n15031), .ZN(n14921) );
  OAI222_X1 U18406 ( .A1(n14834), .A2(n20408), .B1(n14906), .B2(n15192), .C1(
        n14921), .C2(n14899), .ZN(P1_U2845) );
  INV_X1 U18407 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14835) );
  OAI222_X1 U18408 ( .A1(n14835), .A2(n20408), .B1(n14906), .B2(n15199), .C1(
        n15037), .C2(n14899), .ZN(P1_U2846) );
  INV_X1 U18409 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14836) );
  OAI222_X1 U18410 ( .A1(n14836), .A2(n20408), .B1(n14906), .B2(n15213), .C1(
        n14929), .C2(n14899), .ZN(P1_U2847) );
  INV_X1 U18411 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21161) );
  OAI222_X1 U18412 ( .A1(n21161), .A2(n20408), .B1(n14906), .B2(n15220), .C1(
        n14935), .C2(n14899), .ZN(P1_U2848) );
  INV_X1 U18413 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14837) );
  OAI22_X1 U18414 ( .A1(n15230), .A2(n14906), .B1(n14837), .B2(n14905), .ZN(
        n14838) );
  INV_X1 U18415 ( .A(n14838), .ZN(n14839) );
  OAI21_X1 U18416 ( .B1(n14939), .B2(n14899), .A(n14839), .ZN(P1_U2849) );
  AND2_X1 U18417 ( .A1(n14840), .A2(n14841), .ZN(n14842) );
  NOR2_X1 U18418 ( .A1(n14798), .A2(n14842), .ZN(n16216) );
  INV_X1 U18419 ( .A(n16216), .ZN(n14945) );
  INV_X1 U18420 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14846) );
  OR2_X1 U18421 ( .A1(n14851), .A2(n14843), .ZN(n14844) );
  NAND2_X1 U18422 ( .A1(n14845), .A2(n14844), .ZN(n16219) );
  OAI222_X1 U18423 ( .A1(n14899), .A2(n14945), .B1(n14905), .B2(n14846), .C1(
        n16219), .C2(n14906), .ZN(P1_U2850) );
  NAND2_X1 U18424 ( .A1(n10168), .A2(n14847), .ZN(n14848) );
  AND2_X1 U18425 ( .A1(n14840), .A2(n14848), .ZN(n16224) );
  INV_X1 U18426 ( .A(n16224), .ZN(n14951) );
  INV_X1 U18427 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14852) );
  AND2_X1 U18428 ( .A1(n9775), .A2(n14849), .ZN(n14850) );
  OR2_X1 U18429 ( .A1(n14851), .A2(n14850), .ZN(n16222) );
  OAI222_X1 U18430 ( .A1(n14899), .A2(n14951), .B1(n14905), .B2(n14852), .C1(
        n16222), .C2(n14906), .ZN(P1_U2851) );
  INV_X1 U18431 ( .A(n15094), .ZN(n14956) );
  AOI22_X1 U18432 ( .A1(n15267), .A2(n20404), .B1(n13978), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14853) );
  OAI21_X1 U18433 ( .B1(n14956), .B2(n14899), .A(n14853), .ZN(P1_U2852) );
  OR2_X1 U18434 ( .A1(n14854), .A2(n14855), .ZN(n14856) );
  AND2_X1 U18435 ( .A1(n14817), .A2(n14856), .ZN(n16236) );
  INV_X1 U18436 ( .A(n16236), .ZN(n14960) );
  XNOR2_X1 U18437 ( .A(n14867), .B(n14857), .ZN(n16242) );
  OAI22_X1 U18438 ( .A1(n16242), .A2(n14906), .B1(n14858), .B2(n14905), .ZN(
        n14859) );
  INV_X1 U18439 ( .A(n14859), .ZN(n14860) );
  OAI21_X1 U18440 ( .B1(n14960), .B2(n14899), .A(n14860), .ZN(P1_U2853) );
  NOR2_X1 U18441 ( .A1(n14862), .A2(n14863), .ZN(n14864) );
  OR2_X1 U18442 ( .A1(n14854), .A2(n14864), .ZN(n15108) );
  NOR2_X1 U18443 ( .A1(n14875), .A2(n14865), .ZN(n14866) );
  OR2_X1 U18444 ( .A1(n14867), .A2(n14866), .ZN(n16250) );
  OAI22_X1 U18445 ( .A1(n16250), .A2(n14906), .B1(n14868), .B2(n14905), .ZN(
        n14869) );
  INV_X1 U18446 ( .A(n14869), .ZN(n14870) );
  OAI21_X1 U18447 ( .B1(n15108), .B2(n14899), .A(n14870), .ZN(P1_U2854) );
  AND2_X1 U18448 ( .A1(n14871), .A2(n14872), .ZN(n14873) );
  OR2_X1 U18449 ( .A1(n14873), .A2(n14862), .ZN(n15119) );
  AND2_X1 U18450 ( .A1(n14885), .A2(n14874), .ZN(n14876) );
  OR2_X1 U18451 ( .A1(n14876), .A2(n14875), .ZN(n16260) );
  INV_X1 U18452 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14877) );
  OAI22_X1 U18453 ( .A1(n16260), .A2(n14906), .B1(n14877), .B2(n14905), .ZN(
        n14878) );
  INV_X1 U18454 ( .A(n14878), .ZN(n14879) );
  OAI21_X1 U18455 ( .B1(n15119), .B2(n14899), .A(n14879), .ZN(P1_U2855) );
  NAND2_X1 U18456 ( .A1(n14880), .A2(n14881), .ZN(n14882) );
  AND2_X1 U18457 ( .A1(n14871), .A2(n14882), .ZN(n16316) );
  INV_X1 U18458 ( .A(n16316), .ZN(n14976) );
  INV_X1 U18459 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14886) );
  NAND2_X1 U18460 ( .A1(n16269), .A2(n14883), .ZN(n14884) );
  NAND2_X1 U18461 ( .A1(n14885), .A2(n14884), .ZN(n16370) );
  OAI222_X1 U18462 ( .A1(n14899), .A2(n14976), .B1(n14905), .B2(n14886), .C1(
        n16370), .C2(n14906), .ZN(P1_U2856) );
  OAI21_X1 U18463 ( .B1(n9779), .B2(n14888), .A(n14887), .ZN(n21404) );
  INV_X1 U18464 ( .A(n21404), .ZN(n16334) );
  NOR2_X1 U18465 ( .A1(n14897), .A2(n14889), .ZN(n14890) );
  OR2_X1 U18466 ( .A1(n16271), .A2(n14890), .ZN(n21389) );
  OAI22_X1 U18467 ( .A1(n21389), .A2(n14906), .B1(n21392), .B2(n14905), .ZN(
        n14891) );
  AOI21_X1 U18468 ( .B1(n16334), .B2(n20405), .A(n14891), .ZN(n14892) );
  INV_X1 U18469 ( .A(n14892), .ZN(P1_U2858) );
  AND2_X1 U18470 ( .A1(n14603), .A2(n14893), .ZN(n14894) );
  OR2_X1 U18471 ( .A1(n9779), .A2(n14894), .ZN(n16288) );
  AND2_X1 U18472 ( .A1(n14904), .A2(n14895), .ZN(n14896) );
  NOR2_X1 U18473 ( .A1(n14897), .A2(n14896), .ZN(n16405) );
  AOI22_X1 U18474 ( .A1(n16405), .A2(n20404), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n13978), .ZN(n14898) );
  OAI21_X1 U18475 ( .B1(n16288), .B2(n14899), .A(n14898), .ZN(P1_U2859) );
  INV_X1 U18476 ( .A(n14900), .ZN(n16343) );
  NAND2_X1 U18477 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  NAND2_X1 U18478 ( .A1(n14904), .A2(n14903), .ZN(n16415) );
  OAI22_X1 U18479 ( .A1(n16415), .A2(n14906), .B1(n16292), .B2(n14905), .ZN(
        n14907) );
  AOI21_X1 U18480 ( .B1(n16343), .B2(n20405), .A(n14907), .ZN(n14908) );
  INV_X1 U18481 ( .A(n14908), .ZN(P1_U2860) );
  OAI22_X1 U18482 ( .A1(n14969), .A2(n16814), .B1(n14909), .B2(n14985), .ZN(
        n14910) );
  INV_X1 U18483 ( .A(n14910), .ZN(n14912) );
  MUX2_X1 U18484 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14918), .Z(
        n20452) );
  AOI22_X1 U18485 ( .A1(n14973), .A2(n20452), .B1(n14971), .B2(DATAI_29_), 
        .ZN(n14911) );
  OAI211_X1 U18486 ( .C1(n14913), .C2(n14990), .A(n14912), .B(n14911), .ZN(
        P1_U2875) );
  AOI22_X1 U18487 ( .A1(n14964), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14982), .ZN(n14915) );
  AOI22_X1 U18488 ( .A1(n14973), .A2(n20450), .B1(n14971), .B2(DATAI_28_), 
        .ZN(n14914) );
  OAI211_X1 U18489 ( .C1(n15018), .C2(n14990), .A(n14915), .B(n14914), .ZN(
        P1_U2876) );
  OAI22_X1 U18490 ( .A1(n14969), .A2(n16818), .B1(n14916), .B2(n14985), .ZN(
        n14917) );
  INV_X1 U18491 ( .A(n14917), .ZN(n14920) );
  MUX2_X1 U18492 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14918), .Z(
        n20448) );
  AOI22_X1 U18493 ( .A1(n14973), .A2(n20448), .B1(n14971), .B2(DATAI_27_), 
        .ZN(n14919) );
  OAI211_X1 U18494 ( .C1(n14921), .C2(n14990), .A(n14920), .B(n14919), .ZN(
        P1_U2877) );
  OAI22_X1 U18495 ( .A1(n14969), .A2(n16820), .B1(n13603), .B2(n14985), .ZN(
        n14922) );
  INV_X1 U18496 ( .A(n14922), .ZN(n14924) );
  AOI22_X1 U18497 ( .A1(n14973), .A2(n20446), .B1(n14971), .B2(DATAI_26_), 
        .ZN(n14923) );
  OAI211_X1 U18498 ( .C1(n15037), .C2(n14990), .A(n14924), .B(n14923), .ZN(
        P1_U2878) );
  OAI22_X1 U18499 ( .A1(n14969), .A2(n16822), .B1(n14925), .B2(n14985), .ZN(
        n14926) );
  INV_X1 U18500 ( .A(n14926), .ZN(n14928) );
  AOI22_X1 U18501 ( .A1(n14973), .A2(n20444), .B1(n14971), .B2(DATAI_25_), 
        .ZN(n14927) );
  OAI211_X1 U18502 ( .C1(n14929), .C2(n14990), .A(n14928), .B(n14927), .ZN(
        P1_U2879) );
  INV_X1 U18503 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14931) );
  OAI22_X1 U18504 ( .A1(n14969), .A2(n14931), .B1(n14930), .B2(n14985), .ZN(
        n14932) );
  INV_X1 U18505 ( .A(n14932), .ZN(n14934) );
  AOI22_X1 U18506 ( .A1(n14973), .A2(n20442), .B1(n14971), .B2(DATAI_24_), 
        .ZN(n14933) );
  OAI211_X1 U18507 ( .C1(n14935), .C2(n14990), .A(n14934), .B(n14933), .ZN(
        P1_U2880) );
  AOI22_X1 U18508 ( .A1(n14964), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14982), .ZN(n14938) );
  AOI22_X1 U18509 ( .A1(n14973), .A2(n14936), .B1(n14971), .B2(DATAI_23_), 
        .ZN(n14937) );
  OAI211_X1 U18510 ( .C1(n14939), .C2(n14990), .A(n14938), .B(n14937), .ZN(
        P1_U2881) );
  OAI22_X1 U18511 ( .A1(n14969), .A2(n16825), .B1(n14940), .B2(n14985), .ZN(
        n14941) );
  INV_X1 U18512 ( .A(n14941), .ZN(n14944) );
  AOI22_X1 U18513 ( .A1(n14973), .A2(n14942), .B1(n14971), .B2(DATAI_22_), 
        .ZN(n14943) );
  OAI211_X1 U18514 ( .C1(n14945), .C2(n14990), .A(n14944), .B(n14943), .ZN(
        P1_U2882) );
  OAI22_X1 U18515 ( .A1(n14969), .A2(n16828), .B1(n14946), .B2(n14985), .ZN(
        n14947) );
  INV_X1 U18516 ( .A(n14947), .ZN(n14950) );
  AOI22_X1 U18517 ( .A1(n14973), .A2(n14948), .B1(n14971), .B2(DATAI_21_), 
        .ZN(n14949) );
  OAI211_X1 U18518 ( .C1(n14951), .C2(n14990), .A(n14950), .B(n14949), .ZN(
        P1_U2883) );
  OAI22_X1 U18519 ( .A1(n14969), .A2(n21108), .B1(n21072), .B2(n14985), .ZN(
        n14952) );
  INV_X1 U18520 ( .A(n14952), .ZN(n14955) );
  AOI22_X1 U18521 ( .A1(n14973), .A2(n14953), .B1(n14971), .B2(DATAI_20_), 
        .ZN(n14954) );
  OAI211_X1 U18522 ( .C1(n14956), .C2(n14990), .A(n14955), .B(n14954), .ZN(
        P1_U2884) );
  AOI22_X1 U18523 ( .A1(n14964), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14982), .ZN(n14959) );
  AOI22_X1 U18524 ( .A1(n14973), .A2(n14957), .B1(n14971), .B2(DATAI_19_), 
        .ZN(n14958) );
  OAI211_X1 U18525 ( .C1(n14960), .C2(n14990), .A(n14959), .B(n14958), .ZN(
        P1_U2885) );
  AOI22_X1 U18526 ( .A1(n14964), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14982), .ZN(n14963) );
  AOI22_X1 U18527 ( .A1(n14973), .A2(n14961), .B1(n14971), .B2(DATAI_18_), 
        .ZN(n14962) );
  OAI211_X1 U18528 ( .C1(n15108), .C2(n14990), .A(n14963), .B(n14962), .ZN(
        P1_U2886) );
  AOI22_X1 U18529 ( .A1(n14964), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14982), .ZN(n14967) );
  AOI22_X1 U18530 ( .A1(n14973), .A2(n14965), .B1(n14971), .B2(DATAI_17_), 
        .ZN(n14966) );
  OAI211_X1 U18531 ( .C1(n15119), .C2(n14990), .A(n14967), .B(n14966), .ZN(
        P1_U2887) );
  OAI22_X1 U18532 ( .A1(n14969), .A2(n16836), .B1(n14968), .B2(n14985), .ZN(
        n14970) );
  INV_X1 U18533 ( .A(n14970), .ZN(n14975) );
  AOI22_X1 U18534 ( .A1(n14973), .A2(n14972), .B1(n14971), .B2(DATAI_16_), 
        .ZN(n14974) );
  OAI211_X1 U18535 ( .C1(n14976), .C2(n14990), .A(n14975), .B(n14974), .ZN(
        P1_U2888) );
  INV_X1 U18536 ( .A(n14880), .ZN(n14977) );
  AOI21_X1 U18537 ( .B1(n14978), .B2(n14887), .A(n14977), .ZN(n16325) );
  INV_X1 U18538 ( .A(n16325), .ZN(n14980) );
  OAI222_X1 U18539 ( .A1(n14980), .A2(n14990), .B1(n14988), .B2(n14979), .C1(
        n14985), .C2(n13771), .ZN(P1_U2889) );
  AOI22_X1 U18540 ( .A1(n14983), .A2(n20454), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14982), .ZN(n14981) );
  OAI21_X1 U18541 ( .B1(n21404), .B2(n14990), .A(n14981), .ZN(P1_U2890) );
  AOI22_X1 U18542 ( .A1(n14983), .A2(n20452), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14982), .ZN(n14984) );
  OAI21_X1 U18543 ( .B1(n16288), .B2(n14990), .A(n14984), .ZN(P1_U2891) );
  INV_X1 U18544 ( .A(n20448), .ZN(n14987) );
  OAI222_X1 U18545 ( .A1(n14990), .A2(n14989), .B1(n14988), .B2(n14987), .C1(
        n14986), .C2(n14985), .ZN(P1_U2893) );
  NAND2_X1 U18546 ( .A1(n12232), .A2(n15172), .ZN(n14994) );
  NAND2_X1 U18547 ( .A1(n12230), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14992) );
  OAI22_X1 U18548 ( .A1(n14991), .A2(n14994), .B1(n14993), .B2(n14992), .ZN(
        n14995) );
  XNOR2_X1 U18549 ( .A(n14995), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15168) );
  INV_X1 U18550 ( .A(n14996), .ZN(n15001) );
  INV_X1 U18551 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14997) );
  NOR2_X1 U18552 ( .A1(n12460), .A2(n14997), .ZN(n15165) );
  AOI21_X1 U18553 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15165), .ZN(n14998) );
  OAI21_X1 U18554 ( .B1(n20482), .B2(n14999), .A(n14998), .ZN(n15000) );
  OAI21_X1 U18555 ( .B1(n15168), .B2(n20321), .A(n15002), .ZN(P1_U2969) );
  XNOR2_X1 U18556 ( .A(n15063), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15003) );
  XNOR2_X1 U18557 ( .A(n15004), .B(n15003), .ZN(n15178) );
  INV_X1 U18558 ( .A(n15005), .ZN(n15008) );
  NOR2_X1 U18559 ( .A1(n12460), .A2(n15006), .ZN(n15170) );
  AOI21_X1 U18560 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15170), .ZN(n15007) );
  OAI21_X1 U18561 ( .B1(n20482), .B2(n15008), .A(n15007), .ZN(n15009) );
  AOI21_X1 U18562 ( .B1(n15010), .B2(n20477), .A(n15009), .ZN(n15011) );
  OAI21_X1 U18563 ( .B1(n15178), .B2(n20321), .A(n15011), .ZN(P1_U2970) );
  INV_X1 U18564 ( .A(n15014), .ZN(n15013) );
  INV_X1 U18565 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15197) );
  INV_X1 U18566 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15190) );
  NAND4_X1 U18567 ( .A1(n15013), .A2(n15035), .A3(n15197), .A4(n15190), .ZN(
        n15016) );
  NAND3_X1 U18568 ( .A1(n15014), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15015) );
  MUX2_X1 U18569 ( .A(n15016), .B(n15015), .S(n12230), .Z(n15017) );
  XNOR2_X1 U18570 ( .A(n15017), .B(n21118), .ZN(n15185) );
  INV_X1 U18571 ( .A(n15018), .ZN(n15022) );
  NOR2_X1 U18572 ( .A1(n12460), .A2(n21035), .ZN(n15180) );
  AOI21_X1 U18573 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15180), .ZN(n15019) );
  OAI21_X1 U18574 ( .B1(n20482), .B2(n15020), .A(n15019), .ZN(n15021) );
  AOI21_X1 U18575 ( .B1(n15022), .B2(n20477), .A(n15021), .ZN(n15023) );
  OAI21_X1 U18576 ( .B1(n15185), .B2(n20321), .A(n15023), .ZN(P1_U2971) );
  XNOR2_X1 U18577 ( .A(n15025), .B(n15190), .ZN(n15196) );
  INV_X1 U18578 ( .A(n15026), .ZN(n15029) );
  INV_X1 U18579 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15027) );
  NOR2_X1 U18580 ( .A1(n12460), .A2(n15027), .ZN(n15188) );
  AOI21_X1 U18581 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15188), .ZN(n15028) );
  OAI21_X1 U18582 ( .B1(n20482), .B2(n15029), .A(n15028), .ZN(n15030) );
  AOI21_X1 U18583 ( .B1(n15031), .B2(n20477), .A(n15030), .ZN(n15032) );
  OAI21_X1 U18584 ( .B1(n15196), .B2(n20321), .A(n15032), .ZN(P1_U2972) );
  NOR2_X1 U18585 ( .A1(n15065), .A2(n12230), .ZN(n15047) );
  NOR2_X1 U18586 ( .A1(n12232), .A2(n15198), .ZN(n15034) );
  AOI22_X1 U18587 ( .A1(n15047), .A2(n15035), .B1(n15034), .B2(n15044), .ZN(
        n15036) );
  XNOR2_X1 U18588 ( .A(n15036), .B(n15197), .ZN(n15205) );
  INV_X1 U18589 ( .A(n15037), .ZN(n15041) );
  INV_X1 U18590 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21032) );
  NOR2_X1 U18591 ( .A1(n12460), .A2(n21032), .ZN(n15201) );
  AOI21_X1 U18592 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15201), .ZN(n15038) );
  OAI21_X1 U18593 ( .B1(n20482), .B2(n15039), .A(n15038), .ZN(n15040) );
  AOI21_X1 U18594 ( .B1(n15041), .B2(n20477), .A(n15040), .ZN(n15042) );
  OAI21_X1 U18595 ( .B1(n15205), .B2(n20321), .A(n15042), .ZN(P1_U2973) );
  INV_X1 U18596 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15234) );
  INV_X1 U18597 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15043) );
  NOR3_X1 U18598 ( .A1(n12232), .A2(n15234), .A3(n15043), .ZN(n15045) );
  AOI22_X1 U18599 ( .A1(n15047), .A2(n15046), .B1(n15045), .B2(n15044), .ZN(
        n15048) );
  XNOR2_X1 U18600 ( .A(n15048), .B(n15209), .ZN(n15216) );
  NOR2_X1 U18601 ( .A1(n12460), .A2(n15049), .ZN(n15207) );
  AOI21_X1 U18602 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15207), .ZN(n15050) );
  OAI21_X1 U18603 ( .B1(n20482), .B2(n15051), .A(n15050), .ZN(n15052) );
  AOI21_X1 U18604 ( .B1(n15053), .B2(n20477), .A(n15052), .ZN(n15054) );
  OAI21_X1 U18605 ( .B1(n15216), .B2(n20321), .A(n15054), .ZN(P1_U2974) );
  AOI21_X1 U18606 ( .B1(n12232), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15065), .ZN(n15055) );
  AOI21_X1 U18607 ( .B1(n12230), .B2(n15234), .A(n15055), .ZN(n15057) );
  XNOR2_X1 U18608 ( .A(n15063), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15056) );
  XNOR2_X1 U18609 ( .A(n15057), .B(n15056), .ZN(n15226) );
  NOR2_X1 U18610 ( .A1(n12460), .A2(n21028), .ZN(n15223) );
  AOI21_X1 U18611 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15223), .ZN(n15058) );
  OAI21_X1 U18612 ( .B1(n20482), .B2(n15059), .A(n15058), .ZN(n15060) );
  AOI21_X1 U18613 ( .B1(n15061), .B2(n20477), .A(n15060), .ZN(n15062) );
  OAI21_X1 U18614 ( .B1(n15226), .B2(n20321), .A(n15062), .ZN(P1_U2975) );
  XNOR2_X1 U18615 ( .A(n15063), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15064) );
  XNOR2_X1 U18616 ( .A(n15065), .B(n15064), .ZN(n15231) );
  INV_X1 U18617 ( .A(n15066), .ZN(n15069) );
  NOR2_X1 U18618 ( .A1(n12460), .A2(n15067), .ZN(n15227) );
  AOI21_X1 U18619 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15227), .ZN(n15068) );
  OAI21_X1 U18620 ( .B1(n20482), .B2(n15069), .A(n15068), .ZN(n15070) );
  AOI21_X1 U18621 ( .B1(n15071), .B2(n20477), .A(n15070), .ZN(n15072) );
  OAI21_X1 U18622 ( .B1(n15231), .B2(n20321), .A(n15072), .ZN(P1_U2976) );
  NAND2_X1 U18623 ( .A1(n15074), .A2(n15073), .ZN(n15075) );
  XOR2_X1 U18624 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15075), .Z(
        n15251) );
  INV_X1 U18625 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15076) );
  NOR2_X1 U18626 ( .A1(n12460), .A2(n15076), .ZN(n15237) );
  AOI21_X1 U18627 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15237), .ZN(n15077) );
  OAI21_X1 U18628 ( .B1(n20482), .B2(n16211), .A(n15077), .ZN(n15078) );
  AOI21_X1 U18629 ( .B1(n16216), .B2(n20477), .A(n15078), .ZN(n15079) );
  OAI21_X1 U18630 ( .B1(n15251), .B2(n20321), .A(n15079), .ZN(P1_U2977) );
  NAND2_X1 U18631 ( .A1(n15080), .A2(n12230), .ZN(n15088) );
  NAND2_X1 U18632 ( .A1(n15081), .A2(n12232), .ZN(n15089) );
  MUX2_X1 U18633 ( .A(n15088), .B(n15089), .S(n15244), .Z(n15082) );
  XNOR2_X1 U18634 ( .A(n15082), .B(n15256), .ZN(n15260) );
  INV_X1 U18635 ( .A(n16221), .ZN(n15085) );
  INV_X1 U18636 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15083) );
  NOR2_X1 U18637 ( .A1(n12460), .A2(n15083), .ZN(n15252) );
  AOI21_X1 U18638 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15252), .ZN(n15084) );
  OAI21_X1 U18639 ( .B1(n20482), .B2(n15085), .A(n15084), .ZN(n15086) );
  AOI21_X1 U18640 ( .B1(n16224), .B2(n20477), .A(n15086), .ZN(n15087) );
  OAI21_X1 U18641 ( .B1(n15260), .B2(n20321), .A(n15087), .ZN(P1_U2978) );
  NAND2_X1 U18642 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  XNOR2_X1 U18643 ( .A(n15090), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15269) );
  NOR2_X1 U18644 ( .A1(n12460), .A2(n21022), .ZN(n15262) );
  AOI21_X1 U18645 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15262), .ZN(n15091) );
  OAI21_X1 U18646 ( .B1(n20482), .B2(n15092), .A(n15091), .ZN(n15093) );
  AOI21_X1 U18647 ( .B1(n15094), .B2(n20477), .A(n15093), .ZN(n15095) );
  OAI21_X1 U18648 ( .B1(n15269), .B2(n20321), .A(n15095), .ZN(P1_U2979) );
  NAND2_X1 U18650 ( .A1(n15106), .A2(n15280), .ZN(n15097) );
  MUX2_X1 U18651 ( .A(n15106), .B(n15097), .S(n21407), .Z(n15098) );
  XNOR2_X1 U18652 ( .A(n15098), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15270) );
  INV_X1 U18653 ( .A(n15270), .ZN(n15104) );
  INV_X1 U18654 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15099) );
  NOR2_X1 U18655 ( .A1(n12460), .A2(n15099), .ZN(n15274) );
  AOI21_X1 U18656 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15274), .ZN(n15100) );
  OAI21_X1 U18657 ( .B1(n20482), .B2(n15101), .A(n15100), .ZN(n15102) );
  AOI21_X1 U18658 ( .B1(n16236), .B2(n20477), .A(n15102), .ZN(n15103) );
  OAI21_X1 U18659 ( .B1(n15104), .B2(n20321), .A(n15103), .ZN(P1_U2980) );
  OAI21_X1 U18660 ( .B1(n15105), .B2(n15107), .A(n15106), .ZN(n15290) );
  INV_X1 U18661 ( .A(n15108), .ZN(n16248) );
  INV_X1 U18662 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n16238) );
  NOR2_X1 U18663 ( .A1(n12460), .A2(n16238), .ZN(n15285) );
  AOI21_X1 U18664 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15285), .ZN(n15109) );
  OAI21_X1 U18665 ( .B1(n20482), .B2(n16245), .A(n15109), .ZN(n15110) );
  AOI21_X1 U18666 ( .B1(n16248), .B2(n20477), .A(n15110), .ZN(n15111) );
  OAI21_X1 U18667 ( .B1(n15290), .B2(n20321), .A(n15111), .ZN(P1_U2981) );
  OAI21_X1 U18668 ( .B1(n16348), .B2(n9820), .A(n15113), .ZN(n15117) );
  NAND2_X1 U18669 ( .A1(n15117), .A2(n15114), .ZN(n15116) );
  MUX2_X1 U18670 ( .A(n15117), .B(n15116), .S(n21407), .Z(n15118) );
  XNOR2_X1 U18671 ( .A(n15118), .B(n15292), .ZN(n15298) );
  INV_X1 U18672 ( .A(n15119), .ZN(n16255) );
  INV_X1 U18673 ( .A(n16251), .ZN(n15121) );
  NOR2_X1 U18674 ( .A1(n12460), .A2(n21018), .ZN(n15294) );
  AOI21_X1 U18675 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15294), .ZN(n15120) );
  OAI21_X1 U18676 ( .B1(n20482), .B2(n15121), .A(n15120), .ZN(n15122) );
  AOI21_X1 U18677 ( .B1(n16255), .B2(n20477), .A(n15122), .ZN(n15123) );
  OAI21_X1 U18678 ( .B1(n15298), .B2(n20321), .A(n15123), .ZN(P1_U2982) );
  INV_X1 U18679 ( .A(n15124), .ZN(n15125) );
  AOI21_X1 U18680 ( .B1(n16348), .B2(n15126), .A(n15125), .ZN(n16339) );
  AND2_X1 U18681 ( .A1(n15127), .A2(n15128), .ZN(n16338) );
  NAND2_X1 U18682 ( .A1(n16339), .A2(n16338), .ZN(n16337) );
  NAND2_X1 U18683 ( .A1(n16337), .A2(n15128), .ZN(n15129) );
  XOR2_X1 U18684 ( .A(n15130), .B(n15129), .Z(n16406) );
  NAND2_X1 U18685 ( .A1(n16406), .A2(n12479), .ZN(n15135) );
  INV_X1 U18686 ( .A(n20482), .ZN(n16342) );
  INV_X1 U18687 ( .A(n16287), .ZN(n15133) );
  OAI22_X1 U18688 ( .A1(n15131), .A2(n16285), .B1(n12460), .B2(n21387), .ZN(
        n15132) );
  AOI21_X1 U18689 ( .B1(n16342), .B2(n15133), .A(n15132), .ZN(n15134) );
  OAI211_X1 U18690 ( .C1(n15136), .C2(n16288), .A(n15135), .B(n15134), .ZN(
        P1_U2986) );
  MUX2_X1 U18691 ( .A(n16347), .B(n16348), .S(n12230), .Z(n15137) );
  XNOR2_X1 U18692 ( .A(n15137), .B(n16346), .ZN(n16444) );
  INV_X1 U18693 ( .A(n16444), .ZN(n15143) );
  AOI22_X1 U18694 ( .A1(n20474), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15138) );
  OAI21_X1 U18695 ( .B1(n20482), .B2(n15139), .A(n15138), .ZN(n15140) );
  AOI21_X1 U18696 ( .B1(n15141), .B2(n20477), .A(n15140), .ZN(n15142) );
  OAI21_X1 U18697 ( .B1(n15143), .B2(n20321), .A(n15142), .ZN(P1_U2989) );
  INV_X1 U18698 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16453) );
  MUX2_X1 U18699 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n16453), .S(
        n12230), .Z(n15145) );
  XNOR2_X1 U18700 ( .A(n15144), .B(n15145), .ZN(n16450) );
  INV_X1 U18701 ( .A(n16450), .ZN(n15150) );
  AOI22_X1 U18702 ( .A1(n20474), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n15146) );
  OAI21_X1 U18703 ( .B1(n20482), .B2(n15147), .A(n15146), .ZN(n15148) );
  AOI21_X1 U18704 ( .B1(n20348), .B2(n20477), .A(n15148), .ZN(n15149) );
  OAI21_X1 U18705 ( .B1(n15150), .B2(n20321), .A(n15149), .ZN(P1_U2990) );
  XNOR2_X1 U18706 ( .A(n15151), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15152) );
  XNOR2_X1 U18707 ( .A(n15153), .B(n15152), .ZN(n15307) );
  INV_X1 U18708 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15154) );
  NOR2_X1 U18709 ( .A1(n12460), .A2(n15154), .ZN(n15304) );
  AOI21_X1 U18710 ( .B1(n20474), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15304), .ZN(n15155) );
  OAI21_X1 U18711 ( .B1(n20482), .B2(n15156), .A(n15155), .ZN(n15157) );
  AOI21_X1 U18712 ( .B1(n15158), .B2(n20477), .A(n15157), .ZN(n15159) );
  OAI21_X1 U18713 ( .B1(n15307), .B2(n20321), .A(n15159), .ZN(P1_U2991) );
  INV_X1 U18714 ( .A(n15160), .ZN(n15173) );
  AOI21_X1 U18715 ( .B1(n15173), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15163) );
  INV_X1 U18716 ( .A(n15161), .ZN(n15162) );
  NOR2_X1 U18717 ( .A1(n15163), .A2(n15162), .ZN(n15164) );
  OAI21_X1 U18718 ( .B1(n15168), .B2(n16424), .A(n15167), .ZN(P1_U3001) );
  NOR2_X1 U18719 ( .A1(n15169), .A2(n15172), .ZN(n15171) );
  AOI211_X1 U18720 ( .C1(n15173), .C2(n15172), .A(n15171), .B(n15170), .ZN(
        n15177) );
  INV_X1 U18721 ( .A(n15174), .ZN(n15175) );
  NAND2_X1 U18722 ( .A1(n15175), .A2(n20486), .ZN(n15176) );
  OAI211_X1 U18723 ( .C1(n15178), .C2(n16424), .A(n15177), .B(n15176), .ZN(
        P1_U3002) );
  XNOR2_X1 U18724 ( .A(n21118), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15181) );
  INV_X1 U18725 ( .A(n15203), .ZN(n15187) );
  INV_X1 U18726 ( .A(n16436), .ZN(n15186) );
  NOR3_X1 U18727 ( .A1(n15187), .A2(n15186), .A3(n21118), .ZN(n15179) );
  AOI211_X1 U18728 ( .C1(n15191), .C2(n15181), .A(n15180), .B(n15179), .ZN(
        n15184) );
  NAND2_X1 U18729 ( .A1(n15182), .A2(n20486), .ZN(n15183) );
  OAI211_X1 U18730 ( .C1(n15185), .C2(n16424), .A(n15184), .B(n15183), .ZN(
        P1_U3003) );
  NOR3_X1 U18731 ( .A1(n15187), .A2(n15186), .A3(n15190), .ZN(n15189) );
  AOI211_X1 U18732 ( .C1(n15191), .C2(n15190), .A(n15189), .B(n15188), .ZN(
        n15195) );
  INV_X1 U18733 ( .A(n15192), .ZN(n15193) );
  NAND2_X1 U18734 ( .A1(n15193), .A2(n20486), .ZN(n15194) );
  OAI211_X1 U18735 ( .C1(n15196), .C2(n16424), .A(n15195), .B(n15194), .ZN(
        P1_U3004) );
  OAI21_X1 U18736 ( .B1(n15221), .B2(n15198), .A(n15197), .ZN(n15202) );
  NOR2_X1 U18737 ( .A1(n15199), .A2(n20504), .ZN(n15200) );
  AOI211_X1 U18738 ( .C1(n15203), .C2(n15202), .A(n15201), .B(n15200), .ZN(
        n15204) );
  OAI21_X1 U18739 ( .B1(n15205), .B2(n16424), .A(n15204), .ZN(P1_U3005) );
  INV_X1 U18740 ( .A(n15206), .ZN(n15208) );
  AOI21_X1 U18741 ( .B1(n15208), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15207), .ZN(n15212) );
  INV_X1 U18742 ( .A(n15221), .ZN(n15235) );
  NAND3_X1 U18743 ( .A1(n15235), .A2(n15210), .A3(n15209), .ZN(n15211) );
  OAI211_X1 U18744 ( .C1(n15213), .C2(n20504), .A(n15212), .B(n15211), .ZN(
        n15214) );
  INV_X1 U18745 ( .A(n15214), .ZN(n15215) );
  OAI21_X1 U18746 ( .B1(n15216), .B2(n16424), .A(n15215), .ZN(P1_U3006) );
  AOI21_X1 U18747 ( .B1(n15217), .B2(n20502), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15218) );
  OAI21_X1 U18748 ( .B1(n15218), .B2(n15228), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15219) );
  OAI21_X1 U18749 ( .B1(n15220), .B2(n20504), .A(n15219), .ZN(n15224) );
  NOR3_X1 U18750 ( .A1(n15221), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15234), .ZN(n15222) );
  NOR3_X1 U18751 ( .A1(n15224), .A2(n15223), .A3(n15222), .ZN(n15225) );
  OAI21_X1 U18752 ( .B1(n15226), .B2(n16424), .A(n15225), .ZN(P1_U3007) );
  AOI21_X1 U18753 ( .B1(n15228), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15227), .ZN(n15229) );
  OAI21_X1 U18754 ( .B1(n15230), .B2(n20504), .A(n15229), .ZN(n15233) );
  NOR2_X1 U18755 ( .A1(n15231), .A2(n16424), .ZN(n15232) );
  AOI211_X1 U18756 ( .C1(n15235), .C2(n15234), .A(n15233), .B(n15232), .ZN(
        n15236) );
  INV_X1 U18757 ( .A(n15236), .ZN(P1_U3008) );
  INV_X1 U18758 ( .A(n16219), .ZN(n15249) );
  INV_X1 U18759 ( .A(n15237), .ZN(n15247) );
  INV_X1 U18760 ( .A(n15238), .ZN(n15239) );
  NAND2_X1 U18761 ( .A1(n15239), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15240) );
  AOI21_X1 U18762 ( .B1(n15243), .B2(n15241), .A(n15240), .ZN(n15276) );
  INV_X1 U18763 ( .A(n16385), .ZN(n15242) );
  NAND3_X1 U18764 ( .A1(n15242), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n16404), .ZN(n16384) );
  AND2_X1 U18765 ( .A1(n15243), .A2(n16384), .ZN(n16400) );
  NAND2_X1 U18766 ( .A1(n16396), .A2(n16400), .ZN(n15261) );
  NAND3_X1 U18767 ( .A1(n15276), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15261), .ZN(n15265) );
  NOR2_X1 U18768 ( .A1(n15265), .A2(n15244), .ZN(n15253) );
  OAI211_X1 U18769 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15253), .B(n15245), .ZN(
        n15246) );
  OAI211_X1 U18770 ( .C1(n15255), .C2(n9933), .A(n15247), .B(n15246), .ZN(
        n15248) );
  AOI21_X1 U18771 ( .B1(n15249), .B2(n20486), .A(n15248), .ZN(n15250) );
  OAI21_X1 U18772 ( .B1(n15251), .B2(n16424), .A(n15250), .ZN(P1_U3009) );
  INV_X1 U18773 ( .A(n16222), .ZN(n15258) );
  AOI21_X1 U18774 ( .B1(n15253), .B2(n15256), .A(n15252), .ZN(n15254) );
  OAI21_X1 U18775 ( .B1(n15256), .B2(n15255), .A(n15254), .ZN(n15257) );
  AOI21_X1 U18776 ( .B1(n15258), .B2(n20486), .A(n15257), .ZN(n15259) );
  OAI21_X1 U18777 ( .B1(n15260), .B2(n16424), .A(n15259), .ZN(P1_U3010) );
  AND2_X1 U18778 ( .A1(n15261), .A2(n21077), .ZN(n15275) );
  OAI21_X1 U18779 ( .B1(n15271), .B2(n15275), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15264) );
  INV_X1 U18780 ( .A(n15262), .ZN(n15263) );
  OAI211_X1 U18781 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15265), .A(
        n15264), .B(n15263), .ZN(n15266) );
  AOI21_X1 U18782 ( .B1(n15267), .B2(n20486), .A(n15266), .ZN(n15268) );
  OAI21_X1 U18783 ( .B1(n15269), .B2(n16424), .A(n15268), .ZN(P1_U3011) );
  NAND2_X1 U18784 ( .A1(n15270), .A2(n20507), .ZN(n15278) );
  INV_X1 U18785 ( .A(n15271), .ZN(n15272) );
  NOR2_X1 U18786 ( .A1(n15272), .A2(n21077), .ZN(n15273) );
  AOI211_X1 U18787 ( .C1(n15276), .C2(n15275), .A(n15274), .B(n15273), .ZN(
        n15277) );
  OAI211_X1 U18788 ( .C1(n20504), .C2(n16242), .A(n15278), .B(n15277), .ZN(
        P1_U3012) );
  NAND4_X1 U18789 ( .A1(n15291), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        n15287) );
  OAI21_X1 U18790 ( .B1(n20495), .B2(n16397), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15282) );
  NAND2_X1 U18791 ( .A1(n15282), .A2(n15300), .ZN(n15283) );
  AND2_X1 U18792 ( .A1(n16386), .A2(n15283), .ZN(n16369) );
  OAI21_X1 U18793 ( .B1(n16368), .B2(n15292), .A(n15300), .ZN(n15284) );
  NAND2_X1 U18794 ( .A1(n16369), .A2(n15284), .ZN(n15295) );
  AOI21_X1 U18795 ( .B1(n15295), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15285), .ZN(n15286) );
  OAI211_X1 U18796 ( .C1(n20504), .C2(n16250), .A(n15287), .B(n15286), .ZN(
        n15288) );
  INV_X1 U18797 ( .A(n15288), .ZN(n15289) );
  OAI21_X1 U18798 ( .B1(n15290), .B2(n16424), .A(n15289), .ZN(P1_U3013) );
  NAND2_X1 U18799 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15291), .ZN(
        n16379) );
  OAI21_X1 U18800 ( .B1(n16368), .B2(n16379), .A(n15292), .ZN(n15296) );
  NOR2_X1 U18801 ( .A1(n16260), .A2(n20504), .ZN(n15293) );
  AOI211_X1 U18802 ( .C1(n15296), .C2(n15295), .A(n15294), .B(n15293), .ZN(
        n15297) );
  OAI21_X1 U18803 ( .B1(n15298), .B2(n16424), .A(n15297), .ZN(P1_U3014) );
  INV_X1 U18804 ( .A(n15299), .ZN(n15305) );
  INV_X1 U18805 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15301) );
  NOR2_X1 U18806 ( .A1(n15301), .A2(n16432), .ZN(n16454) );
  OAI21_X1 U18807 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16454), .ZN(n15302) );
  AOI21_X1 U18808 ( .B1(n15301), .B2(n15300), .A(n16463), .ZN(n16459) );
  OAI22_X1 U18809 ( .A1(n16439), .A2(n15302), .B1(n16459), .B2(n12358), .ZN(
        n15303) );
  AOI211_X1 U18810 ( .C1(n20486), .C2(n15305), .A(n15304), .B(n15303), .ZN(
        n15306) );
  OAI21_X1 U18811 ( .B1(n15307), .B2(n16424), .A(n15306), .ZN(P1_U3023) );
  NOR2_X1 U18812 ( .A1(n20650), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15308) );
  OAI22_X1 U18813 ( .A1(n20613), .A2(n15308), .B1(n14172), .B2(n15316), .ZN(
        n15309) );
  MUX2_X1 U18814 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15309), .S(
        n20513), .Z(P1_U3477) );
  MUX2_X1 U18815 ( .A(n15310), .B(n20613), .S(n20652), .Z(n15311) );
  OAI21_X1 U18816 ( .B1(n15316), .B2(n9748), .A(n15311), .ZN(n15312) );
  MUX2_X1 U18817 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15312), .S(
        n20513), .Z(P1_U3476) );
  OAI21_X1 U18818 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20515), .A(n20784), 
        .ZN(n15314) );
  OR2_X1 U18819 ( .A1(n20650), .A2(n20683), .ZN(n20779) );
  NOR2_X1 U18820 ( .A1(n15313), .A2(n20779), .ZN(n20909) );
  AOI211_X1 U18821 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n15315), .A(n15314), 
        .B(n20909), .ZN(n15318) );
  INV_X1 U18822 ( .A(n9749), .ZN(n15317) );
  OAI22_X1 U18823 ( .A1(n15318), .A2(n20915), .B1(n15317), .B2(n15316), .ZN(
        n15319) );
  MUX2_X1 U18824 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15319), .S(
        n20513), .Z(P1_U3475) );
  INV_X1 U18825 ( .A(n15320), .ZN(n15323) );
  INV_X1 U18826 ( .A(n15321), .ZN(n15322) );
  NAND2_X1 U18827 ( .A1(n15323), .A2(n15322), .ZN(n15324) );
  NAND2_X1 U18828 ( .A1(n15325), .A2(n15324), .ZN(n15786) );
  AOI21_X1 U18829 ( .B1(n10061), .B2(n10253), .A(n19450), .ZN(n15334) );
  INV_X1 U18830 ( .A(n16493), .ZN(n15333) );
  NOR2_X1 U18831 ( .A1(n9777), .A2(n15326), .ZN(n15327) );
  AOI22_X1 U18832 ( .A1(n15329), .A2(n19422), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n19431), .ZN(n15331) );
  AOI22_X1 U18833 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19444), .ZN(n15330) );
  OAI211_X1 U18834 ( .C1(n15791), .C2(n19442), .A(n15331), .B(n15330), .ZN(
        n15332) );
  OAI21_X1 U18835 ( .B1(n15786), .B2(n19414), .A(n15335), .ZN(P2_U2826) );
  INV_X1 U18836 ( .A(n15336), .ZN(n15339) );
  NAND2_X1 U18837 ( .A1(n15416), .A2(n15337), .ZN(n15338) );
  NAND2_X1 U18838 ( .A1(n15339), .A2(n15338), .ZN(n15805) );
  NAND2_X1 U18839 ( .A1(n15340), .A2(n15341), .ZN(n15342) );
  NAND2_X1 U18840 ( .A1(n15343), .A2(n15342), .ZN(n15802) );
  AOI22_X1 U18841 ( .A1(n15344), .A2(n19422), .B1(P2_REIP_REG_27__SCAN_IN), 
        .B2(n19431), .ZN(n15346) );
  AOI22_X1 U18842 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19444), .ZN(n15345) );
  OAI211_X1 U18843 ( .C1(n15802), .C2(n19442), .A(n15346), .B(n15345), .ZN(
        n15350) );
  AOI211_X1 U18844 ( .C1(n15616), .C2(n15348), .A(n15347), .B(n19450), .ZN(
        n15349) );
  NOR2_X1 U18845 ( .A1(n15350), .A2(n15349), .ZN(n15351) );
  OAI21_X1 U18846 ( .B1(n19414), .B2(n15805), .A(n15351), .ZN(P2_U2828) );
  NAND2_X1 U18847 ( .A1(n15447), .A2(n15352), .ZN(n15353) );
  NAND2_X1 U18848 ( .A1(n9782), .A2(n15353), .ZN(n16561) );
  XNOR2_X1 U18849 ( .A(n15354), .B(n15859), .ZN(n15849) );
  AOI22_X1 U18850 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19431), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19454), .ZN(n15357) );
  AOI22_X1 U18851 ( .A1(n15355), .A2(n19422), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n19444), .ZN(n15356) );
  OAI211_X1 U18852 ( .C1(n15849), .C2(n19442), .A(n15357), .B(n15356), .ZN(
        n15360) );
  AOI211_X1 U18853 ( .C1(n16558), .C2(n10044), .A(n15358), .B(n19450), .ZN(
        n15359) );
  NOR2_X1 U18854 ( .A1(n15360), .A2(n15359), .ZN(n15361) );
  OAI21_X1 U18855 ( .B1(n19414), .B2(n16561), .A(n15361), .ZN(P2_U2832) );
  AOI211_X1 U18856 ( .C1(n15364), .C2(n15363), .A(n15362), .B(n19450), .ZN(
        n15365) );
  INV_X1 U18857 ( .A(n15365), .ZN(n15371) );
  XNOR2_X1 U18858 ( .A(n15565), .B(n9845), .ZN(n15907) );
  INV_X1 U18859 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20229) );
  AOI22_X1 U18860 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19444), .ZN(n15366) );
  OAI211_X1 U18861 ( .C1(n19440), .C2(n20229), .A(n15366), .B(n19272), .ZN(
        n15369) );
  OAI21_X1 U18862 ( .B1(n15474), .B2(n15367), .A(n15463), .ZN(n15904) );
  NOR2_X1 U18863 ( .A1(n15904), .A2(n19414), .ZN(n15368) );
  AOI211_X1 U18864 ( .C1(n19379), .C2(n15907), .A(n15369), .B(n15368), .ZN(
        n15370) );
  OAI211_X1 U18865 ( .C1(n15372), .C2(n19447), .A(n15371), .B(n15370), .ZN(
        P2_U2836) );
  NAND2_X1 U18866 ( .A1(n10049), .A2(n15373), .ZN(n19345) );
  INV_X1 U18867 ( .A(n19345), .ZN(n15374) );
  OAI211_X1 U18868 ( .C1(n15376), .C2(n15375), .A(n19416), .B(n15374), .ZN(
        n15385) );
  NOR2_X1 U18869 ( .A1(n19450), .A2(n10049), .ZN(n19285) );
  AOI22_X1 U18870 ( .A1(n16606), .A2(n19285), .B1(n19444), .B2(
        P2_EBX_REG_11__SCAN_IN), .ZN(n15377) );
  OAI21_X1 U18871 ( .B1(n16614), .B2(n19414), .A(n15377), .ZN(n15382) );
  OAI21_X1 U18872 ( .B1(n15379), .B2(n15378), .A(n15936), .ZN(n19477) );
  AOI22_X1 U18873 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19454), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19431), .ZN(n15380) );
  OAI211_X1 U18874 ( .C1(n19477), .C2(n19442), .A(n15380), .B(n19272), .ZN(
        n15381) );
  AOI211_X1 U18875 ( .C1(n19422), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        n15384) );
  NAND2_X1 U18876 ( .A1(n15385), .A2(n15384), .ZN(P2_U2844) );
  OAI211_X1 U18877 ( .C1(n16006), .C2(n15387), .A(n10049), .B(n15386), .ZN(
        n16013) );
  XNOR2_X1 U18878 ( .A(n15389), .B(n15388), .ZN(n20286) );
  INV_X1 U18879 ( .A(n15390), .ZN(n15392) );
  AOI22_X1 U18880 ( .A1(n19431), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n13043), 
        .B2(n19285), .ZN(n15391) );
  OAI21_X1 U18881 ( .B1(n19447), .B2(n15392), .A(n15391), .ZN(n15394) );
  OAI22_X1 U18882 ( .A1(n19429), .A2(n11396), .B1(n13043), .B2(n19420), .ZN(
        n15393) );
  AOI211_X1 U18883 ( .C1(n19379), .C2(n20286), .A(n15394), .B(n15393), .ZN(
        n15395) );
  OAI21_X1 U18884 ( .B1(n15396), .B2(n19414), .A(n15395), .ZN(n15397) );
  AOI21_X1 U18885 ( .B1(n20284), .B2(n19452), .A(n15397), .ZN(n15398) );
  OAI21_X1 U18886 ( .B1(n16013), .B2(n19450), .A(n15398), .ZN(P2_U2854) );
  INV_X1 U18887 ( .A(n16489), .ZN(n15399) );
  NAND2_X1 U18888 ( .A1(n15399), .A2(n15499), .ZN(n15400) );
  OAI21_X1 U18889 ( .B1(n15499), .B2(n13074), .A(n15400), .ZN(P2_U2856) );
  OR2_X1 U18890 ( .A1(n15402), .A2(n15401), .ZN(n15505) );
  NAND3_X1 U18891 ( .A1(n15505), .A2(n15403), .A3(n15492), .ZN(n15405) );
  NAND2_X1 U18892 ( .A1(n15480), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15404) );
  OAI211_X1 U18893 ( .C1(n15786), .C2(n15480), .A(n15405), .B(n15404), .ZN(
        P2_U2858) );
  NAND2_X1 U18894 ( .A1(n13407), .A2(n15406), .ZN(n15408) );
  XNOR2_X1 U18895 ( .A(n15408), .B(n15407), .ZN(n15511) );
  NAND2_X1 U18896 ( .A1(n15511), .A2(n15492), .ZN(n15410) );
  NAND2_X1 U18897 ( .A1(n15480), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15409) );
  OAI211_X1 U18898 ( .C1(n16496), .C2(n15480), .A(n15410), .B(n15409), .ZN(
        P2_U2859) );
  AOI21_X1 U18899 ( .B1(n15412), .B2(n15411), .A(n9791), .ZN(n15520) );
  NAND2_X1 U18900 ( .A1(n15520), .A2(n15492), .ZN(n15414) );
  NAND2_X1 U18901 ( .A1(n15480), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15413) );
  OAI211_X1 U18902 ( .C1(n15480), .C2(n15805), .A(n15414), .B(n15413), .ZN(
        P2_U2860) );
  OAI21_X1 U18903 ( .B1(n10128), .B2(n10130), .A(n15416), .ZN(n16510) );
  AOI21_X1 U18904 ( .B1(n15419), .B2(n15418), .A(n15417), .ZN(n15527) );
  NAND2_X1 U18905 ( .A1(n15527), .A2(n15492), .ZN(n15421) );
  NAND2_X1 U18906 ( .A1(n15480), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15420) );
  OAI211_X1 U18907 ( .C1(n16510), .C2(n15480), .A(n15421), .B(n15420), .ZN(
        P2_U2861) );
  OAI21_X1 U18908 ( .B1(n15424), .B2(n15423), .A(n15422), .ZN(n15534) );
  OAI21_X1 U18909 ( .B1(n15433), .B2(n15426), .A(n15425), .ZN(n16524) );
  NOR2_X1 U18910 ( .A1(n16524), .A2(n15480), .ZN(n15427) );
  AOI21_X1 U18911 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n13461), .A(n15427), .ZN(
        n15428) );
  OAI21_X1 U18912 ( .B1(n15534), .B2(n15482), .A(n15428), .ZN(P2_U2862) );
  AOI21_X1 U18913 ( .B1(n15429), .B2(n15430), .A(n9824), .ZN(n15431) );
  XOR2_X1 U18914 ( .A(n15432), .B(n15431), .Z(n15542) );
  INV_X1 U18915 ( .A(n15433), .ZN(n15436) );
  NAND2_X1 U18916 ( .A1(n9782), .A2(n15434), .ZN(n15435) );
  NAND2_X1 U18917 ( .A1(n15436), .A2(n15435), .ZN(n16542) );
  NOR2_X1 U18918 ( .A1(n16542), .A2(n15480), .ZN(n15437) );
  AOI21_X1 U18919 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n13461), .A(n15437), .ZN(
        n15438) );
  OAI21_X1 U18920 ( .B1(n15542), .B2(n15482), .A(n15438), .ZN(P2_U2863) );
  AOI21_X1 U18921 ( .B1(n15439), .B2(n15441), .A(n15440), .ZN(n15442) );
  INV_X1 U18922 ( .A(n15442), .ZN(n15548) );
  NOR2_X1 U18923 ( .A1(n16561), .A2(n15480), .ZN(n15443) );
  AOI21_X1 U18924 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n13461), .A(n15443), .ZN(
        n15444) );
  OAI21_X1 U18925 ( .B1(n15548), .B2(n15482), .A(n15444), .ZN(P2_U2864) );
  INV_X1 U18926 ( .A(n15445), .ZN(n15449) );
  INV_X1 U18927 ( .A(n15446), .ZN(n15448) );
  OAI21_X1 U18928 ( .B1(n15449), .B2(n15448), .A(n15447), .ZN(n16131) );
  AOI21_X1 U18929 ( .B1(n15452), .B2(n15450), .A(n15451), .ZN(n16548) );
  NAND2_X1 U18930 ( .A1(n16548), .A2(n15492), .ZN(n15454) );
  NAND2_X1 U18931 ( .A1(n15480), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15453) );
  OAI211_X1 U18932 ( .C1(n16131), .C2(n15480), .A(n15454), .B(n15453), .ZN(
        P2_U2865) );
  INV_X1 U18933 ( .A(n15450), .ZN(n15456) );
  AOI21_X1 U18934 ( .B1(n15457), .B2(n15455), .A(n15456), .ZN(n15549) );
  NAND2_X1 U18935 ( .A1(n15549), .A2(n15492), .ZN(n15459) );
  INV_X1 U18936 ( .A(n15678), .ZN(n15874) );
  NAND2_X1 U18937 ( .A1(n15874), .A2(n15499), .ZN(n15458) );
  OAI211_X1 U18938 ( .C1(n15499), .C2(n11494), .A(n15459), .B(n15458), .ZN(
        P2_U2866) );
  OAI21_X1 U18939 ( .B1(n15461), .B2(n15462), .A(n15455), .ZN(n16553) );
  AOI21_X1 U18940 ( .B1(n15464), .B2(n15463), .A(n9806), .ZN(n19260) );
  INV_X1 U18941 ( .A(n19260), .ZN(n15898) );
  MUX2_X1 U18942 ( .A(n11333), .B(n15898), .S(n15499), .Z(n15465) );
  OAI21_X1 U18943 ( .B1(n16553), .B2(n15482), .A(n15465), .ZN(P2_U2867) );
  INV_X1 U18944 ( .A(n15461), .ZN(n15468) );
  OAI21_X1 U18945 ( .B1(n15472), .B2(n15469), .A(n15468), .ZN(n15555) );
  NOR2_X1 U18946 ( .A1(n15904), .A2(n15480), .ZN(n15470) );
  AOI21_X1 U18947 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n13461), .A(n15470), .ZN(
        n15471) );
  OAI21_X1 U18948 ( .B1(n15555), .B2(n15482), .A(n15471), .ZN(P2_U2868) );
  OAI21_X1 U18949 ( .B1(n9755), .B2(n15473), .A(n15467), .ZN(n15571) );
  INV_X1 U18950 ( .A(n15474), .ZN(n15479) );
  INV_X1 U18951 ( .A(n15485), .ZN(n15477) );
  INV_X1 U18952 ( .A(n15475), .ZN(n15476) );
  NAND2_X1 U18953 ( .A1(n15477), .A2(n15476), .ZN(n15478) );
  NAND2_X1 U18954 ( .A1(n15479), .A2(n15478), .ZN(n19275) );
  MUX2_X1 U18955 ( .A(n19275), .B(n11485), .S(n15480), .Z(n15481) );
  OAI21_X1 U18956 ( .B1(n15571), .B2(n15482), .A(n15481), .ZN(P2_U2869) );
  NOR2_X1 U18957 ( .A1(n15483), .A2(n15493), .ZN(n15484) );
  NOR2_X1 U18958 ( .A1(n15485), .A2(n15484), .ZN(n19290) );
  INV_X1 U18959 ( .A(n19290), .ZN(n16142) );
  AOI21_X1 U18960 ( .B1(n15487), .B2(n10238), .A(n9755), .ZN(n15578) );
  NAND2_X1 U18961 ( .A1(n15578), .A2(n15492), .ZN(n15489) );
  NAND2_X1 U18962 ( .A1(n15480), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15488) );
  OAI211_X1 U18963 ( .C1(n16142), .C2(n15480), .A(n15489), .B(n15488), .ZN(
        P2_U2870) );
  INV_X1 U18964 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15498) );
  AOI21_X1 U18965 ( .B1(n15491), .B2(n15490), .A(n15486), .ZN(n19463) );
  NAND2_X1 U18966 ( .A1(n19463), .A2(n15492), .ZN(n15497) );
  AOI21_X1 U18967 ( .B1(n15495), .B2(n15494), .A(n15493), .ZN(n19303) );
  NAND2_X1 U18968 ( .A1(n15499), .A2(n19303), .ZN(n15496) );
  OAI211_X1 U18969 ( .C1(n15499), .C2(n15498), .A(n15497), .B(n15496), .ZN(
        P2_U2871) );
  INV_X1 U18970 ( .A(n19461), .ZN(n15504) );
  INV_X1 U18971 ( .A(n15500), .ZN(n15501) );
  AOI22_X1 U18972 ( .A1(n15501), .A2(n19523), .B1(P2_EAX_REG_31__SCAN_IN), 
        .B2(n19522), .ZN(n15503) );
  NAND2_X1 U18973 ( .A1(n19460), .A2(BUF2_REG_31__SCAN_IN), .ZN(n15502) );
  OAI211_X1 U18974 ( .C1(n16811), .C2(n15504), .A(n15503), .B(n15502), .ZN(
        P2_U2888) );
  NAND3_X1 U18975 ( .A1(n15505), .A2(n15403), .A3(n19505), .ZN(n15510) );
  INV_X1 U18976 ( .A(n15791), .ZN(n15507) );
  INV_X1 U18977 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19544) );
  OAI22_X1 U18978 ( .A1(n15543), .A2(n19472), .B1(n19489), .B2(n19544), .ZN(
        n15506) );
  AOI21_X1 U18979 ( .B1(n19523), .B2(n15507), .A(n15506), .ZN(n15509) );
  AOI22_X1 U18980 ( .A1(n19461), .A2(BUF1_REG_29__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15508) );
  NAND3_X1 U18981 ( .A1(n15510), .A2(n15509), .A3(n15508), .ZN(P2_U2890) );
  INV_X1 U18982 ( .A(n15511), .ZN(n15515) );
  OAI22_X1 U18983 ( .A1(n15543), .A2(n19474), .B1(n19489), .B2(n19546), .ZN(
        n15512) );
  AOI21_X1 U18984 ( .B1(n19523), .B2(n16497), .A(n15512), .ZN(n15514) );
  AOI22_X1 U18985 ( .A1(n19461), .A2(BUF1_REG_28__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15513) );
  OAI211_X1 U18986 ( .C1(n15515), .C2(n19527), .A(n15514), .B(n15513), .ZN(
        P2_U2891) );
  AOI22_X1 U18987 ( .A1(n19461), .A2(BUF1_REG_27__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U18988 ( .A1(n19459), .A2(n15516), .B1(n19522), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15517) );
  OAI211_X1 U18989 ( .C1(n15576), .C2(n15802), .A(n15518), .B(n15517), .ZN(
        n15519) );
  AOI21_X1 U18990 ( .B1(n15520), .B2(n19505), .A(n15519), .ZN(n15521) );
  INV_X1 U18991 ( .A(n15521), .ZN(P2_U2892) );
  OAI21_X1 U18992 ( .B1(n15523), .B2(n15522), .A(n15340), .ZN(n15811) );
  AOI22_X1 U18993 ( .A1(n19461), .A2(BUF1_REG_26__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U18994 ( .A1(n19459), .A2(n19478), .B1(n19522), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15524) );
  OAI211_X1 U18995 ( .C1(n15576), .C2(n15811), .A(n15525), .B(n15524), .ZN(
        n15526) );
  AOI21_X1 U18996 ( .B1(n15527), .B2(n19505), .A(n15526), .ZN(n15528) );
  INV_X1 U18997 ( .A(n15528), .ZN(P2_U2893) );
  XOR2_X1 U18998 ( .A(n15529), .B(n15538), .Z(n16531) );
  INV_X1 U18999 ( .A(n19481), .ZN(n15530) );
  OAI22_X1 U19000 ( .A1(n15543), .A2(n15530), .B1(n19489), .B2(n19551), .ZN(
        n15531) );
  AOI21_X1 U19001 ( .B1(n19523), .B2(n16531), .A(n15531), .ZN(n15533) );
  AOI22_X1 U19002 ( .A1(n19461), .A2(BUF1_REG_25__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15532) );
  OAI211_X1 U19003 ( .C1(n15534), .C2(n19527), .A(n15533), .B(n15532), .ZN(
        P2_U2894) );
  NAND2_X1 U19004 ( .A1(n15536), .A2(n15535), .ZN(n15537) );
  AND2_X1 U19005 ( .A1(n15538), .A2(n15537), .ZN(n16540) );
  OAI22_X1 U19006 ( .A1(n15543), .A2(n19485), .B1(n19489), .B2(n19553), .ZN(
        n15539) );
  AOI21_X1 U19007 ( .B1(n19523), .B2(n16540), .A(n15539), .ZN(n15541) );
  AOI22_X1 U19008 ( .A1(n19461), .A2(BUF1_REG_24__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15540) );
  OAI211_X1 U19009 ( .C1(n15542), .C2(n19527), .A(n15541), .B(n15540), .ZN(
        P2_U2895) );
  INV_X1 U19010 ( .A(n15849), .ZN(n15545) );
  INV_X1 U19011 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19555) );
  OAI22_X1 U19012 ( .A1(n15543), .A2(n19698), .B1(n19489), .B2(n19555), .ZN(
        n15544) );
  AOI21_X1 U19013 ( .B1(n19523), .B2(n15545), .A(n15544), .ZN(n15547) );
  AOI22_X1 U19014 ( .A1(n19461), .A2(BUF1_REG_23__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15546) );
  OAI211_X1 U19015 ( .C1(n15548), .C2(n19527), .A(n15547), .B(n15546), .ZN(
        P2_U2896) );
  NAND2_X1 U19016 ( .A1(n15549), .A2(n19505), .ZN(n15554) );
  AOI22_X1 U19017 ( .A1(n19459), .A2(n19492), .B1(n19522), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15553) );
  AOI22_X1 U19018 ( .A1(n19461), .A2(BUF1_REG_21__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15552) );
  INV_X1 U19019 ( .A(n15877), .ZN(n15550) );
  NAND2_X1 U19020 ( .A1(n19523), .A2(n15550), .ZN(n15551) );
  NAND4_X1 U19021 ( .A1(n15554), .A2(n15553), .A3(n15552), .A4(n15551), .ZN(
        P2_U2898) );
  OR2_X1 U19022 ( .A1(n15555), .A2(n19527), .ZN(n15560) );
  AOI22_X1 U19023 ( .A1(n19459), .A2(n15556), .B1(n19522), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15559) );
  AOI22_X1 U19024 ( .A1(n19461), .A2(BUF1_REG_19__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15558) );
  NAND2_X1 U19025 ( .A1(n19523), .A2(n15907), .ZN(n15557) );
  NAND4_X1 U19026 ( .A1(n15560), .A2(n15559), .A3(n15558), .A4(n15557), .ZN(
        P2_U2900) );
  INV_X1 U19027 ( .A(n15561), .ZN(n15563) );
  NAND2_X1 U19028 ( .A1(n15572), .A2(n9812), .ZN(n15562) );
  NAND2_X1 U19029 ( .A1(n15563), .A2(n15562), .ZN(n15564) );
  NAND2_X1 U19030 ( .A1(n15565), .A2(n15564), .ZN(n19282) );
  AOI22_X1 U19031 ( .A1(n19461), .A2(BUF1_REG_18__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U19032 ( .A1(n19459), .A2(n15566), .B1(n19522), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15567) );
  OAI211_X1 U19033 ( .C1(n15576), .C2(n19282), .A(n15568), .B(n15567), .ZN(
        n15569) );
  INV_X1 U19034 ( .A(n15569), .ZN(n15570) );
  OAI21_X1 U19035 ( .B1(n15571), .B2(n19527), .A(n15570), .ZN(P2_U2901) );
  XNOR2_X1 U19036 ( .A(n15572), .B(n9812), .ZN(n19288) );
  AOI22_X1 U19037 ( .A1(n19461), .A2(BUF1_REG_17__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n15575) );
  AOI22_X1 U19038 ( .A1(n19459), .A2(n15573), .B1(n19522), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15574) );
  OAI211_X1 U19039 ( .C1(n19288), .C2(n15576), .A(n15575), .B(n15574), .ZN(
        n15577) );
  AOI21_X1 U19040 ( .B1(n15578), .B2(n19505), .A(n15577), .ZN(n15579) );
  INV_X1 U19041 ( .A(n15579), .ZN(P2_U2902) );
  NAND2_X1 U19042 ( .A1(n15580), .A2(n15592), .ZN(n15583) );
  NOR2_X1 U19043 ( .A1(n15581), .A2(n11579), .ZN(n15582) );
  XNOR2_X1 U19044 ( .A(n15583), .B(n15582), .ZN(n15784) );
  XNOR2_X1 U19045 ( .A(n15588), .B(n15779), .ZN(n15782) );
  NAND2_X1 U19046 ( .A1(n16638), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15584) );
  NAND2_X1 U19047 ( .A1(n19643), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15776) );
  OAI211_X1 U19048 ( .C1(n15773), .C2(n14135), .A(n15584), .B(n15776), .ZN(
        n15586) );
  NOR2_X1 U19049 ( .A1(n16492), .A2(n19634), .ZN(n15585) );
  AOI21_X1 U19050 ( .B1(n15782), .B2(n16632), .A(n9790), .ZN(n15587) );
  OAI21_X1 U19051 ( .B1(n15784), .B2(n19619), .A(n15587), .ZN(P2_U2984) );
  INV_X1 U19052 ( .A(n15588), .ZN(n15591) );
  NAND2_X1 U19053 ( .A1(n11597), .A2(n15589), .ZN(n15590) );
  NAND2_X1 U19054 ( .A1(n15591), .A2(n15590), .ZN(n15796) );
  NAND2_X1 U19055 ( .A1(n15593), .A2(n15592), .ZN(n15594) );
  XNOR2_X1 U19056 ( .A(n15595), .B(n15594), .ZN(n15785) );
  NAND2_X1 U19057 ( .A1(n15785), .A2(n12997), .ZN(n15599) );
  NAND2_X1 U19058 ( .A1(n19643), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15790) );
  NAND2_X1 U19059 ( .A1(n16638), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15596) );
  OAI211_X1 U19060 ( .C1(n15786), .C2(n14135), .A(n15790), .B(n15596), .ZN(
        n15597) );
  AOI21_X1 U19061 ( .B1(n10253), .B2(n19613), .A(n15597), .ZN(n15598) );
  OAI211_X1 U19062 ( .C1(n19636), .C2(n15796), .A(n15599), .B(n15598), .ZN(
        P2_U2985) );
  INV_X1 U19063 ( .A(n15600), .ZN(n15606) );
  NOR2_X1 U19064 ( .A1(n16496), .A2(n14135), .ZN(n15601) );
  AOI211_X1 U19065 ( .C1(n16638), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15602), .B(n15601), .ZN(n15603) );
  OAI21_X1 U19066 ( .B1(n15604), .B2(n19634), .A(n15603), .ZN(n15605) );
  AOI21_X1 U19067 ( .B1(n15606), .B2(n16568), .A(n15605), .ZN(n15607) );
  OAI21_X1 U19068 ( .B1(n15608), .B2(n19619), .A(n15607), .ZN(P2_U2986) );
  OR2_X1 U19069 ( .A1(n15609), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15610) );
  NAND2_X1 U19070 ( .A1(n15611), .A2(n15610), .ZN(n15810) );
  OR2_X1 U19071 ( .A1(n15612), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15797) );
  NAND3_X1 U19072 ( .A1(n15797), .A2(n15613), .A3(n12997), .ZN(n15618) );
  INV_X1 U19073 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20243) );
  NOR2_X1 U19074 ( .A1(n19272), .A2(n20243), .ZN(n15798) );
  AOI21_X1 U19075 ( .B1(n16638), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15798), .ZN(n15614) );
  OAI21_X1 U19076 ( .B1(n15805), .B2(n14135), .A(n15614), .ZN(n15615) );
  AOI21_X1 U19077 ( .B1(n15616), .B2(n19613), .A(n15615), .ZN(n15617) );
  OAI211_X1 U19078 ( .C1(n19636), .C2(n15810), .A(n15618), .B(n15617), .ZN(
        P2_U2987) );
  NOR2_X1 U19079 ( .A1(n15619), .A2(n15621), .ZN(n15620) );
  MUX2_X1 U19080 ( .A(n15621), .B(n15620), .S(n15630), .Z(n15623) );
  INV_X1 U19081 ( .A(n15624), .ZN(n15637) );
  NAND2_X1 U19082 ( .A1(n15624), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15831) );
  AOI21_X1 U19083 ( .B1(n15814), .B2(n15831), .A(n15609), .ZN(n15820) );
  INV_X1 U19084 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20240) );
  NOR2_X1 U19085 ( .A1(n19272), .A2(n20240), .ZN(n15816) );
  NOR2_X1 U19086 ( .A1(n16510), .A2(n14135), .ZN(n15625) );
  AOI211_X1 U19087 ( .C1(n16638), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15816), .B(n15625), .ZN(n15626) );
  OAI21_X1 U19088 ( .B1(n19634), .B2(n15627), .A(n15626), .ZN(n15628) );
  AOI21_X1 U19089 ( .B1(n15820), .B2(n16632), .A(n15628), .ZN(n15629) );
  OAI21_X1 U19090 ( .B1(n15822), .B2(n19619), .A(n15629), .ZN(P2_U2988) );
  INV_X1 U19091 ( .A(n15630), .ZN(n15631) );
  NOR2_X1 U19092 ( .A1(n15632), .A2(n15631), .ZN(n15634) );
  XOR2_X1 U19093 ( .A(n15634), .B(n15633), .Z(n15834) );
  INV_X1 U19094 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20238) );
  NOR2_X1 U19095 ( .A1(n19272), .A2(n20238), .ZN(n15826) );
  AOI21_X1 U19096 ( .B1(n16638), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15826), .ZN(n15635) );
  OAI21_X1 U19097 ( .B1(n16524), .B2(n14135), .A(n15635), .ZN(n15636) );
  AOI21_X1 U19098 ( .B1(n16522), .B2(n19613), .A(n15636), .ZN(n15639) );
  NAND2_X1 U19099 ( .A1(n15637), .A2(n15813), .ZN(n15830) );
  NAND3_X1 U19100 ( .A1(n15831), .A2(n16632), .A3(n15830), .ZN(n15638) );
  OAI211_X1 U19101 ( .C1(n15834), .C2(n19619), .A(n15639), .B(n15638), .ZN(
        P2_U2989) );
  NOR2_X1 U19102 ( .A1(n15641), .A2(n10158), .ZN(n15642) );
  XNOR2_X1 U19103 ( .A(n15643), .B(n15642), .ZN(n15842) );
  AOI21_X1 U19104 ( .B1(n15644), .B2(n15844), .A(n15624), .ZN(n15840) );
  INV_X1 U19105 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20236) );
  OAI22_X1 U19106 ( .A1(n20236), .A2(n19272), .B1(n19634), .B2(n15645), .ZN(
        n15648) );
  INV_X1 U19107 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15646) );
  OAI22_X1 U19108 ( .A1(n16542), .A2(n14135), .B1(n15646), .B2(n19642), .ZN(
        n15647) );
  AOI211_X1 U19109 ( .C1(n15840), .C2(n16632), .A(n15648), .B(n15647), .ZN(
        n15649) );
  OAI21_X1 U19110 ( .B1(n15842), .B2(n19619), .A(n15649), .ZN(P2_U2990) );
  NAND2_X1 U19111 ( .A1(n15651), .A2(n15650), .ZN(n15653) );
  XOR2_X1 U19112 ( .A(n15653), .B(n15652), .Z(n15871) );
  NOR2_X1 U19113 ( .A1(n16131), .A2(n14135), .ZN(n15656) );
  INV_X1 U19114 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n21096) );
  OAI22_X1 U19115 ( .A1(n21096), .A2(n19272), .B1(n19634), .B2(n15654), .ZN(
        n15655) );
  AOI211_X1 U19116 ( .C1(n16638), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15656), .B(n15655), .ZN(n15661) );
  INV_X1 U19117 ( .A(n15657), .ZN(n15658) );
  NAND2_X1 U19118 ( .A1(n15658), .A2(n15864), .ZN(n15868) );
  NAND3_X1 U19119 ( .A1(n15868), .A2(n16568), .A3(n15659), .ZN(n15660) );
  OAI211_X1 U19120 ( .C1(n15871), .C2(n19619), .A(n15661), .B(n15660), .ZN(
        P2_U2992) );
  NAND2_X1 U19121 ( .A1(n15663), .A2(n15662), .ZN(n15676) );
  NAND2_X1 U19122 ( .A1(n16586), .A2(n16585), .ZN(n16576) );
  NAND2_X1 U19123 ( .A1(n16576), .A2(n15666), .ZN(n15667) );
  INV_X1 U19124 ( .A(n16121), .ZN(n15668) );
  INV_X1 U19125 ( .A(n15724), .ZN(n15671) );
  INV_X1 U19126 ( .A(n15672), .ZN(n15711) );
  INV_X1 U19127 ( .A(n15673), .ZN(n15674) );
  NAND2_X1 U19128 ( .A1(n15689), .A2(n15684), .ZN(n15675) );
  XOR2_X1 U19129 ( .A(n15676), .B(n15675), .Z(n15884) );
  NOR2_X1 U19130 ( .A1(n19272), .A2(n20232), .ZN(n15873) );
  AOI21_X1 U19131 ( .B1(n16638), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15873), .ZN(n15677) );
  OAI21_X1 U19132 ( .B1(n15678), .B2(n14135), .A(n15677), .ZN(n15681) );
  INV_X1 U19133 ( .A(n15679), .ZN(n15692) );
  NOR2_X1 U19134 ( .A1(n15692), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15878) );
  NOR3_X1 U19135 ( .A1(n15878), .A2(n15657), .A3(n19636), .ZN(n15680) );
  AOI211_X1 U19136 ( .C1(n19613), .C2(n15682), .A(n15681), .B(n15680), .ZN(
        n15683) );
  OAI21_X1 U19137 ( .B1(n15884), .B2(n19619), .A(n15683), .ZN(P2_U2993) );
  INV_X1 U19138 ( .A(n15684), .ZN(n15688) );
  AND2_X1 U19139 ( .A1(n15685), .A2(n15684), .ZN(n15686) );
  OAI22_X1 U19140 ( .A1(n15689), .A2(n15688), .B1(n15687), .B2(n15686), .ZN(
        n15903) );
  AOI21_X1 U19141 ( .B1(n15691), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15693) );
  NOR2_X1 U19142 ( .A1(n15693), .A2(n15692), .ZN(n15901) );
  INV_X1 U19143 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20230) );
  NOR2_X1 U19144 ( .A1(n19272), .A2(n20230), .ZN(n15895) );
  AOI21_X1 U19145 ( .B1(n16638), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15895), .ZN(n15695) );
  NAND2_X1 U19146 ( .A1(n19260), .A2(n19622), .ZN(n15694) );
  OAI211_X1 U19147 ( .C1(n15696), .C2(n19634), .A(n15695), .B(n15694), .ZN(
        n15697) );
  AOI21_X1 U19148 ( .B1(n15901), .B2(n16632), .A(n15697), .ZN(n15698) );
  OAI21_X1 U19149 ( .B1(n15903), .B2(n19619), .A(n15698), .ZN(P2_U2994) );
  NAND2_X1 U19150 ( .A1(n15700), .A2(n15699), .ZN(n15704) );
  INV_X1 U19151 ( .A(n15701), .ZN(n15710) );
  NOR2_X1 U19152 ( .A1(n15702), .A2(n15710), .ZN(n15703) );
  XOR2_X1 U19153 ( .A(n15704), .B(n15703), .Z(n15915) );
  XNOR2_X1 U19154 ( .A(n15690), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15913) );
  NOR2_X1 U19155 ( .A1(n19272), .A2(n20229), .ZN(n15906) );
  NOR2_X1 U19156 ( .A1(n15904), .A2(n14135), .ZN(n15705) );
  AOI211_X1 U19157 ( .C1(n16638), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15906), .B(n15705), .ZN(n15706) );
  OAI21_X1 U19158 ( .B1(n15707), .B2(n19634), .A(n15706), .ZN(n15708) );
  AOI21_X1 U19159 ( .B1(n15913), .B2(n16568), .A(n15708), .ZN(n15709) );
  OAI21_X1 U19160 ( .B1(n15915), .B2(n19619), .A(n15709), .ZN(P2_U2995) );
  NOR2_X1 U19161 ( .A1(n15711), .A2(n15710), .ZN(n15712) );
  XNOR2_X1 U19162 ( .A(n15713), .B(n15712), .ZN(n15928) );
  NOR2_X1 U19163 ( .A1(n19275), .A2(n14135), .ZN(n15716) );
  INV_X1 U19164 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20227) );
  OAI22_X1 U19165 ( .A1(n20227), .A2(n19272), .B1(n19634), .B2(n15714), .ZN(
        n15715) );
  AOI211_X1 U19166 ( .C1(n16638), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15716), .B(n15715), .ZN(n15720) );
  NAND2_X1 U19167 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16146) );
  NOR2_X2 U19168 ( .A1(n16146), .A2(n16583), .ZN(n16567) );
  NAND2_X1 U19169 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16567), .ZN(
        n15725) );
  NAND2_X1 U19170 ( .A1(n15718), .A2(n15725), .ZN(n15925) );
  NAND3_X1 U19171 ( .A1(n15690), .A2(n16568), .A3(n15925), .ZN(n15719) );
  OAI211_X1 U19172 ( .C1(n15928), .C2(n19619), .A(n15720), .B(n15719), .ZN(
        P2_U2996) );
  NOR2_X1 U19173 ( .A1(n15722), .A2(n15721), .ZN(n15723) );
  XNOR2_X1 U19174 ( .A(n15724), .B(n15723), .ZN(n16150) );
  OAI211_X1 U19175 ( .C1(n16567), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16568), .B(n15725), .ZN(n15728) );
  INV_X1 U19176 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20226) );
  NOR2_X1 U19177 ( .A1(n20226), .A2(n19272), .ZN(n16145) );
  INV_X1 U19178 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19283) );
  OAI22_X1 U19179 ( .A1(n19283), .A2(n19642), .B1(n19634), .B2(n19291), .ZN(
        n15726) );
  AOI211_X1 U19180 ( .C1(n19622), .C2(n19290), .A(n16145), .B(n15726), .ZN(
        n15727) );
  OAI211_X1 U19181 ( .C1(n16150), .C2(n19619), .A(n15728), .B(n15727), .ZN(
        P2_U2997) );
  OR2_X1 U19182 ( .A1(n15743), .A2(n15730), .ZN(n16616) );
  INV_X1 U19183 ( .A(n16616), .ZN(n15729) );
  AOI21_X1 U19184 ( .B1(n15730), .B2(n15743), .A(n15729), .ZN(n16699) );
  INV_X1 U19185 ( .A(n15731), .ZN(n15744) );
  OR2_X1 U19186 ( .A1(n15732), .A2(n15744), .ZN(n15736) );
  AND2_X1 U19187 ( .A1(n15734), .A2(n15733), .ZN(n15735) );
  XNOR2_X1 U19188 ( .A(n15736), .B(n15735), .ZN(n16703) );
  AOI22_X1 U19189 ( .A1(n19358), .A2(n19622), .B1(n19613), .B2(n19357), .ZN(
        n15740) );
  INV_X1 U19190 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20215) );
  OAI22_X1 U19191 ( .A1(n20215), .A2(n19272), .B1(n15737), .B2(n19642), .ZN(
        n15738) );
  INV_X1 U19192 ( .A(n15738), .ZN(n15739) );
  OAI211_X1 U19193 ( .C1(n16703), .C2(n19619), .A(n15740), .B(n15739), .ZN(
        n15741) );
  AOI21_X1 U19194 ( .B1(n16699), .B2(n16632), .A(n15741), .ZN(n15742) );
  INV_X1 U19195 ( .A(n15742), .ZN(P2_U3004) );
  OAI21_X1 U19196 ( .B1(n15717), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15743), .ZN(n15953) );
  NOR2_X1 U19197 ( .A1(n15745), .A2(n15744), .ZN(n15746) );
  XNOR2_X1 U19198 ( .A(n15747), .B(n15746), .ZN(n15951) );
  INV_X1 U19199 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19372) );
  OAI22_X1 U19200 ( .A1(n19372), .A2(n19642), .B1(n19634), .B2(n19366), .ZN(
        n15750) );
  INV_X1 U19201 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15748) );
  OAI22_X1 U19202 ( .A1(n19367), .A2(n14135), .B1(n19272), .B2(n15748), .ZN(
        n15749) );
  AOI211_X1 U19203 ( .C1(n15951), .C2(n12997), .A(n15750), .B(n15749), .ZN(
        n15751) );
  OAI21_X1 U19204 ( .B1(n15953), .B2(n19636), .A(n15751), .ZN(P2_U3005) );
  XNOR2_X1 U19205 ( .A(n15752), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15964) );
  INV_X1 U19206 ( .A(n16625), .ZN(n15754) );
  NAND2_X1 U19207 ( .A1(n15754), .A2(n16626), .ZN(n15755) );
  XNOR2_X1 U19208 ( .A(n15753), .B(n15755), .ZN(n15962) );
  INV_X1 U19209 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20211) );
  OAI22_X1 U19210 ( .A1(n20211), .A2(n19272), .B1(n19634), .B2(n19386), .ZN(
        n15758) );
  INV_X1 U19211 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15756) );
  OAI22_X1 U19212 ( .A1(n19390), .A2(n14135), .B1(n19642), .B2(n15756), .ZN(
        n15757) );
  AOI211_X1 U19213 ( .C1(n15962), .C2(n12997), .A(n15758), .B(n15757), .ZN(
        n15759) );
  OAI21_X1 U19214 ( .B1(n15964), .B2(n19636), .A(n15759), .ZN(P2_U3007) );
  AND2_X1 U19215 ( .A1(n15761), .A2(n15760), .ZN(n15763) );
  OAI22_X1 U19216 ( .A1(n9726), .A2(n15764), .B1(n15763), .B2(n15762), .ZN(
        n15991) );
  XOR2_X1 U19217 ( .A(n15766), .B(n15767), .Z(n15993) );
  NAND2_X1 U19218 ( .A1(n15993), .A2(n12997), .ZN(n15772) );
  INV_X1 U19219 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19421) );
  OAI22_X1 U19220 ( .A1(n19421), .A2(n19642), .B1(n19634), .B2(n19412), .ZN(
        n15770) );
  INV_X1 U19221 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15768) );
  OAI22_X1 U19222 ( .A1(n19413), .A2(n14135), .B1(n19272), .B2(n15768), .ZN(
        n15769) );
  NOR2_X1 U19223 ( .A1(n15770), .A2(n15769), .ZN(n15771) );
  OAI211_X1 U19224 ( .C1(n19636), .C2(n15991), .A(n15772), .B(n15771), .ZN(
        P2_U3009) );
  INV_X1 U19225 ( .A(n15773), .ZN(n15778) );
  NAND3_X1 U19226 ( .A1(n15799), .A2(n15774), .A3(n15779), .ZN(n15775) );
  AOI21_X1 U19227 ( .B1(n15782), .B2(n19660), .A(n15781), .ZN(n15783) );
  OAI21_X1 U19228 ( .B1(n15784), .B2(n16702), .A(n15783), .ZN(P2_U3016) );
  NAND2_X1 U19229 ( .A1(n15785), .A2(n19663), .ZN(n15795) );
  NOR2_X1 U19230 ( .A1(n15786), .A2(n16143), .ZN(n15793) );
  OAI211_X1 U19231 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15788), .A(
        n15799), .B(n15787), .ZN(n15789) );
  OAI211_X1 U19232 ( .C1(n19667), .C2(n15791), .A(n15790), .B(n15789), .ZN(
        n15792) );
  AOI211_X1 U19233 ( .C1(n15807), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15793), .B(n15792), .ZN(n15794) );
  OAI211_X1 U19234 ( .C1(n15796), .C2(n19650), .A(n15795), .B(n15794), .ZN(
        P2_U3017) );
  NAND3_X1 U19235 ( .A1(n15797), .A2(n15613), .A3(n19663), .ZN(n15809) );
  INV_X1 U19236 ( .A(n15798), .ZN(n15801) );
  NAND2_X1 U19237 ( .A1(n15799), .A2(n11569), .ZN(n15800) );
  OAI211_X1 U19238 ( .C1(n19667), .C2(n15802), .A(n15801), .B(n15800), .ZN(
        n15803) );
  INV_X1 U19239 ( .A(n15803), .ZN(n15804) );
  OAI21_X1 U19240 ( .B1(n15805), .B2(n16143), .A(n15804), .ZN(n15806) );
  AOI21_X1 U19241 ( .B1(n15807), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15806), .ZN(n15808) );
  OAI211_X1 U19242 ( .C1(n15810), .C2(n19650), .A(n15809), .B(n15808), .ZN(
        P2_U3019) );
  NOR2_X1 U19243 ( .A1(n15823), .A2(n15814), .ZN(n15819) );
  INV_X1 U19244 ( .A(n15811), .ZN(n16511) );
  AOI211_X1 U19245 ( .C1(n15814), .C2(n15813), .A(n15824), .B(n10908), .ZN(
        n15815) );
  AOI211_X1 U19246 ( .C1(n19645), .C2(n16511), .A(n15816), .B(n15815), .ZN(
        n15817) );
  OAI21_X1 U19247 ( .B1(n16510), .B2(n16143), .A(n15817), .ZN(n15818) );
  AOI211_X1 U19248 ( .C1(n15820), .C2(n19660), .A(n15819), .B(n15818), .ZN(
        n15821) );
  OAI21_X1 U19249 ( .B1(n15822), .B2(n16702), .A(n15821), .ZN(P2_U3020) );
  INV_X1 U19250 ( .A(n15823), .ZN(n15829) );
  NOR2_X1 U19251 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15824), .ZN(
        n15825) );
  AOI211_X1 U19252 ( .C1(n19645), .C2(n16531), .A(n15826), .B(n15825), .ZN(
        n15827) );
  OAI21_X1 U19253 ( .B1(n16524), .B2(n16143), .A(n15827), .ZN(n15828) );
  AOI21_X1 U19254 ( .B1(n15829), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15828), .ZN(n15833) );
  NAND3_X1 U19255 ( .A1(n15831), .A2(n19660), .A3(n15830), .ZN(n15832) );
  OAI211_X1 U19256 ( .C1(n15834), .C2(n16702), .A(n15833), .B(n15832), .ZN(
        P2_U3021) );
  OAI21_X1 U19257 ( .B1(n15836), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15835), .ZN(n15838) );
  AOI22_X1 U19258 ( .A1(n19645), .A2(n16540), .B1(n19643), .B2(
        P2_REIP_REG_24__SCAN_IN), .ZN(n15837) );
  OAI211_X1 U19259 ( .C1(n16143), .C2(n16542), .A(n15838), .B(n15837), .ZN(
        n15839) );
  AOI21_X1 U19260 ( .B1(n15840), .B2(n19660), .A(n15839), .ZN(n15841) );
  OAI21_X1 U19261 ( .B1(n15842), .B2(n16702), .A(n15841), .ZN(P2_U3022) );
  NAND2_X1 U19262 ( .A1(n15659), .A2(n15853), .ZN(n15843) );
  AND2_X1 U19263 ( .A1(n15844), .A2(n15843), .ZN(n16563) );
  INV_X1 U19264 ( .A(n16563), .ZN(n15858) );
  OR2_X1 U19265 ( .A1(n15846), .A2(n15845), .ZN(n16559) );
  AND3_X1 U19266 ( .A1(n16559), .A2(n19663), .A3(n15847), .ZN(n15856) );
  AOI211_X1 U19267 ( .C1(n15864), .C2(n15853), .A(n15848), .B(n15865), .ZN(
        n15855) );
  INV_X1 U19268 ( .A(n16561), .ZN(n15851) );
  INV_X1 U19269 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21139) );
  OAI22_X1 U19270 ( .A1(n19667), .A2(n15849), .B1(n21139), .B2(n19272), .ZN(
        n15850) );
  AOI21_X1 U19271 ( .B1(n15851), .B2(n19669), .A(n15850), .ZN(n15852) );
  OAI21_X1 U19272 ( .B1(n15863), .B2(n15853), .A(n15852), .ZN(n15854) );
  NOR3_X1 U19273 ( .A1(n15856), .A2(n15855), .A3(n15854), .ZN(n15857) );
  OAI21_X1 U19274 ( .B1(n15858), .B2(n19650), .A(n15857), .ZN(P2_U3023) );
  AOI21_X1 U19275 ( .B1(n15861), .B2(n15860), .A(n15859), .ZN(n16547) );
  NOR2_X1 U19276 ( .A1(n16131), .A2(n16143), .ZN(n15867) );
  NAND2_X1 U19277 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19643), .ZN(n15862) );
  OAI221_X1 U19278 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15865), 
        .C1(n15864), .C2(n15863), .A(n15862), .ZN(n15866) );
  AOI211_X1 U19279 ( .C1(n19645), .C2(n16547), .A(n15867), .B(n15866), .ZN(
        n15870) );
  NAND3_X1 U19280 ( .A1(n15868), .A2(n19660), .A3(n15659), .ZN(n15869) );
  OAI211_X1 U19281 ( .C1(n15871), .C2(n16702), .A(n15870), .B(n15869), .ZN(
        P2_U3024) );
  NAND3_X1 U19282 ( .A1(n15872), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16115), .ZN(n15876) );
  AOI21_X1 U19283 ( .B1(n15874), .B2(n19669), .A(n15873), .ZN(n15875) );
  OAI211_X1 U19284 ( .C1(n19667), .C2(n15877), .A(n15876), .B(n15875), .ZN(
        n15880) );
  NOR3_X1 U19285 ( .A1(n15878), .A2(n15657), .A3(n19650), .ZN(n15879) );
  AOI211_X1 U19286 ( .C1(n15882), .C2(n15881), .A(n15880), .B(n15879), .ZN(
        n15883) );
  OAI21_X1 U19287 ( .B1(n15884), .B2(n16702), .A(n15883), .ZN(P2_U3025) );
  OAI21_X1 U19288 ( .B1(n15885), .B2(n16681), .A(n16682), .ZN(n15924) );
  NAND2_X1 U19289 ( .A1(n15937), .A2(n16683), .ZN(n16654) );
  NAND2_X1 U19290 ( .A1(n15886), .A2(n16669), .ZN(n16646) );
  NOR2_X1 U19291 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16646), .ZN(
        n15916) );
  NOR2_X1 U19292 ( .A1(n15924), .A2(n15916), .ZN(n15911) );
  AND2_X1 U19293 ( .A1(n15887), .A2(n15910), .ZN(n15888) );
  NAND2_X1 U19294 ( .A1(n16683), .A2(n15888), .ZN(n15908) );
  AOI21_X1 U19295 ( .B1(n15911), .B2(n15908), .A(n15890), .ZN(n15900) );
  INV_X1 U19296 ( .A(n15889), .ZN(n15891) );
  NAND3_X1 U19297 ( .A1(n16683), .A2(n15891), .A3(n15890), .ZN(n15897) );
  AOI21_X1 U19298 ( .B1(n15894), .B2(n15893), .A(n15892), .ZN(n19259) );
  AOI21_X1 U19299 ( .B1(n19645), .B2(n19259), .A(n15895), .ZN(n15896) );
  OAI211_X1 U19300 ( .C1(n15898), .C2(n16143), .A(n15897), .B(n15896), .ZN(
        n15899) );
  AOI211_X1 U19301 ( .C1(n15901), .C2(n19660), .A(n15900), .B(n15899), .ZN(
        n15902) );
  OAI21_X1 U19302 ( .B1(n15903), .B2(n16702), .A(n15902), .ZN(P2_U3026) );
  NOR2_X1 U19303 ( .A1(n16143), .A2(n15904), .ZN(n15905) );
  AOI211_X1 U19304 ( .C1(n19645), .C2(n15907), .A(n15906), .B(n15905), .ZN(
        n15909) );
  OAI211_X1 U19305 ( .C1(n15911), .C2(n15910), .A(n15909), .B(n15908), .ZN(
        n15912) );
  AOI21_X1 U19306 ( .B1(n15913), .B2(n19660), .A(n15912), .ZN(n15914) );
  OAI21_X1 U19307 ( .B1(n15915), .B2(n16702), .A(n15914), .ZN(P2_U3027) );
  INV_X1 U19308 ( .A(n19282), .ZN(n15921) );
  NOR2_X1 U19309 ( .A1(n20227), .A2(n19272), .ZN(n15920) );
  INV_X1 U19310 ( .A(n15916), .ZN(n15918) );
  NOR2_X1 U19311 ( .A1(n15918), .A2(n15917), .ZN(n15919) );
  AOI211_X1 U19312 ( .C1(n19645), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        n15922) );
  OAI21_X1 U19313 ( .B1(n16143), .B2(n19275), .A(n15922), .ZN(n15923) );
  AOI21_X1 U19314 ( .B1(n15924), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15923), .ZN(n15927) );
  NAND3_X1 U19315 ( .A1(n15690), .A2(n19660), .A3(n15925), .ZN(n15926) );
  OAI211_X1 U19316 ( .C1(n15928), .C2(n16702), .A(n15927), .B(n15926), .ZN(
        P2_U3028) );
  NAND2_X1 U19317 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15929), .ZN(
        n16593) );
  OAI21_X1 U19318 ( .B1(n15929), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16593), .ZN(n16602) );
  INV_X1 U19319 ( .A(n15931), .ZN(n15933) );
  NOR2_X1 U19320 ( .A1(n15933), .A2(n15932), .ZN(n15934) );
  XNOR2_X1 U19321 ( .A(n15930), .B(n15934), .ZN(n16601) );
  INV_X1 U19322 ( .A(n16601), .ZN(n15943) );
  XNOR2_X1 U19323 ( .A(n15936), .B(n15935), .ZN(n19475) );
  OAI21_X1 U19324 ( .B1(n15937), .B2(n16726), .A(n16682), .ZN(n16655) );
  INV_X1 U19325 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20217) );
  NOR2_X1 U19326 ( .A1(n20217), .A2(n19272), .ZN(n15938) );
  AOI221_X1 U19327 ( .B1(n16669), .B2(n15939), .C1(n16655), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15938), .ZN(n15941) );
  NAND2_X1 U19328 ( .A1(n19669), .A2(n19347), .ZN(n15940) );
  OAI211_X1 U19329 ( .C1(n19667), .C2(n19475), .A(n15941), .B(n15940), .ZN(
        n15942) );
  AOI21_X1 U19330 ( .B1(n15943), .B2(n19663), .A(n15942), .ZN(n15944) );
  OAI21_X1 U19331 ( .B1(n16602), .B2(n19650), .A(n15944), .ZN(P2_U3034) );
  INV_X1 U19332 ( .A(n16682), .ZN(n15946) );
  NOR2_X1 U19333 ( .A1(n15748), .A2(n19272), .ZN(n15945) );
  AOI221_X1 U19334 ( .B1(n16683), .B2(n11274), .C1(n15946), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15945), .ZN(n15947) );
  INV_X1 U19335 ( .A(n15947), .ZN(n15950) );
  OAI21_X1 U19336 ( .B1(n16704), .B2(n15948), .A(n16694), .ZN(n19483) );
  OAI22_X1 U19337 ( .A1(n19483), .A2(n19667), .B1(n16143), .B2(n19367), .ZN(
        n15949) );
  AOI211_X1 U19338 ( .C1(n15951), .C2(n19663), .A(n15950), .B(n15949), .ZN(
        n15952) );
  OAI21_X1 U19339 ( .B1(n15953), .B2(n19650), .A(n15952), .ZN(P2_U3037) );
  INV_X1 U19340 ( .A(n15954), .ZN(n16711) );
  NOR2_X1 U19341 ( .A1(n20211), .A2(n19272), .ZN(n15955) );
  AOI221_X1 U19342 ( .B1(n16707), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16711), .C2(n11451), .A(n15955), .ZN(n15956) );
  INV_X1 U19343 ( .A(n15956), .ZN(n15961) );
  OR2_X1 U19344 ( .A1(n15958), .A2(n15957), .ZN(n15959) );
  NAND2_X1 U19345 ( .A1(n15959), .A2(n16705), .ZN(n19487) );
  OAI22_X1 U19346 ( .A1(n19487), .A2(n19667), .B1(n16143), .B2(n19390), .ZN(
        n15960) );
  AOI211_X1 U19347 ( .C1(n15962), .C2(n19663), .A(n15961), .B(n15960), .ZN(
        n15963) );
  OAI21_X1 U19348 ( .B1(n15964), .B2(n19650), .A(n15963), .ZN(P2_U3039) );
  XNOR2_X1 U19349 ( .A(n15965), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16640) );
  XNOR2_X1 U19350 ( .A(n15967), .B(n15966), .ZN(n16639) );
  INV_X1 U19351 ( .A(n16639), .ZN(n15976) );
  XNOR2_X1 U19352 ( .A(n15969), .B(n15968), .ZN(n19490) );
  INV_X1 U19353 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20209) );
  NOR2_X1 U19354 ( .A1(n20209), .A2(n19272), .ZN(n15970) );
  AOI221_X1 U19355 ( .B1(n16707), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        n15972), .C2(n15971), .A(n15970), .ZN(n15974) );
  NAND2_X1 U19356 ( .A1(n19669), .A2(n19402), .ZN(n15973) );
  OAI211_X1 U19357 ( .C1(n19667), .C2(n19490), .A(n15974), .B(n15973), .ZN(
        n15975) );
  AOI21_X1 U19358 ( .B1(n15976), .B2(n19663), .A(n15975), .ZN(n15977) );
  OAI21_X1 U19359 ( .B1(n16640), .B2(n19650), .A(n15977), .ZN(P2_U3040) );
  OAI21_X1 U19360 ( .B1(n19425), .B2(n15979), .A(n15978), .ZN(n19500) );
  INV_X1 U19361 ( .A(n19500), .ZN(n15985) );
  NAND2_X1 U19362 ( .A1(n16115), .A2(n15980), .ZN(n19646) );
  INV_X1 U19363 ( .A(n19413), .ZN(n15982) );
  NOR2_X1 U19364 ( .A1(n15768), .A2(n19272), .ZN(n15981) );
  AOI21_X1 U19365 ( .B1(n19669), .B2(n15982), .A(n15981), .ZN(n15983) );
  OAI21_X1 U19366 ( .B1(n19646), .B2(n15987), .A(n15983), .ZN(n15984) );
  AOI21_X1 U19367 ( .B1(n15985), .B2(n19645), .A(n15984), .ZN(n15990) );
  AOI211_X1 U19368 ( .C1(n10787), .C2(n15987), .A(n15986), .B(n19656), .ZN(
        n15988) );
  INV_X1 U19369 ( .A(n15988), .ZN(n15989) );
  OAI211_X1 U19370 ( .C1(n15991), .C2(n19650), .A(n15990), .B(n15989), .ZN(
        n15992) );
  AOI21_X1 U19371 ( .B1(n15993), .B2(n19663), .A(n15992), .ZN(n15994) );
  INV_X1 U19372 ( .A(n15994), .ZN(P2_U3041) );
  OAI211_X1 U19373 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15995), .B(n19670), .ZN(n15998) );
  AOI22_X1 U19374 ( .A1(n16717), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19663), .B2(n15996), .ZN(n15997) );
  AND2_X1 U19375 ( .A1(n15998), .A2(n15997), .ZN(n16005) );
  AOI21_X1 U19376 ( .B1(n19645), .B2(n20286), .A(n15999), .ZN(n16004) );
  NAND2_X1 U19377 ( .A1(n19660), .A2(n16000), .ZN(n16003) );
  NAND2_X1 U19378 ( .A1(n19669), .A2(n16001), .ZN(n16002) );
  NAND4_X1 U19379 ( .A1(n16005), .A2(n16004), .A3(n16003), .A4(n16002), .ZN(
        P2_U3045) );
  INV_X1 U19380 ( .A(n16006), .ZN(n19451) );
  AOI22_X1 U19381 ( .A1(n19410), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19451), .B2(n10049), .ZN(n16012) );
  NAND2_X1 U19382 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16012), .ZN(n16009) );
  NAND2_X1 U19383 ( .A1(n16007), .A2(n20262), .ZN(n16008) );
  OAI211_X1 U19384 ( .C1(n16010), .C2(n16730), .A(n16009), .B(n16008), .ZN(
        n16011) );
  MUX2_X1 U19385 ( .A(n16011), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n16025), .Z(P2_U3601) );
  NOR2_X1 U19386 ( .A1(n16012), .A2(n10591), .ZN(n16018) );
  INV_X1 U19387 ( .A(n16018), .ZN(n16016) );
  OAI21_X1 U19388 ( .B1(n10049), .B2(n16014), .A(n16013), .ZN(n16019) );
  OAI222_X1 U19389 ( .A1(n16730), .A2(n20281), .B1(n16016), .B2(n16019), .C1(
        n16023), .C2(n16015), .ZN(n16017) );
  MUX2_X1 U19390 ( .A(n16017), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16025), .Z(P2_U3600) );
  AOI22_X1 U19391 ( .A1(n16020), .A2(n20262), .B1(n16019), .B2(n16018), .ZN(
        n16021) );
  OAI21_X1 U19392 ( .B1(n20271), .B2(n16730), .A(n16021), .ZN(n16022) );
  MUX2_X1 U19393 ( .A(n16022), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16025), .Z(P2_U3599) );
  OAI22_X1 U19394 ( .A1(n20264), .A2(n16730), .B1(n16024), .B2(n16023), .ZN(
        n16026) );
  MUX2_X1 U19395 ( .A(n16026), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16025), .Z(P2_U3596) );
  NAND2_X1 U19396 ( .A1(n20048), .A2(n20071), .ZN(n20166) );
  NAND2_X1 U19397 ( .A1(n19931), .A2(n19745), .ZN(n19739) );
  OAI21_X1 U19398 ( .B1(n20173), .B2(n19731), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16027) );
  NAND2_X1 U19399 ( .A1(n16027), .A2(n20259), .ZN(n16034) );
  INV_X1 U19400 ( .A(n16034), .ZN(n16030) );
  NAND2_X1 U19401 ( .A1(n21171), .A2(n20278), .ZN(n19771) );
  OR2_X1 U19402 ( .A1(n19771), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19713) );
  NOR2_X1 U19403 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19713), .ZN(
        n19697) );
  INV_X1 U19404 ( .A(n19697), .ZN(n16044) );
  AND2_X1 U19405 ( .A1(n20122), .A2(n16044), .ZN(n16033) );
  AOI211_X1 U19406 ( .C1(n16028), .C2(n19936), .A(n19697), .B(n20259), .ZN(
        n16029) );
  OAI22_X1 U19407 ( .A1(n20135), .A2(n19739), .B1(n19718), .B2(n16044), .ZN(
        n16031) );
  AOI21_X1 U19408 ( .B1(n20173), .B2(n20132), .A(n16031), .ZN(n16036) );
  OAI21_X1 U19409 ( .B1(n16028), .B2(n19697), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16032) );
  NAND2_X1 U19410 ( .A1(n19703), .A2(n14194), .ZN(n16035) );
  OAI211_X1 U19411 ( .C1(n19707), .C2(n16037), .A(n16036), .B(n16035), .ZN(
        P2_U3049) );
  AOI22_X1 U19412 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19693), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19694), .ZN(n20153) );
  INV_X1 U19413 ( .A(n20153), .ZN(n20098) );
  AOI22_X1 U19414 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19693), .ZN(n19951) );
  NAND2_X1 U19415 ( .A1(n16038), .A2(n19686), .ZN(n19725) );
  OAI22_X1 U19416 ( .A1(n19951), .A2(n19739), .B1(n19725), .B2(n16044), .ZN(
        n16039) );
  AOI21_X1 U19417 ( .B1(n20173), .B2(n20098), .A(n16039), .ZN(n16041) );
  INV_X1 U19418 ( .A(n16552), .ZN(n19509) );
  NOR2_X2 U19419 ( .A1(n19509), .A2(n19874), .ZN(n20149) );
  NAND2_X1 U19420 ( .A1(n19703), .A2(n20149), .ZN(n16040) );
  OAI211_X1 U19421 ( .C1(n19707), .C2(n16042), .A(n16041), .B(n16040), .ZN(
        P2_U3052) );
  INV_X1 U19422 ( .A(n19703), .ZN(n16050) );
  NOR2_X2 U19423 ( .A1(n19488), .A2(n19874), .ZN(n20161) );
  INV_X1 U19424 ( .A(n20161), .ZN(n16049) );
  INV_X1 U19425 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18578) );
  OAI22_X2 U19426 ( .A1(n16812), .A2(n19701), .B1(n18578), .B2(n19699), .ZN(
        n20162) );
  NAND2_X1 U19427 ( .A1(n13113), .A2(n19686), .ZN(n19730) );
  INV_X1 U19428 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18581) );
  NAND2_X1 U19429 ( .A1(n20105), .A2(n19731), .ZN(n16043) );
  OAI21_X1 U19430 ( .B1(n16044), .B2(n19730), .A(n16043), .ZN(n16047) );
  NOR2_X1 U19431 ( .A1(n19707), .A2(n16045), .ZN(n16046) );
  AOI211_X1 U19432 ( .C1(n20173), .C2(n20162), .A(n16047), .B(n16046), .ZN(
        n16048) );
  OAI21_X1 U19433 ( .B1(n16050), .B2(n16049), .A(n16048), .ZN(P2_U3054) );
  OAI21_X1 U19434 ( .B1(n19801), .B2(n19830), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16053) );
  INV_X1 U19435 ( .A(n16051), .ZN(n16052) );
  NOR2_X1 U19436 ( .A1(n16052), .A2(n20075), .ZN(n20009) );
  NAND2_X1 U19437 ( .A1(n20009), .A2(n21171), .ZN(n16062) );
  NAND2_X1 U19438 ( .A1(n16053), .A2(n16062), .ZN(n16054) );
  AND2_X1 U19439 ( .A1(n20125), .A2(n16054), .ZN(n16059) );
  NAND2_X1 U19440 ( .A1(n16055), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16056) );
  NAND2_X1 U19441 ( .A1(n16056), .A2(n19936), .ZN(n16057) );
  NOR3_X1 U19442 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19869), .ZN(n19812) );
  INV_X1 U19443 ( .A(n19812), .ZN(n16071) );
  NAND2_X1 U19444 ( .A1(n16057), .A2(n16071), .ZN(n16058) );
  OAI21_X1 U19445 ( .B1(n16060), .B2(n19812), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16061) );
  OAI21_X1 U19446 ( .B1(n16062), .B2(n20261), .A(n16061), .ZN(n19813) );
  AOI22_X1 U19447 ( .A1(n19830), .A2(n20127), .B1(n19801), .B2(n20080), .ZN(
        n16063) );
  OAI21_X1 U19448 ( .B1(n19678), .B2(n16071), .A(n16063), .ZN(n16064) );
  AOI21_X1 U19449 ( .B1(n19813), .B2(n14145), .A(n16064), .ZN(n16065) );
  OAI21_X1 U19450 ( .B1(n19805), .B2(n16066), .A(n16065), .ZN(P2_U3080) );
  AOI22_X1 U19451 ( .A1(n19801), .A2(n20132), .B1(n19830), .B2(n20089), .ZN(
        n16067) );
  OAI21_X1 U19452 ( .B1(n19718), .B2(n16071), .A(n16067), .ZN(n16068) );
  AOI21_X1 U19453 ( .B1(n19813), .B2(n14194), .A(n16068), .ZN(n16069) );
  OAI21_X1 U19454 ( .B1(n19805), .B2(n9985), .A(n16069), .ZN(P2_U3081) );
  AOI22_X1 U19455 ( .A1(n19801), .A2(n20162), .B1(n19830), .B2(n20105), .ZN(
        n16070) );
  OAI21_X1 U19456 ( .B1(n19730), .B2(n16071), .A(n16070), .ZN(n16072) );
  AOI21_X1 U19457 ( .B1(n19813), .B2(n20161), .A(n16072), .ZN(n16073) );
  OAI21_X1 U19458 ( .B1(n19805), .B2(n16074), .A(n16073), .ZN(P2_U3086) );
  NOR2_X1 U19459 ( .A1(n20039), .A2(n16081), .ZN(n19957) );
  AOI21_X1 U19460 ( .B1(n20001), .B2(n19982), .A(n21288), .ZN(n16075) );
  OAI21_X1 U19461 ( .B1(n19957), .B2(n16075), .A(n19936), .ZN(n16076) );
  AOI21_X1 U19462 ( .B1(n16078), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n16076), 
        .ZN(n16077) );
  NOR2_X1 U19463 ( .A1(n20077), .A2(n16081), .ZN(n19977) );
  OAI21_X1 U19464 ( .B1(n16077), .B2(n19977), .A(n20125), .ZN(n19979) );
  INV_X1 U19465 ( .A(n19979), .ZN(n16087) );
  INV_X1 U19466 ( .A(n19742), .ZN(n19838) );
  INV_X1 U19467 ( .A(n16078), .ZN(n16079) );
  OAI21_X1 U19468 ( .B1(n16079), .B2(n19977), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16080) );
  OAI21_X1 U19469 ( .B1(n16081), .B2(n19838), .A(n16080), .ZN(n19978) );
  INV_X1 U19470 ( .A(n19977), .ZN(n16083) );
  AOI22_X1 U19471 ( .A1(n19992), .A2(n20127), .B1(n19974), .B2(n20080), .ZN(
        n16082) );
  OAI21_X1 U19472 ( .B1(n19678), .B2(n16083), .A(n16082), .ZN(n16084) );
  AOI21_X1 U19473 ( .B1(n19978), .B2(n14145), .A(n16084), .ZN(n16085) );
  OAI21_X1 U19474 ( .B1(n16087), .B2(n16086), .A(n16085), .ZN(P2_U3128) );
  OAI21_X1 U19475 ( .B1(n17296), .B2(n16089), .A(n16088), .ZN(n17592) );
  NOR3_X1 U19476 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17300), .A3(n17301), .ZN(
        n16090) );
  AOI21_X1 U19477 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16091), .A(n16090), .ZN(
        n16092) );
  OAI21_X1 U19478 ( .B1(n17592), .B2(n17556), .A(n16092), .ZN(P3_U2675) );
  INV_X1 U19479 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U19480 ( .B1(n19228), .B2(n19179), .A(n19169), .ZN(n19212) );
  NOR2_X1 U19481 ( .A1(n19179), .A2(n16911), .ZN(n18031) );
  NOR2_X1 U19482 ( .A1(n19212), .A2(n18031), .ZN(n16097) );
  NOR2_X1 U19483 ( .A1(n19169), .A2(n19042), .ZN(n18542) );
  NAND2_X1 U19484 ( .A1(n16093), .A2(n10310), .ZN(n18534) );
  NOR2_X1 U19485 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18534), .ZN(n16094) );
  NOR2_X1 U19486 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19221) );
  AOI21_X1 U19487 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n19221), .ZN(n19077) );
  OR2_X1 U19488 ( .A1(n19193), .A2(n19077), .ZN(n18545) );
  OAI21_X1 U19489 ( .B1(n16094), .B2(n19167), .A(n18657), .ZN(n18540) );
  OAI21_X1 U19490 ( .B1(n16097), .B2(n18542), .A(n18540), .ZN(n16098) );
  NOR2_X1 U19491 ( .A1(n19169), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18595) );
  INV_X1 U19492 ( .A(n18595), .ZN(n18728) );
  NAND2_X1 U19493 ( .A1(n18728), .A2(n18540), .ZN(n16096) );
  NAND2_X1 U19494 ( .A1(n19228), .A2(n19169), .ZN(n16908) );
  NOR2_X1 U19495 ( .A1(n16911), .A2(n16908), .ZN(n18913) );
  OAI21_X1 U19496 ( .B1(n16096), .B2(n18913), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16095) );
  OAI21_X1 U19497 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16098), .A(
        n16095), .ZN(P3_U2864) );
  NOR2_X1 U19498 ( .A1(n19044), .A2(n19049), .ZN(n18726) );
  INV_X1 U19499 ( .A(n18726), .ZN(n18541) );
  AOI221_X1 U19500 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18541), .C1(n16097), 
        .C2(n18541), .A(n16096), .ZN(n18539) );
  INV_X1 U19501 ( .A(n16098), .ZN(n16099) );
  AOI22_X1 U19502 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16099), .B1(
        n18913), .B2(n18540), .ZN(n18538) );
  AOI22_X1 U19503 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18539), .B1(
        n18538), .B2(n19049), .ZN(P3_U2865) );
  NAND2_X1 U19504 ( .A1(n16189), .A2(n16190), .ZN(n16102) );
  INV_X1 U19505 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16783) );
  INV_X1 U19506 ( .A(n18521), .ZN(n18526) );
  NOR2_X1 U19507 ( .A1(n16784), .A2(n16783), .ZN(n16760) );
  INV_X1 U19508 ( .A(n16760), .ZN(n16765) );
  NAND2_X1 U19509 ( .A1(n18267), .A2(n18512), .ZN(n18373) );
  INV_X1 U19510 ( .A(n18373), .ZN(n18442) );
  NAND2_X1 U19511 ( .A1(n16758), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16764) );
  AOI22_X1 U19512 ( .A1(n18526), .A2(n16765), .B1(n18442), .B2(n16764), .ZN(
        n16193) );
  NAND2_X1 U19513 ( .A1(n18512), .A2(n16192), .ZN(n16106) );
  NOR2_X1 U19514 ( .A1(n18530), .A2(n18335), .ZN(n18518) );
  INV_X1 U19515 ( .A(n18518), .ZN(n16795) );
  NAND2_X1 U19516 ( .A1(n18513), .A2(n16795), .ZN(n18482) );
  OAI21_X1 U19517 ( .B1(n16104), .B2(n17849), .A(n18482), .ZN(n16105) );
  NAND3_X1 U19518 ( .A1(n16193), .A2(n16106), .A3(n16105), .ZN(n16109) );
  AOI22_X1 U19519 ( .A1(n18267), .A2(n17840), .B1(n18999), .B2(n18211), .ZN(
        n16108) );
  NAND2_X1 U19520 ( .A1(n18203), .A2(n18245), .ZN(n18227) );
  NAND2_X1 U19521 ( .A1(n18203), .A2(n18242), .ZN(n18209) );
  OAI22_X1 U19522 ( .A1(n19031), .A2(n18227), .B1(n18496), .B2(n18209), .ZN(
        n18231) );
  NAND2_X1 U19523 ( .A1(n18205), .A2(n18231), .ZN(n16796) );
  INV_X1 U19524 ( .A(n16775), .ZN(n16107) );
  AOI211_X1 U19525 ( .C1(n16108), .C2(n16796), .A(n18530), .B(n16107), .ZN(
        n16195) );
  AOI22_X1 U19526 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16109), .B1(
        n16195), .B2(n16783), .ZN(n16110) );
  INV_X2 U19527 ( .A(n18529), .ZN(n18523) );
  NAND2_X1 U19528 ( .A1(n18523), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16792) );
  OAI211_X1 U19529 ( .C1(n16779), .C2(n18325), .A(n16110), .B(n16792), .ZN(
        P3_U2833) );
  AOI21_X1 U19530 ( .B1(n16644), .B2(n16111), .A(n9812), .ZN(n19462) );
  AOI22_X1 U19531 ( .A1(n19462), .A2(n19645), .B1(n19669), .B2(n19303), .ZN(
        n16128) );
  AND2_X1 U19532 ( .A1(n19650), .A2(n16112), .ZN(n16113) );
  OR2_X1 U19533 ( .A1(n16567), .A2(n16113), .ZN(n16120) );
  NAND2_X1 U19534 ( .A1(n16115), .A2(n16114), .ZN(n16116) );
  NAND2_X1 U19535 ( .A1(n16682), .A2(n16116), .ZN(n16649) );
  NOR2_X1 U19536 ( .A1(n16117), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16118) );
  NOR2_X1 U19537 ( .A1(n16649), .A2(n16118), .ZN(n16119) );
  NAND2_X1 U19538 ( .A1(n16120), .A2(n16119), .ZN(n16141) );
  NAND2_X1 U19539 ( .A1(n16122), .A2(n16121), .ZN(n16123) );
  AND2_X1 U19540 ( .A1(n16124), .A2(n16123), .ZN(n16566) );
  AOI22_X1 U19541 ( .A1(n16141), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19663), .B2(n16566), .ZN(n16127) );
  OAI21_X1 U19542 ( .B1(n19650), .B2(n16583), .A(n16646), .ZN(n16147) );
  NAND3_X1 U19543 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16125), .A3(
        n16147), .ZN(n16126) );
  NAND2_X1 U19544 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19643), .ZN(n16571) );
  NAND4_X1 U19545 ( .A1(n16128), .A2(n16127), .A3(n16126), .A4(n16571), .ZN(
        P2_U3030) );
  AOI22_X1 U19546 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19431), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19454), .ZN(n16140) );
  INV_X1 U19547 ( .A(n16129), .ZN(n16130) );
  AOI22_X1 U19548 ( .A1(n16130), .A2(n19422), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19444), .ZN(n16139) );
  INV_X1 U19549 ( .A(n16131), .ZN(n16132) );
  AOI22_X1 U19550 ( .A1(n16132), .A2(n19449), .B1(n16547), .B2(n19379), .ZN(
        n16138) );
  AOI21_X1 U19551 ( .B1(n16135), .B2(n16134), .A(n16133), .ZN(n16136) );
  NAND2_X1 U19552 ( .A1(n19416), .A2(n16136), .ZN(n16137) );
  NAND4_X1 U19553 ( .A1(n16140), .A2(n16139), .A3(n16138), .A4(n16137), .ZN(
        P2_U2833) );
  OAI22_X1 U19554 ( .A1(n16143), .A2(n16142), .B1(n19288), .B2(n19667), .ZN(
        n16144) );
  INV_X1 U19555 ( .A(n16146), .ZN(n16149) );
  INV_X1 U19556 ( .A(n16151), .ZN(n16162) );
  INV_X1 U19557 ( .A(n16152), .ZN(n16153) );
  AOI211_X1 U19558 ( .C1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16154), .A(
        n20905), .B(n16153), .ZN(n16158) );
  INV_X1 U19559 ( .A(n16158), .ZN(n16160) );
  INV_X1 U19560 ( .A(n16155), .ZN(n16156) );
  OAI22_X1 U19561 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16158), .B1(
        n16157), .B2(n16156), .ZN(n16159) );
  OAI21_X1 U19562 ( .B1(n16160), .B2(n20870), .A(n16159), .ZN(n16161) );
  AOI222_X1 U19563 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16162), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16161), .C1(n16162), 
        .C2(n16161), .ZN(n16163) );
  AOI222_X1 U19564 ( .A1(n16164), .A2(n16163), .B1(n16164), .B2(n20740), .C1(
        n16163), .C2(n20740), .ZN(n16165) );
  NOR2_X1 U19565 ( .A1(n16165), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16172) );
  NOR2_X1 U19566 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n16167) );
  OAI21_X1 U19567 ( .B1(n16168), .B2(n16167), .A(n16166), .ZN(n16169) );
  NOR4_X1 U19568 ( .A1(n16172), .A2(n16171), .A3(n16170), .A4(n16169), .ZN(
        n16180) );
  AOI21_X1 U19569 ( .B1(n16174), .B2(n20985), .A(n16173), .ZN(n16175) );
  AOI21_X1 U19570 ( .B1(n16177), .B2(n16176), .A(n16175), .ZN(n16479) );
  OAI221_X1 U19571 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16180), 
        .A(n16479), .ZN(n16476) );
  OAI21_X1 U19572 ( .B1(n16180), .B2(n16179), .A(n16178), .ZN(n16181) );
  AOI211_X1 U19573 ( .C1(n20985), .C2(n20913), .A(n16182), .B(n16181), .ZN(
        n16187) );
  NAND2_X1 U19574 ( .A1(n16184), .A2(n16183), .ZN(n16185) );
  AOI21_X1 U19575 ( .B1(n16185), .B2(n16476), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n16186) );
  AOI21_X1 U19576 ( .B1(n16476), .B2(n16187), .A(n16186), .ZN(P1_U3161) );
  INV_X1 U19577 ( .A(n16746), .ZN(n16743) );
  NAND3_X1 U19578 ( .A1(n16190), .A2(n16189), .A3(n16783), .ZN(n16742) );
  NAND2_X1 U19579 ( .A1(n16743), .A2(n16742), .ZN(n16191) );
  INV_X1 U19580 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16798) );
  XOR2_X1 U19581 ( .A(n16191), .B(n16798), .Z(n16778) );
  NOR2_X1 U19582 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16783), .ZN(
        n16774) );
  NAND3_X1 U19583 ( .A1(n16775), .A2(n18512), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16797) );
  AOI22_X1 U19584 ( .A1(n18512), .A2(n16192), .B1(n18482), .B2(n16797), .ZN(
        n16794) );
  AOI21_X1 U19585 ( .B1(n16794), .B2(n16193), .A(n16798), .ZN(n16194) );
  AOI21_X1 U19586 ( .B1(n16774), .B2(n16195), .A(n16194), .ZN(n16196) );
  NAND2_X1 U19587 ( .A1(n18523), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16766) );
  OAI211_X1 U19588 ( .C1(n16778), .C2(n18325), .A(n16196), .B(n16766), .ZN(
        P3_U2832) );
  INV_X1 U19589 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20998) );
  NAND2_X1 U19590 ( .A1(n20998), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20317) );
  INV_X1 U19591 ( .A(HOLD), .ZN(n20981) );
  INV_X1 U19592 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20991) );
  NOR2_X1 U19593 ( .A1(n20992), .A2(n20991), .ZN(n20988) );
  AOI221_X1 U19594 ( .B1(n20998), .B2(n20988), .C1(n20981), .C2(n20988), .A(
        n16197), .ZN(n16198) );
  NAND2_X1 U19595 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20985), .ZN(n20996) );
  OAI211_X1 U19596 ( .C1(n20317), .C2(n20981), .A(n16198), .B(n20996), .ZN(
        P1_U3195) );
  INV_X1 U19597 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16810) );
  NOR2_X1 U19598 ( .A1(n20412), .A2(n16810), .ZN(P1_U2905) );
  NOR3_X1 U19599 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n21192), .A3(n20183), 
        .ZN(n16728) );
  INV_X1 U19600 ( .A(n16201), .ZN(n16729) );
  NOR4_X1 U19601 ( .A1(n16200), .A2(n16199), .A3(n16728), .A4(n16729), .ZN(
        P2_U3178) );
  OAI221_X1 U19602 ( .B1(n16202), .B2(n16201), .C1(n20302), .C2(n16201), .A(
        n19874), .ZN(n20296) );
  NOR2_X1 U19603 ( .A1(n16203), .A2(n20296), .ZN(P2_U3047) );
  INV_X1 U19604 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n21110) );
  NOR3_X1 U19605 ( .A1(n19215), .A2(n17206), .A3(n16204), .ZN(n16205) );
  INV_X1 U19606 ( .A(n16208), .ZN(n16207) );
  INV_X1 U19607 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21141) );
  AOI21_X1 U19608 ( .B1(n18589), .B2(n16207), .A(P3_EAX_REG_0__SCAN_IN), .ZN(
        n16210) );
  OAI222_X1 U19609 ( .A1(n21110), .A2(n17714), .B1(n17720), .B2(n16210), .C1(
        n17711), .C2(n18187), .ZN(P3_U2735) );
  NOR3_X1 U19610 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15083), .A3(n16225), 
        .ZN(n16213) );
  OAI22_X1 U19611 ( .A1(n12789), .A2(n20389), .B1(n16211), .B2(n21398), .ZN(
        n16212) );
  AOI211_X1 U19612 ( .C1(n20353), .C2(P1_EBX_REG_22__SCAN_IN), .A(n16213), .B(
        n16212), .ZN(n16218) );
  OAI21_X1 U19613 ( .B1(n16225), .B2(P1_REIP_REG_21__SCAN_IN), .A(n16214), 
        .ZN(n16215) );
  AOI22_X1 U19614 ( .A1(n16216), .A2(n20368), .B1(P1_REIP_REG_22__SCAN_IN), 
        .B2(n16215), .ZN(n16217) );
  OAI211_X1 U19615 ( .C1(n21390), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        P1_U2818) );
  AOI22_X1 U19616 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n21395), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(n20353), .ZN(n16229) );
  AOI22_X1 U19617 ( .A1(n16221), .A2(n20341), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n16220), .ZN(n16228) );
  NOR2_X1 U19618 ( .A1(n16222), .A2(n21390), .ZN(n16223) );
  AOI21_X1 U19619 ( .B1(n16224), .B2(n20368), .A(n16223), .ZN(n16227) );
  OR2_X1 U19620 ( .A1(n16225), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16226) );
  NAND4_X1 U19621 ( .A1(n16229), .A2(n16228), .A3(n16227), .A4(n16226), .ZN(
        P1_U2819) );
  INV_X1 U19622 ( .A(n16239), .ZN(n16230) );
  NOR3_X1 U19623 ( .A1(n16230), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n16238), 
        .ZN(n16235) );
  AOI22_X1 U19624 ( .A1(n16231), .A2(n20341), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n20378), .ZN(n16232) );
  OAI211_X1 U19625 ( .C1(n16233), .C2(n20389), .A(n16232), .B(n20379), .ZN(
        n16234) );
  AOI211_X1 U19626 ( .C1(n16236), .C2(n20368), .A(n16235), .B(n16234), .ZN(
        n16241) );
  NOR2_X1 U19627 ( .A1(n16281), .A2(n16237), .ZN(n16256) );
  AND2_X1 U19628 ( .A1(n16239), .A2(n16238), .ZN(n16247) );
  OAI21_X1 U19629 ( .B1(n16256), .B2(n16247), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n16240) );
  OAI211_X1 U19630 ( .C1(n16242), .C2(n21390), .A(n16241), .B(n16240), .ZN(
        P1_U2821) );
  AOI22_X1 U19631 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n20378), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n16256), .ZN(n16244) );
  AOI21_X1 U19632 ( .B1(n21395), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21393), .ZN(n16243) );
  OAI211_X1 U19633 ( .C1(n16245), .C2(n21398), .A(n16244), .B(n16243), .ZN(
        n16246) );
  AOI211_X1 U19634 ( .C1(n16248), .C2(n20368), .A(n16247), .B(n16246), .ZN(
        n16249) );
  OAI21_X1 U19635 ( .B1(n21390), .B2(n16250), .A(n16249), .ZN(P1_U2822) );
  AOI22_X1 U19636 ( .A1(n16251), .A2(n20341), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n20353), .ZN(n16252) );
  OAI211_X1 U19637 ( .C1(n16253), .C2(n20389), .A(n16252), .B(n20379), .ZN(
        n16254) );
  AOI21_X1 U19638 ( .B1(n16255), .B2(n20368), .A(n16254), .ZN(n16259) );
  OAI21_X1 U19639 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n16257), .A(n16256), 
        .ZN(n16258) );
  OAI211_X1 U19640 ( .C1(n16260), .C2(n21390), .A(n16259), .B(n16258), .ZN(
        P1_U2823) );
  OAI21_X1 U19641 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n16261), .ZN(n16264) );
  AND2_X1 U19642 ( .A1(n20356), .A2(n16262), .ZN(n21400) );
  AOI22_X1 U19643 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20378), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21400), .ZN(n16263) );
  OAI21_X1 U19644 ( .B1(n16273), .B2(n16264), .A(n16263), .ZN(n16265) );
  AOI211_X1 U19645 ( .C1(n21395), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21393), .B(n16265), .ZN(n16268) );
  AOI22_X1 U19646 ( .A1(n16316), .A2(n20368), .B1(n16266), .B2(n20341), .ZN(
        n16267) );
  OAI211_X1 U19647 ( .C1(n21390), .C2(n16370), .A(n16268), .B(n16267), .ZN(
        P1_U2824) );
  OAI21_X1 U19648 ( .B1(n16271), .B2(n16270), .A(n16269), .ZN(n16272) );
  INV_X1 U19649 ( .A(n16272), .ZN(n16381) );
  INV_X1 U19650 ( .A(n16273), .ZN(n16274) );
  INV_X1 U19651 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21016) );
  AOI22_X1 U19652 ( .A1(n20377), .A2(n16381), .B1(n16274), .B2(n21016), .ZN(
        n16280) );
  OAI22_X1 U19653 ( .A1(n16275), .A2(n20389), .B1(n16308), .B2(n21391), .ZN(
        n16276) );
  AOI211_X1 U19654 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n21400), .A(n21393), 
        .B(n16276), .ZN(n16279) );
  INV_X1 U19655 ( .A(n16277), .ZN(n16324) );
  AOI22_X1 U19656 ( .A1(n16325), .A2(n20368), .B1(n20341), .B2(n16324), .ZN(
        n16278) );
  NAND3_X1 U19657 ( .A1(n16280), .A2(n16279), .A3(n16278), .ZN(P1_U2825) );
  NAND3_X1 U19658 ( .A1(n16304), .A2(P1_REIP_REG_12__SCAN_IN), .A3(
        P1_REIP_REG_11__SCAN_IN), .ZN(n21386) );
  NOR2_X1 U19659 ( .A1(n16412), .A2(n16303), .ZN(n16283) );
  AOI21_X1 U19660 ( .B1(n16283), .B2(n16282), .A(n16281), .ZN(n16294) );
  AOI22_X1 U19661 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20353), .B1(n20377), 
        .B2(n16405), .ZN(n16284) );
  OAI211_X1 U19662 ( .C1(n20389), .C2(n16285), .A(n16284), .B(n20379), .ZN(
        n16286) );
  AOI21_X1 U19663 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n16294), .A(n16286), 
        .ZN(n16291) );
  OAI22_X1 U19664 ( .A1(n16288), .A2(n21403), .B1(n16287), .B2(n21398), .ZN(
        n16289) );
  INV_X1 U19665 ( .A(n16289), .ZN(n16290) );
  OAI211_X1 U19666 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n21386), .A(n16291), 
        .B(n16290), .ZN(P1_U2827) );
  OAI22_X1 U19667 ( .A1(n16292), .A2(n21391), .B1(n21390), .B2(n16415), .ZN(
        n16293) );
  AOI211_X1 U19668 ( .C1(n21395), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21393), .B(n16293), .ZN(n16298) );
  AOI22_X1 U19669 ( .A1(n16343), .A2(n20368), .B1(n20341), .B2(n16341), .ZN(
        n16297) );
  AND2_X1 U19670 ( .A1(n16304), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16295) );
  OAI21_X1 U19671 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n16295), .A(n16294), 
        .ZN(n16296) );
  NAND3_X1 U19672 ( .A1(n16298), .A2(n16297), .A3(n16296), .ZN(P1_U2828) );
  INV_X1 U19673 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16300) );
  AOI22_X1 U19674 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n20378), .B1(n20377), 
        .B2(n16426), .ZN(n16299) );
  OAI211_X1 U19675 ( .C1(n20389), .C2(n16300), .A(n16299), .B(n20379), .ZN(
        n16301) );
  AOI221_X1 U19676 ( .B1(n16304), .B2(n16303), .C1(n16302), .C2(
        P1_REIP_REG_11__SCAN_IN), .A(n16301), .ZN(n16306) );
  NAND2_X1 U19677 ( .A1(n16352), .A2(n20368), .ZN(n16305) );
  OAI211_X1 U19678 ( .C1(n21398), .C2(n16355), .A(n16306), .B(n16305), .ZN(
        P1_U2829) );
  AOI22_X1 U19679 ( .A1(n16325), .A2(n20405), .B1(n20404), .B2(n16381), .ZN(
        n16307) );
  OAI21_X1 U19680 ( .B1(n20408), .B2(n16308), .A(n16307), .ZN(P1_U2857) );
  AOI22_X1 U19681 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16318) );
  INV_X1 U19682 ( .A(n16309), .ZN(n16311) );
  AOI211_X1 U19683 ( .C1(n16348), .C2(n16311), .A(n16310), .B(n16329), .ZN(
        n16322) );
  INV_X1 U19684 ( .A(n16314), .ZN(n16312) );
  NOR2_X1 U19685 ( .A1(n16313), .A2(n16312), .ZN(n16321) );
  NAND2_X1 U19686 ( .A1(n16322), .A2(n16321), .ZN(n16320) );
  NAND2_X1 U19687 ( .A1(n16320), .A2(n16314), .ZN(n16315) );
  AOI22_X1 U19688 ( .A1(n16371), .A2(n12479), .B1(n20477), .B2(n16316), .ZN(
        n16317) );
  OAI211_X1 U19689 ( .C1(n20482), .C2(n16319), .A(n16318), .B(n16317), .ZN(
        P1_U2983) );
  OAI21_X1 U19690 ( .B1(n16322), .B2(n16321), .A(n16320), .ZN(n16323) );
  INV_X1 U19691 ( .A(n16323), .ZN(n16383) );
  AOI22_X1 U19692 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16327) );
  AOI22_X1 U19693 ( .A1(n16325), .A2(n20477), .B1(n16342), .B2(n16324), .ZN(
        n16326) );
  OAI211_X1 U19694 ( .C1(n16383), .C2(n20321), .A(n16327), .B(n16326), .ZN(
        P1_U2984) );
  OAI21_X1 U19695 ( .B1(n16348), .B2(n16329), .A(n16328), .ZN(n16331) );
  NAND2_X1 U19696 ( .A1(n16331), .A2(n16330), .ZN(n16333) );
  MUX2_X1 U19697 ( .A(n12374), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n12230), .Z(n16332) );
  XNOR2_X1 U19698 ( .A(n16333), .B(n16332), .ZN(n16391) );
  AOI22_X1 U19699 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16336) );
  AOI22_X1 U19700 ( .A1(n16334), .A2(n20477), .B1(n16342), .B2(n21388), .ZN(
        n16335) );
  OAI211_X1 U19701 ( .C1(n16391), .C2(n20321), .A(n16336), .B(n16335), .ZN(
        P1_U2985) );
  OAI21_X1 U19702 ( .B1(n16339), .B2(n16338), .A(n16337), .ZN(n16340) );
  INV_X1 U19703 ( .A(n16340), .ZN(n16425) );
  AOI22_X1 U19704 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16345) );
  AOI22_X1 U19705 ( .A1(n16343), .A2(n20477), .B1(n16342), .B2(n16341), .ZN(
        n16344) );
  OAI211_X1 U19706 ( .C1(n16425), .C2(n20321), .A(n16345), .B(n16344), .ZN(
        P1_U2987) );
  AOI22_X1 U19707 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16354) );
  NAND2_X1 U19708 ( .A1(n16347), .A2(n16346), .ZN(n16350) );
  NAND2_X1 U19709 ( .A1(n16348), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16349) );
  MUX2_X1 U19710 ( .A(n16350), .B(n16349), .S(n12230), .Z(n16351) );
  XNOR2_X1 U19711 ( .A(n16351), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16427) );
  AOI22_X1 U19712 ( .A1(n16427), .A2(n12479), .B1(n20477), .B2(n16352), .ZN(
        n16353) );
  OAI211_X1 U19713 ( .C1(n20482), .C2(n16355), .A(n16354), .B(n16353), .ZN(
        P1_U2988) );
  AOI22_X1 U19714 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16361) );
  NAND2_X1 U19715 ( .A1(n9813), .A2(n16356), .ZN(n16357) );
  XNOR2_X1 U19716 ( .A(n16358), .B(n16357), .ZN(n16455) );
  INV_X1 U19717 ( .A(n16359), .ZN(n20358) );
  AOI22_X1 U19718 ( .A1(n16455), .A2(n12479), .B1(n20477), .B2(n20358), .ZN(
        n16360) );
  OAI211_X1 U19719 ( .C1(n20482), .C2(n20361), .A(n16361), .B(n16360), .ZN(
        P1_U2992) );
  AOI22_X1 U19720 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16367) );
  OAI21_X1 U19721 ( .B1(n16364), .B2(n16363), .A(n16362), .ZN(n16365) );
  INV_X1 U19722 ( .A(n16365), .ZN(n16464) );
  AOI22_X1 U19723 ( .A1(n16464), .A2(n12479), .B1(n20477), .B2(n20406), .ZN(
        n16366) );
  OAI211_X1 U19724 ( .C1(n20482), .C2(n20387), .A(n16367), .B(n16366), .ZN(
        P1_U2994) );
  OAI21_X1 U19725 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16368), .ZN(n16375) );
  INV_X1 U19726 ( .A(n16369), .ZN(n16376) );
  INV_X1 U19727 ( .A(n16370), .ZN(n16372) );
  AOI222_X1 U19728 ( .A1(n16376), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .B1(n20486), .B2(n16372), .C1(n20507), .C2(n16371), .ZN(n16374) );
  NAND2_X1 U19729 ( .A1(n20473), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16373) );
  OAI211_X1 U19730 ( .C1(n16379), .C2(n16375), .A(n16374), .B(n16373), .ZN(
        P1_U3015) );
  NAND2_X1 U19731 ( .A1(n16376), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16378) );
  NAND2_X1 U19732 ( .A1(n20473), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16377) );
  OAI211_X1 U19733 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16379), .A(
        n16378), .B(n16377), .ZN(n16380) );
  AOI21_X1 U19734 ( .B1(n16381), .B2(n20486), .A(n16380), .ZN(n16382) );
  OAI21_X1 U19735 ( .B1(n16383), .B2(n16424), .A(n16382), .ZN(P1_U3016) );
  INV_X1 U19736 ( .A(n16384), .ZN(n16389) );
  OAI22_X1 U19737 ( .A1(n16397), .A2(n16396), .B1(n16385), .B2(n16404), .ZN(
        n16388) );
  INV_X1 U19738 ( .A(n16386), .ZN(n16387) );
  AOI211_X1 U19739 ( .C1(n16389), .C2(n16399), .A(n16388), .B(n16387), .ZN(
        n16398) );
  NOR2_X1 U19740 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16390), .ZN(
        n16393) );
  OAI22_X1 U19741 ( .A1(n16391), .A2(n16424), .B1(n20504), .B2(n21389), .ZN(
        n16392) );
  AOI21_X1 U19742 ( .B1(n16393), .B2(n16419), .A(n16392), .ZN(n16395) );
  NAND2_X1 U19743 ( .A1(n20473), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16394) );
  OAI211_X1 U19744 ( .C1(n16398), .C2(n12374), .A(n16395), .B(n16394), .ZN(
        P1_U3017) );
  NOR2_X1 U19745 ( .A1(n16397), .A2(n16396), .ZN(n16403) );
  NOR2_X1 U19746 ( .A1(n12460), .A2(n21387), .ZN(n16402) );
  AOI21_X1 U19747 ( .B1(n16400), .B2(n16399), .A(n16398), .ZN(n16401) );
  AOI211_X1 U19748 ( .C1(n16404), .C2(n16403), .A(n16402), .B(n16401), .ZN(
        n16408) );
  AOI22_X1 U19749 ( .A1(n16406), .A2(n20507), .B1(n20486), .B2(n16405), .ZN(
        n16407) );
  NAND2_X1 U19750 ( .A1(n16408), .A2(n16407), .ZN(P1_U3018) );
  INV_X1 U19751 ( .A(n16409), .ZN(n16421) );
  OAI21_X1 U19752 ( .B1(n16414), .B2(n16433), .A(n16410), .ZN(n16411) );
  OAI211_X1 U19753 ( .C1(n16421), .C2(n20502), .A(n20494), .B(n16411), .ZN(
        n16428) );
  NOR2_X1 U19754 ( .A1(n12460), .A2(n16412), .ZN(n16418) );
  NAND2_X1 U19755 ( .A1(n16413), .A2(n20493), .ZN(n16416) );
  OR2_X1 U19756 ( .A1(n16414), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16431) );
  OAI22_X1 U19757 ( .A1(n16416), .A2(n16431), .B1(n20504), .B2(n16415), .ZN(
        n16417) );
  AOI211_X1 U19758 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16428), .A(
        n16418), .B(n16417), .ZN(n16423) );
  NAND3_X1 U19759 ( .A1(n16421), .A2(n16420), .A3(n16419), .ZN(n16422) );
  OAI211_X1 U19760 ( .C1(n16425), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        P1_U3019) );
  AOI22_X1 U19761 ( .A1(n16426), .A2(n20486), .B1(n20473), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16430) );
  AOI22_X1 U19762 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16428), .B1(
        n20507), .B2(n16427), .ZN(n16429) );
  OAI211_X1 U19763 ( .C1(n16432), .C2(n16431), .A(n16430), .B(n16429), .ZN(
        P1_U3020) );
  NAND3_X1 U19764 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16438) );
  INV_X1 U19765 ( .A(n16433), .ZN(n16435) );
  OAI211_X1 U19766 ( .C1(n16435), .C2(n20495), .A(n16434), .B(n20494), .ZN(
        n16437) );
  OAI21_X1 U19767 ( .B1(n16438), .B2(n16437), .A(n16436), .ZN(n16452) );
  NAND2_X1 U19768 ( .A1(n16439), .A2(n16454), .ZN(n16446) );
  AOI221_X1 U19769 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16346), .C2(n16453), .A(
        n16446), .ZN(n16443) );
  INV_X1 U19770 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16440) );
  OAI22_X1 U19771 ( .A1(n16441), .A2(n20504), .B1(n16440), .B2(n12460), .ZN(
        n16442) );
  AOI211_X1 U19772 ( .C1(n16444), .C2(n20507), .A(n16443), .B(n16442), .ZN(
        n16445) );
  OAI21_X1 U19773 ( .B1(n16346), .B2(n16452), .A(n16445), .ZN(P1_U3021) );
  NOR2_X1 U19774 ( .A1(n16446), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16449) );
  INV_X1 U19775 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21009) );
  OAI22_X1 U19776 ( .A1(n16447), .A2(n20504), .B1(n21009), .B2(n12460), .ZN(
        n16448) );
  AOI211_X1 U19777 ( .C1(n16450), .C2(n20507), .A(n16449), .B(n16448), .ZN(
        n16451) );
  OAI21_X1 U19778 ( .B1(n16453), .B2(n16452), .A(n16451), .ZN(P1_U3022) );
  AOI22_X1 U19779 ( .A1(n20352), .A2(n20486), .B1(n20473), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16457) );
  AOI22_X1 U19780 ( .A1(n16455), .A2(n20507), .B1(n16454), .B2(n16458), .ZN(
        n16456) );
  OAI211_X1 U19781 ( .C1(n16459), .C2(n16458), .A(n16457), .B(n16456), .ZN(
        P1_U3024) );
  AND2_X1 U19782 ( .A1(n16461), .A2(n16460), .ZN(n16462) );
  NOR2_X1 U19783 ( .A1(n9833), .A2(n16462), .ZN(n20403) );
  AOI22_X1 U19784 ( .A1(n20403), .A2(n20486), .B1(n20473), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19785 ( .A1(n16464), .A2(n20507), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16463), .ZN(n16468) );
  NAND3_X1 U19786 ( .A1(n16466), .A2(n20488), .A3(n16465), .ZN(n16467) );
  NAND3_X1 U19787 ( .A1(n16469), .A2(n16468), .A3(n16467), .ZN(P1_U3026) );
  NAND3_X1 U19788 ( .A1(n16472), .A2(n16471), .A3(n16470), .ZN(n16473) );
  OAI21_X1 U19789 ( .B1(n16475), .B2(n16474), .A(n16473), .ZN(P1_U3468) );
  NAND2_X1 U19790 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16476), .ZN(n16483) );
  AOI21_X1 U19791 ( .B1(n20817), .B2(n21066), .A(n21062), .ZN(n16482) );
  NAND4_X1 U19792 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n20913), .A4(n21066), .ZN(n16477) );
  AND2_X1 U19793 ( .A1(n16478), .A2(n16477), .ZN(n20977) );
  AOI21_X1 U19794 ( .B1(n20977), .B2(n16480), .A(n16479), .ZN(n16481) );
  AOI211_X1 U19795 ( .C1(n21247), .C2(n16483), .A(n16482), .B(n16481), .ZN(
        P1_U3162) );
  INV_X1 U19796 ( .A(n16483), .ZN(n16485) );
  OAI21_X1 U19797 ( .B1(n16485), .B2(n20817), .A(n16484), .ZN(P1_U3466) );
  OAI22_X1 U19798 ( .A1(n21234), .A2(n19440), .B1(n16486), .B2(n13074), .ZN(
        n16487) );
  AOI21_X1 U19799 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19454), .A(
        n16487), .ZN(n16488) );
  OAI21_X1 U19800 ( .B1(n16489), .B2(n19414), .A(n16488), .ZN(n16490) );
  AOI21_X1 U19801 ( .B1(n16491), .B2(n19422), .A(n16490), .ZN(n16495) );
  NAND4_X1 U19802 ( .A1(n19416), .A2(n16493), .A3(n16492), .A4(n10049), .ZN(
        n16494) );
  OAI211_X1 U19803 ( .C1(n15500), .C2(n19442), .A(n16495), .B(n16494), .ZN(
        P2_U2824) );
  INV_X1 U19804 ( .A(n16496), .ZN(n16498) );
  AOI22_X1 U19805 ( .A1(n16498), .A2(n19449), .B1(n16497), .B2(n19379), .ZN(
        n16508) );
  AOI211_X1 U19806 ( .C1(n16501), .C2(n16500), .A(n16499), .B(n19450), .ZN(
        n16506) );
  INV_X1 U19807 ( .A(n16502), .ZN(n16504) );
  AOI22_X1 U19808 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19444), .ZN(n16503) );
  OAI21_X1 U19809 ( .B1(n16504), .B2(n19447), .A(n16503), .ZN(n16505) );
  AOI211_X1 U19810 ( .C1(n19431), .C2(P2_REIP_REG_28__SCAN_IN), .A(n16506), 
        .B(n16505), .ZN(n16507) );
  NAND2_X1 U19811 ( .A1(n16508), .A2(n16507), .ZN(P2_U2827) );
  AOI22_X1 U19812 ( .A1(n16509), .A2(n19422), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19454), .ZN(n16519) );
  AOI22_X1 U19813 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19431), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19444), .ZN(n16518) );
  INV_X1 U19814 ( .A(n16510), .ZN(n16512) );
  AOI22_X1 U19815 ( .A1(n16512), .A2(n19449), .B1(n16511), .B2(n19379), .ZN(
        n16517) );
  AOI21_X1 U19816 ( .B1(n16514), .B2(n9804), .A(n16513), .ZN(n16515) );
  NAND2_X1 U19817 ( .A1(n19416), .A2(n16515), .ZN(n16516) );
  NAND4_X1 U19818 ( .A1(n16519), .A2(n16518), .A3(n16517), .A4(n16516), .ZN(
        P2_U2829) );
  AOI211_X1 U19819 ( .C1(n16522), .C2(n16521), .A(n16520), .B(n19450), .ZN(
        n16530) );
  OAI22_X1 U19820 ( .A1(n16523), .A2(n19420), .B1(n19440), .B2(n20238), .ZN(
        n16526) );
  NOR2_X1 U19821 ( .A1(n16524), .A2(n19414), .ZN(n16525) );
  AOI211_X1 U19822 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n19444), .A(n16526), .B(
        n16525), .ZN(n16527) );
  OAI21_X1 U19823 ( .B1(n16528), .B2(n19447), .A(n16527), .ZN(n16529) );
  AOI211_X1 U19824 ( .C1(n19379), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16532) );
  INV_X1 U19825 ( .A(n16532), .ZN(P2_U2830) );
  AOI211_X1 U19826 ( .C1(n16535), .C2(n16534), .A(n16533), .B(n19450), .ZN(
        n16539) );
  AOI22_X1 U19827 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19444), .ZN(n16536) );
  OAI21_X1 U19828 ( .B1(n16537), .B2(n19447), .A(n16536), .ZN(n16538) );
  AOI211_X1 U19829 ( .C1(n19431), .C2(P2_REIP_REG_24__SCAN_IN), .A(n16539), 
        .B(n16538), .ZN(n16545) );
  INV_X1 U19830 ( .A(n16540), .ZN(n16541) );
  OAI22_X1 U19831 ( .A1(n16542), .A2(n19414), .B1(n16541), .B2(n19442), .ZN(
        n16543) );
  INV_X1 U19832 ( .A(n16543), .ZN(n16544) );
  NAND2_X1 U19833 ( .A1(n16545), .A2(n16544), .ZN(P2_U2831) );
  AOI22_X1 U19834 ( .A1(n19459), .A2(n16546), .B1(n19522), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16551) );
  AOI22_X1 U19835 ( .A1(n19461), .A2(BUF1_REG_22__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16550) );
  AOI22_X1 U19836 ( .A1(n16548), .A2(n19505), .B1(n19523), .B2(n16547), .ZN(
        n16549) );
  NAND3_X1 U19837 ( .A1(n16551), .A2(n16550), .A3(n16549), .ZN(P2_U2897) );
  AOI22_X1 U19838 ( .A1(n19459), .A2(n16552), .B1(n19522), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16557) );
  AOI22_X1 U19839 ( .A1(n19461), .A2(BUF1_REG_20__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16556) );
  INV_X1 U19840 ( .A(n16553), .ZN(n16554) );
  AOI22_X1 U19841 ( .A1(n16554), .A2(n19505), .B1(n19523), .B2(n19259), .ZN(
        n16555) );
  NAND3_X1 U19842 ( .A1(n16557), .A2(n16556), .A3(n16555), .ZN(P2_U2899) );
  AOI22_X1 U19843 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16638), .B1(
        n19613), .B2(n16558), .ZN(n16565) );
  NAND3_X1 U19844 ( .A1(n16559), .A2(n12997), .A3(n15847), .ZN(n16560) );
  OAI21_X1 U19845 ( .B1(n14135), .B2(n16561), .A(n16560), .ZN(n16562) );
  AOI21_X1 U19846 ( .B1(n16632), .B2(n16563), .A(n16562), .ZN(n16564) );
  OAI211_X1 U19847 ( .C1(n21139), .C2(n19388), .A(n16565), .B(n16564), .ZN(
        P2_U2991) );
  AOI22_X1 U19848 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16638), .B1(
        n19613), .B2(n19299), .ZN(n16573) );
  AOI22_X1 U19849 ( .A1(n16566), .A2(n12997), .B1(n19622), .B2(n19303), .ZN(
        n16572) );
  INV_X1 U19850 ( .A(n16567), .ZN(n16569) );
  OAI211_X1 U19851 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16579), .A(
        n16569), .B(n16568), .ZN(n16570) );
  NAND4_X1 U19852 ( .A1(n16573), .A2(n16572), .A3(n16571), .A4(n16570), .ZN(
        P2_U2998) );
  AOI22_X1 U19853 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19643), .B1(n19613), 
        .B2(n19312), .ZN(n16582) );
  NAND2_X1 U19854 ( .A1(n16575), .A2(n16574), .ZN(n16578) );
  NAND2_X1 U19855 ( .A1(n16576), .A2(n16584), .ZN(n16577) );
  XOR2_X1 U19856 ( .A(n16578), .B(n16577), .Z(n16653) );
  INV_X1 U19857 ( .A(n16653), .ZN(n16580) );
  INV_X1 U19858 ( .A(n19313), .ZN(n16650) );
  OAI211_X1 U19859 ( .C1(n19318), .C2(n19642), .A(n16582), .B(n16581), .ZN(
        P2_U2999) );
  AOI22_X1 U19860 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19643), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16638), .ZN(n16590) );
  NOR2_X1 U19861 ( .A1(n16656), .A2(n16617), .ZN(n16592) );
  OAI21_X1 U19862 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16592), .A(
        n16583), .ZN(n16668) );
  NAND2_X1 U19863 ( .A1(n16585), .A2(n16584), .ZN(n16587) );
  XOR2_X1 U19864 ( .A(n16587), .B(n16586), .Z(n16664) );
  OAI22_X1 U19865 ( .A1(n16668), .A2(n19636), .B1(n16664), .B2(n19619), .ZN(
        n16588) );
  AOI21_X1 U19866 ( .B1(n19622), .B2(n19326), .A(n16588), .ZN(n16589) );
  OAI211_X1 U19867 ( .C1(n19634), .C2(n16591), .A(n16590), .B(n16589), .ZN(
        P2_U3000) );
  AOI22_X1 U19868 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19643), .B1(n19613), 
        .B2(n19335), .ZN(n16600) );
  AOI21_X1 U19869 ( .B1(n11269), .B2(n16593), .A(n16592), .ZN(n16677) );
  NAND2_X1 U19870 ( .A1(n16595), .A2(n16594), .ZN(n16596) );
  XNOR2_X1 U19871 ( .A(n16597), .B(n16596), .ZN(n16680) );
  INV_X1 U19872 ( .A(n16680), .ZN(n16598) );
  AOI222_X1 U19873 ( .A1(n16677), .A2(n16632), .B1(n12997), .B2(n16598), .C1(
        n19622), .C2(n16676), .ZN(n16599) );
  OAI211_X1 U19874 ( .C1(n21272), .C2(n19642), .A(n16600), .B(n16599), .ZN(
        P2_U3001) );
  AOI22_X1 U19875 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16638), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19643), .ZN(n16605) );
  OAI22_X1 U19876 ( .A1(n16602), .A2(n19636), .B1(n16601), .B2(n19619), .ZN(
        n16603) );
  AOI21_X1 U19877 ( .B1(n19622), .B2(n19347), .A(n16603), .ZN(n16604) );
  OAI211_X1 U19878 ( .C1(n19634), .C2(n19346), .A(n16605), .B(n16604), .ZN(
        P2_U3002) );
  AOI22_X1 U19879 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19643), .B1(n19613), 
        .B2(n16606), .ZN(n16621) );
  INV_X1 U19880 ( .A(n16607), .ZN(n16608) );
  NAND2_X1 U19881 ( .A1(n16609), .A2(n16608), .ZN(n16613) );
  OR2_X1 U19882 ( .A1(n16611), .A2(n16610), .ZN(n16612) );
  XNOR2_X1 U19883 ( .A(n16613), .B(n16612), .ZN(n16689) );
  INV_X1 U19884 ( .A(n16614), .ZN(n16688) );
  NAND2_X1 U19885 ( .A1(n16616), .A2(n16615), .ZN(n16618) );
  NAND2_X1 U19886 ( .A1(n16618), .A2(n16617), .ZN(n16692) );
  INV_X1 U19887 ( .A(n16692), .ZN(n16619) );
  AOI222_X1 U19888 ( .A1(n16689), .A2(n12997), .B1(n19622), .B2(n16688), .C1(
        n16632), .C2(n16619), .ZN(n16620) );
  OAI211_X1 U19889 ( .C1(n16622), .C2(n19642), .A(n16621), .B(n16620), .ZN(
        P2_U3003) );
  AOI22_X1 U19890 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19643), .B1(n19613), 
        .B2(n19375), .ZN(n16636) );
  XOR2_X1 U19891 ( .A(n16623), .B(n16624), .Z(n16708) );
  AOI21_X1 U19892 ( .B1(n15753), .B2(n16626), .A(n16625), .ZN(n16631) );
  INV_X1 U19893 ( .A(n16627), .ZN(n16628) );
  NOR2_X1 U19894 ( .A1(n16629), .A2(n16628), .ZN(n16630) );
  XNOR2_X1 U19895 ( .A(n16631), .B(n16630), .ZN(n16709) );
  AOI22_X1 U19896 ( .A1(n16708), .A2(n16632), .B1(n12997), .B2(n16709), .ZN(
        n16633) );
  INV_X1 U19897 ( .A(n16633), .ZN(n16634) );
  AOI21_X1 U19898 ( .B1(n19622), .B2(n19380), .A(n16634), .ZN(n16635) );
  OAI211_X1 U19899 ( .C1(n16637), .C2(n19642), .A(n16636), .B(n16635), .ZN(
        P2_U3006) );
  AOI22_X1 U19900 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16638), .B1(
        n19613), .B2(n19401), .ZN(n16643) );
  OAI22_X1 U19901 ( .A1(n16640), .A2(n19636), .B1(n19619), .B2(n16639), .ZN(
        n16641) );
  AOI21_X1 U19902 ( .B1(n19622), .B2(n19402), .A(n16641), .ZN(n16642) );
  OAI211_X1 U19903 ( .C1(n20209), .C2(n19388), .A(n16643), .B(n16642), .ZN(
        P2_U3008) );
  INV_X1 U19904 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20222) );
  NOR2_X1 U19905 ( .A1(n20222), .A2(n19272), .ZN(n16648) );
  OAI21_X1 U19906 ( .B1(n16659), .B2(n16645), .A(n16644), .ZN(n19468) );
  OAI22_X1 U19907 ( .A1(n19468), .A2(n19667), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16646), .ZN(n16647) );
  AOI211_X1 U19908 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16649), .A(
        n16648), .B(n16647), .ZN(n16652) );
  AOI22_X1 U19909 ( .A1(n9784), .A2(n19660), .B1(n19669), .B2(n16650), .ZN(
        n16651) );
  OAI211_X1 U19910 ( .C1(n16653), .C2(n16702), .A(n16652), .B(n16651), .ZN(
        P2_U3031) );
  NOR2_X1 U19911 ( .A1(n16656), .A2(n16654), .ZN(n16658) );
  AOI21_X1 U19912 ( .B1(n16669), .B2(n16656), .A(n16655), .ZN(n16674) );
  INV_X1 U19913 ( .A(n16674), .ZN(n16657) );
  MUX2_X1 U19914 ( .A(n16658), .B(n16657), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16663) );
  AOI21_X1 U19915 ( .B1(n16670), .B2(n16660), .A(n16659), .ZN(n19469) );
  NAND2_X1 U19916 ( .A1(n19469), .A2(n19645), .ZN(n16661) );
  OAI21_X1 U19917 ( .B1(n11265), .B2(n19388), .A(n16661), .ZN(n16662) );
  NOR2_X1 U19918 ( .A1(n16663), .A2(n16662), .ZN(n16667) );
  INV_X1 U19919 ( .A(n16664), .ZN(n16665) );
  AOI22_X1 U19920 ( .A1(n16665), .A2(n19663), .B1(n19669), .B2(n19326), .ZN(
        n16666) );
  OAI211_X1 U19921 ( .C1(n19650), .C2(n16668), .A(n16667), .B(n16666), .ZN(
        P2_U3032) );
  AOI21_X1 U19922 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16669), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16673) );
  OAI21_X1 U19923 ( .B1(n16672), .B2(n16671), .A(n16670), .ZN(n19473) );
  OAI22_X1 U19924 ( .A1(n16674), .A2(n16673), .B1(n19473), .B2(n19667), .ZN(
        n16675) );
  AOI21_X1 U19925 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19643), .A(n16675), 
        .ZN(n16679) );
  AOI22_X1 U19926 ( .A1(n16677), .A2(n19660), .B1(n19669), .B2(n16676), .ZN(
        n16678) );
  OAI211_X1 U19927 ( .C1(n16702), .C2(n16680), .A(n16679), .B(n16678), .ZN(
        P2_U3033) );
  AOI21_X1 U19928 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16682), .A(
        n16681), .ZN(n16698) );
  INV_X1 U19929 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n21297) );
  NOR2_X1 U19930 ( .A1(n21297), .A2(n19272), .ZN(n16687) );
  NAND2_X1 U19931 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16683), .ZN(
        n16695) );
  OAI21_X1 U19932 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16684), .ZN(n16685) );
  OAI22_X1 U19933 ( .A1(n19477), .A2(n19667), .B1(n16695), .B2(n16685), .ZN(
        n16686) );
  AOI211_X1 U19934 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16698), .A(
        n16687), .B(n16686), .ZN(n16691) );
  AOI22_X1 U19935 ( .A1(n16689), .A2(n19663), .B1(n19669), .B2(n16688), .ZN(
        n16690) );
  OAI211_X1 U19936 ( .C1(n19650), .C2(n16692), .A(n16691), .B(n16690), .ZN(
        P2_U3035) );
  NOR2_X1 U19937 ( .A1(n20215), .A2(n19272), .ZN(n16697) );
  XNOR2_X1 U19938 ( .A(n16694), .B(n16693), .ZN(n19480) );
  OAI22_X1 U19939 ( .A1(n19480), .A2(n19667), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16695), .ZN(n16696) );
  AOI211_X1 U19940 ( .C1(n16698), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16697), .B(n16696), .ZN(n16701) );
  AOI22_X1 U19941 ( .A1(n16699), .A2(n19660), .B1(n19669), .B2(n19358), .ZN(
        n16700) );
  OAI211_X1 U19942 ( .C1(n16703), .C2(n16702), .A(n16701), .B(n16700), .ZN(
        P2_U3036) );
  AOI21_X1 U19943 ( .B1(n16706), .B2(n16705), .A(n16704), .ZN(n19484) );
  AOI22_X1 U19944 ( .A1(n16707), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19645), .B2(n19484), .ZN(n16715) );
  AOI222_X1 U19945 ( .A1(n16709), .A2(n19663), .B1(n19669), .B2(n19380), .C1(
        n16708), .C2(n19660), .ZN(n16714) );
  NAND2_X1 U19946 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19643), .ZN(n16713) );
  OAI211_X1 U19947 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16711), .B(n16710), .ZN(n16712) );
  NAND4_X1 U19948 ( .A1(n16715), .A2(n16714), .A3(n16713), .A4(n16712), .ZN(
        P2_U3038) );
  AOI22_X1 U19949 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16717), .B1(
        n19663), .B2(n16716), .ZN(n16725) );
  AOI21_X1 U19950 ( .B1(n19669), .B2(n13096), .A(n16718), .ZN(n16723) );
  NAND2_X1 U19951 ( .A1(n19660), .A2(n16719), .ZN(n16722) );
  NAND2_X1 U19952 ( .A1(n19645), .A2(n16720), .ZN(n16721) );
  AND3_X1 U19953 ( .A1(n16723), .A2(n16722), .A3(n16721), .ZN(n16724) );
  OAI211_X1 U19954 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16726), .A(
        n16725), .B(n16724), .ZN(P2_U3046) );
  AOI211_X1 U19955 ( .C1(n20302), .C2(n16729), .A(n16728), .B(n16727), .ZN(
        n16739) );
  OAI21_X1 U19956 ( .B1(n16731), .B2(n16730), .A(n21192), .ZN(n16733) );
  INV_X1 U19957 ( .A(n16735), .ZN(n16732) );
  NAND2_X1 U19958 ( .A1(n16733), .A2(n16732), .ZN(n16737) );
  NAND3_X1 U19959 ( .A1(n16735), .A2(n16734), .A3(n21192), .ZN(n16736) );
  NAND2_X1 U19960 ( .A1(n16737), .A2(n16736), .ZN(n16738) );
  OAI211_X1 U19961 ( .C1(n16740), .C2(n19533), .A(n16739), .B(n16738), .ZN(
        P2_U3176) );
  NAND2_X1 U19962 ( .A1(n18107), .A2(n16742), .ZN(n16747) );
  OAI211_X1 U19963 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16798), .A(
        n16743), .B(n16747), .ZN(n16745) );
  INV_X1 U19964 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19180) );
  AOI22_X1 U19965 ( .A1(n18109), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n19180), .B2(n18107), .ZN(n16749) );
  NOR2_X1 U19966 ( .A1(n19180), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16744) );
  OAI21_X1 U19967 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16746), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16748) );
  NAND3_X1 U19968 ( .A1(n16749), .A2(n16748), .A3(n16747), .ZN(n16750) );
  NOR2_X1 U19969 ( .A1(n18529), .A2(n21249), .ZN(n16800) );
  NAND2_X1 U19970 ( .A1(n9844), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16753) );
  NAND2_X1 U19971 ( .A1(n19218), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19080) );
  OR2_X1 U19972 ( .A1(n16753), .A2(n18028), .ZN(n16769) );
  XNOR2_X1 U19973 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16756) );
  INV_X1 U19974 ( .A(n17980), .ZN(n17950) );
  NOR2_X1 U19975 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17950), .ZN(
        n16788) );
  INV_X1 U19976 ( .A(n19080), .ZN(n17921) );
  AOI22_X1 U19977 ( .A1(n18585), .A2(n16753), .B1(n17921), .B2(n16752), .ZN(
        n16754) );
  NAND2_X1 U19978 ( .A1(n16754), .A2(n9733), .ZN(n16789) );
  NOR2_X1 U19979 ( .A1(n16788), .A2(n16789), .ZN(n16767) );
  OAI22_X1 U19980 ( .A1(n16769), .A2(n16756), .B1(n16767), .B2(n16755), .ZN(
        n16757) );
  AOI211_X1 U19981 ( .C1(n18050), .C2(n9958), .A(n16800), .B(n16757), .ZN(
        n16763) );
  NAND2_X1 U19982 ( .A1(n17691), .A2(n18191), .ZN(n18072) );
  INV_X1 U19983 ( .A(n18072), .ZN(n18111) );
  NAND3_X1 U19984 ( .A1(n16758), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16759) );
  XOR2_X1 U19985 ( .A(n16759), .B(n19180), .Z(n16803) );
  NAND2_X1 U19986 ( .A1(n16760), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16761) );
  XOR2_X1 U19987 ( .A(n16761), .B(n19180), .Z(n16802) );
  AOI22_X1 U19988 ( .A1(n18111), .A2(n16803), .B1(n18143), .B2(n16802), .ZN(
        n16762) );
  OAI211_X1 U19989 ( .C1(n17979), .C2(n16806), .A(n16763), .B(n16762), .ZN(
        P3_U2799) );
  NAND2_X1 U19990 ( .A1(n18111), .A2(n16764), .ZN(n16780) );
  NAND2_X1 U19991 ( .A1(n18143), .A2(n16765), .ZN(n16782) );
  AOI21_X1 U19992 ( .B1(n16780), .B2(n16782), .A(n16798), .ZN(n16771) );
  OAI221_X1 U19993 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16769), .C1(
        n16768), .C2(n16767), .A(n16766), .ZN(n16770) );
  AOI211_X1 U19994 ( .C1(n18050), .C2(n16772), .A(n16771), .B(n16770), .ZN(
        n16777) );
  INV_X1 U19995 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18212) );
  OAI22_X1 U19996 ( .A1(n18039), .A2(n18072), .B1(n18202), .B2(n18021), .ZN(
        n18058) );
  NAND2_X1 U19997 ( .A1(n18058), .A2(n16773), .ZN(n18001) );
  NAND4_X1 U19998 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n18251), .A4(n17976), .ZN(
        n17865) );
  NOR2_X1 U19999 ( .A1(n18212), .A2(n17865), .ZN(n17859) );
  NAND3_X1 U20000 ( .A1(n16775), .A2(n17859), .A3(n16774), .ZN(n16776) );
  OAI211_X1 U20001 ( .C1(n16778), .C2(n17979), .A(n16777), .B(n16776), .ZN(
        P3_U2800) );
  INV_X1 U20002 ( .A(n16779), .ZN(n16787) );
  AOI21_X1 U20003 ( .B1(n16781), .B2(n16783), .A(n16780), .ZN(n16786) );
  AOI21_X1 U20004 ( .B1(n16784), .B2(n16783), .A(n16782), .ZN(n16785) );
  OAI21_X1 U20005 ( .B1(n16788), .B2(n18050), .A(n16933), .ZN(n16791) );
  OAI221_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9844), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18585), .A(n16789), .ZN(
        n16790) );
  NAND4_X1 U20007 ( .A1(n16793), .A2(n16792), .A3(n16791), .A4(n16790), .ZN(
        P3_U2801) );
  OAI21_X1 U20008 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16795), .A(
        n16794), .ZN(n16801) );
  NOR4_X1 U20009 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16798), .A3(
        n16797), .A4(n16796), .ZN(n16799) );
  AOI211_X1 U20010 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16801), .A(
        n16800), .B(n16799), .ZN(n16805) );
  AOI22_X1 U20011 ( .A1(n16803), .A2(n18442), .B1(n16802), .B2(n18526), .ZN(
        n16804) );
  OAI211_X1 U20012 ( .C1(n18325), .C2(n16806), .A(n16805), .B(n16804), .ZN(
        P3_U2831) );
  NOR3_X1 U20013 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16808) );
  NOR4_X1 U20014 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16807) );
  INV_X2 U20015 ( .A(n16900), .ZN(U215) );
  NAND4_X1 U20016 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16808), .A3(n16807), .A4(
        U215), .ZN(U213) );
  INV_X1 U20017 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19538) );
  OAI222_X1 U20018 ( .A1(U212), .A2(n19538), .B1(n16866), .B2(n16811), .C1(
        U214), .C2(n16810), .ZN(U216) );
  INV_X1 U20019 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19542) );
  INV_X1 U20020 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n20413) );
  OAI222_X1 U20021 ( .A1(U212), .A2(n19542), .B1(n16866), .B2(n16812), .C1(
        U214), .C2(n20413), .ZN(U217) );
  INV_X2 U20022 ( .A(U212), .ZN(n16864) );
  AOI22_X1 U20023 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16863), .ZN(n16813) );
  OAI21_X1 U20024 ( .B1(n16814), .B2(n16866), .A(n16813), .ZN(U218) );
  AOI22_X1 U20025 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16863), .ZN(n16815) );
  OAI21_X1 U20026 ( .B1(n16816), .B2(n16866), .A(n16815), .ZN(U219) );
  AOI22_X1 U20027 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16863), .ZN(n16817) );
  OAI21_X1 U20028 ( .B1(n16818), .B2(n16866), .A(n16817), .ZN(U220) );
  AOI22_X1 U20029 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16863), .ZN(n16819) );
  OAI21_X1 U20030 ( .B1(n16820), .B2(n16866), .A(n16819), .ZN(U221) );
  AOI22_X1 U20031 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16863), .ZN(n16821) );
  OAI21_X1 U20032 ( .B1(n16822), .B2(n16866), .A(n16821), .ZN(U222) );
  AOI22_X1 U20033 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16863), .ZN(n16823) );
  OAI21_X1 U20034 ( .B1(n14931), .B2(n16866), .A(n16823), .ZN(U223) );
  AOI22_X1 U20035 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16863), .ZN(n16824) );
  OAI21_X1 U20036 ( .B1(n19702), .B2(n16866), .A(n16824), .ZN(U224) );
  INV_X1 U20037 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n16826) );
  INV_X1 U20038 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21122) );
  OAI222_X1 U20039 ( .A1(U214), .A2(n16826), .B1(n16866), .B2(n16825), .C1(
        U212), .C2(n21122), .ZN(U225) );
  AOI22_X1 U20040 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16863), .ZN(n16827) );
  OAI21_X1 U20041 ( .B1(n16828), .B2(n16866), .A(n16827), .ZN(U226) );
  AOI22_X1 U20042 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16863), .ZN(n16829) );
  OAI21_X1 U20043 ( .B1(n21108), .B2(n16866), .A(n16829), .ZN(U227) );
  AOI22_X1 U20044 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16863), .ZN(n16830) );
  OAI21_X1 U20045 ( .B1(n21087), .B2(n16866), .A(n16830), .ZN(U228) );
  AOI22_X1 U20046 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16863), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16864), .ZN(n16831) );
  OAI21_X1 U20047 ( .B1(n16832), .B2(n16866), .A(n16831), .ZN(U229) );
  AOI22_X1 U20048 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16863), .ZN(n16833) );
  OAI21_X1 U20049 ( .B1(n16834), .B2(n16866), .A(n16833), .ZN(U230) );
  AOI22_X1 U20050 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16863), .ZN(n16835) );
  OAI21_X1 U20051 ( .B1(n16836), .B2(n16866), .A(n16835), .ZN(U231) );
  AOI22_X1 U20052 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16863), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16864), .ZN(n16837) );
  OAI21_X1 U20053 ( .B1(n13766), .B2(n16866), .A(n16837), .ZN(U232) );
  AOI22_X1 U20054 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16863), .ZN(n16838) );
  OAI21_X1 U20055 ( .B1(n14687), .B2(n16866), .A(n16838), .ZN(U233) );
  AOI22_X1 U20056 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16863), .ZN(n16839) );
  OAI21_X1 U20057 ( .B1(n13708), .B2(n16866), .A(n16839), .ZN(U234) );
  INV_X1 U20058 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U20059 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16863), .ZN(n16840) );
  OAI21_X1 U20060 ( .B1(n16841), .B2(n16866), .A(n16840), .ZN(U235) );
  AOI22_X1 U20061 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16863), .ZN(n16842) );
  OAI21_X1 U20062 ( .B1(n16843), .B2(n16866), .A(n16842), .ZN(U236) );
  AOI22_X1 U20063 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16863), .ZN(n16844) );
  OAI21_X1 U20064 ( .B1(n16845), .B2(n16866), .A(n16844), .ZN(U237) );
  AOI22_X1 U20065 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16863), .ZN(n16846) );
  OAI21_X1 U20066 ( .B1(n16847), .B2(n16866), .A(n16846), .ZN(U238) );
  INV_X1 U20067 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U20068 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16863), .ZN(n16848) );
  OAI21_X1 U20069 ( .B1(n16849), .B2(n16866), .A(n16848), .ZN(U239) );
  INV_X1 U20070 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16851) );
  AOI22_X1 U20071 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16863), .ZN(n16850) );
  OAI21_X1 U20072 ( .B1(n16851), .B2(n16866), .A(n16850), .ZN(U240) );
  INV_X1 U20073 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16853) );
  AOI22_X1 U20074 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16863), .ZN(n16852) );
  OAI21_X1 U20075 ( .B1(n16853), .B2(n16866), .A(n16852), .ZN(U241) );
  INV_X1 U20076 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U20077 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16863), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16864), .ZN(n16854) );
  OAI21_X1 U20078 ( .B1(n16855), .B2(n16866), .A(n16854), .ZN(U242) );
  AOI22_X1 U20079 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16863), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16864), .ZN(n16856) );
  OAI21_X1 U20080 ( .B1(n16857), .B2(n16866), .A(n16856), .ZN(U243) );
  INV_X1 U20081 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20082 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16863), .ZN(n16858) );
  OAI21_X1 U20083 ( .B1(n16859), .B2(n16866), .A(n16858), .ZN(U244) );
  INV_X1 U20084 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20085 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16863), .ZN(n16860) );
  OAI21_X1 U20086 ( .B1(n16861), .B2(n16866), .A(n16860), .ZN(U245) );
  INV_X1 U20087 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n21264) );
  AOI22_X1 U20088 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16863), .ZN(n16862) );
  OAI21_X1 U20089 ( .B1(n21264), .B2(n16866), .A(n16862), .ZN(U246) );
  INV_X1 U20090 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20091 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16864), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16863), .ZN(n16865) );
  OAI21_X1 U20092 ( .B1(n16867), .B2(n16866), .A(n16865), .ZN(U247) );
  OAI22_X1 U20093 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16900), .ZN(n16868) );
  INV_X1 U20094 ( .A(n16868), .ZN(U251) );
  OAI22_X1 U20095 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16900), .ZN(n16869) );
  INV_X1 U20096 ( .A(n16869), .ZN(U252) );
  OAI22_X1 U20097 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16900), .ZN(n16870) );
  INV_X1 U20098 ( .A(n16870), .ZN(U253) );
  OAI22_X1 U20099 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16900), .ZN(n16871) );
  INV_X1 U20100 ( .A(n16871), .ZN(U254) );
  OAI22_X1 U20101 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16900), .ZN(n16872) );
  INV_X1 U20102 ( .A(n16872), .ZN(U255) );
  OAI22_X1 U20103 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16900), .ZN(n16873) );
  INV_X1 U20104 ( .A(n16873), .ZN(U256) );
  OAI22_X1 U20105 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16900), .ZN(n16874) );
  INV_X1 U20106 ( .A(n16874), .ZN(U257) );
  OAI22_X1 U20107 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16900), .ZN(n16875) );
  INV_X1 U20108 ( .A(n16875), .ZN(U258) );
  OAI22_X1 U20109 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16900), .ZN(n16876) );
  INV_X1 U20110 ( .A(n16876), .ZN(U259) );
  OAI22_X1 U20111 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16890), .ZN(n16877) );
  INV_X1 U20112 ( .A(n16877), .ZN(U260) );
  OAI22_X1 U20113 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16890), .ZN(n16878) );
  INV_X1 U20114 ( .A(n16878), .ZN(U261) );
  OAI22_X1 U20115 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16900), .ZN(n16879) );
  INV_X1 U20116 ( .A(n16879), .ZN(U262) );
  OAI22_X1 U20117 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16890), .ZN(n16880) );
  INV_X1 U20118 ( .A(n16880), .ZN(U263) );
  OAI22_X1 U20119 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16900), .ZN(n16881) );
  INV_X1 U20120 ( .A(n16881), .ZN(U264) );
  OAI22_X1 U20121 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16900), .ZN(n16882) );
  INV_X1 U20122 ( .A(n16882), .ZN(U265) );
  OAI22_X1 U20123 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16890), .ZN(n16883) );
  INV_X1 U20124 ( .A(n16883), .ZN(U266) );
  OAI22_X1 U20125 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16890), .ZN(n16884) );
  INV_X1 U20126 ( .A(n16884), .ZN(U267) );
  OAI22_X1 U20127 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16890), .ZN(n16885) );
  INV_X1 U20128 ( .A(n16885), .ZN(U268) );
  OAI22_X1 U20129 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16890), .ZN(n16886) );
  INV_X1 U20130 ( .A(n16886), .ZN(U269) );
  OAI22_X1 U20131 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16890), .ZN(n16887) );
  INV_X1 U20132 ( .A(n16887), .ZN(U270) );
  OAI22_X1 U20133 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16890), .ZN(n16888) );
  INV_X1 U20134 ( .A(n16888), .ZN(U271) );
  OAI22_X1 U20135 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16900), .ZN(n16889) );
  INV_X1 U20136 ( .A(n16889), .ZN(U272) );
  AOI22_X1 U20137 ( .A1(n16900), .A2(n21122), .B1(n18581), .B2(U215), .ZN(U273) );
  OAI22_X1 U20138 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16890), .ZN(n16891) );
  INV_X1 U20139 ( .A(n16891), .ZN(U274) );
  OAI22_X1 U20140 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16900), .ZN(n16892) );
  INV_X1 U20141 ( .A(n16892), .ZN(U275) );
  OAI22_X1 U20142 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16900), .ZN(n16893) );
  INV_X1 U20143 ( .A(n16893), .ZN(U276) );
  OAI22_X1 U20144 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16900), .ZN(n16894) );
  INV_X1 U20145 ( .A(n16894), .ZN(U277) );
  OAI22_X1 U20146 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16900), .ZN(n16895) );
  INV_X1 U20147 ( .A(n16895), .ZN(U278) );
  OAI22_X1 U20148 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16900), .ZN(n16896) );
  INV_X1 U20149 ( .A(n16896), .ZN(U279) );
  OAI22_X1 U20150 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16900), .ZN(n16897) );
  INV_X1 U20151 ( .A(n16897), .ZN(U280) );
  AOI22_X1 U20152 ( .A1(n16900), .A2(n19542), .B1(n18578), .B2(U215), .ZN(U281) );
  INV_X1 U20153 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20154 ( .A1(n16900), .A2(n19538), .B1(n16899), .B2(U215), .ZN(U282) );
  INV_X1 U20155 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16901) );
  OAI222_X1 U20156 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n20413), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n19542), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16901), .ZN(n16903) );
  INV_X2 U20157 ( .A(n16904), .ZN(n16902) );
  INV_X1 U20158 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19117) );
  INV_X1 U20159 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U20160 ( .A1(n16902), .A2(n19117), .B1(n20216), .B2(n16904), .ZN(
        U347) );
  INV_X1 U20161 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19115) );
  INV_X1 U20162 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20214) );
  AOI22_X1 U20163 ( .A1(n16902), .A2(n19115), .B1(n20214), .B2(n16904), .ZN(
        U348) );
  INV_X1 U20164 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19112) );
  INV_X1 U20165 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20213) );
  AOI22_X1 U20166 ( .A1(n16902), .A2(n19112), .B1(n20213), .B2(n16904), .ZN(
        U349) );
  INV_X1 U20167 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19111) );
  INV_X1 U20168 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n21080) );
  AOI22_X1 U20169 ( .A1(n16902), .A2(n19111), .B1(n21080), .B2(n16904), .ZN(
        U350) );
  INV_X1 U20170 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19108) );
  INV_X1 U20171 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U20172 ( .A1(n16902), .A2(n19108), .B1(n20210), .B2(n16904), .ZN(
        U351) );
  INV_X1 U20173 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19107) );
  INV_X1 U20174 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U20175 ( .A1(n16902), .A2(n19107), .B1(n20208), .B2(n16904), .ZN(
        U352) );
  INV_X1 U20176 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19105) );
  AOI22_X1 U20177 ( .A1(n16902), .A2(n19105), .B1(n20207), .B2(n16904), .ZN(
        U353) );
  INV_X1 U20178 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19103) );
  INV_X1 U20179 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n21237) );
  AOI22_X1 U20180 ( .A1(n16902), .A2(n19103), .B1(n21237), .B2(n16904), .ZN(
        U354) );
  INV_X1 U20181 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19158) );
  INV_X1 U20182 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20248) );
  AOI22_X1 U20183 ( .A1(n16902), .A2(n19158), .B1(n20248), .B2(n16903), .ZN(
        U355) );
  INV_X1 U20184 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19154) );
  INV_X1 U20185 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20246) );
  AOI22_X1 U20186 ( .A1(n16902), .A2(n19154), .B1(n20246), .B2(n16904), .ZN(
        U356) );
  INV_X1 U20187 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19152) );
  INV_X1 U20188 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20244) );
  AOI22_X1 U20189 ( .A1(n16902), .A2(n19152), .B1(n20244), .B2(n16904), .ZN(
        U357) );
  INV_X1 U20190 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19149) );
  INV_X1 U20191 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20242) );
  AOI22_X1 U20192 ( .A1(n16902), .A2(n19149), .B1(n20242), .B2(n16903), .ZN(
        U358) );
  INV_X1 U20193 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19148) );
  INV_X1 U20194 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20241) );
  AOI22_X1 U20195 ( .A1(n16902), .A2(n19148), .B1(n20241), .B2(n16903), .ZN(
        U359) );
  INV_X1 U20196 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19146) );
  INV_X1 U20197 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20239) );
  AOI22_X1 U20198 ( .A1(n16902), .A2(n19146), .B1(n20239), .B2(n16903), .ZN(
        U360) );
  INV_X1 U20199 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19143) );
  INV_X1 U20200 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20237) );
  AOI22_X1 U20201 ( .A1(n16902), .A2(n19143), .B1(n20237), .B2(n16903), .ZN(
        U361) );
  INV_X1 U20202 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19141) );
  INV_X1 U20203 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20235) );
  AOI22_X1 U20204 ( .A1(n16902), .A2(n19141), .B1(n20235), .B2(n16904), .ZN(
        U362) );
  INV_X1 U20205 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19140) );
  INV_X1 U20206 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20234) );
  AOI22_X1 U20207 ( .A1(n16902), .A2(n19140), .B1(n20234), .B2(n16904), .ZN(
        U363) );
  INV_X1 U20208 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19139) );
  INV_X1 U20209 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20233) );
  AOI22_X1 U20210 ( .A1(n16902), .A2(n19139), .B1(n20233), .B2(n16904), .ZN(
        U364) );
  INV_X1 U20211 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19101) );
  INV_X1 U20212 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20203) );
  AOI22_X1 U20213 ( .A1(n16902), .A2(n19101), .B1(n20203), .B2(n16904), .ZN(
        U365) );
  INV_X1 U20214 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19137) );
  INV_X1 U20215 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20231) );
  AOI22_X1 U20216 ( .A1(n16902), .A2(n19137), .B1(n20231), .B2(n16904), .ZN(
        U366) );
  INV_X1 U20217 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19135) );
  INV_X1 U20218 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21280) );
  AOI22_X1 U20219 ( .A1(n16902), .A2(n19135), .B1(n21280), .B2(n16904), .ZN(
        U367) );
  INV_X1 U20220 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19133) );
  INV_X1 U20221 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20228) );
  AOI22_X1 U20222 ( .A1(n16902), .A2(n19133), .B1(n20228), .B2(n16904), .ZN(
        U368) );
  INV_X1 U20223 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19131) );
  INV_X1 U20224 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21202) );
  AOI22_X1 U20225 ( .A1(n16902), .A2(n19131), .B1(n21202), .B2(n16904), .ZN(
        U369) );
  INV_X1 U20226 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19129) );
  INV_X1 U20227 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U20228 ( .A1(n16902), .A2(n19129), .B1(n20225), .B2(n16904), .ZN(
        U370) );
  INV_X1 U20229 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19126) );
  INV_X1 U20230 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20223) );
  AOI22_X1 U20231 ( .A1(n16902), .A2(n19126), .B1(n20223), .B2(n16904), .ZN(
        U371) );
  INV_X1 U20232 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19125) );
  INV_X1 U20233 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20221) );
  AOI22_X1 U20234 ( .A1(n16902), .A2(n19125), .B1(n20221), .B2(n16903), .ZN(
        U372) );
  INV_X1 U20235 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19123) );
  INV_X1 U20236 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20220) );
  AOI22_X1 U20237 ( .A1(n16902), .A2(n19123), .B1(n20220), .B2(n16904), .ZN(
        U373) );
  INV_X1 U20238 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19121) );
  INV_X1 U20239 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U20240 ( .A1(n16902), .A2(n19121), .B1(n20218), .B2(n16903), .ZN(
        U374) );
  INV_X1 U20241 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19119) );
  INV_X1 U20242 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n21227) );
  AOI22_X1 U20243 ( .A1(n16902), .A2(n19119), .B1(n21227), .B2(n16903), .ZN(
        U375) );
  INV_X1 U20244 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19100) );
  INV_X1 U20245 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20201) );
  AOI22_X1 U20246 ( .A1(n16902), .A2(n19100), .B1(n20201), .B2(n16904), .ZN(
        U376) );
  INV_X1 U20247 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19098) );
  NAND2_X1 U20248 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19098), .ZN(n16905) );
  AOI22_X1 U20249 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n16905), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19096), .ZN(n19166) );
  AOI21_X1 U20250 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19166), .ZN(n16906) );
  INV_X1 U20251 ( .A(n16906), .ZN(P3_U2633) );
  INV_X1 U20252 ( .A(n18198), .ZN(n19071) );
  OAI21_X1 U20253 ( .B1(n16914), .B2(n17784), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16907) );
  OAI21_X1 U20254 ( .B1(n16908), .B2(n19071), .A(n16907), .ZN(P3_U2634) );
  AOI21_X1 U20255 ( .B1(n19096), .B2(n19098), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16909) );
  AOI22_X1 U20256 ( .A1(n19225), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16909), 
        .B2(n19226), .ZN(P3_U2635) );
  INV_X1 U20257 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19083) );
  NAND2_X1 U20258 ( .A1(n19083), .A2(n19098), .ZN(n19082) );
  INV_X1 U20259 ( .A(n19082), .ZN(n16910) );
  OAI21_X1 U20260 ( .B1(n16910), .B2(BS16), .A(n19166), .ZN(n19164) );
  OAI21_X1 U20261 ( .B1(n19166), .B2(n16911), .A(n19164), .ZN(P3_U2636) );
  NOR3_X1 U20262 ( .A1(n16914), .A2(n16913), .A3(n16912), .ZN(n19006) );
  NOR2_X1 U20263 ( .A1(n19006), .A2(n19068), .ZN(n19208) );
  OAI21_X1 U20264 ( .B1(n19208), .B2(n18535), .A(n16915), .ZN(P3_U2637) );
  NOR4_X1 U20265 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16919) );
  NOR4_X1 U20266 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16918) );
  NOR4_X1 U20267 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16917) );
  NOR4_X1 U20268 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16916) );
  NAND4_X1 U20269 ( .A1(n16919), .A2(n16918), .A3(n16917), .A4(n16916), .ZN(
        n16925) );
  NOR4_X1 U20270 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16923) );
  AOI211_X1 U20271 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_9__SCAN_IN), .B(
        P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n16922) );
  NOR4_X1 U20272 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16921) );
  NOR4_X1 U20273 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16920) );
  NAND4_X1 U20274 ( .A1(n16923), .A2(n16922), .A3(n16921), .A4(n16920), .ZN(
        n16924) );
  NOR2_X1 U20275 ( .A1(n16925), .A2(n16924), .ZN(n19206) );
  INV_X1 U20276 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16927) );
  NOR3_X1 U20277 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16928) );
  OAI21_X1 U20278 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16928), .A(n19206), .ZN(
        n16926) );
  OAI21_X1 U20279 ( .B1(n19206), .B2(n16927), .A(n16926), .ZN(P3_U2638) );
  INV_X1 U20280 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19165) );
  AOI21_X1 U20281 ( .B1(n19099), .B2(n19165), .A(n16928), .ZN(n16930) );
  INV_X1 U20282 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16929) );
  INV_X1 U20283 ( .A(n19206), .ZN(n19203) );
  AOI22_X1 U20284 ( .A1(n19206), .A2(n16930), .B1(n16929), .B2(n19203), .ZN(
        P3_U2639) );
  INV_X1 U20285 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19153) );
  NAND3_X1 U20286 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16941), .ZN(n16935) );
  OAI22_X1 U20287 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16935), .B1(n16934), 
        .B2(n17254), .ZN(n16936) );
  INV_X1 U20288 ( .A(n16937), .ZN(n16938) );
  OAI21_X1 U20289 ( .B1(n16942), .B2(n17275), .A(n16938), .ZN(n16939) );
  NAND2_X1 U20290 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16941), .ZN(n16951) );
  AOI22_X1 U20291 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17244), .B1(
        n17266), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16950) );
  INV_X1 U20292 ( .A(n16941), .ZN(n16953) );
  OAI21_X1 U20293 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16953), .A(n16969), 
        .ZN(n16948) );
  AOI211_X1 U20294 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16956), .A(n16942), .B(
        n17258), .ZN(n16947) );
  AOI211_X1 U20295 ( .C1(n16945), .C2(n16944), .A(n16943), .B(n19076), .ZN(
        n16946) );
  AOI211_X1 U20296 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16948), .A(n16947), 
        .B(n16946), .ZN(n16949) );
  OAI211_X1 U20297 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16951), .A(n16950), 
        .B(n16949), .ZN(P3_U2643) );
  INV_X1 U20298 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19150) );
  AOI211_X1 U20299 ( .C1(n17853), .C2(n16952), .A(n9951), .B(n19076), .ZN(
        n16955) );
  OAI22_X1 U20300 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16953), .B1(n17857), 
        .B2(n17254), .ZN(n16954) );
  AOI211_X1 U20301 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17266), .A(n16955), .B(
        n16954), .ZN(n16958) );
  OAI211_X1 U20302 ( .C1(n16960), .C2(n17300), .A(n17265), .B(n16956), .ZN(
        n16957) );
  OAI211_X1 U20303 ( .C1(n16969), .C2(n19150), .A(n16958), .B(n16957), .ZN(
        P3_U2644) );
  INV_X1 U20304 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19145) );
  INV_X1 U20305 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19147) );
  OAI21_X1 U20306 ( .B1(n19145), .B2(n16974), .A(n19147), .ZN(n16959) );
  INV_X1 U20307 ( .A(n16959), .ZN(n16968) );
  AOI22_X1 U20308 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17244), .B1(
        n17266), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16967) );
  AOI211_X1 U20309 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16961), .A(n16960), .B(
        n17258), .ZN(n16965) );
  AOI211_X1 U20310 ( .C1(n17867), .C2(n16963), .A(n16962), .B(n19076), .ZN(
        n16964) );
  NOR2_X1 U20311 ( .A1(n16965), .A2(n16964), .ZN(n16966) );
  OAI211_X1 U20312 ( .C1(n16969), .C2(n16968), .A(n16967), .B(n16966), .ZN(
        P3_U2645) );
  OR2_X1 U20313 ( .A1(n17258), .A2(n16970), .ZN(n16983) );
  AOI21_X1 U20314 ( .B1(n17265), .B2(n16970), .A(n17266), .ZN(n16979) );
  INV_X1 U20315 ( .A(n16989), .ZN(n17001) );
  OAI21_X1 U20316 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17245), .A(n17001), 
        .ZN(n16977) );
  AOI211_X1 U20317 ( .C1(n17877), .C2(n16971), .A(n16972), .B(n19076), .ZN(
        n16976) );
  OAI22_X1 U20318 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16974), .B1(n16973), 
        .B2(n17254), .ZN(n16975) );
  AOI211_X1 U20319 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16977), .A(n16976), 
        .B(n16975), .ZN(n16978) );
  OAI221_X1 U20320 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16983), .C1(n16980), 
        .C2(n16979), .A(n16978), .ZN(P3_U2646) );
  NOR2_X1 U20321 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17245), .ZN(n16981) );
  AOI22_X1 U20322 ( .A1(n17266), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16982), 
        .B2(n16981), .ZN(n16991) );
  AOI21_X1 U20323 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16998), .A(n16983), .ZN(
        n16988) );
  AOI211_X1 U20324 ( .C1(n16986), .C2(n16985), .A(n16984), .B(n19076), .ZN(
        n16987) );
  AOI211_X1 U20325 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16989), .A(n16988), 
        .B(n16987), .ZN(n16990) );
  OAI211_X1 U20326 ( .C1(n21279), .C2(n17254), .A(n16991), .B(n16990), .ZN(
        P3_U2647) );
  AOI211_X1 U20327 ( .C1(n17903), .C2(n16992), .A(n16993), .B(n19076), .ZN(
        n16997) );
  NAND2_X1 U20328 ( .A1(n17247), .A2(n19142), .ZN(n16994) );
  OAI22_X1 U20329 ( .A1(n17897), .A2(n17254), .B1(n16995), .B2(n16994), .ZN(
        n16996) );
  AOI211_X1 U20330 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n17266), .A(n16997), .B(
        n16996), .ZN(n17000) );
  OAI211_X1 U20331 ( .C1(n17002), .C2(n17274), .A(n17265), .B(n16998), .ZN(
        n16999) );
  OAI211_X1 U20332 ( .C1(n17001), .C2(n19142), .A(n17000), .B(n16999), .ZN(
        P3_U2648) );
  AOI22_X1 U20333 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17244), .B1(
        n17266), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n17010) );
  OAI221_X1 U20334 ( .B1(n17245), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17245), 
        .C2(n17020), .A(n17268), .ZN(n17007) );
  AOI211_X1 U20335 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17014), .A(n17002), .B(
        n17258), .ZN(n17006) );
  AOI211_X1 U20336 ( .C1(n17929), .C2(n17003), .A(n17004), .B(n19076), .ZN(
        n17005) );
  AOI211_X1 U20337 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17007), .A(n17006), 
        .B(n17005), .ZN(n17009) );
  INV_X1 U20338 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21123) );
  NAND4_X1 U20339 ( .A1(n17247), .A2(P3_REIP_REG_21__SCAN_IN), .A3(n17020), 
        .A4(n21123), .ZN(n17008) );
  NAND3_X1 U20340 ( .A1(n17010), .A2(n17009), .A3(n17008), .ZN(P3_U2649) );
  AOI22_X1 U20341 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17244), .B1(
        n17266), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n17018) );
  OAI21_X1 U20342 ( .B1(n17020), .B2(n17245), .A(n17268), .ZN(n17019) );
  AOI211_X1 U20343 ( .C1(n17936), .C2(n17011), .A(n17012), .B(n19076), .ZN(
        n17013) );
  AOI21_X1 U20344 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n17019), .A(n17013), 
        .ZN(n17017) );
  INV_X1 U20345 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19138) );
  NAND3_X1 U20346 ( .A1(n17247), .A2(n17020), .A3(n19138), .ZN(n17016) );
  OAI211_X1 U20347 ( .C1(n17024), .C2(n17348), .A(n17265), .B(n17014), .ZN(
        n17015) );
  NAND4_X1 U20348 ( .A1(n17018), .A2(n17017), .A3(n17016), .A4(n17015), .ZN(
        P3_U2650) );
  INV_X1 U20349 ( .A(n17019), .ZN(n17031) );
  AOI22_X1 U20350 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17244), .B1(
        n17266), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n17030) );
  NOR2_X1 U20351 ( .A1(n17020), .A2(n17245), .ZN(n17028) );
  INV_X1 U20352 ( .A(n17021), .ZN(n17027) );
  AOI211_X1 U20353 ( .C1(n17951), .C2(n17023), .A(n17022), .B(n19076), .ZN(
        n17026) );
  AOI211_X1 U20354 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17039), .A(n17024), .B(
        n17258), .ZN(n17025) );
  AOI211_X1 U20355 ( .C1(n17028), .C2(n17027), .A(n17026), .B(n17025), .ZN(
        n17029) );
  OAI211_X1 U20356 ( .C1(n17031), .C2(n19136), .A(n17030), .B(n17029), .ZN(
        P3_U2651) );
  OAI221_X1 U20357 ( .B1(n17245), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n17245), 
        .C2(n17043), .A(n17268), .ZN(n17038) );
  AOI211_X1 U20358 ( .C1(n17957), .C2(n17032), .A(n17033), .B(n19076), .ZN(
        n17037) );
  INV_X1 U20359 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19134) );
  NAND4_X1 U20360 ( .A1(n17247), .A2(P3_REIP_REG_18__SCAN_IN), .A3(n17043), 
        .A4(n19134), .ZN(n17034) );
  OAI211_X1 U20361 ( .C1(n17035), .C2(n17254), .A(n18529), .B(n17034), .ZN(
        n17036) );
  AOI211_X1 U20362 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17038), .A(n17037), 
        .B(n17036), .ZN(n17041) );
  OAI211_X1 U20363 ( .C1(n17047), .C2(n17042), .A(n17265), .B(n17039), .ZN(
        n17040) );
  OAI211_X1 U20364 ( .C1(n17042), .C2(n17259), .A(n17041), .B(n17040), .ZN(
        P3_U2652) );
  INV_X1 U20365 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19132) );
  OAI21_X1 U20366 ( .B1(n17245), .B2(n17043), .A(n17268), .ZN(n17061) );
  INV_X1 U20367 ( .A(n17061), .ZN(n17052) );
  NAND2_X1 U20368 ( .A1(n17247), .A2(n17043), .ZN(n17044) );
  NOR2_X1 U20369 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17044), .ZN(n17045) );
  AOI211_X1 U20370 ( .C1(n17266), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18523), .B(
        n17045), .ZN(n17051) );
  AOI211_X1 U20371 ( .C1(n17970), .C2(n9842), .A(n17046), .B(n19076), .ZN(
        n17049) );
  AOI211_X1 U20372 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17056), .A(n17047), .B(
        n17258), .ZN(n17048) );
  AOI211_X1 U20373 ( .C1(n17244), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17049), .B(n17048), .ZN(n17050) );
  OAI211_X1 U20374 ( .C1(n19132), .C2(n17052), .A(n17051), .B(n17050), .ZN(
        P3_U2653) );
  OAI21_X1 U20375 ( .B1(n17245), .B2(n17053), .A(n19130), .ZN(n17060) );
  AOI211_X1 U20376 ( .C1(n17984), .C2(n17055), .A(n17054), .B(n19076), .ZN(
        n17059) );
  OAI211_X1 U20377 ( .C1(n17067), .C2(n17401), .A(n17265), .B(n17056), .ZN(
        n17057) );
  OAI21_X1 U20378 ( .B1(n17254), .B2(n9977), .A(n17057), .ZN(n17058) );
  AOI211_X1 U20379 ( .C1(n17061), .C2(n17060), .A(n17059), .B(n17058), .ZN(
        n17062) );
  OAI211_X1 U20380 ( .C1(n17259), .C2(n17401), .A(n17062), .B(n18529), .ZN(
        P3_U2654) );
  NOR2_X1 U20381 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17245), .ZN(n17063) );
  AOI22_X1 U20382 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17244), .B1(
        n17064), .B2(n17063), .ZN(n17074) );
  AOI211_X1 U20383 ( .C1(n17993), .C2(n17066), .A(n17065), .B(n19076), .ZN(
        n17069) );
  AOI211_X1 U20384 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17082), .A(n17067), .B(
        n17258), .ZN(n17068) );
  AOI211_X1 U20385 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17266), .A(n17069), .B(
        n17068), .ZN(n17073) );
  NOR2_X1 U20386 ( .A1(n17246), .A2(n17071), .ZN(n17092) );
  NOR2_X1 U20387 ( .A1(n17070), .A2(n17092), .ZN(n17094) );
  NOR3_X1 U20388 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17245), .A3(n17071), 
        .ZN(n17078) );
  OAI21_X1 U20389 ( .B1(n17094), .B2(n17078), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n17072) );
  NAND4_X1 U20390 ( .A1(n17074), .A2(n17073), .A3(n18418), .A4(n17072), .ZN(
        P3_U2655) );
  OAI21_X1 U20391 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17992), .A(
        n17075), .ZN(n18002) );
  NAND2_X1 U20392 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17256), .ZN(
        n17213) );
  OAI21_X1 U20393 ( .B1(n17994), .B2(n17213), .A(n9958), .ZN(n17077) );
  OAI21_X1 U20394 ( .B1(n18002), .B2(n17077), .A(n17229), .ZN(n17076) );
  AOI21_X1 U20395 ( .B1(n18002), .B2(n17077), .A(n17076), .ZN(n17081) );
  AOI211_X1 U20396 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17244), .A(
        n18523), .B(n17078), .ZN(n17079) );
  INV_X1 U20397 ( .A(n17079), .ZN(n17080) );
  AOI211_X1 U20398 ( .C1(n17094), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17081), 
        .B(n17080), .ZN(n17084) );
  OAI211_X1 U20399 ( .C1(n17088), .C2(n17085), .A(n17265), .B(n17082), .ZN(
        n17083) );
  OAI211_X1 U20400 ( .C1(n17259), .C2(n17085), .A(n17084), .B(n17083), .ZN(
        P3_U2656) );
  INV_X1 U20401 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17086) );
  INV_X1 U20402 ( .A(n18064), .ZN(n18102) );
  NAND2_X1 U20403 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18102), .ZN(
        n17186) );
  NOR2_X1 U20404 ( .A1(n18014), .A2(n17186), .ZN(n18032) );
  NAND2_X1 U20405 ( .A1(n18030), .A2(n18032), .ZN(n17100) );
  AOI21_X1 U20406 ( .B1(n17086), .B2(n17100), .A(n17992), .ZN(n18015) );
  OAI21_X1 U20407 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17100), .A(
        n9958), .ZN(n17087) );
  XOR2_X1 U20408 ( .A(n18015), .B(n17087), .Z(n17097) );
  AOI211_X1 U20409 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17107), .A(n17088), .B(
        n17258), .ZN(n17089) );
  AOI21_X1 U20410 ( .B1(n17244), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17089), .ZN(n17096) );
  NAND2_X1 U20411 ( .A1(n17247), .A2(n17090), .ZN(n17091) );
  INV_X1 U20412 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17444) );
  OAI22_X1 U20413 ( .A1(n17092), .A2(n17091), .B1(n17259), .B2(n17444), .ZN(
        n17093) );
  AOI211_X1 U20414 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n17094), .A(n18523), 
        .B(n17093), .ZN(n17095) );
  OAI211_X1 U20415 ( .C1(n19076), .C2(n17097), .A(n17096), .B(n17095), .ZN(
        P3_U2657) );
  NOR3_X1 U20416 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17245), .A3(n17098), 
        .ZN(n17106) );
  OAI21_X1 U20417 ( .B1(n17117), .B2(n17245), .A(n17268), .ZN(n17133) );
  NOR2_X1 U20418 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17245), .ZN(n17116) );
  OAI21_X1 U20419 ( .B1(n17133), .B2(n17116), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n17104) );
  INV_X1 U20420 ( .A(n18032), .ZN(n17114) );
  NOR2_X1 U20421 ( .A1(n18046), .A2(n17114), .ZN(n17113) );
  OAI21_X1 U20422 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17113), .A(
        n17100), .ZN(n18034) );
  OAI211_X1 U20423 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n17100), .A(
        n17099), .B(n18034), .ZN(n17103) );
  INV_X1 U20424 ( .A(n18034), .ZN(n17101) );
  AOI21_X1 U20425 ( .B1(n9958), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19076), .ZN(n17262) );
  OAI211_X1 U20426 ( .C1(n18036), .C2(n9968), .A(n17101), .B(n17262), .ZN(
        n17102) );
  NAND4_X1 U20427 ( .A1(n18418), .A2(n17104), .A3(n17103), .A4(n17102), .ZN(
        n17105) );
  AOI211_X1 U20428 ( .C1(n17244), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17106), .B(n17105), .ZN(n17109) );
  OAI211_X1 U20429 ( .C1(n17111), .C2(n17110), .A(n17265), .B(n17107), .ZN(
        n17108) );
  OAI211_X1 U20430 ( .C1(n17110), .C2(n17259), .A(n17109), .B(n17108), .ZN(
        P3_U2658) );
  INV_X1 U20431 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19120) );
  INV_X1 U20432 ( .A(n17133), .ZN(n17123) );
  AOI211_X1 U20433 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17128), .A(n17111), .B(
        n17258), .ZN(n17121) );
  INV_X1 U20434 ( .A(n17213), .ZN(n17239) );
  AOI21_X1 U20435 ( .B1(n18046), .B2(n17114), .A(n17113), .ZN(n18049) );
  AOI211_X1 U20436 ( .C1(n17112), .C2(n17239), .A(n18049), .B(n17255), .ZN(
        n17115) );
  AOI211_X1 U20437 ( .C1(n17117), .C2(n17116), .A(n18523), .B(n17115), .ZN(
        n17119) );
  OAI211_X1 U20438 ( .C1(n18046), .C2(n9968), .A(n18049), .B(n17262), .ZN(
        n17118) );
  OAI211_X1 U20439 ( .C1(n17254), .C2(n18046), .A(n17119), .B(n17118), .ZN(
        n17120) );
  AOI211_X1 U20440 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17266), .A(n17121), .B(
        n17120), .ZN(n17122) );
  OAI21_X1 U20441 ( .B1(n19120), .B2(n17123), .A(n17122), .ZN(P3_U2659) );
  OAI21_X1 U20442 ( .B1(n17245), .B2(n17124), .A(n19118), .ZN(n17132) );
  OR2_X1 U20443 ( .A1(n18101), .A2(n17186), .ZN(n17159) );
  OR2_X1 U20444 ( .A1(n18066), .A2(n17159), .ZN(n17137) );
  AOI21_X1 U20445 ( .B1(n9946), .B2(n17137), .A(n18032), .ZN(n17127) );
  OAI21_X1 U20446 ( .B1(n17186), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n9958), .ZN(n17187) );
  OAI21_X1 U20447 ( .B1(n9968), .B2(n17125), .A(n17187), .ZN(n17126) );
  INV_X1 U20448 ( .A(n17127), .ZN(n18067) );
  INV_X1 U20449 ( .A(n17126), .ZN(n17138) );
  OAI221_X1 U20450 ( .B1(n17127), .B2(n17126), .C1(n18067), .C2(n17138), .A(
        n17229), .ZN(n17130) );
  OAI211_X1 U20451 ( .C1(n17146), .C2(n17135), .A(n17265), .B(n17128), .ZN(
        n17129) );
  OAI211_X1 U20452 ( .C1(n17254), .C2(n9946), .A(n17130), .B(n17129), .ZN(
        n17131) );
  AOI21_X1 U20453 ( .B1(n17133), .B2(n17132), .A(n17131), .ZN(n17134) );
  OAI211_X1 U20454 ( .C1(n17259), .C2(n17135), .A(n17134), .B(n18418), .ZN(
        P3_U2660) );
  AOI21_X1 U20455 ( .B1(n17148), .B2(P3_EBX_REG_10__SCAN_IN), .A(n17258), .ZN(
        n17136) );
  AOI21_X1 U20456 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17266), .A(n17136), .ZN(
        n17145) );
  NOR2_X1 U20457 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17159), .ZN(
        n17152) );
  AOI21_X1 U20458 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17152), .A(
        n9968), .ZN(n17150) );
  INV_X1 U20459 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18087) );
  NOR2_X1 U20460 ( .A1(n18087), .A2(n17159), .ZN(n17147) );
  OAI21_X1 U20461 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17147), .A(
        n17137), .ZN(n18085) );
  INV_X1 U20462 ( .A(n18085), .ZN(n17139) );
  AOI221_X1 U20463 ( .B1(n17150), .B2(n17139), .C1(n17138), .C2(n18085), .A(
        n19076), .ZN(n17140) );
  AOI211_X1 U20464 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n17244), .A(
        n18523), .B(n17140), .ZN(n17144) );
  OAI21_X1 U20465 ( .B1(n17141), .B2(n17245), .A(n17268), .ZN(n17163) );
  INV_X1 U20466 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19116) );
  INV_X1 U20467 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19114) );
  NOR3_X1 U20468 ( .A1(n17245), .A2(n19110), .A3(n17176), .ZN(n17164) );
  NAND2_X1 U20469 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17164), .ZN(n17158) );
  AOI221_X1 U20470 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n19116), .C2(n19114), .A(n17158), .ZN(n17142) );
  AOI21_X1 U20471 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17163), .A(n17142), 
        .ZN(n17143) );
  OAI211_X1 U20472 ( .C1(n17146), .C2(n17145), .A(n17144), .B(n17143), .ZN(
        P3_U2661) );
  INV_X1 U20473 ( .A(n17163), .ZN(n17157) );
  AOI21_X1 U20474 ( .B1(n18087), .B2(n17159), .A(n17147), .ZN(n18091) );
  NOR2_X1 U20475 ( .A1(n9958), .A2(n19076), .ZN(n17236) );
  OAI211_X1 U20476 ( .C1(n17162), .C2(n17430), .A(n17265), .B(n17148), .ZN(
        n17149) );
  OAI21_X1 U20477 ( .B1(n17254), .B2(n18087), .A(n17149), .ZN(n17155) );
  INV_X1 U20478 ( .A(n18091), .ZN(n17151) );
  OAI211_X1 U20479 ( .C1(n17152), .C2(n17151), .A(n17229), .B(n17150), .ZN(
        n17153) );
  OAI211_X1 U20480 ( .C1(n17430), .C2(n17259), .A(n18529), .B(n17153), .ZN(
        n17154) );
  AOI211_X1 U20481 ( .C1(n18091), .C2(n17236), .A(n17155), .B(n17154), .ZN(
        n17156) );
  OAI221_X1 U20482 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n17158), .C1(n19114), 
        .C2(n17157), .A(n17156), .ZN(P3_U2662) );
  NOR2_X1 U20483 ( .A1(n18118), .A2(n17186), .ZN(n17173) );
  OAI21_X1 U20484 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17173), .A(
        n17159), .ZN(n18104) );
  NOR2_X1 U20485 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17186), .ZN(
        n17160) );
  AOI21_X1 U20486 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17160), .A(
        n9968), .ZN(n17161) );
  XOR2_X1 U20487 ( .A(n18104), .B(n17161), .Z(n17170) );
  AOI211_X1 U20488 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17181), .A(n17162), .B(
        n17258), .ZN(n17168) );
  OAI21_X1 U20489 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n17164), .A(n17163), .ZN(
        n17165) );
  OAI211_X1 U20490 ( .C1(n17166), .C2(n17254), .A(n18529), .B(n17165), .ZN(
        n17167) );
  AOI211_X1 U20491 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17266), .A(n17168), .B(
        n17167), .ZN(n17169) );
  OAI21_X1 U20492 ( .B1(n19076), .B2(n17170), .A(n17169), .ZN(P3_U2663) );
  OAI21_X1 U20493 ( .B1(n17245), .B2(n17172), .A(n17268), .ZN(n17171) );
  INV_X1 U20494 ( .A(n17171), .ZN(n17196) );
  INV_X1 U20495 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19109) );
  NAND3_X1 U20496 ( .A1(n17247), .A2(n17172), .A3(n19109), .ZN(n17193) );
  AOI21_X1 U20497 ( .B1(n17196), .B2(n17193), .A(n19110), .ZN(n17180) );
  AOI21_X1 U20498 ( .B1(n18118), .B2(n17186), .A(n17173), .ZN(n18124) );
  INV_X1 U20499 ( .A(n17187), .ZN(n17175) );
  INV_X1 U20500 ( .A(n18124), .ZN(n17174) );
  AOI221_X1 U20501 ( .B1(n18124), .B2(n17175), .C1(n17174), .C2(n17187), .A(
        n19076), .ZN(n17179) );
  OR2_X1 U20502 ( .A1(n17245), .A2(n17176), .ZN(n17177) );
  OAI22_X1 U20503 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17177), .B1(n17259), 
        .B2(n17542), .ZN(n17178) );
  NOR4_X1 U20504 ( .A1(n18523), .A2(n17180), .A3(n17179), .A4(n17178), .ZN(
        n17183) );
  OAI211_X1 U20505 ( .C1(n17184), .C2(n17542), .A(n17265), .B(n17181), .ZN(
        n17182) );
  OAI211_X1 U20506 ( .C1(n17254), .C2(n18118), .A(n17183), .B(n17182), .ZN(
        P3_U2664) );
  AOI211_X1 U20507 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17198), .A(n17184), .B(
        n17258), .ZN(n17192) );
  NAND3_X1 U20508 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17185), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17208) );
  NOR2_X1 U20509 ( .A1(n18144), .A2(n17208), .ZN(n17195) );
  OAI21_X1 U20510 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17195), .A(
        n17186), .ZN(n18132) );
  AOI21_X1 U20511 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9958), .A(
        n18132), .ZN(n17189) );
  NOR2_X1 U20512 ( .A1(n19076), .A2(n17187), .ZN(n17188) );
  AOI22_X1 U20513 ( .A1(n17189), .A2(n17262), .B1(n17188), .B2(n18132), .ZN(
        n17190) );
  OAI211_X1 U20514 ( .C1(n17196), .C2(n19109), .A(n17190), .B(n18529), .ZN(
        n17191) );
  AOI211_X1 U20515 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17266), .A(n17192), .B(
        n17191), .ZN(n17194) );
  OAI211_X1 U20516 ( .C1(n17254), .C2(n9948), .A(n17194), .B(n17193), .ZN(
        P3_U2665) );
  AOI21_X1 U20517 ( .B1(n18144), .B2(n17208), .A(n17195), .ZN(n18146) );
  OAI21_X1 U20518 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17208), .A(
        n9958), .ZN(n17214) );
  XNOR2_X1 U20519 ( .A(n18146), .B(n17214), .ZN(n17202) );
  AOI221_X1 U20520 ( .B1(n17245), .B2(n19106), .C1(n17197), .C2(n19106), .A(
        n17196), .ZN(n17201) );
  OAI211_X1 U20521 ( .C1(n17207), .C2(n17204), .A(n17265), .B(n17198), .ZN(
        n17199) );
  OAI21_X1 U20522 ( .B1(n17254), .B2(n18144), .A(n17199), .ZN(n17200) );
  AOI211_X1 U20523 ( .C1(n17202), .C2(n17229), .A(n17201), .B(n17200), .ZN(
        n17203) );
  OAI211_X1 U20524 ( .C1(n17259), .C2(n17204), .A(n17203), .B(n18529), .ZN(
        P3_U2666) );
  NOR2_X1 U20525 ( .A1(n17206), .A2(n17205), .ZN(n19233) );
  AOI221_X1 U20526 ( .B1(n10308), .B2(n19233), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19233), .A(n18523), .ZN(
        n17221) );
  AOI211_X1 U20527 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17230), .A(n17207), .B(
        n17258), .ZN(n17211) );
  INV_X1 U20528 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17212) );
  AND2_X1 U20529 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17185), .ZN(
        n17223) );
  OAI21_X1 U20530 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17223), .A(
        n17208), .ZN(n18163) );
  INV_X1 U20531 ( .A(n17236), .ZN(n17209) );
  OAI22_X1 U20532 ( .A1(n17212), .A2(n17254), .B1(n18163), .B2(n17209), .ZN(
        n17210) );
  AOI211_X1 U20533 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17266), .A(n17211), .B(
        n17210), .ZN(n17220) );
  INV_X1 U20534 ( .A(n18163), .ZN(n17215) );
  NAND2_X1 U20535 ( .A1(n17185), .A2(n17212), .ZN(n18155) );
  OAI22_X1 U20536 ( .A1(n17215), .A2(n17214), .B1(n17213), .B2(n18155), .ZN(
        n17216) );
  OAI21_X1 U20537 ( .B1(n17217), .B2(n17245), .A(n17268), .ZN(n17227) );
  AOI22_X1 U20538 ( .A1(n17229), .A2(n17216), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n17227), .ZN(n17219) );
  INV_X1 U20539 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19104) );
  NAND3_X1 U20540 ( .A1(n17247), .A2(n17217), .A3(n19104), .ZN(n17218) );
  NAND4_X1 U20541 ( .A1(n17221), .A2(n17220), .A3(n17219), .A4(n17218), .ZN(
        P3_U2667) );
  AOI22_X1 U20542 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17244), .B1(
        n17266), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17235) );
  NAND2_X1 U20543 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17240) );
  AOI21_X1 U20544 ( .B1(n17222), .B2(n17240), .A(n17223), .ZN(n18170) );
  OAI21_X1 U20545 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17240), .A(
        n9958), .ZN(n17224) );
  XNOR2_X1 U20546 ( .A(n18170), .B(n17224), .ZN(n17228) );
  NAND2_X1 U20547 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n17225) );
  OAI21_X1 U20548 ( .B1(n17245), .B2(n17225), .A(n19102), .ZN(n17226) );
  AOI22_X1 U20549 ( .A1(n17229), .A2(n17228), .B1(n17227), .B2(n17226), .ZN(
        n17234) );
  OAI211_X1 U20550 ( .C1(n17238), .C2(n17552), .A(n17265), .B(n17230), .ZN(
        n17233) );
  INV_X1 U20551 ( .A(n19012), .ZN(n19027) );
  NOR2_X1 U20552 ( .A1(n19198), .A2(n19027), .ZN(n19018) );
  INV_X1 U20553 ( .A(n19018), .ZN(n17231) );
  AOI21_X1 U20554 ( .B1(n19175), .B2(n17231), .A(n10308), .ZN(n19170) );
  NAND2_X1 U20555 ( .A1(n19170), .A2(n19233), .ZN(n17232) );
  NAND4_X1 U20556 ( .A1(n17235), .A2(n17234), .A3(n17233), .A4(n17232), .ZN(
        P3_U2668) );
  AOI21_X1 U20557 ( .B1(n19186), .B2(n19033), .A(n19018), .ZN(n19182) );
  OAI21_X1 U20558 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17240), .ZN(n18181) );
  INV_X1 U20559 ( .A(n18181), .ZN(n17237) );
  AOI22_X1 U20560 ( .A1(n19182), .A2(n19233), .B1(n17237), .B2(n17236), .ZN(
        n17251) );
  INV_X1 U20561 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17571) );
  INV_X1 U20562 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17565) );
  NAND2_X1 U20563 ( .A1(n17571), .A2(n17565), .ZN(n17257) );
  AOI211_X1 U20564 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17257), .A(n17238), .B(
        n17258), .ZN(n17243) );
  OAI22_X1 U20565 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17240), .B1(
        n17239), .B2(n18181), .ZN(n17241) );
  OAI22_X1 U20566 ( .A1(n17259), .A2(n17559), .B1(n17255), .B2(n17241), .ZN(
        n17242) );
  AOI211_X1 U20567 ( .C1(n17244), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17243), .B(n17242), .ZN(n17250) );
  NOR2_X1 U20568 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17245), .ZN(n17253) );
  OAI21_X1 U20569 ( .B1(n17246), .B2(n17253), .A(P3_REIP_REG_2__SCAN_IN), .ZN(
        n17249) );
  NAND3_X1 U20570 ( .A1(n17247), .A2(P3_REIP_REG_1__SCAN_IN), .A3(n21303), 
        .ZN(n17248) );
  NAND4_X1 U20571 ( .A1(n17251), .A2(n17250), .A3(n17249), .A4(n17248), .ZN(
        P3_U2669) );
  NAND2_X1 U20572 ( .A1(n19033), .A2(n17252), .ZN(n19040) );
  INV_X1 U20573 ( .A(n19040), .ZN(n19189) );
  AOI21_X1 U20574 ( .B1(n19233), .B2(n19189), .A(n17253), .ZN(n17264) );
  OAI21_X1 U20575 ( .B1(n17256), .B2(n17255), .A(n17254), .ZN(n17261) );
  NAND2_X1 U20576 ( .A1(n17257), .A2(n17561), .ZN(n17567) );
  OAI22_X1 U20577 ( .A1(n17259), .A2(n17565), .B1(n17258), .B2(n17567), .ZN(
        n17260) );
  AOI221_X1 U20578 ( .B1(n17262), .B2(n9961), .C1(n17261), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17260), .ZN(n17263) );
  OAI211_X1 U20579 ( .C1(n17268), .C2(n19099), .A(n17264), .B(n17263), .ZN(
        P3_U2670) );
  NOR2_X1 U20580 ( .A1(n17266), .A2(n17265), .ZN(n17271) );
  AOI22_X1 U20581 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17267), .B1(n19233), 
        .B2(n19198), .ZN(n17270) );
  NAND3_X1 U20582 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19173), .A3(
        n17268), .ZN(n17269) );
  OAI211_X1 U20583 ( .C1(n17271), .C2(n17571), .A(n17270), .B(n17269), .ZN(
        P3_U2671) );
  INV_X1 U20584 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17272) );
  NOR2_X1 U20585 ( .A1(n17272), .A2(n17374), .ZN(n17347) );
  NOR4_X1 U20586 ( .A1(n17275), .A2(n17274), .A3(n17333), .A4(n17273), .ZN(
        n17276) );
  NAND4_X1 U20587 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17347), .A4(n17276), .ZN(n17279) );
  NOR2_X1 U20588 ( .A1(n17280), .A2(n17279), .ZN(n17295) );
  NAND2_X1 U20589 ( .A1(n17556), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17278) );
  NAND2_X1 U20590 ( .A1(n17295), .A2(n18589), .ZN(n17277) );
  OAI22_X1 U20591 ( .A1(n17295), .A2(n17278), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17277), .ZN(P3_U2672) );
  NAND2_X1 U20592 ( .A1(n17280), .A2(n17279), .ZN(n17281) );
  NAND2_X1 U20593 ( .A1(n17281), .A2(n17556), .ZN(n17294) );
  AOI22_X1 U20594 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20595 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17505), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U20596 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20597 ( .A1(n11673), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17282) );
  NAND4_X1 U20598 ( .A1(n17285), .A2(n17284), .A3(n17283), .A4(n17282), .ZN(
        n17291) );
  AOI22_X1 U20599 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U20600 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U20601 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20602 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17286) );
  NAND4_X1 U20603 ( .A1(n17289), .A2(n17288), .A3(n17287), .A4(n17286), .ZN(
        n17290) );
  NOR2_X1 U20604 ( .A1(n17291), .A2(n17290), .ZN(n17292) );
  XOR2_X1 U20605 ( .A(n17293), .B(n17292), .Z(n17583) );
  OAI22_X1 U20606 ( .A1(n17295), .A2(n17294), .B1(n17583), .B2(n17556), .ZN(
        P3_U2673) );
  AOI21_X1 U20607 ( .B1(n17297), .B2(n17302), .A(n17296), .ZN(n17593) );
  NAND2_X1 U20608 ( .A1(n17593), .A2(n17569), .ZN(n17298) );
  OAI221_X1 U20609 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17301), .C1(n17300), 
        .C2(n17299), .A(n17298), .ZN(P3_U2676) );
  INV_X1 U20610 ( .A(n17301), .ZN(n17305) );
  AOI21_X1 U20611 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17556), .A(n17310), .ZN(
        n17304) );
  OAI21_X1 U20612 ( .B1(n17306), .B2(n17303), .A(n17302), .ZN(n17601) );
  OAI22_X1 U20613 ( .A1(n17305), .A2(n17304), .B1(n17601), .B2(n17556), .ZN(
        P3_U2677) );
  AOI21_X1 U20614 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17556), .A(n17314), .ZN(
        n17309) );
  AOI21_X1 U20615 ( .B1(n17307), .B2(n17311), .A(n17306), .ZN(n17602) );
  INV_X1 U20616 ( .A(n17602), .ZN(n17308) );
  OAI22_X1 U20617 ( .A1(n17310), .A2(n17309), .B1(n17556), .B2(n17308), .ZN(
        P3_U2678) );
  AOI21_X1 U20618 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17556), .A(n17320), .ZN(
        n17313) );
  OAI21_X1 U20619 ( .B1(n17315), .B2(n17312), .A(n17311), .ZN(n17611) );
  OAI22_X1 U20620 ( .A1(n17314), .A2(n17313), .B1(n17556), .B2(n17611), .ZN(
        P3_U2679) );
  NOR2_X1 U20621 ( .A1(n17333), .A2(n17332), .ZN(n17336) );
  AOI21_X1 U20622 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17556), .A(n17336), .ZN(
        n17319) );
  AOI21_X1 U20623 ( .B1(n17317), .B2(n17316), .A(n17315), .ZN(n17612) );
  INV_X1 U20624 ( .A(n17612), .ZN(n17318) );
  OAI22_X1 U20625 ( .A1(n17320), .A2(n17319), .B1(n17556), .B2(n17318), .ZN(
        P3_U2680) );
  AOI22_X1 U20626 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9719), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n14519), .ZN(n17324) );
  AOI22_X1 U20627 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20628 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14517), .B1(
        n17504), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U20629 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11673), .B1(
        P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n10308), .ZN(n17321) );
  NAND4_X1 U20630 ( .A1(n17324), .A2(n17323), .A3(n17322), .A4(n17321), .ZN(
        n17331) );
  AOI22_X1 U20631 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20632 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17526), .B1(
        P3_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n17523), .ZN(n17328) );
  AOI22_X1 U20633 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n17503), .ZN(n17327) );
  AOI22_X1 U20634 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n14480), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17326) );
  NAND4_X1 U20635 ( .A1(n17329), .A2(n17328), .A3(n17327), .A4(n17326), .ZN(
        n17330) );
  NOR2_X1 U20636 ( .A1(n17331), .A2(n17330), .ZN(n17619) );
  OAI21_X1 U20637 ( .B1(n17333), .B2(n17569), .A(n17332), .ZN(n17334) );
  INV_X1 U20638 ( .A(n17334), .ZN(n17335) );
  OAI22_X1 U20639 ( .A1(n17619), .A2(n17556), .B1(n17336), .B2(n17335), .ZN(
        P3_U2681) );
  AOI22_X1 U20640 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17340) );
  AOI22_X1 U20641 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U20642 ( .A1(n9719), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20643 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17337) );
  NAND4_X1 U20644 ( .A1(n17340), .A2(n17339), .A3(n17338), .A4(n17337), .ZN(
        n17346) );
  AOI22_X1 U20645 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U20646 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20647 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20648 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17341) );
  NAND4_X1 U20649 ( .A1(n17344), .A2(n17343), .A3(n17342), .A4(n17341), .ZN(
        n17345) );
  NOR2_X1 U20650 ( .A1(n17346), .A2(n17345), .ZN(n17627) );
  NOR2_X1 U20651 ( .A1(n17569), .A2(n17347), .ZN(n17361) );
  AOI22_X1 U20652 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17361), .B1(n17349), 
        .B2(n17348), .ZN(n17350) );
  OAI21_X1 U20653 ( .B1(n17627), .B2(n17556), .A(n17350), .ZN(P3_U2682) );
  AOI22_X1 U20654 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U20655 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20656 ( .A1(n11704), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9731), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20657 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17351) );
  NAND4_X1 U20658 ( .A1(n17354), .A2(n17353), .A3(n17352), .A4(n17351), .ZN(
        n17360) );
  AOI22_X1 U20659 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U20660 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20661 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20662 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17355) );
  NAND4_X1 U20663 ( .A1(n17358), .A2(n17357), .A3(n17356), .A4(n17355), .ZN(
        n17359) );
  NOR2_X1 U20664 ( .A1(n17360), .A2(n17359), .ZN(n17631) );
  OAI21_X1 U20665 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17362), .A(n17361), .ZN(
        n17363) );
  OAI21_X1 U20666 ( .B1(n17631), .B2(n17556), .A(n17363), .ZN(P3_U2683) );
  AOI22_X1 U20667 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20668 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20669 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20670 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17364) );
  NAND4_X1 U20671 ( .A1(n17367), .A2(n17366), .A3(n17365), .A4(n17364), .ZN(
        n17373) );
  AOI22_X1 U20672 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U20673 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U20674 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20675 ( .A1(n14517), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17368) );
  NAND4_X1 U20676 ( .A1(n17371), .A2(n17370), .A3(n17369), .A4(n17368), .ZN(
        n17372) );
  NOR2_X1 U20677 ( .A1(n17373), .A2(n17372), .ZN(n17636) );
  OAI21_X1 U20678 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17375), .A(n17374), .ZN(
        n17376) );
  AOI22_X1 U20679 ( .A1(n17569), .A2(n17636), .B1(n17376), .B2(n17556), .ZN(
        P3_U2684) );
  NAND2_X1 U20680 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17377), .ZN(n17389) );
  AOI22_X1 U20681 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20682 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20683 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20684 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17378) );
  NAND4_X1 U20685 ( .A1(n17381), .A2(n17380), .A3(n17379), .A4(n17378), .ZN(
        n17387) );
  AOI22_X1 U20686 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9719), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20687 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20688 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20689 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17382) );
  NAND4_X1 U20690 ( .A1(n17385), .A2(n17384), .A3(n17383), .A4(n17382), .ZN(
        n17386) );
  NOR2_X1 U20691 ( .A1(n17387), .A2(n17386), .ZN(n17641) );
  OR4_X1 U20692 ( .A1(n17659), .A2(n17401), .A3(n17402), .A4(
        P3_EBX_REG_18__SCAN_IN), .ZN(n17388) );
  OAI221_X1 U20693 ( .B1(n17569), .B2(n17389), .C1(n17556), .C2(n17641), .A(
        n17388), .ZN(P3_U2685) );
  AOI22_X1 U20694 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U20695 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20696 ( .A1(n9719), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20697 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17390) );
  NAND4_X1 U20698 ( .A1(n17393), .A2(n17392), .A3(n17391), .A4(n17390), .ZN(
        n17399) );
  AOI22_X1 U20699 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20700 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20701 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20702 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17394) );
  NAND4_X1 U20703 ( .A1(n17397), .A2(n17396), .A3(n17395), .A4(n17394), .ZN(
        n17398) );
  NOR2_X1 U20704 ( .A1(n17399), .A2(n17398), .ZN(n17646) );
  OAI33_X1 U20705 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17659), .A3(n17402), 
        .B1(n17401), .B2(n17569), .B3(n17400), .ZN(n17403) );
  INV_X1 U20706 ( .A(n17403), .ZN(n17404) );
  OAI21_X1 U20707 ( .B1(n17646), .B2(n17556), .A(n17404), .ZN(P3_U2686) );
  AOI22_X1 U20708 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9719), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20709 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20710 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20711 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17405) );
  NAND4_X1 U20712 ( .A1(n17408), .A2(n17407), .A3(n17406), .A4(n17405), .ZN(
        n17414) );
  AOI22_X1 U20713 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20714 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20715 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20716 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17409) );
  NAND4_X1 U20717 ( .A1(n17412), .A2(n17411), .A3(n17410), .A4(n17409), .ZN(
        n17413) );
  NOR2_X1 U20718 ( .A1(n17414), .A2(n17413), .ZN(n17652) );
  INV_X1 U20719 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17416) );
  OAI33_X1 U20720 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17659), .A3(n17432), 
        .B1(n17416), .B2(n17569), .B3(n17415), .ZN(n17417) );
  INV_X1 U20721 ( .A(n17417), .ZN(n17418) );
  OAI21_X1 U20722 ( .B1(n17652), .B2(n17556), .A(n17418), .ZN(P3_U2687) );
  AOI22_X1 U20723 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20724 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U20725 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20726 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17419) );
  NAND4_X1 U20727 ( .A1(n17422), .A2(n17421), .A3(n17420), .A4(n17419), .ZN(
        n17429) );
  AOI22_X1 U20728 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20729 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9719), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20730 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U20731 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17424) );
  NAND4_X1 U20732 ( .A1(n17427), .A2(n17426), .A3(n17425), .A4(n17424), .ZN(
        n17428) );
  NOR2_X1 U20733 ( .A1(n17429), .A2(n17428), .ZN(n17657) );
  INV_X1 U20734 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17431) );
  NOR2_X1 U20735 ( .A1(n17430), .A2(n17539), .ZN(n17490) );
  NAND3_X1 U20736 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n17490), .ZN(n17471) );
  NOR2_X1 U20737 ( .A1(n17431), .A2(n17471), .ZN(n17472) );
  NAND2_X1 U20738 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17472), .ZN(n17459) );
  NOR2_X1 U20739 ( .A1(n17444), .A2(n17459), .ZN(n17447) );
  OAI211_X1 U20740 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17447), .A(n17432), .B(
        n17556), .ZN(n17433) );
  OAI21_X1 U20741 ( .B1(n17657), .B2(n17556), .A(n17433), .ZN(P3_U2688) );
  AOI22_X1 U20742 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n10331), .ZN(n17437) );
  AOI22_X1 U20743 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20744 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n17503), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20745 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n14519), .B1(
        P3_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n11673), .ZN(n17434) );
  NAND4_X1 U20746 ( .A1(n17437), .A2(n17436), .A3(n17435), .A4(n17434), .ZN(
        n17443) );
  AOI22_X1 U20747 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17504), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U20748 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17523), .B1(
        n9732), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20749 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14517), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n10308), .ZN(n17439) );
  AOI22_X1 U20750 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17438) );
  NAND4_X1 U20751 ( .A1(n17441), .A2(n17440), .A3(n17439), .A4(n17438), .ZN(
        n17442) );
  NOR2_X1 U20752 ( .A1(n17443), .A2(n17442), .ZN(n17664) );
  AOI21_X1 U20753 ( .B1(n17444), .B2(n17459), .A(n17569), .ZN(n17445) );
  INV_X1 U20754 ( .A(n17445), .ZN(n17446) );
  OAI22_X1 U20755 ( .A1(n17664), .A2(n17556), .B1(n17447), .B2(n17446), .ZN(
        P3_U2689) );
  AOI22_X1 U20756 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9732), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20757 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U20758 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U20759 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17449) );
  NAND4_X1 U20760 ( .A1(n17452), .A2(n17451), .A3(n17450), .A4(n17449), .ZN(
        n17458) );
  AOI22_X1 U20761 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20762 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20763 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17533), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20764 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17453) );
  NAND4_X1 U20765 ( .A1(n17456), .A2(n17455), .A3(n17454), .A4(n17453), .ZN(
        n17457) );
  NOR2_X1 U20766 ( .A1(n17458), .A2(n17457), .ZN(n17666) );
  OAI21_X1 U20767 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17472), .A(n17459), .ZN(
        n17460) );
  AOI22_X1 U20768 ( .A1(n17569), .A2(n17666), .B1(n17460), .B2(n17556), .ZN(
        P3_U2690) );
  AOI22_X1 U20769 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U20770 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17463) );
  AOI22_X1 U20771 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20772 ( .A1(n11656), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17461) );
  NAND4_X1 U20773 ( .A1(n17464), .A2(n17463), .A3(n17462), .A4(n17461), .ZN(
        n17470) );
  AOI22_X1 U20774 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9731), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20775 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U20776 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U20777 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17465) );
  NAND4_X1 U20778 ( .A1(n17468), .A2(n17467), .A3(n17466), .A4(n17465), .ZN(
        n17469) );
  NOR2_X1 U20779 ( .A1(n17470), .A2(n17469), .ZN(n17670) );
  NAND2_X1 U20780 ( .A1(n17556), .A2(n17471), .ZN(n17487) );
  NAND2_X1 U20781 ( .A1(n18589), .A2(n17472), .ZN(n17473) );
  OAI21_X1 U20782 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17487), .A(n17473), .ZN(
        n17474) );
  AOI21_X1 U20783 ( .B1(n17569), .B2(n17670), .A(n17474), .ZN(P3_U2691) );
  AOI22_X1 U20784 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14480), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U20785 ( .A1(n17504), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U20786 ( .A1(n17503), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20787 ( .B1(n17476), .B2(n21246), .A(n17475), .ZN(n17483) );
  AOI22_X1 U20788 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17477), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U20789 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17480) );
  AOI22_X1 U20790 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U20791 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17478) );
  NAND4_X1 U20792 ( .A1(n17481), .A2(n17480), .A3(n17479), .A4(n17478), .ZN(
        n17482) );
  AOI211_X1 U20793 ( .C1(n9718), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17483), .B(n17482), .ZN(n17484) );
  NAND3_X1 U20794 ( .A1(n17486), .A2(n17485), .A3(n17484), .ZN(n17673) );
  INV_X1 U20795 ( .A(n17673), .ZN(n17489) );
  AOI21_X1 U20796 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17490), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n17488) );
  OAI22_X1 U20797 ( .A1(n17489), .A2(n17556), .B1(n17488), .B2(n17487), .ZN(
        P3_U2692) );
  NAND2_X1 U20798 ( .A1(n18589), .A2(n17490), .ZN(n17502) );
  NOR2_X1 U20799 ( .A1(n17569), .A2(n17490), .ZN(n17518) );
  AOI22_X1 U20800 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U20801 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17504), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U20802 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U20803 ( .B1(n10309), .B2(n21174), .A(n17491), .ZN(n17497) );
  AOI22_X1 U20804 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U20805 ( .A1(n11671), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20806 ( .A1(n14517), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U20807 ( .A1(n9732), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17523), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17492) );
  NAND4_X1 U20808 ( .A1(n17495), .A2(n17494), .A3(n17493), .A4(n17492), .ZN(
        n17496) );
  AOI211_X1 U20809 ( .C1(n17325), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17497), .B(n17496), .ZN(n17498) );
  NAND3_X1 U20810 ( .A1(n17500), .A2(n17499), .A3(n17498), .ZN(n17676) );
  AOI22_X1 U20811 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17518), .B1(n17569), 
        .B2(n17676), .ZN(n17501) );
  OAI21_X1 U20812 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17502), .A(n17501), .ZN(
        P3_U2693) );
  AOI22_X1 U20813 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U20814 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17504), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U20815 ( .A1(n14480), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14519), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U20816 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17506) );
  NAND4_X1 U20817 ( .A1(n17509), .A2(n17508), .A3(n17507), .A4(n17506), .ZN(
        n17517) );
  AOI22_X1 U20818 ( .A1(n11671), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17515) );
  AOI22_X1 U20819 ( .A1(n11704), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17510), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U20820 ( .A1(n14517), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20821 ( .A1(n17511), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17512) );
  NAND4_X1 U20822 ( .A1(n17515), .A2(n17514), .A3(n17513), .A4(n17512), .ZN(
        n17516) );
  NOR2_X1 U20823 ( .A1(n17517), .A2(n17516), .ZN(n17681) );
  INV_X1 U20824 ( .A(n17539), .ZN(n17519) );
  OAI21_X1 U20825 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17519), .A(n17518), .ZN(
        n17520) );
  OAI21_X1 U20826 ( .B1(n17681), .B2(n17556), .A(n17520), .ZN(P3_U2694) );
  AOI22_X1 U20827 ( .A1(n17522), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17536) );
  AOI22_X1 U20828 ( .A1(n9731), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17535) );
  INV_X1 U20829 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21155) );
  AOI22_X1 U20830 ( .A1(n17523), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14517), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U20831 ( .B1(n17525), .B2(n21155), .A(n17524), .ZN(n17532) );
  AOI22_X1 U20832 ( .A1(n11671), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17526), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U20833 ( .A1(n17505), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10308), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17529) );
  AOI22_X1 U20834 ( .A1(n14520), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17528) );
  AOI22_X1 U20835 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11673), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17527) );
  NAND4_X1 U20836 ( .A1(n17530), .A2(n17529), .A3(n17528), .A4(n17527), .ZN(
        n17531) );
  AOI211_X1 U20837 ( .C1(n10331), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17532), .B(n17531), .ZN(n17534) );
  NAND3_X1 U20838 ( .A1(n17536), .A2(n17535), .A3(n17534), .ZN(n17684) );
  INV_X1 U20839 ( .A(n17684), .ZN(n17541) );
  NOR2_X1 U20840 ( .A1(n17537), .A2(n17566), .ZN(n17554) );
  NAND2_X1 U20841 ( .A1(n17538), .A2(n17554), .ZN(n17546) );
  NOR2_X1 U20842 ( .A1(n17542), .A2(n17546), .ZN(n17545) );
  OAI21_X1 U20843 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17545), .A(n17539), .ZN(
        n17540) );
  AOI22_X1 U20844 ( .A1(n17569), .A2(n17541), .B1(n17540), .B2(n17556), .ZN(
        P3_U2695) );
  OAI21_X1 U20845 ( .B1(n17542), .B2(n17569), .A(n17546), .ZN(n17543) );
  INV_X1 U20846 ( .A(n17543), .ZN(n17544) );
  INV_X1 U20847 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18593) );
  OAI22_X1 U20848 ( .A1(n17545), .A2(n17544), .B1(n18593), .B2(n17556), .ZN(
        P3_U2696) );
  AND2_X1 U20849 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17548), .ZN(n17550) );
  OAI21_X1 U20850 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17550), .A(n17546), .ZN(
        n17547) );
  AOI22_X1 U20851 ( .A1(n17569), .A2(n18584), .B1(n17547), .B2(n17556), .ZN(
        P3_U2697) );
  OAI21_X1 U20852 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17548), .A(n17556), .ZN(
        n17549) );
  OAI22_X1 U20853 ( .A1(n17550), .A2(n17549), .B1(n18577), .B2(n17556), .ZN(
        P3_U2698) );
  NAND2_X1 U20854 ( .A1(n17551), .A2(n17568), .ZN(n17555) );
  NOR2_X1 U20855 ( .A1(n17552), .A2(n17555), .ZN(n17558) );
  AOI21_X1 U20856 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17556), .A(n17558), .ZN(
        n17553) );
  INV_X1 U20857 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18571) );
  OAI22_X1 U20858 ( .A1(n17554), .A2(n17553), .B1(n18571), .B2(n17556), .ZN(
        P3_U2699) );
  INV_X1 U20859 ( .A(n17555), .ZN(n17563) );
  AOI21_X1 U20860 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17556), .A(n17563), .ZN(
        n17557) );
  OAI22_X1 U20861 ( .A1(n17558), .A2(n17557), .B1(n21246), .B2(n17556), .ZN(
        P3_U2700) );
  INV_X1 U20862 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18561) );
  OAI221_X1 U20863 ( .B1(n17561), .B2(n17560), .C1(n18589), .C2(n17560), .A(
        n17559), .ZN(n17562) );
  INV_X1 U20864 ( .A(n17562), .ZN(n17564) );
  AOI211_X1 U20865 ( .C1(n17569), .C2(n18561), .A(n17564), .B(n17563), .ZN(
        P3_U2701) );
  OAI222_X1 U20866 ( .A1(n17567), .A2(n17566), .B1(n17565), .B2(n17572), .C1(
        n21310), .C2(n17556), .ZN(P3_U2702) );
  AOI22_X1 U20867 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17569), .B1(
        n17568), .B2(n17571), .ZN(n17570) );
  OAI21_X1 U20868 ( .B1(n17572), .B2(n17571), .A(n17570), .ZN(P3_U2703) );
  INV_X1 U20869 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17727) );
  INV_X1 U20870 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17732) );
  INV_X1 U20871 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17834) );
  INV_X1 U20872 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17763) );
  INV_X1 U20873 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17765) );
  NAND4_X1 U20874 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n17690) );
  OR3_X1 U20875 ( .A1(n17763), .A2(n17765), .A3(n17690), .ZN(n17689) );
  INV_X1 U20876 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17829) );
  INV_X1 U20877 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17820) );
  INV_X1 U20878 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17814) );
  NAND2_X1 U20879 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17660) );
  NOR4_X1 U20880 ( .A1(n17829), .A2(n17820), .A3(n17814), .A4(n17660), .ZN(
        n17573) );
  NAND3_X1 U20881 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .ZN(n17617) );
  NAND3_X1 U20882 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .ZN(n17574) );
  NAND2_X1 U20883 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17614), .ZN(n17613) );
  NAND2_X1 U20884 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17580), .ZN(n17579) );
  NAND2_X1 U20885 ( .A1(n17579), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17577) );
  NAND2_X1 U20886 ( .A1(n17575), .A2(n17654), .ZN(n17618) );
  NAND2_X1 U20887 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17647), .ZN(n17576) );
  OAI221_X1 U20888 ( .B1(n17579), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17577), 
        .C2(n17654), .A(n17576), .ZN(P3_U2704) );
  NOR2_X2 U20889 ( .A1(n17578), .A2(n17719), .ZN(n17648) );
  AOI22_X1 U20890 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17647), .ZN(n17582) );
  OAI211_X1 U20891 ( .C1(n17580), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17719), .B(
        n17579), .ZN(n17581) );
  INV_X1 U20892 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18572) );
  AOI22_X1 U20893 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17648), .B1(n17716), .B2(
        n17584), .ZN(n17587) );
  OAI211_X1 U20894 ( .C1(n17588), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17719), .B(
        n17585), .ZN(n17586) );
  OAI211_X1 U20895 ( .C1(n17618), .C2(n18572), .A(n17587), .B(n17586), .ZN(
        P3_U2706) );
  AOI22_X1 U20896 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17647), .ZN(n17591) );
  AOI211_X1 U20897 ( .C1(n17727), .C2(n17594), .A(n17588), .B(n17654), .ZN(
        n17589) );
  INV_X1 U20898 ( .A(n17589), .ZN(n17590) );
  OAI211_X1 U20899 ( .C1(n17592), .C2(n17711), .A(n17591), .B(n17590), .ZN(
        P3_U2707) );
  INV_X1 U20900 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21126) );
  AOI22_X1 U20901 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17648), .B1(n17716), .B2(
        n17593), .ZN(n17597) );
  OAI211_X1 U20902 ( .C1(n17595), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17719), .B(
        n17594), .ZN(n17596) );
  OAI211_X1 U20903 ( .C1(n17618), .C2(n21126), .A(n17597), .B(n17596), .ZN(
        P3_U2708) );
  AOI22_X1 U20904 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17647), .ZN(n17600) );
  OAI211_X1 U20905 ( .C1(n17603), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17719), .B(
        n17598), .ZN(n17599) );
  OAI211_X1 U20906 ( .C1(n17601), .C2(n17711), .A(n17600), .B(n17599), .ZN(
        P3_U2709) );
  AOI22_X1 U20907 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17648), .B1(n17716), .B2(
        n17602), .ZN(n17606) );
  AOI211_X1 U20908 ( .C1(n17732), .C2(n17607), .A(n17603), .B(n17654), .ZN(
        n17604) );
  INV_X1 U20909 ( .A(n17604), .ZN(n17605) );
  OAI211_X1 U20910 ( .C1(n17618), .C2(n18551), .A(n17606), .B(n17605), .ZN(
        P3_U2710) );
  AOI22_X1 U20911 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17647), .ZN(n17610) );
  OAI211_X1 U20912 ( .C1(n17608), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17719), .B(
        n17607), .ZN(n17609) );
  OAI211_X1 U20913 ( .C1(n17611), .C2(n17711), .A(n17610), .B(n17609), .ZN(
        P3_U2711) );
  INV_X1 U20914 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19700) );
  AOI22_X1 U20915 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17648), .B1(n17716), .B2(
        n17612), .ZN(n17616) );
  OAI211_X1 U20916 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17614), .A(n17719), .B(
        n17613), .ZN(n17615) );
  OAI211_X1 U20917 ( .C1(n17618), .C2(n19700), .A(n17616), .B(n17615), .ZN(
        P3_U2712) );
  NOR3_X1 U20918 ( .A1(n17659), .A2(n17649), .A3(n17617), .ZN(n17632) );
  NAND2_X1 U20919 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17632), .ZN(n17628) );
  INV_X1 U20920 ( .A(n17628), .ZN(n17624) );
  NAND2_X1 U20921 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17624), .ZN(n17623) );
  NAND2_X1 U20922 ( .A1(n17623), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17622) );
  OAI22_X1 U20923 ( .A1(n17619), .A2(n17711), .B1(n18581), .B2(n17618), .ZN(
        n17620) );
  AOI21_X1 U20924 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17648), .A(n17620), .ZN(
        n17621) );
  OAI221_X1 U20925 ( .B1(n17623), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17622), 
        .C2(n17654), .A(n17621), .ZN(P3_U2713) );
  AOI22_X1 U20926 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17647), .ZN(n17626) );
  OAI211_X1 U20927 ( .C1(n17624), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17719), .B(
        n17623), .ZN(n17625) );
  OAI211_X1 U20928 ( .C1(n17627), .C2(n17711), .A(n17626), .B(n17625), .ZN(
        P3_U2714) );
  AOI22_X1 U20929 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17647), .ZN(n17630) );
  OAI211_X1 U20930 ( .C1(n17632), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17719), .B(
        n17628), .ZN(n17629) );
  OAI211_X1 U20931 ( .C1(n17631), .C2(n17711), .A(n17630), .B(n17629), .ZN(
        P3_U2715) );
  AOI22_X1 U20932 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17647), .ZN(n17635) );
  INV_X1 U20933 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17743) );
  INV_X1 U20934 ( .A(n17649), .ZN(n17643) );
  NAND2_X1 U20935 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17643), .ZN(n17642) );
  NAND2_X1 U20936 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17638), .ZN(n17637) );
  AOI211_X1 U20937 ( .C1(n17743), .C2(n17637), .A(n17632), .B(n17654), .ZN(
        n17633) );
  INV_X1 U20938 ( .A(n17633), .ZN(n17634) );
  OAI211_X1 U20939 ( .C1(n17636), .C2(n17711), .A(n17635), .B(n17634), .ZN(
        P3_U2716) );
  AOI22_X1 U20940 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17647), .ZN(n17640) );
  OAI211_X1 U20941 ( .C1(n17638), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17719), .B(
        n17637), .ZN(n17639) );
  OAI211_X1 U20942 ( .C1(n17641), .C2(n17711), .A(n17640), .B(n17639), .ZN(
        P3_U2717) );
  AOI22_X1 U20943 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17647), .ZN(n17645) );
  OAI211_X1 U20944 ( .C1(n17643), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17719), .B(
        n17642), .ZN(n17644) );
  OAI211_X1 U20945 ( .C1(n17646), .C2(n17711), .A(n17645), .B(n17644), .ZN(
        P3_U2718) );
  AOI22_X1 U20946 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17648), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17647), .ZN(n17651) );
  OAI211_X1 U20947 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17653), .A(n17719), .B(
        n17649), .ZN(n17650) );
  OAI211_X1 U20948 ( .C1(n17652), .C2(n17711), .A(n17651), .B(n17650), .ZN(
        P3_U2719) );
  AOI211_X1 U20949 ( .C1(n17834), .C2(n17661), .A(n17654), .B(n17653), .ZN(
        n17655) );
  AOI21_X1 U20950 ( .B1(n17717), .B2(BUF2_REG_15__SCAN_IN), .A(n17655), .ZN(
        n17656) );
  OAI21_X1 U20951 ( .B1(n17657), .B2(n17711), .A(n17656), .ZN(P3_U2720) );
  NOR3_X1 U20952 ( .A1(n17689), .A2(n17814), .A3(n17718), .ZN(n17680) );
  NAND2_X1 U20953 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17680), .ZN(n17678) );
  INV_X1 U20954 ( .A(n17678), .ZN(n17683) );
  NAND2_X1 U20955 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17683), .ZN(n17675) );
  NOR2_X1 U20956 ( .A1(n17820), .A2(n17675), .ZN(n17669) );
  INV_X1 U20957 ( .A(n17669), .ZN(n17665) );
  NOR2_X1 U20958 ( .A1(n17660), .A2(n17665), .ZN(n17667) );
  AOI22_X1 U20959 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17717), .B1(n17667), .B2(
        n17829), .ZN(n17663) );
  NAND3_X1 U20960 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17719), .A3(n17661), 
        .ZN(n17662) );
  OAI211_X1 U20961 ( .C1(n17664), .C2(n17711), .A(n17663), .B(n17662), .ZN(
        P3_U2721) );
  INV_X1 U20962 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17827) );
  INV_X1 U20963 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17755) );
  NOR2_X1 U20964 ( .A1(n17755), .A2(n17665), .ZN(n17672) );
  AOI21_X1 U20965 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17719), .A(n17672), .ZN(
        n17668) );
  OAI222_X1 U20966 ( .A1(n17714), .A2(n17827), .B1(n17668), .B2(n17667), .C1(
        n17711), .C2(n17666), .ZN(P3_U2722) );
  INV_X1 U20967 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17823) );
  AOI21_X1 U20968 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17719), .A(n17669), .ZN(
        n17671) );
  OAI222_X1 U20969 ( .A1(n17714), .A2(n17823), .B1(n17672), .B2(n17671), .C1(
        n17711), .C2(n17670), .ZN(P3_U2723) );
  NAND2_X1 U20970 ( .A1(n17719), .A2(n17675), .ZN(n17679) );
  AOI22_X1 U20971 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17717), .B1(n17716), .B2(
        n17673), .ZN(n17674) );
  OAI221_X1 U20972 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17675), .C1(n17820), 
        .C2(n17679), .A(n17674), .ZN(P3_U2724) );
  INV_X1 U20973 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17758) );
  AOI22_X1 U20974 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17717), .B1(n17716), .B2(
        n17676), .ZN(n17677) );
  OAI221_X1 U20975 ( .B1(n17679), .B2(n17758), .C1(n17679), .C2(n17678), .A(
        n17677), .ZN(P3_U2725) );
  INV_X1 U20976 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17816) );
  AOI21_X1 U20977 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17719), .A(n17680), .ZN(
        n17682) );
  OAI222_X1 U20978 ( .A1(n17714), .A2(n17816), .B1(n17683), .B2(n17682), .C1(
        n17711), .C2(n17681), .ZN(P3_U2726) );
  AOI22_X1 U20979 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17717), .B1(n17716), .B2(
        n17684), .ZN(n17688) );
  INV_X1 U20980 ( .A(n17686), .ZN(n17685) );
  OAI221_X1 U20981 ( .B1(n17686), .B2(P3_EAX_REG_8__SCAN_IN), .C1(n17685), 
        .C2(n17814), .A(n17719), .ZN(n17687) );
  NAND2_X1 U20982 ( .A1(n17688), .A2(n17687), .ZN(P3_U2727) );
  INV_X1 U20983 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18586) );
  NOR2_X1 U20984 ( .A1(n17689), .A2(n17718), .ZN(n17693) );
  NOR2_X1 U20985 ( .A1(n17690), .A2(n17718), .ZN(n17699) );
  AOI22_X1 U20986 ( .A1(n17699), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17719), .ZN(n17692) );
  OAI222_X1 U20987 ( .A1(n17714), .A2(n18586), .B1(n17693), .B2(n17692), .C1(
        n17711), .C2(n17691), .ZN(P3_U2728) );
  INV_X1 U20988 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18579) );
  AND2_X1 U20989 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17699), .ZN(n17696) );
  AOI21_X1 U20990 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17719), .A(n17699), .ZN(
        n17695) );
  OAI222_X1 U20991 ( .A1(n18579), .A2(n17714), .B1(n17696), .B2(n17695), .C1(
        n17711), .C2(n17694), .ZN(P3_U2729) );
  INV_X1 U20992 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18573) );
  INV_X1 U20993 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17769) );
  INV_X1 U20994 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17775) );
  NOR2_X1 U20995 ( .A1(n17775), .A2(n17718), .ZN(n17713) );
  NAND2_X1 U20996 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17713), .ZN(n17700) );
  NOR2_X1 U20997 ( .A1(n17769), .A2(n17700), .ZN(n17704) );
  AOI21_X1 U20998 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17719), .A(n17704), .ZN(
        n17698) );
  OAI222_X1 U20999 ( .A1(n18573), .A2(n17714), .B1(n17699), .B2(n17698), .C1(
        n17711), .C2(n17697), .ZN(P3_U2730) );
  INV_X1 U21000 ( .A(n17700), .ZN(n17707) );
  AOI21_X1 U21001 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17719), .A(n17707), .ZN(
        n17703) );
  INV_X1 U21002 ( .A(n17701), .ZN(n17702) );
  OAI222_X1 U21003 ( .A1(n18567), .A2(n17714), .B1(n17704), .B2(n17703), .C1(
        n17711), .C2(n17702), .ZN(P3_U2731) );
  INV_X1 U21004 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18562) );
  AOI21_X1 U21005 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17719), .A(n17713), .ZN(
        n17706) );
  OAI222_X1 U21006 ( .A1(n18562), .A2(n17714), .B1(n17707), .B2(n17706), .C1(
        n17711), .C2(n17705), .ZN(P3_U2732) );
  INV_X1 U21007 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18555) );
  AOI21_X1 U21008 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17719), .A(n17708), .ZN(
        n17712) );
  INV_X1 U21009 ( .A(n17709), .ZN(n17710) );
  OAI222_X1 U21010 ( .A1(n18555), .A2(n17714), .B1(n17713), .B2(n17712), .C1(
        n17711), .C2(n17710), .ZN(P3_U2733) );
  AOI22_X1 U21011 ( .A1(n17717), .A2(BUF2_REG_1__SCAN_IN), .B1(n17716), .B2(
        n17715), .ZN(n17722) );
  OAI211_X1 U21012 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17720), .A(n17719), .B(
        n17718), .ZN(n17721) );
  NAND2_X1 U21013 ( .A1(n17722), .A2(n17721), .ZN(P3_U2734) );
  NAND2_X1 U21014 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17921), .ZN(n17772) );
  INV_X2 U21015 ( .A(n17772), .ZN(n17778) );
  AND2_X1 U21016 ( .A1(n17773), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21017 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17803) );
  NOR2_X1 U21018 ( .A1(n17780), .A2(n18547), .ZN(n17729) );
  AOI22_X1 U21019 ( .A1(n17778), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17724) );
  OAI21_X1 U21020 ( .B1(n17803), .B2(n17748), .A(n17724), .ZN(P3_U2737) );
  AOI22_X1 U21021 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(n17777), .B1(n17778), 
        .B2(P3_UWORD_REG_13__SCAN_IN), .ZN(n17725) );
  OAI21_X1 U21022 ( .B1(n9862), .B2(n17748), .A(n17725), .ZN(P3_U2738) );
  AOI22_X1 U21023 ( .A1(n17778), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17726) );
  OAI21_X1 U21024 ( .B1(n17727), .B2(n17748), .A(n17726), .ZN(P3_U2739) );
  INV_X1 U21025 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U21026 ( .A1(n17778), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17728) );
  OAI21_X1 U21027 ( .B1(n17799), .B2(n17748), .A(n17728), .ZN(P3_U2740) );
  INV_X1 U21028 ( .A(P3_UWORD_REG_10__SCAN_IN), .ZN(n21184) );
  AOI22_X1 U21029 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17729), .B1(n17773), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17730) );
  OAI21_X1 U21030 ( .B1(n21184), .B2(n17772), .A(n17730), .ZN(P3_U2741) );
  AOI22_X1 U21031 ( .A1(n17778), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17731) );
  OAI21_X1 U21032 ( .B1(n17732), .B2(n17748), .A(n17731), .ZN(P3_U2742) );
  INV_X1 U21033 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17795) );
  AOI22_X1 U21034 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(n17777), .B1(n17778), 
        .B2(P3_UWORD_REG_8__SCAN_IN), .ZN(n17733) );
  OAI21_X1 U21035 ( .B1(n17795), .B2(n17748), .A(n17733), .ZN(P3_U2743) );
  INV_X1 U21036 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U21037 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(n17777), .B1(n17778), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n17734) );
  OAI21_X1 U21038 ( .B1(n17735), .B2(n17748), .A(n17734), .ZN(P3_U2744) );
  INV_X1 U21039 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17737) );
  AOI22_X1 U21040 ( .A1(n17778), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17736) );
  OAI21_X1 U21041 ( .B1(n17737), .B2(n17748), .A(n17736), .ZN(P3_U2745) );
  INV_X1 U21042 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U21043 ( .A1(n17778), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17738) );
  OAI21_X1 U21044 ( .B1(n17739), .B2(n17748), .A(n17738), .ZN(P3_U2746) );
  INV_X1 U21045 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U21046 ( .A1(n17778), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17740) );
  OAI21_X1 U21047 ( .B1(n17741), .B2(n17748), .A(n17740), .ZN(P3_U2747) );
  AOI22_X1 U21048 ( .A1(n17778), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17742) );
  OAI21_X1 U21049 ( .B1(n17743), .B2(n17748), .A(n17742), .ZN(P3_U2748) );
  INV_X1 U21050 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17745) );
  AOI22_X1 U21051 ( .A1(n17778), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17744) );
  OAI21_X1 U21052 ( .B1(n17745), .B2(n17748), .A(n17744), .ZN(P3_U2749) );
  INV_X1 U21053 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U21054 ( .A1(n17778), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17746) );
  OAI21_X1 U21055 ( .B1(n17787), .B2(n17748), .A(n17746), .ZN(P3_U2750) );
  INV_X1 U21056 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U21057 ( .A1(n17778), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17747) );
  OAI21_X1 U21058 ( .B1(n17749), .B2(n17748), .A(n17747), .ZN(P3_U2751) );
  AOI22_X1 U21059 ( .A1(n17778), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17750) );
  OAI21_X1 U21060 ( .B1(n17834), .B2(n17780), .A(n17750), .ZN(P3_U2752) );
  AOI22_X1 U21061 ( .A1(n17778), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17751) );
  OAI21_X1 U21062 ( .B1(n17829), .B2(n17780), .A(n17751), .ZN(P3_U2753) );
  INV_X1 U21063 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17753) );
  AOI22_X1 U21064 ( .A1(n17778), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17752) );
  OAI21_X1 U21065 ( .B1(n17753), .B2(n17780), .A(n17752), .ZN(P3_U2754) );
  AOI22_X1 U21066 ( .A1(n17778), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17754) );
  OAI21_X1 U21067 ( .B1(n17755), .B2(n17780), .A(n17754), .ZN(P3_U2755) );
  AOI22_X1 U21068 ( .A1(n17778), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17756) );
  OAI21_X1 U21069 ( .B1(n17820), .B2(n17780), .A(n17756), .ZN(P3_U2756) );
  AOI22_X1 U21070 ( .A1(n17778), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17757) );
  OAI21_X1 U21071 ( .B1(n17758), .B2(n17780), .A(n17757), .ZN(P3_U2757) );
  INV_X1 U21072 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17760) );
  AOI22_X1 U21073 ( .A1(n17778), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17759) );
  OAI21_X1 U21074 ( .B1(n17760), .B2(n17780), .A(n17759), .ZN(P3_U2758) );
  AOI22_X1 U21075 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(n17777), .B1(n17778), 
        .B2(P3_LWORD_REG_8__SCAN_IN), .ZN(n17761) );
  OAI21_X1 U21076 ( .B1(n17814), .B2(n17780), .A(n17761), .ZN(P3_U2759) );
  AOI22_X1 U21077 ( .A1(n17778), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17762) );
  OAI21_X1 U21078 ( .B1(n17763), .B2(n17780), .A(n17762), .ZN(P3_U2760) );
  AOI22_X1 U21079 ( .A1(n17778), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17764) );
  OAI21_X1 U21080 ( .B1(n17765), .B2(n17780), .A(n17764), .ZN(P3_U2761) );
  INV_X1 U21081 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U21082 ( .A1(n17778), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17766) );
  OAI21_X1 U21083 ( .B1(n17767), .B2(n17780), .A(n17766), .ZN(P3_U2762) );
  AOI22_X1 U21084 ( .A1(n17778), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17768) );
  OAI21_X1 U21085 ( .B1(n17769), .B2(n17780), .A(n17768), .ZN(P3_U2763) );
  INV_X1 U21086 ( .A(P3_LWORD_REG_3__SCAN_IN), .ZN(n21111) );
  AOI22_X1 U21087 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17770), .B1(n17777), .B2(
        P3_DATAO_REG_3__SCAN_IN), .ZN(n17771) );
  OAI21_X1 U21088 ( .B1(n21111), .B2(n17772), .A(n17771), .ZN(P3_U2764) );
  AOI22_X1 U21089 ( .A1(n17778), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17773), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17774) );
  OAI21_X1 U21090 ( .B1(n17775), .B2(n17780), .A(n17774), .ZN(P3_U2765) );
  INV_X1 U21091 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17806) );
  AOI22_X1 U21092 ( .A1(n17778), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17776) );
  OAI21_X1 U21093 ( .B1(n17806), .B2(n17780), .A(n17776), .ZN(P3_U2766) );
  AOI22_X1 U21094 ( .A1(n17778), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17777), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17779) );
  OAI21_X1 U21095 ( .B1(n21141), .B2(n17780), .A(n17779), .ZN(P3_U2767) );
  AOI211_X1 U21096 ( .C1(n19216), .C2(n19215), .A(n17781), .B(n17784), .ZN(
        n17782) );
  INV_X2 U21097 ( .A(n17782), .ZN(n17830) );
  INV_X1 U21098 ( .A(n17783), .ZN(n19062) );
  AOI22_X1 U21099 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17824), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17830), .ZN(n17785) );
  OAI21_X1 U21100 ( .B1(n21110), .B2(n17826), .A(n17785), .ZN(P3_U2768) );
  INV_X1 U21101 ( .A(n17824), .ZN(n17833) );
  AOI22_X1 U21102 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17831), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17830), .ZN(n17786) );
  OAI21_X1 U21103 ( .B1(n17787), .B2(n17833), .A(n17786), .ZN(P3_U2769) );
  AOI22_X1 U21104 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17830), .ZN(n17788) );
  OAI21_X1 U21105 ( .B1(n18555), .B2(n17826), .A(n17788), .ZN(P3_U2770) );
  AOI22_X1 U21106 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17824), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17830), .ZN(n17789) );
  OAI21_X1 U21107 ( .B1(n18562), .B2(n17826), .A(n17789), .ZN(P3_U2771) );
  AOI22_X1 U21108 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17824), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17830), .ZN(n17790) );
  OAI21_X1 U21109 ( .B1(n18567), .B2(n17826), .A(n17790), .ZN(P3_U2772) );
  AOI22_X1 U21110 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17830), .ZN(n17791) );
  OAI21_X1 U21111 ( .B1(n18573), .B2(n17826), .A(n17791), .ZN(P3_U2773) );
  AOI22_X1 U21112 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17824), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17830), .ZN(n17792) );
  OAI21_X1 U21113 ( .B1(n18579), .B2(n17826), .A(n17792), .ZN(P3_U2774) );
  AOI22_X1 U21114 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17824), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17830), .ZN(n17793) );
  OAI21_X1 U21115 ( .B1(n18586), .B2(n17826), .A(n17793), .ZN(P3_U2775) );
  AOI22_X1 U21116 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17831), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17830), .ZN(n17794) );
  OAI21_X1 U21117 ( .B1(n17795), .B2(n17833), .A(n17794), .ZN(P3_U2776) );
  AOI22_X1 U21118 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17830), .ZN(n17796) );
  OAI21_X1 U21119 ( .B1(n17816), .B2(n17826), .A(n17796), .ZN(P3_U2777) );
  INV_X1 U21120 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17818) );
  AOI22_X1 U21121 ( .A1(P3_UWORD_REG_10__SCAN_IN), .A2(n17830), .B1(
        P3_EAX_REG_26__SCAN_IN), .B2(n17821), .ZN(n17797) );
  OAI21_X1 U21122 ( .B1(n17818), .B2(n17826), .A(n17797), .ZN(P3_U2778) );
  AOI22_X1 U21123 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17831), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17830), .ZN(n17798) );
  OAI21_X1 U21124 ( .B1(n17799), .B2(n17833), .A(n17798), .ZN(P3_U2779) );
  AOI22_X1 U21125 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17824), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17830), .ZN(n17800) );
  OAI21_X1 U21126 ( .B1(n17823), .B2(n17826), .A(n17800), .ZN(P3_U2780) );
  AOI22_X1 U21127 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17830), .ZN(n17801) );
  OAI21_X1 U21128 ( .B1(n17827), .B2(n17826), .A(n17801), .ZN(P3_U2781) );
  AOI22_X1 U21129 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17831), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17830), .ZN(n17802) );
  OAI21_X1 U21130 ( .B1(n17803), .B2(n17833), .A(n17802), .ZN(P3_U2782) );
  AOI22_X1 U21131 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17824), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17830), .ZN(n17804) );
  OAI21_X1 U21132 ( .B1(n21110), .B2(n17826), .A(n17804), .ZN(P3_U2783) );
  AOI22_X1 U21133 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17831), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17830), .ZN(n17805) );
  OAI21_X1 U21134 ( .B1(n17806), .B2(n17833), .A(n17805), .ZN(P3_U2784) );
  AOI22_X1 U21135 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17824), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17830), .ZN(n17807) );
  OAI21_X1 U21136 ( .B1(n18555), .B2(n17826), .A(n17807), .ZN(P3_U2785) );
  AOI22_X1 U21137 ( .A1(P3_LWORD_REG_3__SCAN_IN), .A2(n17830), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n17821), .ZN(n17808) );
  OAI21_X1 U21138 ( .B1(n18562), .B2(n17826), .A(n17808), .ZN(P3_U2786) );
  AOI22_X1 U21139 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17830), .ZN(n17809) );
  OAI21_X1 U21140 ( .B1(n18567), .B2(n17826), .A(n17809), .ZN(P3_U2787) );
  AOI22_X1 U21141 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17830), .ZN(n17810) );
  OAI21_X1 U21142 ( .B1(n18573), .B2(n17826), .A(n17810), .ZN(P3_U2788) );
  AOI22_X1 U21143 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17830), .ZN(n17811) );
  OAI21_X1 U21144 ( .B1(n18579), .B2(n17826), .A(n17811), .ZN(P3_U2789) );
  AOI22_X1 U21145 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17830), .ZN(n17812) );
  OAI21_X1 U21146 ( .B1(n18586), .B2(n17826), .A(n17812), .ZN(P3_U2790) );
  AOI22_X1 U21147 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17831), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17830), .ZN(n17813) );
  OAI21_X1 U21148 ( .B1(n17814), .B2(n17833), .A(n17813), .ZN(P3_U2791) );
  AOI22_X1 U21149 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17824), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17830), .ZN(n17815) );
  OAI21_X1 U21150 ( .B1(n17816), .B2(n17826), .A(n17815), .ZN(P3_U2792) );
  AOI22_X1 U21151 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17830), .ZN(n17817) );
  OAI21_X1 U21152 ( .B1(n17818), .B2(n17826), .A(n17817), .ZN(P3_U2793) );
  AOI22_X1 U21153 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17831), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17830), .ZN(n17819) );
  OAI21_X1 U21154 ( .B1(n17820), .B2(n17833), .A(n17819), .ZN(P3_U2794) );
  AOI22_X1 U21155 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17830), .ZN(n17822) );
  OAI21_X1 U21156 ( .B1(n17823), .B2(n17826), .A(n17822), .ZN(P3_U2795) );
  AOI22_X1 U21157 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17824), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17830), .ZN(n17825) );
  OAI21_X1 U21158 ( .B1(n17827), .B2(n17826), .A(n17825), .ZN(P3_U2796) );
  AOI22_X1 U21159 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17831), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17830), .ZN(n17828) );
  OAI21_X1 U21160 ( .B1(n17829), .B2(n17833), .A(n17828), .ZN(P3_U2797) );
  AOI22_X1 U21161 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17831), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17830), .ZN(n17832) );
  OAI21_X1 U21162 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(P3_U2798) );
  OAI21_X1 U21163 ( .B1(n17837), .B2(n17836), .A(n17835), .ZN(n17852) );
  OAI21_X1 U21164 ( .B1(n17838), .B2(n19080), .A(n9733), .ZN(n17839) );
  AOI21_X1 U21165 ( .B1(n18031), .B2(n17842), .A(n17839), .ZN(n17870) );
  OAI21_X1 U21166 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17950), .A(
        n17870), .ZN(n17854) );
  NOR2_X1 U21167 ( .A1(n18111), .A2(n18143), .ZN(n17943) );
  OAI22_X1 U21168 ( .A1(n18211), .A2(n18202), .B1(n17840), .B2(n18072), .ZN(
        n17872) );
  NOR2_X1 U21169 ( .A1(n21186), .A2(n17872), .ZN(n17841) );
  NOR3_X1 U21170 ( .A1(n17943), .A2(n17841), .A3(n17849), .ZN(n17848) );
  NOR2_X1 U21171 ( .A1(n18028), .A2(n17842), .ZN(n17858) );
  OAI211_X1 U21172 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17858), .B(n17843), .ZN(n17844) );
  OAI211_X1 U21173 ( .C1(n18035), .C2(n17846), .A(n17845), .B(n17844), .ZN(
        n17847) );
  AOI211_X1 U21174 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17854), .A(
        n17848), .B(n17847), .ZN(n17851) );
  NAND3_X1 U21175 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17859), .A3(
        n17849), .ZN(n17850) );
  OAI211_X1 U21176 ( .C1(n17979), .C2(n17852), .A(n17851), .B(n17850), .ZN(
        P3_U2802) );
  AOI22_X1 U21177 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17854), .B1(
        n18050), .B2(n17853), .ZN(n17862) );
  OAI21_X1 U21178 ( .B1(n18109), .B2(n17856), .A(n17855), .ZN(n18216) );
  AOI22_X1 U21179 ( .A1(n18110), .A2(n18216), .B1(n17858), .B2(n17857), .ZN(
        n17861) );
  AOI22_X1 U21180 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17872), .B1(
        n17859), .B2(n21186), .ZN(n17860) );
  NAND2_X1 U21181 ( .A1(n18523), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18218) );
  NAND4_X1 U21182 ( .A1(n17862), .A2(n17861), .A3(n17860), .A4(n18218), .ZN(
        P3_U2803) );
  AOI21_X1 U21183 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17864), .A(
        n17863), .ZN(n18226) );
  INV_X1 U21184 ( .A(n17865), .ZN(n17873) );
  AOI21_X1 U21185 ( .B1(n18585), .B2(n17866), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17869) );
  OAI21_X1 U21186 ( .B1(n18050), .B2(n17980), .A(n17867), .ZN(n17868) );
  NAND2_X1 U21187 ( .A1(n18523), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18224) );
  OAI211_X1 U21188 ( .C1(n17870), .C2(n17869), .A(n17868), .B(n18224), .ZN(
        n17871) );
  AOI221_X1 U21189 ( .B1(n17873), .B2(n18212), .C1(n17872), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17871), .ZN(n17874) );
  OAI21_X1 U21190 ( .B1(n18226), .B2(n17979), .A(n17874), .ZN(P3_U2804) );
  NAND2_X1 U21191 ( .A1(n18585), .A2(n17875), .ZN(n17896) );
  OAI211_X1 U21192 ( .C1(n17876), .C2(n19080), .A(n9733), .B(n17896), .ZN(
        n17900) );
  AOI22_X1 U21193 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17900), .B1(
        n18050), .B2(n17877), .ZN(n17887) );
  XOR2_X1 U21194 ( .A(n17878), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18238) );
  XOR2_X1 U21195 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17879), .Z(
        n18234) );
  OAI21_X1 U21196 ( .B1(n18107), .B2(n17881), .A(n17880), .ZN(n17882) );
  XOR2_X1 U21197 ( .A(n17882), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18235) );
  OAI22_X1 U21198 ( .A1(n18202), .A2(n18234), .B1(n17979), .B2(n18235), .ZN(
        n17883) );
  AOI21_X1 U21199 ( .B1(n18111), .B2(n18238), .A(n17883), .ZN(n17886) );
  NAND2_X1 U21200 ( .A1(n18523), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18233) );
  NOR2_X1 U21201 ( .A1(n18028), .A2(n17875), .ZN(n17888) );
  OAI211_X1 U21202 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17888), .B(n17884), .ZN(n17885) );
  NAND4_X1 U21203 ( .A1(n17887), .A2(n17886), .A3(n18233), .A4(n17885), .ZN(
        P3_U2805) );
  NOR2_X1 U21204 ( .A1(n18529), .A2(n19144), .ZN(n18248) );
  AOI221_X1 U21205 ( .B1(n17888), .B2(n21279), .C1(n17900), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18248), .ZN(n17894) );
  AOI21_X1 U21206 ( .B1(n18263), .B2(n18251), .A(n18072), .ZN(n17910) );
  AOI21_X1 U21207 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18240), .A(
        n18202), .ZN(n17911) );
  NAND2_X1 U21208 ( .A1(n18251), .A2(n17976), .ZN(n17891) );
  AOI21_X1 U21209 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17890), .A(
        n17889), .ZN(n18254) );
  OAI22_X1 U21210 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17891), .B1(
        n18254), .B2(n17979), .ZN(n17892) );
  AOI221_X1 U21211 ( .B1(n17910), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), 
        .C1(n17911), .C2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n17892), .ZN(
        n17893) );
  OAI211_X1 U21212 ( .C1(n18035), .C2(n17895), .A(n17894), .B(n17893), .ZN(
        P3_U2806) );
  INV_X1 U21213 ( .A(n17896), .ZN(n17901) );
  OAI21_X1 U21214 ( .B1(n17950), .B2(n17898), .A(n17897), .ZN(n17899) );
  AOI22_X1 U21215 ( .A1(n17902), .A2(n17901), .B1(n17900), .B2(n17899), .ZN(
        n17915) );
  AOI22_X1 U21216 ( .A1(n18523), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18050), 
        .B2(n17903), .ZN(n17914) );
  AOI22_X1 U21217 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18107), .B1(
        n17904), .B2(n17916), .ZN(n17905) );
  NAND2_X1 U21218 ( .A1(n17944), .A2(n17905), .ZN(n17906) );
  XOR2_X1 U21219 ( .A(n17906), .B(n17908), .Z(n18256) );
  NAND2_X1 U21220 ( .A1(n17908), .A2(n17907), .ZN(n17909) );
  AOI22_X1 U21221 ( .A1(n18110), .A2(n18256), .B1(n17910), .B2(n17909), .ZN(
        n17913) );
  OAI21_X1 U21222 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18240), .A(
        n17911), .ZN(n17912) );
  NAND4_X1 U21223 ( .A1(n17915), .A2(n17914), .A3(n17913), .A4(n17912), .ZN(
        P3_U2807) );
  INV_X1 U21224 ( .A(n17916), .ZN(n17918) );
  NAND2_X1 U21225 ( .A1(n18317), .A2(n17917), .ZN(n18261) );
  INV_X1 U21226 ( .A(n18261), .ZN(n18269) );
  OAI221_X1 U21227 ( .B1(n17918), .B2(n18269), .C1(n17918), .C2(n17990), .A(
        n17944), .ZN(n17919) );
  XOR2_X1 U21228 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17919), .Z(
        n18278) );
  NOR2_X1 U21229 ( .A1(n18529), .A2(n21123), .ZN(n18260) );
  AOI22_X1 U21230 ( .A1(n17921), .A2(n17920), .B1(n18031), .B2(n17924), .ZN(
        n17922) );
  NAND2_X1 U21231 ( .A1(n17922), .A2(n9733), .ZN(n17948) );
  AOI21_X1 U21232 ( .B1(n17980), .B2(n17923), .A(n17948), .ZN(n17932) );
  OR2_X1 U21233 ( .A1(n17924), .A2(n18028), .ZN(n17934) );
  OAI21_X1 U21234 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17925), .ZN(n17926) );
  OAI22_X1 U21235 ( .A1(n17932), .A2(n17927), .B1(n17934), .B2(n17926), .ZN(
        n17928) );
  AOI211_X1 U21236 ( .C1(n17929), .C2(n18050), .A(n18260), .B(n17928), .ZN(
        n17931) );
  INV_X1 U21237 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18270) );
  NOR2_X1 U21238 ( .A1(n18263), .A2(n18072), .ZN(n18009) );
  AOI21_X1 U21239 ( .B1(n18143), .B2(n18348), .A(n18009), .ZN(n18000) );
  OAI21_X1 U21240 ( .B1(n17943), .B2(n18269), .A(n18000), .ZN(n17940) );
  OAI222_X1 U21241 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17976), 
        .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18269), .C1(n18270), 
        .C2(n17940), .ZN(n17930) );
  OAI211_X1 U21242 ( .C1(n17979), .C2(n18278), .A(n17931), .B(n17930), .ZN(
        P3_U2808) );
  NAND2_X1 U21243 ( .A1(n18287), .A2(n18280), .ZN(n18293) );
  NOR2_X1 U21244 ( .A1(n17975), .A2(n18320), .ZN(n18281) );
  NAND2_X1 U21245 ( .A1(n17976), .A2(n18281), .ZN(n17960) );
  NAND2_X1 U21246 ( .A1(n18523), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18291) );
  OAI221_X1 U21247 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17934), .C1(
        n17933), .C2(n17932), .A(n18291), .ZN(n17935) );
  AOI21_X1 U21248 ( .B1(n18050), .B2(n17936), .A(n17935), .ZN(n17942) );
  NOR3_X1 U21249 ( .A1(n18107), .A2(n18320), .A3(n17937), .ZN(n17958) );
  AOI22_X1 U21250 ( .A1(n18287), .A2(n17958), .B1(n17969), .B2(n17938), .ZN(
        n17939) );
  XOR2_X1 U21251 ( .A(n18280), .B(n17939), .Z(n18290) );
  AOI22_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17940), .B1(
        n18110), .B2(n18290), .ZN(n17941) );
  OAI211_X1 U21253 ( .C1(n18293), .C2(n17960), .A(n17942), .B(n17941), .ZN(
        P3_U2809) );
  NAND2_X1 U21254 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18281), .ZN(
        n18264) );
  INV_X1 U21255 ( .A(n18264), .ZN(n18295) );
  OAI21_X1 U21256 ( .B1(n17943), .B2(n18295), .A(n18000), .ZN(n17962) );
  OAI221_X1 U21257 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17967), 
        .C1(n18307), .C2(n17958), .A(n17944), .ZN(n17945) );
  XOR2_X1 U21258 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17945), .Z(
        n18299) );
  NAND2_X1 U21259 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17946), .ZN(
        n18304) );
  OAI22_X1 U21260 ( .A1(n17979), .A2(n18299), .B1(n17960), .B2(n18304), .ZN(
        n17947) );
  AOI21_X1 U21261 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n17962), .A(
        n17947), .ZN(n17954) );
  NAND2_X1 U21262 ( .A1(n18523), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18302) );
  OAI221_X1 U21263 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17949), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18585), .A(n17948), .ZN(
        n17953) );
  OAI21_X1 U21264 ( .B1(n18050), .B2(n17980), .A(n17951), .ZN(n17952) );
  NAND4_X1 U21265 ( .A1(n17954), .A2(n18302), .A3(n17953), .A4(n17952), .ZN(
        P3_U2810) );
  AOI21_X1 U21266 ( .B1(n18031), .B2(n17955), .A(n18183), .ZN(n17981) );
  OAI21_X1 U21267 ( .B1(n17956), .B2(n19080), .A(n17981), .ZN(n17972) );
  AOI22_X1 U21268 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17972), .B1(
        n18050), .B2(n17957), .ZN(n17966) );
  AOI21_X1 U21269 ( .B1(n17969), .B2(n17967), .A(n17958), .ZN(n17959) );
  XOR2_X1 U21270 ( .A(n17959), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18311) );
  OAI22_X1 U21271 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17960), .B1(
        n18311), .B2(n17979), .ZN(n17961) );
  AOI21_X1 U21272 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17962), .A(
        n17961), .ZN(n17965) );
  NAND2_X1 U21273 ( .A1(n18523), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18310) );
  NOR2_X1 U21274 ( .A1(n18028), .A2(n17955), .ZN(n17974) );
  OAI211_X1 U21275 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17974), .B(n17963), .ZN(n17964) );
  NAND4_X1 U21276 ( .A1(n17966), .A2(n17965), .A3(n18310), .A4(n17964), .ZN(
        P3_U2811) );
  AOI21_X1 U21277 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18109), .A(
        n17967), .ZN(n17968) );
  XNOR2_X1 U21278 ( .A(n17969), .B(n17968), .ZN(n18326) );
  OAI22_X1 U21279 ( .A1(n18529), .A2(n19132), .B1(n18035), .B2(n9966), .ZN(
        n17971) );
  AOI221_X1 U21280 ( .B1(n17974), .B2(n17973), .C1(n17972), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17971), .ZN(n17978) );
  OAI21_X1 U21281 ( .B1(n18317), .B2(n18001), .A(n18000), .ZN(n17987) );
  NOR2_X1 U21282 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17975), .ZN(
        n18322) );
  AOI22_X1 U21283 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17987), .B1(
        n17976), .B2(n18322), .ZN(n17977) );
  OAI211_X1 U21284 ( .C1(n17979), .C2(n18326), .A(n17978), .B(n17977), .ZN(
        P3_U2812) );
  NAND2_X1 U21285 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18327), .ZN(
        n18333) );
  AOI21_X1 U21286 ( .B1(n10281), .B2(n18585), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17982) );
  OAI22_X1 U21287 ( .A1(n17982), .A2(n17981), .B1(n18418), .B2(n19130), .ZN(
        n17983) );
  AOI21_X1 U21288 ( .B1(n17984), .B2(n18169), .A(n17983), .ZN(n17989) );
  OAI21_X1 U21289 ( .B1(n17986), .B2(n18327), .A(n17985), .ZN(n18331) );
  AOI22_X1 U21290 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17987), .B1(
        n18110), .B2(n18331), .ZN(n17988) );
  OAI211_X1 U21291 ( .C1(n18001), .C2(n18333), .A(n17989), .B(n17988), .ZN(
        P3_U2813) );
  NOR2_X1 U21292 ( .A1(n18107), .A2(n18039), .ZN(n18051) );
  INV_X1 U21293 ( .A(n18051), .ZN(n18093) );
  OAI22_X1 U21294 ( .A1(n18109), .A2(n17990), .B1(n18093), .B2(n18314), .ZN(
        n17991) );
  XOR2_X1 U21295 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17991), .Z(
        n18343) );
  INV_X1 U21296 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19128) );
  AOI21_X1 U21297 ( .B1(n18031), .B2(n17994), .A(n18183), .ZN(n18026) );
  OAI21_X1 U21298 ( .B1(n17992), .B2(n19080), .A(n18026), .ZN(n18004) );
  AOI22_X1 U21299 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18004), .B1(
        n18050), .B2(n17993), .ZN(n17997) );
  NOR2_X1 U21300 ( .A1(n18028), .A2(n17994), .ZN(n18006) );
  OAI211_X1 U21301 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18006), .B(n17995), .ZN(n17996) );
  OAI211_X1 U21302 ( .C1(n19128), .C2(n18418), .A(n17997), .B(n17996), .ZN(
        n17998) );
  AOI21_X1 U21303 ( .B1(n18110), .B2(n18343), .A(n17998), .ZN(n17999) );
  OAI221_X1 U21304 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18001), 
        .C1(n18341), .C2(n18000), .A(n17999), .ZN(P3_U2814) );
  INV_X1 U21305 ( .A(n18360), .ZN(n18362) );
  NAND4_X1 U21306 ( .A1(n18362), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n18396), .ZN(n18022) );
  NAND2_X1 U21307 ( .A1(n11731), .A2(n18022), .ZN(n18350) );
  INV_X1 U21308 ( .A(n18350), .ZN(n18013) );
  NAND2_X1 U21309 ( .A1(n18143), .A2(n18348), .ZN(n18012) );
  INV_X1 U21310 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18005) );
  NAND2_X1 U21311 ( .A1(n18523), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18356) );
  OAI21_X1 U21312 ( .B1(n18035), .B2(n18002), .A(n18356), .ZN(n18003) );
  AOI221_X1 U21313 ( .B1(n18006), .B2(n18005), .C1(n18004), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18003), .ZN(n18011) );
  NAND2_X1 U21314 ( .A1(n18362), .A2(n18051), .ZN(n18018) );
  NAND2_X1 U21315 ( .A1(n18359), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18044) );
  INV_X1 U21316 ( .A(n18044), .ZN(n18384) );
  AOI221_X1 U21317 ( .B1(n18363), .B2(n18007), .C1(n18018), .C2(n18007), .A(
        n18384), .ZN(n18008) );
  XOR2_X1 U21318 ( .A(n18008), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n18355) );
  NAND2_X1 U21319 ( .A1(n11731), .A2(n18020), .ZN(n18352) );
  AOI22_X1 U21320 ( .A1(n18110), .A2(n18355), .B1(n18009), .B2(n18352), .ZN(
        n18010) );
  OAI211_X1 U21321 ( .C1(n18013), .C2(n18012), .A(n18011), .B(n18010), .ZN(
        P3_U2815) );
  NOR3_X1 U21322 ( .A1(n18557), .A2(n18064), .A3(n18014), .ZN(n18069) );
  AOI21_X1 U21323 ( .B1(n18030), .B2(n18069), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18027) );
  AOI22_X1 U21324 ( .A1(n18523), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18015), 
        .B2(n18169), .ZN(n18025) );
  INV_X1 U21325 ( .A(n18016), .ZN(n18017) );
  AOI21_X1 U21326 ( .B1(n18018), .B2(n18017), .A(n18384), .ZN(n18019) );
  XOR2_X1 U21327 ( .A(n18019), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18375) );
  OAI221_X1 U21328 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18399), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18368), .A(n18020), .ZN(
        n18372) );
  NOR2_X1 U21329 ( .A1(n18021), .A2(n18360), .ZN(n18379) );
  OAI221_X1 U21330 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18379), .A(n18022), .ZN(
        n18371) );
  OAI22_X1 U21331 ( .A1(n18072), .A2(n18372), .B1(n18202), .B2(n18371), .ZN(
        n18023) );
  AOI21_X1 U21332 ( .B1(n18110), .B2(n18375), .A(n18023), .ZN(n18024) );
  OAI211_X1 U21333 ( .C1(n18027), .C2(n18026), .A(n18025), .B(n18024), .ZN(
        P3_U2816) );
  NAND2_X1 U21334 ( .A1(n18408), .A2(n18058), .ZN(n18057) );
  INV_X1 U21335 ( .A(n18028), .ZN(n18029) );
  NAND2_X1 U21336 ( .A1(n17112), .A2(n18029), .ZN(n18047) );
  AOI211_X1 U21337 ( .C1(n18046), .C2(n18036), .A(n18030), .B(n18047), .ZN(
        n18038) );
  INV_X1 U21338 ( .A(n18031), .ZN(n18160) );
  OAI22_X1 U21339 ( .A1(n17112), .A2(n18160), .B1(n18032), .B2(n19080), .ZN(
        n18033) );
  NOR2_X1 U21340 ( .A1(n18183), .A2(n18033), .ZN(n18045) );
  OAI22_X1 U21341 ( .A1(n18045), .A2(n18036), .B1(n18035), .B2(n18034), .ZN(
        n18037) );
  AOI211_X1 U21342 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18523), .A(n18038), 
        .B(n18037), .ZN(n18043) );
  NOR2_X1 U21343 ( .A1(n18039), .A2(n18360), .ZN(n18378) );
  OAI22_X1 U21344 ( .A1(n18379), .A2(n18202), .B1(n18378), .B2(n18072), .ZN(
        n18054) );
  AOI22_X1 U21345 ( .A1(n18399), .A2(n18362), .B1(n18107), .B2(n11732), .ZN(
        n18040) );
  AOI21_X1 U21346 ( .B1(n18107), .B2(n18052), .A(n18040), .ZN(n18041) );
  XNOR2_X1 U21347 ( .A(n18359), .B(n18041), .ZN(n18385) );
  AOI22_X1 U21348 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18054), .B1(
        n18110), .B2(n18385), .ZN(n18042) );
  OAI211_X1 U21349 ( .C1(n18044), .C2(n18057), .A(n18043), .B(n18042), .ZN(
        P3_U2817) );
  NAND2_X1 U21350 ( .A1(n18523), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18393) );
  OAI221_X1 U21351 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18047), .C1(
        n18046), .C2(n18045), .A(n18393), .ZN(n18048) );
  AOI21_X1 U21352 ( .B1(n18050), .B2(n18049), .A(n18048), .ZN(n18056) );
  NAND2_X1 U21353 ( .A1(n18406), .A2(n18051), .ZN(n18059) );
  OAI21_X1 U21354 ( .B1(n18063), .B2(n18059), .A(n18052), .ZN(n18053) );
  XOR2_X1 U21355 ( .A(n18053), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18392) );
  AOI22_X1 U21356 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18054), .B1(
        n18110), .B2(n18392), .ZN(n18055) );
  OAI211_X1 U21357 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18057), .A(
        n18056), .B(n18055), .ZN(P3_U2818) );
  INV_X1 U21358 ( .A(n18058), .ZN(n18098) );
  NAND2_X1 U21359 ( .A1(n18406), .A2(n18063), .ZN(n18412) );
  INV_X1 U21360 ( .A(n18059), .ZN(n18060) );
  NOR2_X1 U21361 ( .A1(n18061), .A2(n18060), .ZN(n18062) );
  XOR2_X1 U21362 ( .A(n18063), .B(n18062), .Z(n18395) );
  NOR2_X1 U21363 ( .A1(n18529), .A2(n19118), .ZN(n18071) );
  INV_X1 U21364 ( .A(n18193), .ZN(n18077) );
  NOR2_X1 U21365 ( .A1(n18557), .A2(n18064), .ZN(n18119) );
  NAND2_X1 U21366 ( .A1(n18065), .A2(n18119), .ZN(n18088) );
  NOR2_X1 U21367 ( .A1(n18066), .A2(n18088), .ZN(n18079) );
  AOI21_X1 U21368 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18077), .A(
        n18079), .ZN(n18068) );
  OAI22_X1 U21369 ( .A1(n18069), .A2(n18068), .B1(n18194), .B2(n18067), .ZN(
        n18070) );
  AOI211_X1 U21370 ( .C1(n18110), .C2(n18395), .A(n18071), .B(n18070), .ZN(
        n18074) );
  NOR2_X1 U21371 ( .A1(n18406), .A2(n18098), .ZN(n18076) );
  OAI22_X1 U21372 ( .A1(n18399), .A2(n18072), .B1(n18202), .B2(n18396), .ZN(
        n18095) );
  OAI21_X1 U21373 ( .B1(n18076), .B2(n18095), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18073) );
  OAI211_X1 U21374 ( .C1(n18098), .C2(n18412), .A(n18074), .B(n18073), .ZN(
        P3_U2819) );
  INV_X1 U21375 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18428) );
  AOI22_X1 U21376 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18093), .B1(
        n18092), .B2(n18428), .ZN(n18075) );
  XOR2_X1 U21377 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18075), .Z(
        n18416) );
  NOR2_X1 U21378 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18081) );
  AOI21_X1 U21379 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18095), .A(
        n18076), .ZN(n18080) );
  NOR2_X1 U21380 ( .A1(n18087), .A2(n18088), .ZN(n18086) );
  AOI21_X1 U21381 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18077), .A(
        n18086), .ZN(n18078) );
  OAI22_X1 U21382 ( .A1(n18081), .A2(n18080), .B1(n18079), .B2(n18078), .ZN(
        n18082) );
  AOI21_X1 U21383 ( .B1(n18110), .B2(n18416), .A(n18082), .ZN(n18084) );
  NAND2_X1 U21384 ( .A1(n18523), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18083) );
  OAI211_X1 U21385 ( .C1(n18194), .C2(n18085), .A(n18084), .B(n18083), .ZN(
        P3_U2820) );
  AOI211_X1 U21386 ( .C1(n18088), .C2(n18087), .A(n18193), .B(n18086), .ZN(
        n18090) );
  NOR2_X1 U21387 ( .A1(n18529), .A2(n19114), .ZN(n18089) );
  AOI211_X1 U21388 ( .C1(n18091), .C2(n18169), .A(n18090), .B(n18089), .ZN(
        n18097) );
  NAND2_X1 U21389 ( .A1(n18093), .A2(n18092), .ZN(n18094) );
  XOR2_X1 U21390 ( .A(n18094), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18425) );
  AOI22_X1 U21391 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18095), .B1(
        n18110), .B2(n18425), .ZN(n18096) );
  OAI211_X1 U21392 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18098), .A(
        n18097), .B(n18096), .ZN(P3_U2821) );
  OAI21_X1 U21393 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18100), .A(
        n18099), .ZN(n18446) );
  OAI21_X1 U21394 ( .B1(n18102), .B2(n18160), .A(n9733), .ZN(n18120) );
  NOR2_X1 U21395 ( .A1(n18529), .A2(n19113), .ZN(n18437) );
  OAI211_X1 U21396 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18102), .B(n18101), .ZN(n18103)
         );
  OAI22_X1 U21397 ( .A1(n18194), .A2(n18104), .B1(n18557), .B2(n18103), .ZN(
        n18105) );
  AOI211_X1 U21398 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18120), .A(
        n18437), .B(n18105), .ZN(n18113) );
  INV_X1 U21399 ( .A(n18443), .ZN(n18108) );
  AOI22_X1 U21400 ( .A1(n18109), .A2(n18108), .B1(n18443), .B2(n18107), .ZN(
        n18440) );
  AOI22_X1 U21401 ( .A1(n18443), .A2(n18111), .B1(n18110), .B2(n18440), .ZN(
        n18112) );
  OAI211_X1 U21402 ( .C1(n18202), .C2(n18446), .A(n18113), .B(n18112), .ZN(
        P3_U2822) );
  OAI21_X1 U21403 ( .B1(n18116), .B2(n18115), .A(n18114), .ZN(n18117) );
  XOR2_X1 U21404 ( .A(n18117), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18456) );
  NOR2_X1 U21405 ( .A1(n18529), .A2(n19110), .ZN(n18450) );
  AOI221_X1 U21406 ( .B1(n18120), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18119), .C2(n18118), .A(n18450), .ZN(n18126) );
  AOI21_X1 U21407 ( .B1(n18123), .B2(n18122), .A(n18121), .ZN(n18453) );
  AOI22_X1 U21408 ( .A1(n18191), .A2(n18453), .B1(n18124), .B2(n18169), .ZN(
        n18125) );
  OAI211_X1 U21409 ( .C1(n18202), .C2(n18456), .A(n18126), .B(n18125), .ZN(
        P3_U2823) );
  NAND2_X1 U21410 ( .A1(n18585), .A2(n18129), .ZN(n18136) );
  AOI21_X1 U21411 ( .B1(n18128), .B2(n18127), .A(n9839), .ZN(n18463) );
  AOI22_X1 U21412 ( .A1(n18523), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18191), 
        .B2(n18463), .ZN(n18135) );
  AOI21_X1 U21413 ( .B1(n18129), .B2(n18585), .A(n18193), .ZN(n18148) );
  OAI21_X1 U21414 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18131), .A(
        n18130), .ZN(n18465) );
  OAI22_X1 U21415 ( .A1(n18194), .A2(n18132), .B1(n18202), .B2(n18465), .ZN(
        n18133) );
  AOI21_X1 U21416 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18148), .A(
        n18133), .ZN(n18134) );
  OAI211_X1 U21417 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18136), .A(
        n18135), .B(n18134), .ZN(P3_U2824) );
  OAI21_X1 U21418 ( .B1(n18139), .B2(n18138), .A(n18137), .ZN(n18140) );
  XOR2_X1 U21419 ( .A(n18140), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18474) );
  XOR2_X1 U21420 ( .A(n18142), .B(n18141), .Z(n18472) );
  AOI22_X1 U21421 ( .A1(n18523), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18143), 
        .B2(n18472), .ZN(n18150) );
  OAI21_X1 U21422 ( .B1(n18183), .B2(n18145), .A(n18144), .ZN(n18147) );
  AOI22_X1 U21423 ( .A1(n18148), .A2(n18147), .B1(n18146), .B2(n18169), .ZN(
        n18149) );
  OAI211_X1 U21424 ( .C1(n18201), .C2(n18474), .A(n18150), .B(n18149), .ZN(
        P3_U2825) );
  OAI21_X1 U21425 ( .B1(n18153), .B2(n18152), .A(n18151), .ZN(n18154) );
  XOR2_X1 U21426 ( .A(n18154), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18486) );
  OAI22_X1 U21427 ( .A1(n18202), .A2(n18486), .B1(n18557), .B2(n18155), .ZN(
        n18156) );
  AOI21_X1 U21428 ( .B1(n18523), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18156), .ZN(
        n18162) );
  AOI21_X1 U21429 ( .B1(n18159), .B2(n18158), .A(n18157), .ZN(n18475) );
  OAI21_X1 U21430 ( .B1(n17185), .B2(n18160), .A(n9733), .ZN(n18172) );
  AOI22_X1 U21431 ( .A1(n18191), .A2(n18475), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18172), .ZN(n18161) );
  OAI211_X1 U21432 ( .C1(n18194), .C2(n18163), .A(n18162), .B(n18161), .ZN(
        P3_U2826) );
  OAI21_X1 U21433 ( .B1(n18166), .B2(n18165), .A(n18164), .ZN(n18494) );
  AOI21_X1 U21434 ( .B1(n18489), .B2(n18168), .A(n18167), .ZN(n18492) );
  AOI22_X1 U21435 ( .A1(n18523), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18191), 
        .B2(n18492), .ZN(n18174) );
  OAI21_X1 U21436 ( .B1(n18183), .B2(n18184), .A(n17222), .ZN(n18171) );
  AOI22_X1 U21437 ( .A1(n18172), .A2(n18171), .B1(n18170), .B2(n18169), .ZN(
        n18173) );
  OAI211_X1 U21438 ( .C1(n18202), .C2(n18494), .A(n18174), .B(n18173), .ZN(
        P3_U2827) );
  OAI21_X1 U21439 ( .B1(n18177), .B2(n18176), .A(n18175), .ZN(n18504) );
  XNOR2_X1 U21440 ( .A(n18180), .B(n18179), .ZN(n18502) );
  OAI22_X1 U21441 ( .A1(n18194), .A2(n18181), .B1(n18201), .B2(n18502), .ZN(
        n18182) );
  AOI221_X1 U21442 ( .B1(n18585), .B2(n18184), .C1(n18183), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18182), .ZN(n18185) );
  NAND2_X1 U21443 ( .A1(n18523), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18508) );
  OAI211_X1 U21444 ( .C1(n18202), .C2(n18504), .A(n18185), .B(n18508), .ZN(
        P3_U2828) );
  AOI21_X1 U21445 ( .B1(n18195), .B2(n18188), .A(n18186), .ZN(n18516) );
  NAND2_X1 U21446 ( .A1(n19195), .A2(n18187), .ZN(n18189) );
  XNOR2_X1 U21447 ( .A(n18189), .B(n18188), .ZN(n18522) );
  OAI22_X1 U21448 ( .A1(n18522), .A2(n18202), .B1(n18418), .B2(n19099), .ZN(
        n18190) );
  AOI21_X1 U21449 ( .B1(n18191), .B2(n18516), .A(n18190), .ZN(n18192) );
  OAI221_X1 U21450 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18194), .C1(
        n9961), .C2(n18193), .A(n18192), .ZN(P3_U2829) );
  OAI21_X1 U21451 ( .B1(n18196), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18195), .ZN(n18525) );
  INV_X1 U21452 ( .A(n18525), .ZN(n18527) );
  OAI21_X1 U21453 ( .B1(n18198), .B2(n19221), .A(n9733), .ZN(n18199) );
  AOI22_X1 U21454 ( .A1(n18523), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18199), .ZN(n18200) );
  OAI221_X1 U21455 ( .B1(n18527), .B2(n18202), .C1(n18525), .C2(n18201), .A(
        n18200), .ZN(P3_U2830) );
  NOR3_X1 U21456 ( .A1(n18270), .A2(n18262), .A3(n18261), .ZN(n18255) );
  NAND2_X1 U21457 ( .A1(n18203), .A2(n18255), .ZN(n18220) );
  NOR2_X1 U21458 ( .A1(n18204), .A2(n18220), .ZN(n18215) );
  OAI22_X1 U21459 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19038), .B1(
        n18205), .B2(n19024), .ZN(n18206) );
  AOI211_X1 U21460 ( .C1(n18267), .C2(n18208), .A(n18207), .B(n18206), .ZN(
        n18210) );
  NOR2_X1 U21461 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19024), .ZN(
        n18476) );
  OAI21_X1 U21462 ( .B1(n18476), .B2(n18209), .A(n18477), .ZN(n18228) );
  OAI211_X1 U21463 ( .C1(n18211), .C2(n18397), .A(n18210), .B(n18228), .ZN(
        n18221) );
  AOI21_X1 U21464 ( .B1(n18212), .B2(n19020), .A(n18221), .ZN(n18213) );
  INV_X1 U21465 ( .A(n18213), .ZN(n18214) );
  MUX2_X1 U21466 ( .A(n18215), .B(n18214), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18217) );
  AOI22_X1 U21467 ( .A1(n18512), .A2(n18217), .B1(n18441), .B2(n18216), .ZN(
        n18219) );
  OAI211_X1 U21468 ( .C1(n18513), .C2(n21186), .A(n18219), .B(n18218), .ZN(
        P3_U2835) );
  NOR2_X1 U21469 ( .A1(n21104), .A2(n18220), .ZN(n18222) );
  MUX2_X1 U21470 ( .A(n18222), .B(n18221), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n18223) );
  AOI22_X1 U21471 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18458), .B1(
        n18512), .B2(n18223), .ZN(n18225) );
  OAI211_X1 U21472 ( .C1(n18226), .C2(n18325), .A(n18225), .B(n18224), .ZN(
        P3_U2836) );
  INV_X1 U21473 ( .A(n18227), .ZN(n18229) );
  OAI21_X1 U21474 ( .B1(n18229), .B2(n19031), .A(n18228), .ZN(n18230) );
  OAI221_X1 U21475 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18231), 
        .C1(n21104), .C2(n18230), .A(n18512), .ZN(n18232) );
  OAI211_X1 U21476 ( .C1(n18513), .C2(n21104), .A(n18233), .B(n18232), .ZN(
        n18237) );
  OAI22_X1 U21477 ( .A1(n18325), .A2(n18235), .B1(n18521), .B2(n18234), .ZN(
        n18236) );
  AOI211_X1 U21478 ( .C1(n18442), .C2(n18238), .A(n18237), .B(n18236), .ZN(
        n18239) );
  INV_X1 U21479 ( .A(n18239), .ZN(P3_U2837) );
  AOI21_X1 U21480 ( .B1(n18263), .B2(n18251), .A(n18398), .ZN(n18244) );
  AND2_X1 U21481 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18240), .ZN(
        n18241) );
  OAI22_X1 U21482 ( .A1(n18242), .A2(n18431), .B1(n18241), .B2(n18397), .ZN(
        n18243) );
  OAI211_X1 U21483 ( .C1(n18245), .C2(n19031), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18247), .ZN(n18246) );
  NAND2_X1 U21484 ( .A1(n18418), .A2(n18246), .ZN(n18258) );
  AOI21_X1 U21485 ( .B1(n18335), .B2(n18247), .A(n18258), .ZN(n18249) );
  AOI21_X1 U21486 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18249), .A(
        n18248), .ZN(n18253) );
  NAND3_X1 U21487 ( .A1(n18251), .A2(n18279), .A3(n18250), .ZN(n18252) );
  OAI211_X1 U21488 ( .C1(n18254), .C2(n18325), .A(n18253), .B(n18252), .ZN(
        P3_U2838) );
  AOI21_X1 U21489 ( .B1(n18255), .B2(n18513), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U21490 ( .A1(n18523), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18441), 
        .B2(n18256), .ZN(n18257) );
  OAI21_X1 U21491 ( .B1(n18259), .B2(n18258), .A(n18257), .ZN(P3_U2839) );
  AOI21_X1 U21492 ( .B1(n18458), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n18260), .ZN(n18277) );
  NOR2_X1 U21493 ( .A1(n18262), .A2(n18261), .ZN(n18275) );
  NOR2_X1 U21494 ( .A1(n18263), .A2(n18398), .ZN(n18351) );
  AOI21_X1 U21495 ( .B1(n18999), .B2(n18348), .A(n18351), .ZN(n18283) );
  OAI21_X1 U21496 ( .B1(n18315), .B2(n18264), .A(n19020), .ZN(n18265) );
  OAI221_X1 U21497 ( .B1(n19031), .B2(n18266), .C1(n19031), .C2(n18281), .A(
        n18265), .ZN(n18297) );
  NOR2_X1 U21498 ( .A1(n18267), .A2(n18999), .ZN(n18405) );
  OAI22_X1 U21499 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19038), .B1(
        n18269), .B2(n18405), .ZN(n18268) );
  NOR2_X1 U21500 ( .A1(n18297), .A2(n18268), .ZN(n18285) );
  AOI21_X1 U21501 ( .B1(n18282), .B2(n18269), .A(n19024), .ZN(n18271) );
  AOI211_X1 U21502 ( .C1(n18272), .C2(n18413), .A(n18271), .B(n18270), .ZN(
        n18273) );
  NAND3_X1 U21503 ( .A1(n18283), .A2(n18285), .A3(n18273), .ZN(n18274) );
  OAI211_X1 U21504 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18275), .A(
        n18512), .B(n18274), .ZN(n18276) );
  OAI211_X1 U21505 ( .C1(n18278), .C2(n18325), .A(n18277), .B(n18276), .ZN(
        P3_U2840) );
  NAND2_X1 U21506 ( .A1(n18279), .A2(n18281), .ZN(n18305) );
  NOR2_X1 U21507 ( .A1(n18523), .A2(n18280), .ZN(n18289) );
  NAND2_X1 U21508 ( .A1(n19031), .A2(n19024), .ZN(n18511) );
  INV_X1 U21509 ( .A(n18511), .ZN(n18286) );
  AOI21_X1 U21510 ( .B1(n18282), .B2(n18281), .A(n19024), .ZN(n18284) );
  NAND2_X1 U21511 ( .A1(n18512), .A2(n18283), .ZN(n18340) );
  NOR2_X1 U21512 ( .A1(n18284), .A2(n18340), .ZN(n18294) );
  OAI211_X1 U21513 ( .C1(n18287), .C2(n18286), .A(n18285), .B(n18294), .ZN(
        n18288) );
  AOI22_X1 U21514 ( .A1(n18441), .A2(n18290), .B1(n18289), .B2(n18288), .ZN(
        n18292) );
  OAI211_X1 U21515 ( .C1(n18293), .C2(n18305), .A(n18292), .B(n18291), .ZN(
        P3_U2841) );
  OAI21_X1 U21516 ( .B1(n18295), .B2(n18405), .A(n18294), .ZN(n18296) );
  OAI21_X1 U21517 ( .B1(n18297), .B2(n18296), .A(n18529), .ZN(n18306) );
  NAND3_X1 U21518 ( .A1(n18511), .A2(n18307), .A3(P3_STATE2_REG_2__SCAN_IN), 
        .ZN(n18298) );
  NAND2_X1 U21519 ( .A1(n18306), .A2(n18298), .ZN(n18301) );
  INV_X1 U21520 ( .A(n18299), .ZN(n18300) );
  AOI22_X1 U21521 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18301), .B1(
        n18441), .B2(n18300), .ZN(n18303) );
  OAI211_X1 U21522 ( .C1(n18304), .C2(n18305), .A(n18303), .B(n18302), .ZN(
        P3_U2842) );
  OAI22_X1 U21523 ( .A1(n18307), .A2(n18306), .B1(n18305), .B2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18308) );
  INV_X1 U21524 ( .A(n18308), .ZN(n18309) );
  OAI211_X1 U21525 ( .C1(n18311), .C2(n18325), .A(n18310), .B(n18309), .ZN(
        P3_U2843) );
  OAI22_X1 U21526 ( .A1(n18495), .A2(n19031), .B1(n18478), .B2(n18496), .ZN(
        n18430) );
  INV_X1 U21527 ( .A(n18430), .ZN(n18488) );
  NOR3_X1 U21528 ( .A1(n18438), .A2(n18436), .A3(n18447), .ZN(n18367) );
  OAI21_X1 U21529 ( .B1(n18367), .B2(n18313), .A(n18512), .ZN(n18429) );
  NOR2_X1 U21530 ( .A1(n18314), .A2(n18429), .ZN(n18342) );
  NOR3_X1 U21531 ( .A1(n18476), .A2(n18315), .A3(n18341), .ZN(n18316) );
  OAI22_X1 U21532 ( .A1(n18317), .A2(n18405), .B1(n18431), .B2(n18316), .ZN(
        n18318) );
  AOI211_X1 U21533 ( .C1(n19010), .C2(n18319), .A(n18340), .B(n18318), .ZN(
        n18328) );
  AOI221_X1 U21534 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18328), 
        .C1(n18431), .C2(n18328), .A(n18320), .ZN(n18321) );
  AOI22_X1 U21535 ( .A1(n18342), .A2(n18322), .B1(n18321), .B2(n18529), .ZN(
        n18324) );
  NAND2_X1 U21536 ( .A1(n18523), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18323) );
  OAI211_X1 U21537 ( .C1(n18326), .C2(n18325), .A(n18324), .B(n18323), .ZN(
        P3_U2844) );
  INV_X1 U21538 ( .A(n18342), .ZN(n18334) );
  NOR2_X1 U21539 ( .A1(n18529), .A2(n19130), .ZN(n18330) );
  NOR3_X1 U21540 ( .A1(n18523), .A2(n18328), .A3(n18327), .ZN(n18329) );
  AOI211_X1 U21541 ( .C1(n18441), .C2(n18331), .A(n18330), .B(n18329), .ZN(
        n18332) );
  OAI21_X1 U21542 ( .B1(n18334), .B2(n18333), .A(n18332), .ZN(P3_U2845) );
  INV_X1 U21543 ( .A(n18335), .ZN(n18339) );
  AOI21_X1 U21544 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18336), .A(
        n19038), .ZN(n18402) );
  AOI21_X1 U21545 ( .B1(n19010), .B2(n18401), .A(n18402), .ZN(n18361) );
  OAI21_X1 U21546 ( .B1(n19036), .B2(n11731), .A(n18337), .ZN(n18338) );
  OAI211_X1 U21547 ( .C1(n18346), .C2(n18407), .A(n18361), .B(n18338), .ZN(
        n18353) );
  OAI221_X1 U21548 ( .B1(n18340), .B2(n18339), .C1(n18340), .C2(n18353), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U21549 ( .A1(n18441), .A2(n18343), .B1(n18342), .B2(n18341), .ZN(
        n18344) );
  OAI221_X1 U21550 ( .B1(n18523), .B2(n18345), .C1(n18418), .C2(n19128), .A(
        n18344), .ZN(P3_U2846) );
  AOI21_X1 U21551 ( .B1(n18346), .B2(n18367), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18347) );
  INV_X1 U21552 ( .A(n18347), .ZN(n18354) );
  AND2_X1 U21553 ( .A1(n18348), .A2(n18999), .ZN(n18349) );
  AOI222_X1 U21554 ( .A1(n18354), .A2(n18353), .B1(n18352), .B2(n18351), .C1(
        n18350), .C2(n18349), .ZN(n18358) );
  AOI22_X1 U21555 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18458), .B1(
        n18441), .B2(n18355), .ZN(n18357) );
  OAI211_X1 U21556 ( .C1(n18358), .C2(n18530), .A(n18357), .B(n18356), .ZN(
        P3_U2847) );
  INV_X1 U21557 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19124) );
  AOI22_X1 U21558 ( .A1(n19010), .A2(n18360), .B1(n18359), .B2(n18511), .ZN(
        n18366) );
  OAI221_X1 U21559 ( .B1(n19024), .B2(n18362), .C1(n19024), .C2(n18422), .A(
        n18361), .ZN(n18381) );
  AOI211_X1 U21560 ( .C1(n18364), .C2(n19020), .A(n18363), .B(n18381), .ZN(
        n18365) );
  AOI21_X1 U21561 ( .B1(n18366), .B2(n18365), .A(n18530), .ZN(n18370) );
  AND2_X1 U21562 ( .A1(n18368), .A2(n18367), .ZN(n18369) );
  AOI222_X1 U21563 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18370), 
        .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18458), .C1(n18370), 
        .C2(n18369), .ZN(n18377) );
  OAI22_X1 U21564 ( .A1(n18373), .A2(n18372), .B1(n18521), .B2(n18371), .ZN(
        n18374) );
  AOI21_X1 U21565 ( .B1(n18441), .B2(n18375), .A(n18374), .ZN(n18376) );
  OAI211_X1 U21566 ( .C1(n18418), .C2(n19124), .A(n18377), .B(n18376), .ZN(
        P3_U2848) );
  OAI22_X1 U21567 ( .A1(n18379), .A2(n18397), .B1(n18378), .B2(n18398), .ZN(
        n18380) );
  AOI211_X1 U21568 ( .C1(n18383), .C2(n18413), .A(n18381), .B(n18380), .ZN(
        n18390) );
  OAI211_X1 U21569 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18407), .A(
        n18512), .B(n18390), .ZN(n18382) );
  NAND2_X1 U21570 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18382), .ZN(
        n18387) );
  NOR2_X1 U21571 ( .A1(n18383), .A2(n18429), .ZN(n18388) );
  AOI22_X1 U21572 ( .A1(n18441), .A2(n18385), .B1(n18384), .B2(n18388), .ZN(
        n18386) );
  OAI221_X1 U21573 ( .B1(n18523), .B2(n18387), .C1(n18418), .C2(n19122), .A(
        n18386), .ZN(P3_U2849) );
  AOI21_X1 U21574 ( .B1(n18512), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18388), .ZN(n18389) );
  AOI21_X1 U21575 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18390), .A(
        n18389), .ZN(n18391) );
  AOI21_X1 U21576 ( .B1(n18441), .B2(n18392), .A(n18391), .ZN(n18394) );
  OAI211_X1 U21577 ( .C1(n18513), .C2(n11732), .A(n18394), .B(n18393), .ZN(
        P3_U2850) );
  AOI22_X1 U21578 ( .A1(n18523), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18441), 
        .B2(n18395), .ZN(n18411) );
  OAI22_X1 U21579 ( .A1(n18399), .A2(n18398), .B1(n18397), .B2(n18396), .ZN(
        n18400) );
  AOI211_X1 U21580 ( .C1(n19010), .C2(n18401), .A(n18530), .B(n18400), .ZN(
        n18420) );
  AOI221_X1 U21581 ( .B1(n18428), .B2(n19036), .C1(n18403), .C2(n19036), .A(
        n18402), .ZN(n18404) );
  OAI211_X1 U21582 ( .C1(n18406), .C2(n18405), .A(n18420), .B(n18404), .ZN(
        n18414) );
  OAI22_X1 U21583 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n19024), .B1(
        n18408), .B2(n18407), .ZN(n18409) );
  OAI211_X1 U21584 ( .C1(n18414), .C2(n18409), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18418), .ZN(n18410) );
  OAI211_X1 U21585 ( .C1(n18412), .C2(n18429), .A(n18411), .B(n18410), .ZN(
        P3_U2851) );
  OAI221_X1 U21586 ( .B1(n18414), .B2(n18428), .C1(n18414), .C2(n18413), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18419) );
  NOR3_X1 U21587 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18428), .A3(
        n18429), .ZN(n18415) );
  AOI21_X1 U21588 ( .B1(n18441), .B2(n18416), .A(n18415), .ZN(n18417) );
  OAI221_X1 U21589 ( .B1(n18523), .B2(n18419), .C1(n18418), .C2(n19116), .A(
        n18417), .ZN(P3_U2852) );
  NAND2_X1 U21590 ( .A1(n18438), .A2(n19020), .ZN(n18421) );
  OAI211_X1 U21591 ( .C1(n18422), .C2(n19024), .A(n18421), .B(n18420), .ZN(
        n18424) );
  OAI221_X1 U21592 ( .B1(n18424), .B2(n19020), .C1(n18424), .C2(n18423), .A(
        n18529), .ZN(n18427) );
  AOI22_X1 U21593 ( .A1(n18523), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18441), 
        .B2(n18425), .ZN(n18426) );
  OAI221_X1 U21594 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18429), .C1(
        n18428), .C2(n18427), .A(n18426), .ZN(P3_U2853) );
  NAND3_X1 U21595 ( .A1(n18430), .A2(n18512), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18466) );
  INV_X1 U21596 ( .A(n18466), .ZN(n18481) );
  NAND3_X1 U21597 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n18481), .ZN(n18461) );
  NOR2_X1 U21598 ( .A1(n18436), .A2(n18461), .ZN(n18439) );
  OAI22_X1 U21599 ( .A1(n18433), .A2(n19031), .B1(n18432), .B2(n18431), .ZN(
        n18434) );
  NOR2_X1 U21600 ( .A1(n18476), .A2(n18434), .ZN(n18435) );
  NOR2_X1 U21601 ( .A1(n18530), .A2(n18435), .ZN(n18457) );
  AOI21_X1 U21602 ( .B1(n18518), .B2(n18436), .A(n18457), .ZN(n18448) );
  NAND2_X1 U21603 ( .A1(n18448), .A2(n18513), .ZN(n18451) );
  AOI221_X1 U21604 ( .B1(n18439), .B2(n18438), .C1(n18451), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18437), .ZN(n18445) );
  AOI22_X1 U21605 ( .A1(n18443), .A2(n18442), .B1(n18441), .B2(n18440), .ZN(
        n18444) );
  OAI211_X1 U21606 ( .C1(n18521), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2854) );
  NOR3_X1 U21607 ( .A1(n18448), .A2(n18447), .A3(n18460), .ZN(n18449) );
  AOI211_X1 U21608 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18451), .A(
        n18450), .B(n18449), .ZN(n18455) );
  NAND2_X1 U21609 ( .A1(n18452), .A2(n18512), .ZN(n18503) );
  INV_X1 U21610 ( .A(n18503), .ZN(n18528) );
  NAND2_X1 U21611 ( .A1(n18453), .A2(n18528), .ZN(n18454) );
  OAI211_X1 U21612 ( .C1(n18456), .C2(n18521), .A(n18455), .B(n18454), .ZN(
        P3_U2855) );
  NOR2_X1 U21613 ( .A1(n18458), .A2(n18457), .ZN(n18467) );
  NAND2_X1 U21614 ( .A1(n18523), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18459) );
  OAI221_X1 U21615 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18461), .C1(
        n18460), .C2(n18467), .A(n18459), .ZN(n18462) );
  AOI21_X1 U21616 ( .B1(n18528), .B2(n18463), .A(n18462), .ZN(n18464) );
  OAI21_X1 U21617 ( .B1(n18521), .B2(n18465), .A(n18464), .ZN(P3_U2856) );
  NOR2_X1 U21618 ( .A1(n18529), .A2(n19106), .ZN(n18471) );
  NOR2_X1 U21619 ( .A1(n18480), .A2(n18466), .ZN(n18469) );
  INV_X1 U21620 ( .A(n18467), .ZN(n18468) );
  MUX2_X1 U21621 ( .A(n18469), .B(n18468), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18470) );
  AOI211_X1 U21622 ( .C1(n18526), .C2(n18472), .A(n18471), .B(n18470), .ZN(
        n18473) );
  OAI21_X1 U21623 ( .B1(n18503), .B2(n18474), .A(n18473), .ZN(P3_U2857) );
  AOI22_X1 U21624 ( .A1(n18523), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18528), 
        .B2(n18475), .ZN(n18485) );
  AOI21_X1 U21625 ( .B1(n18478), .B2(n18477), .A(n18476), .ZN(n18479) );
  INV_X1 U21626 ( .A(n18479), .ZN(n18497) );
  AOI211_X1 U21627 ( .C1(n18495), .C2(n19010), .A(n18489), .B(n18497), .ZN(
        n18487) );
  AOI21_X1 U21628 ( .B1(n18512), .B2(n18487), .A(n18480), .ZN(n18483) );
  AOI22_X1 U21629 ( .A1(n18483), .A2(n18482), .B1(n18481), .B2(n18480), .ZN(
        n18484) );
  OAI211_X1 U21630 ( .C1(n18521), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P3_U2858) );
  AOI211_X1 U21631 ( .C1(n18488), .C2(n18489), .A(n18487), .B(n18530), .ZN(
        n18491) );
  OAI22_X1 U21632 ( .A1(n18529), .A2(n19102), .B1(n18489), .B2(n18513), .ZN(
        n18490) );
  AOI211_X1 U21633 ( .C1(n18492), .C2(n18528), .A(n18491), .B(n18490), .ZN(
        n18493) );
  OAI21_X1 U21634 ( .B1(n18521), .B2(n18494), .A(n18493), .ZN(P3_U2859) );
  AND2_X1 U21635 ( .A1(n19010), .A2(n18495), .ZN(n18507) );
  NOR2_X1 U21636 ( .A1(n19181), .A2(n18496), .ZN(n18501) );
  NOR2_X1 U21637 ( .A1(n19181), .A2(n19195), .ZN(n18498) );
  AOI21_X1 U21638 ( .B1(n19010), .B2(n18498), .A(n18497), .ZN(n18499) );
  INV_X1 U21639 ( .A(n18499), .ZN(n18500) );
  MUX2_X1 U21640 ( .A(n18501), .B(n18500), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18506) );
  OAI22_X1 U21641 ( .A1(n18521), .A2(n18504), .B1(n18503), .B2(n18502), .ZN(
        n18505) );
  AOI221_X1 U21642 ( .B1(n18507), .B2(n18512), .C1(n18506), .C2(n18512), .A(
        n18505), .ZN(n18509) );
  OAI211_X1 U21643 ( .C1(n18513), .C2(n18510), .A(n18509), .B(n18508), .ZN(
        P3_U2860) );
  NOR2_X1 U21644 ( .A1(n18529), .A2(n19099), .ZN(n18515) );
  NAND3_X1 U21645 ( .A1(n18512), .A2(n19195), .A3(n18511), .ZN(n18532) );
  AOI21_X1 U21646 ( .B1(n18513), .B2(n18532), .A(n19181), .ZN(n18514) );
  AOI211_X1 U21647 ( .C1(n18516), .C2(n18528), .A(n18515), .B(n18514), .ZN(
        n18520) );
  NAND3_X1 U21648 ( .A1(n18518), .A2(n19181), .A3(n18517), .ZN(n18519) );
  OAI211_X1 U21649 ( .C1(n18522), .C2(n18521), .A(n18520), .B(n18519), .ZN(
        P3_U2861) );
  AND2_X1 U21650 ( .A1(n18523), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18524) );
  AOI221_X1 U21651 ( .B1(n18528), .B2(n18527), .C1(n18526), .C2(n18525), .A(
        n18524), .ZN(n18533) );
  OAI211_X1 U21652 ( .C1(n19020), .C2(n18530), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18529), .ZN(n18531) );
  NAND3_X1 U21653 ( .A1(n18533), .A2(n18532), .A3(n18531), .ZN(P3_U2862) );
  AOI211_X1 U21654 ( .C1(n18535), .C2(n18534), .A(n19179), .B(n19228), .ZN(
        n19063) );
  OAI21_X1 U21655 ( .B1(n19063), .B2(n18595), .A(n18540), .ZN(n18536) );
  OAI221_X1 U21656 ( .B1(n19042), .B2(n19212), .C1(n19042), .C2(n18540), .A(
        n18536), .ZN(P3_U2863) );
  INV_X1 U21657 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19052) );
  NAND2_X1 U21658 ( .A1(n19049), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18800) );
  INV_X1 U21659 ( .A(n18800), .ZN(n18846) );
  NAND2_X1 U21660 ( .A1(n19052), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18703) );
  INV_X1 U21661 ( .A(n18703), .ZN(n18729) );
  NOR2_X1 U21662 ( .A1(n18846), .A2(n18729), .ZN(n18537) );
  OAI22_X1 U21663 ( .A1(n18539), .A2(n19052), .B1(n18538), .B2(n18537), .ZN(
        P3_U2866) );
  NOR2_X1 U21664 ( .A1(n19053), .A2(n18540), .ZN(P3_U2867) );
  NOR2_X1 U21665 ( .A1(n19052), .A2(n18541), .ZN(n18943) );
  NAND2_X1 U21666 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18943), .ZN(
        n18996) );
  NOR2_X1 U21667 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18656) );
  NOR2_X1 U21668 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18635) );
  NAND2_X1 U21669 ( .A1(n18656), .A2(n18635), .ZN(n18650) );
  NOR2_X1 U21670 ( .A1(n18969), .A2(n18652), .ZN(n18615) );
  NOR2_X1 U21671 ( .A1(n18657), .A2(n18542), .ZN(n18911) );
  INV_X1 U21672 ( .A(n18911), .ZN(n18750) );
  NAND2_X1 U21673 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18544) );
  NAND2_X1 U21674 ( .A1(n19042), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18796) );
  INV_X1 U21675 ( .A(n18796), .ZN(n18614) );
  NOR2_X1 U21676 ( .A1(n19042), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18773) );
  NOR2_X1 U21677 ( .A1(n18614), .A2(n18773), .ZN(n18848) );
  NOR2_X1 U21678 ( .A1(n18544), .A2(n18848), .ZN(n18914) );
  INV_X1 U21679 ( .A(n18914), .ZN(n18909) );
  OAI22_X1 U21680 ( .A1(n18615), .A2(n18750), .B1(n18557), .B2(n18909), .ZN(
        n18592) );
  NOR2_X2 U21681 ( .A1(n18657), .A2(n21110), .ZN(n18941) );
  NOR2_X1 U21682 ( .A1(n19072), .A2(n18615), .ZN(n18587) );
  AND2_X1 U21683 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18585), .ZN(n18940) );
  NOR2_X1 U21684 ( .A1(n18544), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18944) );
  NAND2_X1 U21685 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18944), .ZN(
        n18973) );
  INV_X1 U21686 ( .A(n18973), .ZN(n18991) );
  AOI22_X1 U21687 ( .A1(n18941), .A2(n18587), .B1(n18940), .B2(n18991), .ZN(
        n18549) );
  INV_X1 U21688 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18543) );
  NOR2_X2 U21689 ( .A1(n18557), .A2(n18543), .ZN(n18945) );
  NOR2_X2 U21690 ( .A1(n18796), .A2(n18544), .ZN(n18917) );
  NAND2_X1 U21691 ( .A1(n18546), .A2(n18545), .ZN(n18588) );
  NOR2_X1 U21692 ( .A1(n18547), .A2(n18588), .ZN(n18878) );
  AOI22_X1 U21693 ( .A1(n18945), .A2(n18917), .B1(n18878), .B2(n18652), .ZN(
        n18548) );
  OAI211_X1 U21694 ( .C1(n18550), .C2(n18592), .A(n18549), .B(n18548), .ZN(
        P3_U2868) );
  INV_X1 U21695 ( .A(n18657), .ZN(n18849) );
  AND2_X1 U21696 ( .A1(n18849), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18950) );
  NOR2_X2 U21697 ( .A1(n18551), .A2(n18557), .ZN(n18949) );
  AOI22_X1 U21698 ( .A1(n18950), .A2(n18587), .B1(n18949), .B2(n18991), .ZN(
        n18554) );
  NAND2_X1 U21699 ( .A1(n18585), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18954) );
  INV_X1 U21700 ( .A(n18954), .ZN(n18881) );
  NOR2_X1 U21701 ( .A1(n18552), .A2(n18588), .ZN(n18951) );
  AOI22_X1 U21702 ( .A1(n18881), .A2(n18917), .B1(n18951), .B2(n18652), .ZN(
        n18553) );
  OAI211_X1 U21703 ( .C1(n21310), .C2(n18592), .A(n18554), .B(n18553), .ZN(
        P3_U2869) );
  NOR2_X2 U21704 ( .A1(n18657), .A2(n18555), .ZN(n18955) );
  AND2_X1 U21705 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18585), .ZN(n18957) );
  AOI22_X1 U21706 ( .A1(n18955), .A2(n18587), .B1(n18957), .B2(n18991), .ZN(
        n18560) );
  INV_X1 U21707 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18556) );
  NOR2_X1 U21708 ( .A1(n18557), .A2(n18556), .ZN(n18956) );
  NOR2_X1 U21709 ( .A1(n18558), .A2(n18588), .ZN(n18885) );
  AOI22_X1 U21710 ( .A1(n18956), .A2(n18917), .B1(n18885), .B2(n18652), .ZN(
        n18559) );
  OAI211_X1 U21711 ( .C1(n18561), .C2(n18592), .A(n18560), .B(n18559), .ZN(
        P3_U2870) );
  NOR2_X2 U21712 ( .A1(n18657), .A2(n18562), .ZN(n18961) );
  NOR2_X2 U21713 ( .A1(n21126), .A2(n18557), .ZN(n18963) );
  AOI22_X1 U21714 ( .A1(n18961), .A2(n18587), .B1(n18963), .B2(n18991), .ZN(
        n18565) );
  NAND2_X1 U21715 ( .A1(n18585), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18861) );
  INV_X1 U21716 ( .A(n18861), .ZN(n18962) );
  NOR2_X1 U21717 ( .A1(n18563), .A2(n18588), .ZN(n18889) );
  AOI22_X1 U21718 ( .A1(n18962), .A2(n18917), .B1(n18889), .B2(n18652), .ZN(
        n18564) );
  OAI211_X1 U21719 ( .C1(n21246), .C2(n18592), .A(n18565), .B(n18564), .ZN(
        P3_U2871) );
  INV_X1 U21720 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18566) );
  NOR2_X1 U21721 ( .A1(n18557), .A2(n18566), .ZN(n18925) );
  NOR2_X2 U21722 ( .A1(n18657), .A2(n18567), .ZN(n18967) );
  AOI22_X1 U21723 ( .A1(n18925), .A2(n18917), .B1(n18967), .B2(n18587), .ZN(
        n18570) );
  NOR2_X1 U21724 ( .A1(n18568), .A2(n18588), .ZN(n18970) );
  AND2_X1 U21725 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18585), .ZN(n18968) );
  AOI22_X1 U21726 ( .A1(n18970), .A2(n18652), .B1(n18968), .B2(n18991), .ZN(
        n18569) );
  OAI211_X1 U21727 ( .C1(n18571), .C2(n18592), .A(n18570), .B(n18569), .ZN(
        P3_U2872) );
  NOR2_X2 U21728 ( .A1(n18657), .A2(n18573), .ZN(n18975) );
  AOI22_X1 U21729 ( .A1(n18976), .A2(n18991), .B1(n18975), .B2(n18587), .ZN(
        n18576) );
  NOR2_X1 U21730 ( .A1(n18574), .A2(n18588), .ZN(n18864) );
  AND2_X1 U21731 ( .A1(n18585), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18977) );
  AOI22_X1 U21732 ( .A1(n18864), .A2(n18652), .B1(n18977), .B2(n18917), .ZN(
        n18575) );
  OAI211_X1 U21733 ( .C1(n18577), .C2(n18592), .A(n18576), .B(n18575), .ZN(
        P3_U2873) );
  NOR2_X2 U21734 ( .A1(n18657), .A2(n18579), .ZN(n18981) );
  AOI22_X1 U21735 ( .A1(n18982), .A2(n18991), .B1(n18981), .B2(n18587), .ZN(
        n18583) );
  NOR2_X1 U21736 ( .A1(n18580), .A2(n18588), .ZN(n18899) );
  NOR2_X2 U21737 ( .A1(n18557), .A2(n18581), .ZN(n18983) );
  AOI22_X1 U21738 ( .A1(n18899), .A2(n18652), .B1(n18983), .B2(n18917), .ZN(
        n18582) );
  OAI211_X1 U21739 ( .C1(n18584), .C2(n18592), .A(n18583), .B(n18582), .ZN(
        P3_U2874) );
  NAND2_X1 U21740 ( .A1(n18585), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18823) );
  INV_X1 U21741 ( .A(n18823), .ZN(n18990) );
  NOR2_X2 U21742 ( .A1(n18586), .A2(n18657), .ZN(n18988) );
  AOI22_X1 U21743 ( .A1(n18990), .A2(n18991), .B1(n18988), .B2(n18587), .ZN(
        n18591) );
  NOR2_X1 U21744 ( .A1(n18589), .A2(n18588), .ZN(n18819) );
  NOR2_X2 U21745 ( .A1(n19700), .A2(n18557), .ZN(n18992) );
  AOI22_X1 U21746 ( .A1(n18819), .A2(n18652), .B1(n18992), .B2(n18917), .ZN(
        n18590) );
  OAI211_X1 U21747 ( .C1(n18593), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U2875) );
  NAND2_X1 U21748 ( .A1(n18773), .A2(n18635), .ZN(n18680) );
  INV_X1 U21749 ( .A(n18635), .ZN(n18594) );
  AOI22_X1 U21750 ( .A1(n18941), .A2(n18610), .B1(n18940), .B2(n18917), .ZN(
        n18597) );
  NOR2_X1 U21751 ( .A1(n18657), .A2(n18595), .ZN(n18942) );
  AND2_X1 U21752 ( .A1(n19044), .A2(n18942), .ZN(n18682) );
  AOI22_X1 U21753 ( .A1(n18585), .A2(n18943), .B1(n18635), .B2(n18682), .ZN(
        n18611) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18611), .B1(
        n18945), .B2(n18969), .ZN(n18596) );
  OAI211_X1 U21755 ( .C1(n18948), .C2(n18680), .A(n18597), .B(n18596), .ZN(
        P3_U2876) );
  INV_X1 U21756 ( .A(n18951), .ZN(n18855) );
  AOI22_X1 U21757 ( .A1(n18881), .A2(n18969), .B1(n18950), .B2(n18610), .ZN(
        n18599) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18611), .B1(
        n18949), .B2(n18917), .ZN(n18598) );
  OAI211_X1 U21759 ( .C1(n18855), .C2(n18680), .A(n18599), .B(n18598), .ZN(
        P3_U2877) );
  INV_X1 U21760 ( .A(n18885), .ZN(n18960) );
  AOI22_X1 U21761 ( .A1(n18956), .A2(n18969), .B1(n18955), .B2(n18610), .ZN(
        n18601) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18611), .B1(
        n18957), .B2(n18917), .ZN(n18600) );
  OAI211_X1 U21763 ( .C1(n18960), .C2(n18680), .A(n18601), .B(n18600), .ZN(
        P3_U2878) );
  INV_X1 U21764 ( .A(n18889), .ZN(n18966) );
  AOI22_X1 U21765 ( .A1(n18962), .A2(n18969), .B1(n18961), .B2(n18610), .ZN(
        n18603) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18611), .B1(
        n18963), .B2(n18917), .ZN(n18602) );
  OAI211_X1 U21767 ( .C1(n18966), .C2(n18680), .A(n18603), .B(n18602), .ZN(
        P3_U2879) );
  INV_X1 U21768 ( .A(n18970), .ZN(n18928) );
  AOI22_X1 U21769 ( .A1(n18925), .A2(n18969), .B1(n18967), .B2(n18610), .ZN(
        n18605) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18611), .B1(
        n18968), .B2(n18917), .ZN(n18604) );
  OAI211_X1 U21771 ( .C1(n18928), .C2(n18680), .A(n18605), .B(n18604), .ZN(
        P3_U2880) );
  AOI22_X1 U21772 ( .A1(n18977), .A2(n18969), .B1(n18975), .B2(n18610), .ZN(
        n18607) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18611), .B1(
        n18976), .B2(n18917), .ZN(n18606) );
  OAI211_X1 U21774 ( .C1(n18980), .C2(n18680), .A(n18607), .B(n18606), .ZN(
        P3_U2881) );
  INV_X1 U21775 ( .A(n18899), .ZN(n18986) );
  AOI22_X1 U21776 ( .A1(n18982), .A2(n18917), .B1(n18981), .B2(n18610), .ZN(
        n18609) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18611), .B1(
        n18983), .B2(n18969), .ZN(n18608) );
  OAI211_X1 U21778 ( .C1(n18986), .C2(n18680), .A(n18609), .B(n18608), .ZN(
        P3_U2882) );
  INV_X1 U21779 ( .A(n18819), .ZN(n18997) );
  AOI22_X1 U21780 ( .A1(n18990), .A2(n18917), .B1(n18988), .B2(n18610), .ZN(
        n18613) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18611), .B1(
        n18992), .B2(n18969), .ZN(n18612) );
  OAI211_X1 U21782 ( .C1(n18997), .C2(n18680), .A(n18613), .B(n18612), .ZN(
        P3_U2883) );
  INV_X1 U21783 ( .A(n18680), .ZN(n18673) );
  NAND2_X1 U21784 ( .A1(n18614), .A2(n18635), .ZN(n18668) );
  NOR2_X1 U21785 ( .A1(n18673), .A2(n18699), .ZN(n18658) );
  AOI221_X1 U21786 ( .B1(n18615), .B2(n18658), .C1(n18798), .C2(n18658), .A(
        n18750), .ZN(n18618) );
  NOR2_X1 U21787 ( .A1(n19072), .A2(n18658), .ZN(n18631) );
  AOI22_X1 U21788 ( .A1(n18945), .A2(n18652), .B1(n18941), .B2(n18631), .ZN(
        n18617) );
  AOI22_X1 U21789 ( .A1(n18878), .A2(n18699), .B1(n18940), .B2(n18969), .ZN(
        n18616) );
  OAI211_X1 U21790 ( .C1(n18618), .C2(n21155), .A(n18617), .B(n18616), .ZN(
        P3_U2884) );
  AOI22_X1 U21791 ( .A1(n18950), .A2(n18631), .B1(n18949), .B2(n18969), .ZN(
        n18620) );
  INV_X1 U21792 ( .A(n18618), .ZN(n18632) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18632), .B1(
        n18951), .B2(n18699), .ZN(n18619) );
  OAI211_X1 U21794 ( .C1(n18954), .C2(n18650), .A(n18620), .B(n18619), .ZN(
        P3_U2885) );
  INV_X1 U21795 ( .A(n18956), .ZN(n18858) );
  AOI22_X1 U21796 ( .A1(n18955), .A2(n18631), .B1(n18957), .B2(n18969), .ZN(
        n18622) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18632), .B1(
        n18885), .B2(n18699), .ZN(n18621) );
  OAI211_X1 U21798 ( .C1(n18858), .C2(n18650), .A(n18622), .B(n18621), .ZN(
        P3_U2886) );
  AOI22_X1 U21799 ( .A1(n18961), .A2(n18631), .B1(n18963), .B2(n18969), .ZN(
        n18624) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18632), .B1(
        n18889), .B2(n18699), .ZN(n18623) );
  OAI211_X1 U21801 ( .C1(n18861), .C2(n18650), .A(n18624), .B(n18623), .ZN(
        P3_U2887) );
  INV_X1 U21802 ( .A(n18925), .ZN(n18974) );
  AOI22_X1 U21803 ( .A1(n18968), .A2(n18969), .B1(n18967), .B2(n18631), .ZN(
        n18626) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18632), .B1(
        n18970), .B2(n18699), .ZN(n18625) );
  OAI211_X1 U21805 ( .C1(n18974), .C2(n18650), .A(n18626), .B(n18625), .ZN(
        P3_U2888) );
  INV_X1 U21806 ( .A(n18976), .ZN(n18867) );
  AOI22_X1 U21807 ( .A1(n18977), .A2(n18652), .B1(n18975), .B2(n18631), .ZN(
        n18628) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18632), .B1(
        n18864), .B2(n18699), .ZN(n18627) );
  OAI211_X1 U21809 ( .C1(n18867), .C2(n18996), .A(n18628), .B(n18627), .ZN(
        P3_U2889) );
  AOI22_X1 U21810 ( .A1(n18982), .A2(n18969), .B1(n18981), .B2(n18631), .ZN(
        n18630) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18632), .B1(
        n18983), .B2(n18652), .ZN(n18629) );
  OAI211_X1 U21812 ( .C1(n18986), .C2(n18668), .A(n18630), .B(n18629), .ZN(
        P3_U2890) );
  AOI22_X1 U21813 ( .A1(n18992), .A2(n18652), .B1(n18988), .B2(n18631), .ZN(
        n18634) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18632), .B1(
        n18819), .B2(n18699), .ZN(n18633) );
  OAI211_X1 U21815 ( .C1(n18823), .C2(n18996), .A(n18634), .B(n18633), .ZN(
        P3_U2891) );
  NAND2_X1 U21816 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18635), .ZN(
        n18681) );
  INV_X1 U21817 ( .A(n9709), .ZN(n18720) );
  NOR2_X1 U21818 ( .A1(n19072), .A2(n18681), .ZN(n18651) );
  AOI22_X1 U21819 ( .A1(n18941), .A2(n18651), .B1(n18940), .B2(n18652), .ZN(
        n18637) );
  AOI21_X1 U21820 ( .B1(n19044), .B2(n18798), .A(n18657), .ZN(n18727) );
  OAI211_X1 U21821 ( .C1(n9709), .C2(n19169), .A(n18635), .B(n18727), .ZN(
        n18653) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18653), .B1(
        n18945), .B2(n18673), .ZN(n18636) );
  OAI211_X1 U21823 ( .C1(n18948), .C2(n18720), .A(n18637), .B(n18636), .ZN(
        P3_U2892) );
  AOI22_X1 U21824 ( .A1(n18950), .A2(n18651), .B1(n18949), .B2(n18652), .ZN(
        n18639) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18653), .B1(
        n18951), .B2(n9709), .ZN(n18638) );
  OAI211_X1 U21826 ( .C1(n18954), .C2(n18680), .A(n18639), .B(n18638), .ZN(
        P3_U2893) );
  AOI22_X1 U21827 ( .A1(n18956), .A2(n18673), .B1(n18955), .B2(n18651), .ZN(
        n18641) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18653), .B1(
        n18957), .B2(n18652), .ZN(n18640) );
  OAI211_X1 U21829 ( .C1(n18960), .C2(n18720), .A(n18641), .B(n18640), .ZN(
        P3_U2894) );
  AOI22_X1 U21830 ( .A1(n18962), .A2(n18673), .B1(n18961), .B2(n18651), .ZN(
        n18643) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18653), .B1(
        n18963), .B2(n18652), .ZN(n18642) );
  OAI211_X1 U21832 ( .C1(n18966), .C2(n18720), .A(n18643), .B(n18642), .ZN(
        P3_U2895) );
  AOI22_X1 U21833 ( .A1(n18968), .A2(n18652), .B1(n18967), .B2(n18651), .ZN(
        n18645) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18653), .B1(
        n18970), .B2(n9709), .ZN(n18644) );
  OAI211_X1 U21835 ( .C1(n18974), .C2(n18680), .A(n18645), .B(n18644), .ZN(
        P3_U2896) );
  AOI22_X1 U21836 ( .A1(n18977), .A2(n18673), .B1(n18975), .B2(n18651), .ZN(
        n18647) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18653), .B1(
        n18864), .B2(n9709), .ZN(n18646) );
  OAI211_X1 U21838 ( .C1(n18867), .C2(n18650), .A(n18647), .B(n18646), .ZN(
        P3_U2897) );
  INV_X1 U21839 ( .A(n18982), .ZN(n18902) );
  AOI22_X1 U21840 ( .A1(n18983), .A2(n18673), .B1(n18981), .B2(n18651), .ZN(
        n18649) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18653), .B1(
        n18899), .B2(n9709), .ZN(n18648) );
  OAI211_X1 U21842 ( .C1(n18902), .C2(n18650), .A(n18649), .B(n18648), .ZN(
        P3_U2898) );
  AOI22_X1 U21843 ( .A1(n18990), .A2(n18652), .B1(n18988), .B2(n18651), .ZN(
        n18655) );
  AOI22_X1 U21844 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18653), .B1(
        n18992), .B2(n18673), .ZN(n18654) );
  OAI211_X1 U21845 ( .C1(n18997), .C2(n18720), .A(n18655), .B(n18654), .ZN(
        P3_U2899) );
  INV_X1 U21846 ( .A(n18656), .ZN(n19045) );
  INV_X1 U21847 ( .A(n18740), .ZN(n18749) );
  NOR2_X1 U21848 ( .A1(n9709), .A2(n18740), .ZN(n18704) );
  NOR2_X1 U21849 ( .A1(n19072), .A2(n18704), .ZN(n18676) );
  AOI22_X1 U21850 ( .A1(n18941), .A2(n18676), .B1(n18940), .B2(n18673), .ZN(
        n18661) );
  OAI22_X1 U21851 ( .A1(n18658), .A2(n18557), .B1(n18704), .B2(n18657), .ZN(
        n18659) );
  OAI21_X1 U21852 ( .B1(n18740), .B2(n19169), .A(n18659), .ZN(n18677) );
  AOI22_X1 U21853 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18677), .B1(
        n18945), .B2(n18699), .ZN(n18660) );
  OAI211_X1 U21854 ( .C1(n18948), .C2(n18749), .A(n18661), .B(n18660), .ZN(
        P3_U2900) );
  AOI22_X1 U21855 ( .A1(n18881), .A2(n18699), .B1(n18950), .B2(n18676), .ZN(
        n18663) );
  AOI22_X1 U21856 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18677), .B1(
        n18949), .B2(n18673), .ZN(n18662) );
  OAI211_X1 U21857 ( .C1(n18855), .C2(n18749), .A(n18663), .B(n18662), .ZN(
        P3_U2901) );
  AOI22_X1 U21858 ( .A1(n18955), .A2(n18676), .B1(n18957), .B2(n18673), .ZN(
        n18665) );
  AOI22_X1 U21859 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18677), .B1(
        n18885), .B2(n18740), .ZN(n18664) );
  OAI211_X1 U21860 ( .C1(n18858), .C2(n18668), .A(n18665), .B(n18664), .ZN(
        P3_U2902) );
  AOI22_X1 U21861 ( .A1(n18961), .A2(n18676), .B1(n18963), .B2(n18673), .ZN(
        n18667) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18677), .B1(
        n18889), .B2(n18740), .ZN(n18666) );
  OAI211_X1 U21863 ( .C1(n18861), .C2(n18668), .A(n18667), .B(n18666), .ZN(
        P3_U2903) );
  AOI22_X1 U21864 ( .A1(n18925), .A2(n18699), .B1(n18967), .B2(n18676), .ZN(
        n18670) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18677), .B1(
        n18968), .B2(n18673), .ZN(n18669) );
  OAI211_X1 U21866 ( .C1(n18928), .C2(n18749), .A(n18670), .B(n18669), .ZN(
        P3_U2904) );
  AOI22_X1 U21867 ( .A1(n18976), .A2(n18673), .B1(n18975), .B2(n18676), .ZN(
        n18672) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18677), .B1(
        n18977), .B2(n18699), .ZN(n18671) );
  OAI211_X1 U21869 ( .C1(n18980), .C2(n18749), .A(n18672), .B(n18671), .ZN(
        P3_U2905) );
  AOI22_X1 U21870 ( .A1(n18982), .A2(n18673), .B1(n18981), .B2(n18676), .ZN(
        n18675) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18677), .B1(
        n18983), .B2(n18699), .ZN(n18674) );
  OAI211_X1 U21872 ( .C1(n18986), .C2(n18749), .A(n18675), .B(n18674), .ZN(
        P3_U2906) );
  AOI22_X1 U21873 ( .A1(n18992), .A2(n18699), .B1(n18988), .B2(n18676), .ZN(
        n18679) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18677), .B1(
        n18819), .B2(n18740), .ZN(n18678) );
  OAI211_X1 U21875 ( .C1(n18823), .C2(n18680), .A(n18679), .B(n18678), .ZN(
        P3_U2907) );
  NAND2_X1 U21876 ( .A1(n18773), .A2(n18729), .ZN(n18772) );
  AOI22_X1 U21877 ( .A1(n18945), .A2(n9709), .B1(n18941), .B2(n18698), .ZN(
        n18685) );
  INV_X1 U21878 ( .A(n18681), .ZN(n18683) );
  AOI22_X1 U21879 ( .A1(n18585), .A2(n18683), .B1(n18729), .B2(n18682), .ZN(
        n18700) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18700), .B1(
        n18940), .B2(n18699), .ZN(n18684) );
  OAI211_X1 U21881 ( .C1(n18948), .C2(n18772), .A(n18685), .B(n18684), .ZN(
        P3_U2908) );
  AOI22_X1 U21882 ( .A1(n18950), .A2(n18698), .B1(n18949), .B2(n18699), .ZN(
        n18687) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18700), .B1(
        n18881), .B2(n9709), .ZN(n18686) );
  OAI211_X1 U21884 ( .C1(n18855), .C2(n18772), .A(n18687), .B(n18686), .ZN(
        P3_U2909) );
  AOI22_X1 U21885 ( .A1(n18955), .A2(n18698), .B1(n18957), .B2(n18699), .ZN(
        n18689) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18700), .B1(
        n18956), .B2(n9709), .ZN(n18688) );
  OAI211_X1 U21887 ( .C1(n18960), .C2(n18772), .A(n18689), .B(n18688), .ZN(
        P3_U2910) );
  AOI22_X1 U21888 ( .A1(n18961), .A2(n18698), .B1(n18963), .B2(n18699), .ZN(
        n18691) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18700), .B1(
        n18962), .B2(n9709), .ZN(n18690) );
  OAI211_X1 U21890 ( .C1(n18966), .C2(n18772), .A(n18691), .B(n18690), .ZN(
        P3_U2911) );
  AOI22_X1 U21891 ( .A1(n18968), .A2(n18699), .B1(n18967), .B2(n18698), .ZN(
        n18693) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18700), .B1(
        n18925), .B2(n9709), .ZN(n18692) );
  OAI211_X1 U21893 ( .C1(n18928), .C2(n18772), .A(n18693), .B(n18692), .ZN(
        P3_U2912) );
  AOI22_X1 U21894 ( .A1(n18976), .A2(n18699), .B1(n18975), .B2(n18698), .ZN(
        n18695) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18700), .B1(
        n18977), .B2(n9709), .ZN(n18694) );
  OAI211_X1 U21896 ( .C1(n18980), .C2(n18772), .A(n18695), .B(n18694), .ZN(
        P3_U2913) );
  AOI22_X1 U21897 ( .A1(n18982), .A2(n18699), .B1(n18981), .B2(n18698), .ZN(
        n18697) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18700), .B1(
        n18983), .B2(n9709), .ZN(n18696) );
  OAI211_X1 U21899 ( .C1(n18986), .C2(n18772), .A(n18697), .B(n18696), .ZN(
        P3_U2914) );
  AOI22_X1 U21900 ( .A1(n18992), .A2(n9709), .B1(n18988), .B2(n18698), .ZN(
        n18702) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18700), .B1(
        n18990), .B2(n18699), .ZN(n18701) );
  OAI211_X1 U21902 ( .C1(n18997), .C2(n18772), .A(n18702), .B(n18701), .ZN(
        P3_U2915) );
  NOR2_X2 U21903 ( .A1(n18796), .A2(n18703), .ZN(n18788) );
  INV_X1 U21904 ( .A(n18788), .ZN(n18795) );
  INV_X1 U21905 ( .A(n18772), .ZN(n18765) );
  NOR2_X1 U21906 ( .A1(n18765), .A2(n18788), .ZN(n18751) );
  NOR2_X1 U21907 ( .A1(n19072), .A2(n18751), .ZN(n18721) );
  AOI22_X1 U21908 ( .A1(n18941), .A2(n18721), .B1(n18940), .B2(n9709), .ZN(
        n18707) );
  AOI221_X1 U21909 ( .B1(n18751), .B2(n18798), .C1(n18751), .C2(n18704), .A(
        n18750), .ZN(n18705) );
  INV_X1 U21910 ( .A(n18705), .ZN(n18723) );
  AOI22_X1 U21911 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18723), .B1(
        n18945), .B2(n18740), .ZN(n18706) );
  OAI211_X1 U21912 ( .C1(n18948), .C2(n18795), .A(n18707), .B(n18706), .ZN(
        P3_U2916) );
  AOI22_X1 U21913 ( .A1(n18881), .A2(n18740), .B1(n18950), .B2(n18721), .ZN(
        n18709) );
  AOI22_X1 U21914 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18723), .B1(
        n18949), .B2(n9709), .ZN(n18708) );
  OAI211_X1 U21915 ( .C1(n18855), .C2(n18795), .A(n18709), .B(n18708), .ZN(
        P3_U2917) );
  AOI22_X1 U21916 ( .A1(n18956), .A2(n18740), .B1(n18955), .B2(n18721), .ZN(
        n18711) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18723), .B1(
        n18957), .B2(n9709), .ZN(n18710) );
  OAI211_X1 U21918 ( .C1(n18960), .C2(n18795), .A(n18711), .B(n18710), .ZN(
        P3_U2918) );
  AOI22_X1 U21919 ( .A1(n18962), .A2(n18740), .B1(n18961), .B2(n18721), .ZN(
        n18713) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18723), .B1(
        n18963), .B2(n9709), .ZN(n18712) );
  OAI211_X1 U21921 ( .C1(n18966), .C2(n18795), .A(n18713), .B(n18712), .ZN(
        P3_U2919) );
  AOI22_X1 U21922 ( .A1(n18925), .A2(n18740), .B1(n18967), .B2(n18721), .ZN(
        n18715) );
  AOI22_X1 U21923 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18723), .B1(
        n18968), .B2(n9709), .ZN(n18714) );
  OAI211_X1 U21924 ( .C1(n18928), .C2(n18795), .A(n18715), .B(n18714), .ZN(
        P3_U2920) );
  AOI22_X1 U21925 ( .A1(n18976), .A2(n9709), .B1(n18975), .B2(n18721), .ZN(
        n18717) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18723), .B1(
        n18977), .B2(n18740), .ZN(n18716) );
  OAI211_X1 U21927 ( .C1(n18980), .C2(n18795), .A(n18717), .B(n18716), .ZN(
        P3_U2921) );
  AOI22_X1 U21928 ( .A1(n18983), .A2(n18740), .B1(n18981), .B2(n18721), .ZN(
        n18719) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18723), .B1(
        n18899), .B2(n18788), .ZN(n18718) );
  OAI211_X1 U21930 ( .C1(n18902), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2922) );
  AOI22_X1 U21931 ( .A1(n18990), .A2(n9709), .B1(n18988), .B2(n18721), .ZN(
        n18725) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18723), .B1(
        n18992), .B2(n18740), .ZN(n18724) );
  OAI211_X1 U21933 ( .C1(n18997), .C2(n18795), .A(n18725), .B(n18724), .ZN(
        P3_U2923) );
  NAND2_X1 U21934 ( .A1(n19052), .A2(n18726), .ZN(n18774) );
  NOR2_X2 U21935 ( .A1(n19042), .A2(n18774), .ZN(n18810) );
  INV_X1 U21936 ( .A(n18810), .ZN(n18824) );
  NOR2_X1 U21937 ( .A1(n19072), .A2(n18774), .ZN(n18745) );
  AOI22_X1 U21938 ( .A1(n18941), .A2(n18745), .B1(n18940), .B2(n18740), .ZN(
        n18731) );
  NAND3_X1 U21939 ( .A1(n18729), .A2(n18728), .A3(n18727), .ZN(n18746) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18746), .B1(
        n18945), .B2(n18765), .ZN(n18730) );
  OAI211_X1 U21941 ( .C1(n18824), .C2(n18948), .A(n18731), .B(n18730), .ZN(
        P3_U2924) );
  AOI22_X1 U21942 ( .A1(n18881), .A2(n18765), .B1(n18950), .B2(n18745), .ZN(
        n18733) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18746), .B1(
        n18949), .B2(n18740), .ZN(n18732) );
  OAI211_X1 U21944 ( .C1(n18824), .C2(n18855), .A(n18733), .B(n18732), .ZN(
        P3_U2925) );
  AOI22_X1 U21945 ( .A1(n18956), .A2(n18765), .B1(n18955), .B2(n18745), .ZN(
        n18735) );
  AOI22_X1 U21946 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18746), .B1(
        n18957), .B2(n18740), .ZN(n18734) );
  OAI211_X1 U21947 ( .C1(n18824), .C2(n18960), .A(n18735), .B(n18734), .ZN(
        P3_U2926) );
  AOI22_X1 U21948 ( .A1(n18961), .A2(n18745), .B1(n18963), .B2(n18740), .ZN(
        n18737) );
  AOI22_X1 U21949 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18746), .B1(
        n18810), .B2(n18889), .ZN(n18736) );
  OAI211_X1 U21950 ( .C1(n18861), .C2(n18772), .A(n18737), .B(n18736), .ZN(
        P3_U2927) );
  AOI22_X1 U21951 ( .A1(n18925), .A2(n18765), .B1(n18967), .B2(n18745), .ZN(
        n18739) );
  AOI22_X1 U21952 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18746), .B1(
        n18968), .B2(n18740), .ZN(n18738) );
  OAI211_X1 U21953 ( .C1(n18824), .C2(n18928), .A(n18739), .B(n18738), .ZN(
        P3_U2928) );
  AOI22_X1 U21954 ( .A1(n18976), .A2(n18740), .B1(n18975), .B2(n18745), .ZN(
        n18742) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18746), .B1(
        n18977), .B2(n18765), .ZN(n18741) );
  OAI211_X1 U21956 ( .C1(n18824), .C2(n18980), .A(n18742), .B(n18741), .ZN(
        P3_U2929) );
  AOI22_X1 U21957 ( .A1(n18982), .A2(n18740), .B1(n18981), .B2(n18745), .ZN(
        n18744) );
  AOI22_X1 U21958 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18746), .B1(
        n18983), .B2(n18765), .ZN(n18743) );
  OAI211_X1 U21959 ( .C1(n18824), .C2(n18986), .A(n18744), .B(n18743), .ZN(
        P3_U2930) );
  AOI22_X1 U21960 ( .A1(n18992), .A2(n18765), .B1(n18988), .B2(n18745), .ZN(
        n18748) );
  AOI22_X1 U21961 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18746), .B1(
        n18810), .B2(n18819), .ZN(n18747) );
  OAI211_X1 U21962 ( .C1(n18823), .C2(n18749), .A(n18748), .B(n18747), .ZN(
        P3_U2931) );
  NOR2_X2 U21963 ( .A1(n19045), .A2(n18800), .ZN(n18842) );
  INV_X1 U21964 ( .A(n18842), .ZN(n18813) );
  NOR2_X1 U21965 ( .A1(n18842), .A2(n18810), .ZN(n18797) );
  NOR2_X1 U21966 ( .A1(n19072), .A2(n18797), .ZN(n18768) );
  AOI22_X1 U21967 ( .A1(n18941), .A2(n18768), .B1(n18940), .B2(n18765), .ZN(
        n18754) );
  AOI221_X1 U21968 ( .B1(n18797), .B2(n18798), .C1(n18797), .C2(n18751), .A(
        n18750), .ZN(n18752) );
  INV_X1 U21969 ( .A(n18752), .ZN(n18769) );
  AOI22_X1 U21970 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18769), .B1(
        n18945), .B2(n18788), .ZN(n18753) );
  OAI211_X1 U21971 ( .C1(n18813), .C2(n18948), .A(n18754), .B(n18753), .ZN(
        P3_U2932) );
  AOI22_X1 U21972 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18769), .B1(
        n18950), .B2(n18768), .ZN(n18756) );
  AOI22_X1 U21973 ( .A1(n18842), .A2(n18951), .B1(n18949), .B2(n18765), .ZN(
        n18755) );
  OAI211_X1 U21974 ( .C1(n18954), .C2(n18795), .A(n18756), .B(n18755), .ZN(
        P3_U2933) );
  AOI22_X1 U21975 ( .A1(n18955), .A2(n18768), .B1(n18957), .B2(n18765), .ZN(
        n18758) );
  AOI22_X1 U21976 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18769), .B1(
        n18842), .B2(n18885), .ZN(n18757) );
  OAI211_X1 U21977 ( .C1(n18858), .C2(n18795), .A(n18758), .B(n18757), .ZN(
        P3_U2934) );
  AOI22_X1 U21978 ( .A1(n18961), .A2(n18768), .B1(n18963), .B2(n18765), .ZN(
        n18760) );
  AOI22_X1 U21979 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18769), .B1(
        n18842), .B2(n18889), .ZN(n18759) );
  OAI211_X1 U21980 ( .C1(n18861), .C2(n18795), .A(n18760), .B(n18759), .ZN(
        P3_U2935) );
  AOI22_X1 U21981 ( .A1(n18925), .A2(n18788), .B1(n18967), .B2(n18768), .ZN(
        n18762) );
  AOI22_X1 U21982 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18769), .B1(
        n18968), .B2(n18765), .ZN(n18761) );
  OAI211_X1 U21983 ( .C1(n18813), .C2(n18928), .A(n18762), .B(n18761), .ZN(
        P3_U2936) );
  AOI22_X1 U21984 ( .A1(n18977), .A2(n18788), .B1(n18975), .B2(n18768), .ZN(
        n18764) );
  AOI22_X1 U21985 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18769), .B1(
        n18842), .B2(n18864), .ZN(n18763) );
  OAI211_X1 U21986 ( .C1(n18867), .C2(n18772), .A(n18764), .B(n18763), .ZN(
        P3_U2937) );
  AOI22_X1 U21987 ( .A1(n18982), .A2(n18765), .B1(n18981), .B2(n18768), .ZN(
        n18767) );
  AOI22_X1 U21988 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18769), .B1(
        n18983), .B2(n18788), .ZN(n18766) );
  OAI211_X1 U21989 ( .C1(n18813), .C2(n18986), .A(n18767), .B(n18766), .ZN(
        P3_U2938) );
  AOI22_X1 U21990 ( .A1(n18992), .A2(n18788), .B1(n18988), .B2(n18768), .ZN(
        n18771) );
  AOI22_X1 U21991 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18769), .B1(
        n18842), .B2(n18819), .ZN(n18770) );
  OAI211_X1 U21992 ( .C1(n18823), .C2(n18772), .A(n18771), .B(n18770), .ZN(
        P3_U2939) );
  NAND2_X1 U21993 ( .A1(n18846), .A2(n18773), .ZN(n18870) );
  AOI22_X1 U21994 ( .A1(n18945), .A2(n18810), .B1(n18941), .B2(n18791), .ZN(
        n18777) );
  INV_X1 U21995 ( .A(n18774), .ZN(n18775) );
  NOR2_X1 U21996 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18800), .ZN(
        n18826) );
  AOI22_X1 U21997 ( .A1(n18585), .A2(n18775), .B1(n18942), .B2(n18826), .ZN(
        n18792) );
  AOI22_X1 U21998 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18792), .B1(
        n18940), .B2(n18788), .ZN(n18776) );
  OAI211_X1 U21999 ( .C1(n18870), .C2(n18948), .A(n18777), .B(n18776), .ZN(
        P3_U2940) );
  AOI22_X1 U22000 ( .A1(n18950), .A2(n18791), .B1(n18949), .B2(n18788), .ZN(
        n18779) );
  INV_X1 U22001 ( .A(n18870), .ZN(n18872) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18792), .B1(
        n18872), .B2(n18951), .ZN(n18778) );
  OAI211_X1 U22003 ( .C1(n18824), .C2(n18954), .A(n18779), .B(n18778), .ZN(
        P3_U2941) );
  AOI22_X1 U22004 ( .A1(n18955), .A2(n18791), .B1(n18957), .B2(n18788), .ZN(
        n18781) );
  AOI22_X1 U22005 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18792), .B1(
        n18872), .B2(n18885), .ZN(n18780) );
  OAI211_X1 U22006 ( .C1(n18824), .C2(n18858), .A(n18781), .B(n18780), .ZN(
        P3_U2942) );
  AOI22_X1 U22007 ( .A1(n18810), .A2(n18962), .B1(n18961), .B2(n18791), .ZN(
        n18783) );
  AOI22_X1 U22008 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18792), .B1(
        n18963), .B2(n18788), .ZN(n18782) );
  OAI211_X1 U22009 ( .C1(n18870), .C2(n18966), .A(n18783), .B(n18782), .ZN(
        P3_U2943) );
  AOI22_X1 U22010 ( .A1(n18968), .A2(n18788), .B1(n18967), .B2(n18791), .ZN(
        n18785) );
  AOI22_X1 U22011 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18792), .B1(
        n18872), .B2(n18970), .ZN(n18784) );
  OAI211_X1 U22012 ( .C1(n18824), .C2(n18974), .A(n18785), .B(n18784), .ZN(
        P3_U2944) );
  AOI22_X1 U22013 ( .A1(n18976), .A2(n18788), .B1(n18975), .B2(n18791), .ZN(
        n18787) );
  AOI22_X1 U22014 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18792), .B1(
        n18810), .B2(n18977), .ZN(n18786) );
  OAI211_X1 U22015 ( .C1(n18870), .C2(n18980), .A(n18787), .B(n18786), .ZN(
        P3_U2945) );
  AOI22_X1 U22016 ( .A1(n18982), .A2(n18788), .B1(n18981), .B2(n18791), .ZN(
        n18790) );
  AOI22_X1 U22017 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18792), .B1(
        n18810), .B2(n18983), .ZN(n18789) );
  OAI211_X1 U22018 ( .C1(n18870), .C2(n18986), .A(n18790), .B(n18789), .ZN(
        P3_U2946) );
  AOI22_X1 U22019 ( .A1(n18810), .A2(n18992), .B1(n18988), .B2(n18791), .ZN(
        n18794) );
  AOI22_X1 U22020 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18792), .B1(
        n18872), .B2(n18819), .ZN(n18793) );
  OAI211_X1 U22021 ( .C1(n18823), .C2(n18795), .A(n18794), .B(n18793), .ZN(
        P3_U2947) );
  NOR2_X1 U22022 ( .A1(n18800), .A2(n18796), .ZN(n18905) );
  CLKBUF_X1 U22023 ( .A(n18905), .Z(n18894) );
  AOI221_X1 U22024 ( .B1(n18870), .B2(n18798), .C1(n18870), .C2(n18797), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18799) );
  OAI21_X1 U22025 ( .B1(n18894), .B2(n18799), .A(n18849), .ZN(n18820) );
  INV_X1 U22026 ( .A(n18820), .ZN(n18803) );
  INV_X1 U22027 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21086) );
  AOI22_X1 U22028 ( .A1(n18810), .A2(n18940), .B1(n18941), .B2(n18818), .ZN(
        n18802) );
  AOI22_X1 U22029 ( .A1(n18945), .A2(n18842), .B1(n18894), .B2(n18878), .ZN(
        n18801) );
  OAI211_X1 U22030 ( .C1(n18803), .C2(n21086), .A(n18802), .B(n18801), .ZN(
        P3_U2948) );
  AOI22_X1 U22031 ( .A1(n18810), .A2(n18949), .B1(n18818), .B2(n18950), .ZN(
        n18805) );
  AOI22_X1 U22032 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18820), .B1(
        n18905), .B2(n18951), .ZN(n18804) );
  OAI211_X1 U22033 ( .C1(n18813), .C2(n18954), .A(n18805), .B(n18804), .ZN(
        P3_U2949) );
  AOI22_X1 U22034 ( .A1(n18810), .A2(n18957), .B1(n18818), .B2(n18955), .ZN(
        n18807) );
  AOI22_X1 U22035 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18820), .B1(
        n18894), .B2(n18885), .ZN(n18806) );
  OAI211_X1 U22036 ( .C1(n18813), .C2(n18858), .A(n18807), .B(n18806), .ZN(
        P3_U2950) );
  AOI22_X1 U22037 ( .A1(n18810), .A2(n18963), .B1(n18818), .B2(n18961), .ZN(
        n18809) );
  AOI22_X1 U22038 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18820), .B1(
        n18894), .B2(n18889), .ZN(n18808) );
  OAI211_X1 U22039 ( .C1(n18813), .C2(n18861), .A(n18809), .B(n18808), .ZN(
        P3_U2951) );
  AOI22_X1 U22040 ( .A1(n18810), .A2(n18968), .B1(n18818), .B2(n18967), .ZN(
        n18812) );
  AOI22_X1 U22041 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18820), .B1(
        n18905), .B2(n18970), .ZN(n18811) );
  OAI211_X1 U22042 ( .C1(n18813), .C2(n18974), .A(n18812), .B(n18811), .ZN(
        P3_U2952) );
  AOI22_X1 U22043 ( .A1(n18842), .A2(n18977), .B1(n18818), .B2(n18975), .ZN(
        n18815) );
  AOI22_X1 U22044 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18820), .B1(
        n18894), .B2(n18864), .ZN(n18814) );
  OAI211_X1 U22045 ( .C1(n18824), .C2(n18867), .A(n18815), .B(n18814), .ZN(
        P3_U2953) );
  AOI22_X1 U22046 ( .A1(n18842), .A2(n18983), .B1(n18818), .B2(n18981), .ZN(
        n18817) );
  AOI22_X1 U22047 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18820), .B1(
        n18894), .B2(n18899), .ZN(n18816) );
  OAI211_X1 U22048 ( .C1(n18824), .C2(n18902), .A(n18817), .B(n18816), .ZN(
        P3_U2954) );
  AOI22_X1 U22049 ( .A1(n18842), .A2(n18992), .B1(n18818), .B2(n18988), .ZN(
        n18822) );
  AOI22_X1 U22050 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18820), .B1(
        n18894), .B2(n18819), .ZN(n18821) );
  OAI211_X1 U22051 ( .C1(n18824), .C2(n18823), .A(n18822), .B(n18821), .ZN(
        P3_U2955) );
  NAND2_X1 U22052 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18846), .ZN(
        n18825) );
  NOR2_X2 U22053 ( .A1(n19042), .A2(n18825), .ZN(n18934) );
  NOR2_X1 U22054 ( .A1(n19072), .A2(n18825), .ZN(n18841) );
  AOI22_X1 U22055 ( .A1(n18945), .A2(n18872), .B1(n18941), .B2(n18841), .ZN(
        n18828) );
  INV_X1 U22056 ( .A(n18825), .ZN(n18876) );
  AOI22_X1 U22057 ( .A1(n18585), .A2(n18826), .B1(n18942), .B2(n18876), .ZN(
        n18843) );
  AOI22_X1 U22058 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18843), .B1(
        n18842), .B2(n18940), .ZN(n18827) );
  OAI211_X1 U22059 ( .C1(n18948), .C2(n18910), .A(n18828), .B(n18827), .ZN(
        P3_U2956) );
  AOI22_X1 U22060 ( .A1(n18842), .A2(n18949), .B1(n18950), .B2(n18841), .ZN(
        n18830) );
  AOI22_X1 U22061 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18843), .B1(
        n18872), .B2(n18881), .ZN(n18829) );
  OAI211_X1 U22062 ( .C1(n18855), .C2(n18910), .A(n18830), .B(n18829), .ZN(
        P3_U2957) );
  AOI22_X1 U22063 ( .A1(n18842), .A2(n18957), .B1(n18955), .B2(n18841), .ZN(
        n18832) );
  AOI22_X1 U22064 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18843), .B1(
        n18872), .B2(n18956), .ZN(n18831) );
  OAI211_X1 U22065 ( .C1(n18960), .C2(n18910), .A(n18832), .B(n18831), .ZN(
        P3_U2958) );
  AOI22_X1 U22066 ( .A1(n18872), .A2(n18962), .B1(n18961), .B2(n18841), .ZN(
        n18834) );
  AOI22_X1 U22067 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18843), .B1(
        n18842), .B2(n18963), .ZN(n18833) );
  OAI211_X1 U22068 ( .C1(n18966), .C2(n18910), .A(n18834), .B(n18833), .ZN(
        P3_U2959) );
  AOI22_X1 U22069 ( .A1(n18842), .A2(n18968), .B1(n18967), .B2(n18841), .ZN(
        n18836) );
  AOI22_X1 U22070 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18843), .B1(
        n18872), .B2(n18925), .ZN(n18835) );
  OAI211_X1 U22071 ( .C1(n18928), .C2(n18910), .A(n18836), .B(n18835), .ZN(
        P3_U2960) );
  AOI22_X1 U22072 ( .A1(n18842), .A2(n18976), .B1(n18975), .B2(n18841), .ZN(
        n18838) );
  AOI22_X1 U22073 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18843), .B1(
        n18872), .B2(n18977), .ZN(n18837) );
  OAI211_X1 U22074 ( .C1(n18980), .C2(n18910), .A(n18838), .B(n18837), .ZN(
        P3_U2961) );
  AOI22_X1 U22075 ( .A1(n18872), .A2(n18983), .B1(n18981), .B2(n18841), .ZN(
        n18840) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18843), .B1(
        n18842), .B2(n18982), .ZN(n18839) );
  OAI211_X1 U22077 ( .C1(n18986), .C2(n18910), .A(n18840), .B(n18839), .ZN(
        P3_U2962) );
  AOI22_X1 U22078 ( .A1(n18872), .A2(n18992), .B1(n18988), .B2(n18841), .ZN(
        n18845) );
  AOI22_X1 U22079 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18843), .B1(
        n18842), .B2(n18990), .ZN(n18844) );
  OAI211_X1 U22080 ( .C1(n18997), .C2(n18910), .A(n18845), .B(n18844), .ZN(
        P3_U2963) );
  INV_X1 U22081 ( .A(n18944), .ZN(n18877) );
  INV_X1 U22082 ( .A(n9711), .ZN(n18920) );
  AOI21_X1 U22083 ( .B1(n18910), .B2(n18920), .A(n19072), .ZN(n18871) );
  AOI22_X1 U22084 ( .A1(n18945), .A2(n18894), .B1(n18941), .B2(n18871), .ZN(
        n18852) );
  NAND2_X1 U22085 ( .A1(n18913), .A2(n18846), .ZN(n18847) );
  AOI221_X1 U22086 ( .B1(n18848), .B2(n18910), .C1(n18847), .C2(n18910), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18850) );
  OAI21_X1 U22087 ( .B1(n9711), .B2(n18850), .A(n18849), .ZN(n18873) );
  AOI22_X1 U22088 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18873), .B1(
        n18872), .B2(n18940), .ZN(n18851) );
  OAI211_X1 U22089 ( .C1(n18948), .C2(n18920), .A(n18852), .B(n18851), .ZN(
        P3_U2964) );
  AOI22_X1 U22090 ( .A1(n18905), .A2(n18881), .B1(n18950), .B2(n18871), .ZN(
        n18854) );
  AOI22_X1 U22091 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18873), .B1(
        n18872), .B2(n18949), .ZN(n18853) );
  OAI211_X1 U22092 ( .C1(n18855), .C2(n18920), .A(n18854), .B(n18853), .ZN(
        P3_U2965) );
  INV_X1 U22093 ( .A(n18905), .ZN(n18903) );
  AOI22_X1 U22094 ( .A1(n18872), .A2(n18957), .B1(n18955), .B2(n18871), .ZN(
        n18857) );
  AOI22_X1 U22095 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18873), .B1(
        n18885), .B2(n9711), .ZN(n18856) );
  OAI211_X1 U22096 ( .C1(n18903), .C2(n18858), .A(n18857), .B(n18856), .ZN(
        P3_U2966) );
  AOI22_X1 U22097 ( .A1(n18872), .A2(n18963), .B1(n18961), .B2(n18871), .ZN(
        n18860) );
  AOI22_X1 U22098 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18873), .B1(
        n18889), .B2(n9711), .ZN(n18859) );
  OAI211_X1 U22099 ( .C1(n18903), .C2(n18861), .A(n18860), .B(n18859), .ZN(
        P3_U2967) );
  AOI22_X1 U22100 ( .A1(n18872), .A2(n18968), .B1(n18967), .B2(n18871), .ZN(
        n18863) );
  AOI22_X1 U22101 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18873), .B1(
        n18970), .B2(n9711), .ZN(n18862) );
  OAI211_X1 U22102 ( .C1(n18903), .C2(n18974), .A(n18863), .B(n18862), .ZN(
        P3_U2968) );
  AOI22_X1 U22103 ( .A1(n18905), .A2(n18977), .B1(n18975), .B2(n18871), .ZN(
        n18866) );
  AOI22_X1 U22104 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18873), .B1(
        n18864), .B2(n9711), .ZN(n18865) );
  OAI211_X1 U22105 ( .C1(n18870), .C2(n18867), .A(n18866), .B(n18865), .ZN(
        P3_U2969) );
  AOI22_X1 U22106 ( .A1(n18894), .A2(n18983), .B1(n18981), .B2(n18871), .ZN(
        n18869) );
  AOI22_X1 U22107 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18873), .B1(
        n18899), .B2(n9711), .ZN(n18868) );
  OAI211_X1 U22108 ( .C1(n18870), .C2(n18902), .A(n18869), .B(n18868), .ZN(
        P3_U2970) );
  AOI22_X1 U22109 ( .A1(n18872), .A2(n18990), .B1(n18988), .B2(n18871), .ZN(
        n18875) );
  AOI22_X1 U22110 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18873), .B1(
        n18905), .B2(n18992), .ZN(n18874) );
  OAI211_X1 U22111 ( .C1(n18997), .C2(n18920), .A(n18875), .B(n18874), .ZN(
        P3_U2971) );
  AOI22_X1 U22112 ( .A1(n18585), .A2(n18876), .B1(n18944), .B2(n18942), .ZN(
        n18906) );
  INV_X1 U22113 ( .A(n18906), .ZN(n18892) );
  NOR2_X1 U22114 ( .A1(n19072), .A2(n18877), .ZN(n18904) );
  AOI22_X1 U22115 ( .A1(n18945), .A2(n18934), .B1(n18941), .B2(n18904), .ZN(
        n18880) );
  AOI22_X1 U22116 ( .A1(n18894), .A2(n18940), .B1(n18878), .B2(n18991), .ZN(
        n18879) );
  OAI211_X1 U22117 ( .C1(n21295), .C2(n18892), .A(n18880), .B(n18879), .ZN(
        P3_U2972) );
  INV_X1 U22118 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18884) );
  AOI22_X1 U22119 ( .A1(n18881), .A2(n18934), .B1(n18950), .B2(n18904), .ZN(
        n18883) );
  AOI22_X1 U22120 ( .A1(n18905), .A2(n18949), .B1(n18951), .B2(n18991), .ZN(
        n18882) );
  OAI211_X1 U22121 ( .C1(n18884), .C2(n18892), .A(n18883), .B(n18882), .ZN(
        P3_U2973) );
  INV_X1 U22122 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18888) );
  AOI22_X1 U22123 ( .A1(n18956), .A2(n18934), .B1(n18955), .B2(n18904), .ZN(
        n18887) );
  AOI22_X1 U22124 ( .A1(n18905), .A2(n18957), .B1(n18885), .B2(n18991), .ZN(
        n18886) );
  OAI211_X1 U22125 ( .C1(n18888), .C2(n18892), .A(n18887), .B(n18886), .ZN(
        P3_U2974) );
  INV_X1 U22126 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18893) );
  AOI22_X1 U22127 ( .A1(n18962), .A2(n18934), .B1(n18961), .B2(n18904), .ZN(
        n18891) );
  AOI22_X1 U22128 ( .A1(n18894), .A2(n18963), .B1(n18889), .B2(n18991), .ZN(
        n18890) );
  OAI211_X1 U22129 ( .C1(n18893), .C2(n18892), .A(n18891), .B(n18890), .ZN(
        P3_U2975) );
  AOI22_X1 U22130 ( .A1(n18894), .A2(n18968), .B1(n18967), .B2(n18904), .ZN(
        n18896) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18906), .B1(
        n18970), .B2(n18991), .ZN(n18895) );
  OAI211_X1 U22132 ( .C1(n18974), .C2(n18910), .A(n18896), .B(n18895), .ZN(
        P3_U2976) );
  AOI22_X1 U22133 ( .A1(n18905), .A2(n18976), .B1(n18975), .B2(n18904), .ZN(
        n18898) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18906), .B1(
        n18977), .B2(n18934), .ZN(n18897) );
  OAI211_X1 U22135 ( .C1(n18980), .C2(n18973), .A(n18898), .B(n18897), .ZN(
        P3_U2977) );
  AOI22_X1 U22136 ( .A1(n18983), .A2(n18934), .B1(n18981), .B2(n18904), .ZN(
        n18901) );
  AOI22_X1 U22137 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18906), .B1(
        n18899), .B2(n18991), .ZN(n18900) );
  OAI211_X1 U22138 ( .C1(n18903), .C2(n18902), .A(n18901), .B(n18900), .ZN(
        P3_U2978) );
  AOI22_X1 U22139 ( .A1(n18905), .A2(n18990), .B1(n18988), .B2(n18904), .ZN(
        n18908) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18906), .B1(
        n18992), .B2(n18934), .ZN(n18907) );
  OAI211_X1 U22141 ( .C1(n18997), .C2(n18973), .A(n18908), .B(n18907), .ZN(
        P3_U2979) );
  INV_X1 U22142 ( .A(n18917), .ZN(n18938) );
  NOR2_X1 U22143 ( .A1(n19072), .A2(n18909), .ZN(n18933) );
  AOI22_X1 U22144 ( .A1(n18945), .A2(n9711), .B1(n18941), .B2(n18933), .ZN(
        n18916) );
  NAND2_X1 U22145 ( .A1(n18910), .A2(n18920), .ZN(n18912) );
  OAI221_X1 U22146 ( .B1(n18914), .B2(n18913), .C1(n18914), .C2(n18912), .A(
        n18911), .ZN(n18935) );
  AOI22_X1 U22147 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18935), .B1(
        n18940), .B2(n18934), .ZN(n18915) );
  OAI211_X1 U22148 ( .C1(n18948), .C2(n18938), .A(n18916), .B(n18915), .ZN(
        P3_U2980) );
  AOI22_X1 U22149 ( .A1(n18950), .A2(n18933), .B1(n18949), .B2(n18934), .ZN(
        n18919) );
  AOI22_X1 U22150 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18935), .B1(
        n18951), .B2(n18917), .ZN(n18918) );
  OAI211_X1 U22151 ( .C1(n18954), .C2(n18920), .A(n18919), .B(n18918), .ZN(
        P3_U2981) );
  AOI22_X1 U22152 ( .A1(n18956), .A2(n9711), .B1(n18955), .B2(n18933), .ZN(
        n18922) );
  AOI22_X1 U22153 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18935), .B1(
        n18957), .B2(n18934), .ZN(n18921) );
  OAI211_X1 U22154 ( .C1(n18960), .C2(n18938), .A(n18922), .B(n18921), .ZN(
        P3_U2982) );
  AOI22_X1 U22155 ( .A1(n18962), .A2(n9711), .B1(n18961), .B2(n18933), .ZN(
        n18924) );
  AOI22_X1 U22156 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18935), .B1(
        n18963), .B2(n18934), .ZN(n18923) );
  OAI211_X1 U22157 ( .C1(n18966), .C2(n18938), .A(n18924), .B(n18923), .ZN(
        P3_U2983) );
  AOI22_X1 U22158 ( .A1(n18925), .A2(n9711), .B1(n18967), .B2(n18933), .ZN(
        n18927) );
  AOI22_X1 U22159 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18935), .B1(
        n18968), .B2(n18934), .ZN(n18926) );
  OAI211_X1 U22160 ( .C1(n18928), .C2(n18938), .A(n18927), .B(n18926), .ZN(
        P3_U2984) );
  AOI22_X1 U22161 ( .A1(n18976), .A2(n18934), .B1(n18975), .B2(n18933), .ZN(
        n18930) );
  AOI22_X1 U22162 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18935), .B1(
        n18977), .B2(n9711), .ZN(n18929) );
  OAI211_X1 U22163 ( .C1(n18980), .C2(n18938), .A(n18930), .B(n18929), .ZN(
        P3_U2985) );
  AOI22_X1 U22164 ( .A1(n18982), .A2(n18934), .B1(n18981), .B2(n18933), .ZN(
        n18932) );
  AOI22_X1 U22165 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18935), .B1(
        n18983), .B2(n9711), .ZN(n18931) );
  OAI211_X1 U22166 ( .C1(n18986), .C2(n18938), .A(n18932), .B(n18931), .ZN(
        P3_U2986) );
  AOI22_X1 U22167 ( .A1(n18990), .A2(n18934), .B1(n18988), .B2(n18933), .ZN(
        n18937) );
  AOI22_X1 U22168 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18935), .B1(
        n18992), .B2(n9711), .ZN(n18936) );
  OAI211_X1 U22169 ( .C1(n18997), .C2(n18938), .A(n18937), .B(n18936), .ZN(
        P3_U2987) );
  INV_X1 U22170 ( .A(n18943), .ZN(n18939) );
  NOR2_X1 U22171 ( .A1(n19072), .A2(n18939), .ZN(n18987) );
  AOI22_X1 U22172 ( .A1(n18941), .A2(n18987), .B1(n18940), .B2(n9711), .ZN(
        n18947) );
  AOI22_X1 U22173 ( .A1(n18585), .A2(n18944), .B1(n18943), .B2(n18942), .ZN(
        n18993) );
  AOI22_X1 U22174 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18993), .B1(
        n18945), .B2(n18991), .ZN(n18946) );
  OAI211_X1 U22175 ( .C1(n18948), .C2(n18996), .A(n18947), .B(n18946), .ZN(
        P3_U2988) );
  AOI22_X1 U22176 ( .A1(n18950), .A2(n18987), .B1(n18949), .B2(n9711), .ZN(
        n18953) );
  AOI22_X1 U22177 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18993), .B1(
        n18951), .B2(n18969), .ZN(n18952) );
  OAI211_X1 U22178 ( .C1(n18954), .C2(n18973), .A(n18953), .B(n18952), .ZN(
        P3_U2989) );
  AOI22_X1 U22179 ( .A1(n18956), .A2(n18991), .B1(n18955), .B2(n18987), .ZN(
        n18959) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18993), .B1(
        n18957), .B2(n9711), .ZN(n18958) );
  OAI211_X1 U22181 ( .C1(n18960), .C2(n18996), .A(n18959), .B(n18958), .ZN(
        P3_U2990) );
  AOI22_X1 U22182 ( .A1(n18962), .A2(n18991), .B1(n18961), .B2(n18987), .ZN(
        n18965) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18993), .B1(
        n18963), .B2(n9711), .ZN(n18964) );
  OAI211_X1 U22184 ( .C1(n18966), .C2(n18996), .A(n18965), .B(n18964), .ZN(
        P3_U2991) );
  AOI22_X1 U22185 ( .A1(n18968), .A2(n9711), .B1(n18967), .B2(n18987), .ZN(
        n18972) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18993), .B1(
        n18970), .B2(n18969), .ZN(n18971) );
  OAI211_X1 U22187 ( .C1(n18974), .C2(n18973), .A(n18972), .B(n18971), .ZN(
        P3_U2992) );
  AOI22_X1 U22188 ( .A1(n18976), .A2(n9711), .B1(n18975), .B2(n18987), .ZN(
        n18979) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18993), .B1(
        n18977), .B2(n18991), .ZN(n18978) );
  OAI211_X1 U22190 ( .C1(n18980), .C2(n18996), .A(n18979), .B(n18978), .ZN(
        P3_U2993) );
  AOI22_X1 U22191 ( .A1(n18982), .A2(n9711), .B1(n18981), .B2(n18987), .ZN(
        n18985) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18993), .B1(
        n18983), .B2(n18991), .ZN(n18984) );
  OAI211_X1 U22193 ( .C1(n18986), .C2(n18996), .A(n18985), .B(n18984), .ZN(
        P3_U2994) );
  AOI22_X1 U22194 ( .A1(n18990), .A2(n9711), .B1(n18988), .B2(n18987), .ZN(
        n18995) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18993), .B1(
        n18992), .B2(n18991), .ZN(n18994) );
  OAI211_X1 U22196 ( .C1(n18997), .C2(n18996), .A(n18995), .B(n18994), .ZN(
        P3_U2995) );
  INV_X1 U22197 ( .A(n18998), .ZN(n19005) );
  NOR2_X1 U22198 ( .A1(n19010), .A2(n18999), .ZN(n19002) );
  OAI222_X1 U22199 ( .A1(n19005), .A2(n19004), .B1(n19003), .B2(n19002), .C1(
        n19001), .C2(n19000), .ZN(n19209) );
  INV_X1 U22200 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U22201 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n19006), .ZN(n19008) );
  OAI211_X1 U22202 ( .C1(n19035), .C2(n19009), .A(n19008), .B(n19007), .ZN(
        n19058) );
  NOR2_X1 U22203 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19020), .ZN(
        n19039) );
  INV_X1 U22204 ( .A(n19039), .ZN(n19011) );
  NAND2_X1 U22205 ( .A1(n19186), .A2(n19033), .ZN(n19017) );
  AOI22_X1 U22206 ( .A1(n19012), .A2(n19011), .B1(n19010), .B2(n19017), .ZN(
        n19013) );
  NOR2_X1 U22207 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19013), .ZN(
        n19171) );
  AOI21_X1 U22208 ( .B1(n19016), .B2(n19015), .A(n19014), .ZN(n19023) );
  OAI21_X1 U22209 ( .B1(n19023), .B2(n19018), .A(n19017), .ZN(n19019) );
  AOI21_X1 U22210 ( .B1(n19027), .B2(n19020), .A(n19019), .ZN(n19172) );
  AOI21_X1 U22211 ( .B1(n19172), .B2(n19035), .A(n19175), .ZN(n19021) );
  AOI21_X1 U22212 ( .B1(n19035), .B2(n19171), .A(n19021), .ZN(n19056) );
  INV_X1 U22213 ( .A(n19035), .ZN(n19047) );
  AOI221_X1 U22214 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19023), 
        .C1(n19022), .C2(n19023), .A(n19186), .ZN(n19034) );
  NOR2_X1 U22215 ( .A1(n19024), .A2(n19198), .ZN(n19026) );
  OAI211_X1 U22216 ( .C1(n19026), .C2(n19025), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n19186), .ZN(n19030) );
  OAI211_X1 U22217 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n19028), .B(n19027), .ZN(
        n19029) );
  OAI211_X1 U22218 ( .C1(n19182), .C2(n19031), .A(n19030), .B(n19029), .ZN(
        n19032) );
  AOI21_X1 U22219 ( .B1(n19034), .B2(n19033), .A(n19032), .ZN(n19178) );
  AOI22_X1 U22220 ( .A1(n19047), .A2(n19186), .B1(n19178), .B2(n19035), .ZN(
        n19051) );
  NOR2_X1 U22221 ( .A1(n19037), .A2(n19036), .ZN(n19041) );
  AOI22_X1 U22222 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19038), .B1(
        n19041), .B2(n19198), .ZN(n19194) );
  OAI22_X1 U22223 ( .A1(n19041), .A2(n19040), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19039), .ZN(n19190) );
  OR3_X1 U22224 ( .A1(n19194), .A2(n19044), .A3(n19042), .ZN(n19043) );
  AOI22_X1 U22225 ( .A1(n19194), .A2(n19044), .B1(n19190), .B2(n19043), .ZN(
        n19046) );
  OAI21_X1 U22226 ( .B1(n19047), .B2(n19046), .A(n19045), .ZN(n19050) );
  AND2_X1 U22227 ( .A1(n19051), .A2(n19050), .ZN(n19048) );
  OAI221_X1 U22228 ( .B1(n19051), .B2(n19050), .C1(n19049), .C2(n19048), .A(
        n19053), .ZN(n19055) );
  AOI21_X1 U22229 ( .B1(n19053), .B2(n19052), .A(n19051), .ZN(n19054) );
  AOI222_X1 U22230 ( .A1(n19056), .A2(n19055), .B1(n19056), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19055), .C2(n19054), .ZN(
        n19057) );
  NOR4_X1 U22231 ( .A1(n19059), .A2(n19209), .A3(n19058), .A4(n19057), .ZN(
        n19069) );
  AOI22_X1 U22232 ( .A1(n19216), .A2(n17778), .B1(n19193), .B2(n19221), .ZN(
        n19060) );
  INV_X1 U22233 ( .A(n19060), .ZN(n19065) );
  OAI211_X1 U22234 ( .C1(n19062), .C2(n19061), .A(n19213), .B(n19069), .ZN(
        n19168) );
  OAI21_X1 U22235 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19210), .A(n19168), 
        .ZN(n19070) );
  NOR2_X1 U22236 ( .A1(n19063), .A2(n19070), .ZN(n19064) );
  MUX2_X1 U22237 ( .A(n19065), .B(n19064), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19067) );
  OAI211_X1 U22238 ( .C1(n19069), .C2(n19068), .A(n19067), .B(n19066), .ZN(
        P3_U2996) );
  NAND2_X1 U22239 ( .A1(n19216), .A2(n17778), .ZN(n19075) );
  NOR4_X1 U22240 ( .A1(n19218), .A2(n19179), .A3(n19210), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19078) );
  INV_X1 U22241 ( .A(n19078), .ZN(n19074) );
  OR3_X1 U22242 ( .A1(n19072), .A2(n19071), .A3(n19070), .ZN(n19073) );
  NAND4_X1 U22243 ( .A1(n19076), .A2(n19075), .A3(n19074), .A4(n19073), .ZN(
        P3_U2997) );
  OAI21_X1 U22244 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19077), .ZN(n19079) );
  AOI21_X1 U22245 ( .B1(n19080), .B2(n19079), .A(n19078), .ZN(P3_U2998) );
  AND2_X1 U22246 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19081), .ZN(
        P3_U2999) );
  AND2_X1 U22247 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19081), .ZN(
        P3_U3000) );
  AND2_X1 U22248 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19081), .ZN(
        P3_U3001) );
  AND2_X1 U22249 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19081), .ZN(
        P3_U3002) );
  AND2_X1 U22250 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19081), .ZN(
        P3_U3003) );
  AND2_X1 U22251 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19081), .ZN(
        P3_U3004) );
  INV_X1 U22252 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21300) );
  NOR2_X1 U22253 ( .A1(n21300), .A2(n19166), .ZN(P3_U3005) );
  AND2_X1 U22254 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19081), .ZN(
        P3_U3006) );
  AND2_X1 U22255 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19081), .ZN(
        P3_U3007) );
  AND2_X1 U22256 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19081), .ZN(
        P3_U3008) );
  AND2_X1 U22257 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19081), .ZN(
        P3_U3009) );
  AND2_X1 U22258 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19081), .ZN(
        P3_U3010) );
  AND2_X1 U22259 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19081), .ZN(
        P3_U3011) );
  AND2_X1 U22260 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19081), .ZN(
        P3_U3012) );
  AND2_X1 U22261 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19081), .ZN(
        P3_U3013) );
  AND2_X1 U22262 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19081), .ZN(
        P3_U3014) );
  AND2_X1 U22263 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19081), .ZN(
        P3_U3015) );
  AND2_X1 U22264 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19081), .ZN(
        P3_U3016) );
  AND2_X1 U22265 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19081), .ZN(
        P3_U3017) );
  AND2_X1 U22266 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19081), .ZN(
        P3_U3018) );
  AND2_X1 U22267 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19081), .ZN(
        P3_U3019) );
  AND2_X1 U22268 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19081), .ZN(
        P3_U3020) );
  AND2_X1 U22269 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19081), .ZN(P3_U3021) );
  AND2_X1 U22270 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19081), .ZN(P3_U3022) );
  AND2_X1 U22271 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19081), .ZN(P3_U3023) );
  AND2_X1 U22272 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19081), .ZN(P3_U3024) );
  AND2_X1 U22273 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19081), .ZN(P3_U3025) );
  AND2_X1 U22274 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19081), .ZN(P3_U3026) );
  AND2_X1 U22275 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19081), .ZN(P3_U3027) );
  AND2_X1 U22276 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19081), .ZN(P3_U3028) );
  INV_X1 U22277 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19223) );
  AOI21_X1 U22278 ( .B1(HOLD), .B2(n19082), .A(n19223), .ZN(n19085) );
  NOR2_X1 U22279 ( .A1(n19210), .A2(n19083), .ZN(n19091) );
  OAI21_X1 U22280 ( .B1(n19091), .B2(n19096), .A(n19098), .ZN(n19084) );
  NAND3_X1 U22281 ( .A1(NA), .A2(n19096), .A3(n19083), .ZN(n19090) );
  OAI211_X1 U22282 ( .C1(n19225), .C2(n19085), .A(n19084), .B(n19090), .ZN(
        P3_U3029) );
  AOI21_X1 U22283 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19086) );
  AOI21_X1 U22284 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n19086), .ZN(
        n19087) );
  AOI22_X1 U22285 ( .A1(n19216), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19087), .ZN(n19089) );
  NAND2_X1 U22286 ( .A1(n19089), .A2(n19088), .ZN(P3_U3030) );
  AOI21_X1 U22287 ( .B1(n19096), .B2(n19090), .A(n19091), .ZN(n19097) );
  NOR2_X1 U22288 ( .A1(n19098), .A2(n20981), .ZN(n19094) );
  INV_X1 U22289 ( .A(n19091), .ZN(n19092) );
  OAI22_X1 U22290 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19092), .ZN(n19093) );
  OAI22_X1 U22291 ( .A1(n19094), .A2(n19093), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19095) );
  OAI22_X1 U22292 ( .A1(n19097), .A2(n19098), .B1(n19096), .B2(n19095), .ZN(
        P3_U3031) );
  OAI222_X1 U22293 ( .A1(n19155), .A2(n21303), .B1(n19100), .B2(n19225), .C1(
        n19099), .C2(n19156), .ZN(P3_U3032) );
  OAI222_X1 U22294 ( .A1(n21303), .A2(n19156), .B1(n19101), .B2(n19225), .C1(
        n19102), .C2(n19155), .ZN(P3_U3033) );
  OAI222_X1 U22295 ( .A1(n19155), .A2(n19104), .B1(n19103), .B2(n19225), .C1(
        n19102), .C2(n19156), .ZN(P3_U3034) );
  OAI222_X1 U22296 ( .A1(n19155), .A2(n19106), .B1(n19105), .B2(n19225), .C1(
        n19104), .C2(n19156), .ZN(P3_U3035) );
  OAI222_X1 U22297 ( .A1(n19155), .A2(n19109), .B1(n19107), .B2(n19225), .C1(
        n19106), .C2(n19156), .ZN(P3_U3036) );
  OAI222_X1 U22298 ( .A1(n19109), .A2(n19156), .B1(n19108), .B2(n19225), .C1(
        n19110), .C2(n19155), .ZN(P3_U3037) );
  OAI222_X1 U22299 ( .A1(n19155), .A2(n19113), .B1(n19111), .B2(n19225), .C1(
        n19110), .C2(n19156), .ZN(P3_U3038) );
  OAI222_X1 U22300 ( .A1(n19113), .A2(n19156), .B1(n19112), .B2(n19225), .C1(
        n19114), .C2(n19155), .ZN(P3_U3039) );
  OAI222_X1 U22301 ( .A1(n19155), .A2(n19116), .B1(n19115), .B2(n19225), .C1(
        n19114), .C2(n19156), .ZN(P3_U3040) );
  OAI222_X1 U22302 ( .A1(n19155), .A2(n19118), .B1(n19117), .B2(n19225), .C1(
        n19116), .C2(n19156), .ZN(P3_U3041) );
  OAI222_X1 U22303 ( .A1(n19155), .A2(n19120), .B1(n19119), .B2(n19225), .C1(
        n19118), .C2(n19156), .ZN(P3_U3042) );
  OAI222_X1 U22304 ( .A1(n19155), .A2(n19122), .B1(n19121), .B2(n19225), .C1(
        n19120), .C2(n19156), .ZN(P3_U3043) );
  OAI222_X1 U22305 ( .A1(n19155), .A2(n19124), .B1(n19123), .B2(n19225), .C1(
        n19122), .C2(n19156), .ZN(P3_U3044) );
  OAI222_X1 U22306 ( .A1(n19155), .A2(n19127), .B1(n19125), .B2(n19225), .C1(
        n19124), .C2(n19156), .ZN(P3_U3045) );
  OAI222_X1 U22307 ( .A1(n19127), .A2(n19156), .B1(n19126), .B2(n19225), .C1(
        n19128), .C2(n19155), .ZN(P3_U3046) );
  OAI222_X1 U22308 ( .A1(n19155), .A2(n19130), .B1(n19129), .B2(n19225), .C1(
        n19128), .C2(n19156), .ZN(P3_U3047) );
  OAI222_X1 U22309 ( .A1(n19155), .A2(n19132), .B1(n19131), .B2(n19225), .C1(
        n19130), .C2(n19156), .ZN(P3_U3048) );
  OAI222_X1 U22310 ( .A1(n19155), .A2(n19134), .B1(n19133), .B2(n19225), .C1(
        n19132), .C2(n19156), .ZN(P3_U3049) );
  OAI222_X1 U22311 ( .A1(n19155), .A2(n19136), .B1(n19135), .B2(n19225), .C1(
        n19134), .C2(n19156), .ZN(P3_U3050) );
  OAI222_X1 U22312 ( .A1(n19155), .A2(n19138), .B1(n19137), .B2(n19225), .C1(
        n19136), .C2(n19156), .ZN(P3_U3051) );
  OAI222_X1 U22313 ( .A1(n19155), .A2(n21123), .B1(n19139), .B2(n19225), .C1(
        n19138), .C2(n19156), .ZN(P3_U3052) );
  OAI222_X1 U22314 ( .A1(n21123), .A2(n19156), .B1(n19140), .B2(n19225), .C1(
        n19142), .C2(n19155), .ZN(P3_U3053) );
  OAI222_X1 U22315 ( .A1(n19142), .A2(n19156), .B1(n19141), .B2(n19225), .C1(
        n19144), .C2(n19155), .ZN(P3_U3054) );
  OAI222_X1 U22316 ( .A1(n19144), .A2(n19156), .B1(n19143), .B2(n19225), .C1(
        n19145), .C2(n19155), .ZN(P3_U3055) );
  OAI222_X1 U22317 ( .A1(n19155), .A2(n19147), .B1(n19146), .B2(n19225), .C1(
        n19145), .C2(n19156), .ZN(P3_U3056) );
  OAI222_X1 U22318 ( .A1(n19155), .A2(n19150), .B1(n19148), .B2(n19225), .C1(
        n19147), .C2(n19156), .ZN(P3_U3057) );
  INV_X1 U22319 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19151) );
  OAI222_X1 U22320 ( .A1(n19156), .A2(n19150), .B1(n19149), .B2(n19225), .C1(
        n19151), .C2(n19155), .ZN(P3_U3058) );
  OAI222_X1 U22321 ( .A1(n19155), .A2(n19153), .B1(n19152), .B2(n19225), .C1(
        n19151), .C2(n19156), .ZN(P3_U3059) );
  OAI222_X1 U22322 ( .A1(n19155), .A2(n19157), .B1(n19154), .B2(n19225), .C1(
        n19153), .C2(n19156), .ZN(P3_U3060) );
  OAI222_X1 U22323 ( .A1(n19155), .A2(n21249), .B1(n19158), .B2(n19225), .C1(
        n19157), .C2(n19156), .ZN(P3_U3061) );
  OAI22_X1 U22324 ( .A1(n19226), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19225), .ZN(n19159) );
  INV_X1 U22325 ( .A(n19159), .ZN(P3_U3274) );
  OAI22_X1 U22326 ( .A1(n19226), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19225), .ZN(n19160) );
  INV_X1 U22327 ( .A(n19160), .ZN(P3_U3275) );
  OAI22_X1 U22328 ( .A1(n19226), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19225), .ZN(n19161) );
  INV_X1 U22329 ( .A(n19161), .ZN(P3_U3276) );
  OAI22_X1 U22330 ( .A1(n19226), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19225), .ZN(n19162) );
  INV_X1 U22331 ( .A(n19162), .ZN(P3_U3277) );
  OAI21_X1 U22332 ( .B1(n19166), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19164), 
        .ZN(n19163) );
  INV_X1 U22333 ( .A(n19163), .ZN(P3_U3280) );
  OAI21_X1 U22334 ( .B1(n19166), .B2(n19165), .A(n19164), .ZN(P3_U3281) );
  OAI221_X1 U22335 ( .B1(n19169), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19169), 
        .C2(n19168), .A(n19167), .ZN(P3_U3282) );
  AOI22_X1 U22336 ( .A1(n19229), .A2(n19171), .B1(n19193), .B2(n19170), .ZN(
        n19177) );
  INV_X1 U22337 ( .A(n19199), .ZN(n19196) );
  OAI21_X1 U22338 ( .B1(n19173), .B2(n19172), .A(n19196), .ZN(n19174) );
  INV_X1 U22339 ( .A(n19174), .ZN(n19176) );
  OAI22_X1 U22340 ( .A1(n19199), .A2(n19177), .B1(n19176), .B2(n19175), .ZN(
        P3_U3285) );
  INV_X1 U22341 ( .A(n19178), .ZN(n19184) );
  NOR2_X1 U22342 ( .A1(n19179), .A2(n19195), .ZN(n19187) );
  OAI22_X1 U22343 ( .A1(n19181), .A2(n19180), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19188) );
  INV_X1 U22344 ( .A(n19188), .ZN(n19183) );
  AOI222_X1 U22345 ( .A1(n19184), .A2(n19229), .B1(n19187), .B2(n19183), .C1(
        n19193), .C2(n19182), .ZN(n19185) );
  AOI22_X1 U22346 ( .A1(n19199), .A2(n19186), .B1(n19185), .B2(n19196), .ZN(
        P3_U3288) );
  AOI222_X1 U22347 ( .A1(n19190), .A2(n19229), .B1(n19193), .B2(n19189), .C1(
        n19188), .C2(n19187), .ZN(n19191) );
  AOI22_X1 U22348 ( .A1(n19199), .A2(n19192), .B1(n19191), .B2(n19196), .ZN(
        P3_U3289) );
  AOI222_X1 U22349 ( .A1(n19195), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19229), 
        .B2(n19194), .C1(n19198), .C2(n19193), .ZN(n19197) );
  AOI22_X1 U22350 ( .A1(n19199), .A2(n19198), .B1(n19197), .B2(n19196), .ZN(
        P3_U3290) );
  AOI211_X1 U22351 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19200) );
  AOI21_X1 U22352 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19200), .ZN(n19202) );
  INV_X1 U22353 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19201) );
  AOI22_X1 U22354 ( .A1(n19206), .A2(n19202), .B1(n19201), .B2(n19203), .ZN(
        P3_U3292) );
  NOR2_X1 U22355 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19205) );
  INV_X1 U22356 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19204) );
  AOI22_X1 U22357 ( .A1(n19206), .A2(n19205), .B1(n19204), .B2(n19203), .ZN(
        P3_U3293) );
  INV_X1 U22358 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19232) );
  OAI22_X1 U22359 ( .A1(n19226), .A2(n19232), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n19225), .ZN(n19207) );
  INV_X1 U22360 ( .A(n19207), .ZN(P3_U3294) );
  MUX2_X1 U22361 ( .A(P3_MORE_REG_SCAN_IN), .B(n19209), .S(n19208), .Z(
        P3_U3295) );
  AOI21_X1 U22362 ( .B1(n17778), .B2(n19210), .A(n19231), .ZN(n19211) );
  OAI21_X1 U22363 ( .B1(n19213), .B2(n19212), .A(n19211), .ZN(n19224) );
  OAI21_X1 U22364 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19215), .A(n19214), 
        .ZN(n19217) );
  AOI211_X1 U22365 ( .C1(n19230), .C2(n19217), .A(n19216), .B(n19228), .ZN(
        n19219) );
  NOR2_X1 U22366 ( .A1(n19219), .A2(n19218), .ZN(n19220) );
  OAI21_X1 U22367 ( .B1(n19221), .B2(n19220), .A(n19224), .ZN(n19222) );
  OAI21_X1 U22368 ( .B1(n19224), .B2(n19223), .A(n19222), .ZN(P3_U3296) );
  OAI22_X1 U22369 ( .A1(n19226), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19225), .ZN(n19227) );
  INV_X1 U22370 ( .A(n19227), .ZN(P3_U3297) );
  AOI21_X1 U22371 ( .B1(n19229), .B2(n19228), .A(n19231), .ZN(n19235) );
  AOI22_X1 U22372 ( .A1(n19235), .A2(n19232), .B1(n19231), .B2(n19230), .ZN(
        P3_U3298) );
  INV_X1 U22373 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19234) );
  AOI21_X1 U22374 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(P3_U3299) );
  NAND2_X1 U22375 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20200), .ZN(n20193) );
  NAND2_X1 U22376 ( .A1(n20189), .A2(n20182), .ZN(n20190) );
  OAI21_X1 U22377 ( .B1(n20189), .B2(n20193), .A(n20190), .ZN(n20256) );
  AOI21_X1 U22378 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20256), .ZN(n19236) );
  INV_X1 U22379 ( .A(n19236), .ZN(P2_U2815) );
  AOI21_X1 U22380 ( .B1(n20189), .B2(n20200), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19237) );
  AOI22_X1 U22381 ( .A1(n20314), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19237), 
        .B2(n20315), .ZN(P2_U2817) );
  INV_X1 U22382 ( .A(n20194), .ZN(n20181) );
  OAI21_X1 U22383 ( .B1(n20181), .B2(BS16), .A(n20256), .ZN(n20254) );
  OAI21_X1 U22384 ( .B1(n20256), .B2(n21288), .A(n20254), .ZN(P2_U2818) );
  NOR4_X1 U22385 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19247) );
  NOR4_X1 U22386 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19246) );
  AOI211_X1 U22387 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_8__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19238) );
  INV_X1 U22388 ( .A(P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21090) );
  INV_X1 U22389 ( .A(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20180) );
  NAND3_X1 U22390 ( .A1(n19238), .A2(n21090), .A3(n20180), .ZN(n19244) );
  NOR4_X1 U22391 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19242) );
  NOR4_X1 U22392 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_14__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n19241) );
  NOR4_X1 U22393 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19240) );
  NOR4_X1 U22394 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19239) );
  NAND4_X1 U22395 ( .A1(n19242), .A2(n19241), .A3(n19240), .A4(n19239), .ZN(
        n19243) );
  NOR4_X1 U22396 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(n19244), .A4(n19243), .ZN(n19245)
         );
  NAND3_X1 U22397 ( .A1(n19247), .A2(n19246), .A3(n19245), .ZN(n19255) );
  NOR2_X1 U22398 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19255), .ZN(n19250) );
  INV_X1 U22399 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19248) );
  AOI22_X1 U22400 ( .A1(n19250), .A2(n19439), .B1(n19255), .B2(n19248), .ZN(
        P2_U2820) );
  OR3_X1 U22401 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19254) );
  INV_X1 U22402 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19249) );
  AOI22_X1 U22403 ( .A1(n19250), .A2(n19254), .B1(n19255), .B2(n19249), .ZN(
        P2_U2821) );
  INV_X1 U22404 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20255) );
  NAND2_X1 U22405 ( .A1(n19250), .A2(n20255), .ZN(n19253) );
  INV_X1 U22406 ( .A(n19255), .ZN(n19257) );
  OAI21_X1 U22407 ( .B1(n19439), .B2(n20202), .A(n19257), .ZN(n19251) );
  OAI21_X1 U22408 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19257), .A(n19251), 
        .ZN(n19252) );
  OAI221_X1 U22409 ( .B1(n19253), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19253), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19252), .ZN(P2_U2822) );
  INV_X1 U22410 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19256) );
  OAI221_X1 U22411 ( .B1(n19257), .B2(n19256), .C1(n19255), .C2(n19254), .A(
        n19253), .ZN(P2_U2823) );
  AOI22_X1 U22412 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19454), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19431), .ZN(n19268) );
  AOI22_X1 U22413 ( .A1(n19258), .A2(n19422), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19444), .ZN(n19267) );
  AOI22_X1 U22414 ( .A1(n19260), .A2(n19449), .B1(n19259), .B2(n19379), .ZN(
        n19266) );
  AOI21_X1 U22415 ( .B1(n19263), .B2(n19262), .A(n19261), .ZN(n19264) );
  NAND2_X1 U22416 ( .A1(n19416), .A2(n19264), .ZN(n19265) );
  NAND4_X1 U22417 ( .A1(n19268), .A2(n19267), .A3(n19266), .A4(n19265), .ZN(
        P2_U2835) );
  AOI211_X1 U22418 ( .C1(n19270), .C2(n9834), .A(n19269), .B(n19450), .ZN(
        n19280) );
  AOI22_X1 U22419 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19444), .ZN(n19271) );
  NAND2_X1 U22420 ( .A1(n19272), .A2(n19271), .ZN(n19273) );
  AOI21_X1 U22421 ( .B1(n19431), .B2(P2_REIP_REG_18__SCAN_IN), .A(n19273), 
        .ZN(n19274) );
  OAI21_X1 U22422 ( .B1(n19275), .B2(n19414), .A(n19274), .ZN(n19276) );
  INV_X1 U22423 ( .A(n19276), .ZN(n19277) );
  OAI21_X1 U22424 ( .B1(n19278), .B2(n19447), .A(n19277), .ZN(n19279) );
  NOR2_X1 U22425 ( .A1(n19280), .A2(n19279), .ZN(n19281) );
  OAI21_X1 U22426 ( .B1(n19282), .B2(n19442), .A(n19281), .ZN(P2_U2837) );
  INV_X1 U22427 ( .A(n19291), .ZN(n19286) );
  OAI22_X1 U22428 ( .A1(n19283), .A2(n19420), .B1(n20226), .B2(n19440), .ZN(
        n19284) );
  AOI211_X1 U22429 ( .C1(n19286), .C2(n19285), .A(n19643), .B(n19284), .ZN(
        n19296) );
  AOI22_X1 U22430 ( .A1(n19287), .A2(n19422), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n19444), .ZN(n19295) );
  INV_X1 U22431 ( .A(n19288), .ZN(n19289) );
  AOI22_X1 U22432 ( .A1(n19290), .A2(n19449), .B1(n19379), .B2(n19289), .ZN(
        n19294) );
  OAI211_X1 U22433 ( .C1(n19292), .C2(n19291), .A(n19416), .B(n9834), .ZN(
        n19293) );
  NAND4_X1 U22434 ( .A1(n19296), .A2(n19295), .A3(n19294), .A4(n19293), .ZN(
        P2_U2838) );
  NAND2_X1 U22435 ( .A1(n10049), .A2(n19297), .ZN(n19298) );
  XOR2_X1 U22436 ( .A(n19299), .B(n19298), .Z(n19306) );
  AOI22_X1 U22437 ( .A1(n19300), .A2(n19422), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19444), .ZN(n19301) );
  OAI21_X1 U22438 ( .B1(n21240), .B2(n19420), .A(n19301), .ZN(n19302) );
  AOI211_X1 U22439 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19431), .A(n19643), 
        .B(n19302), .ZN(n19305) );
  AOI22_X1 U22440 ( .A1(n19462), .A2(n19379), .B1(n19449), .B2(n19303), .ZN(
        n19304) );
  OAI211_X1 U22441 ( .C1(n19450), .C2(n19306), .A(n19305), .B(n19304), .ZN(
        P2_U2839) );
  OAI22_X1 U22442 ( .A1(n19308), .A2(n19447), .B1(n19307), .B2(n19429), .ZN(
        n19309) );
  AOI211_X1 U22443 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19431), .A(n19643), 
        .B(n19309), .ZN(n19317) );
  NOR2_X1 U22444 ( .A1(n19410), .A2(n19310), .ZN(n19311) );
  XOR2_X1 U22445 ( .A(n19312), .B(n19311), .Z(n19315) );
  OAI22_X1 U22446 ( .A1(n19468), .A2(n19442), .B1(n19414), .B2(n19313), .ZN(
        n19314) );
  AOI21_X1 U22447 ( .B1(n19315), .B2(n19416), .A(n19314), .ZN(n19316) );
  OAI211_X1 U22448 ( .C1(n19318), .C2(n19420), .A(n19317), .B(n19316), .ZN(
        P2_U2840) );
  NAND2_X1 U22449 ( .A1(n10049), .A2(n19319), .ZN(n19320) );
  XOR2_X1 U22450 ( .A(n19321), .B(n19320), .Z(n19329) );
  INV_X1 U22451 ( .A(n19322), .ZN(n19324) );
  AOI22_X1 U22452 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19444), .ZN(n19323) );
  OAI21_X1 U22453 ( .B1(n19324), .B2(n19447), .A(n19323), .ZN(n19325) );
  AOI211_X1 U22454 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19431), .A(n19643), 
        .B(n19325), .ZN(n19328) );
  AOI22_X1 U22455 ( .A1(n19469), .A2(n19379), .B1(n19449), .B2(n19326), .ZN(
        n19327) );
  OAI211_X1 U22456 ( .C1(n19450), .C2(n19329), .A(n19328), .B(n19327), .ZN(
        P2_U2841) );
  INV_X1 U22457 ( .A(n19330), .ZN(n19331) );
  OAI22_X1 U22458 ( .A1(n19331), .A2(n19447), .B1(n21151), .B2(n19429), .ZN(
        n19332) );
  AOI211_X1 U22459 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19431), .A(n19643), 
        .B(n19332), .ZN(n19340) );
  NOR2_X1 U22460 ( .A1(n19410), .A2(n19333), .ZN(n19334) );
  XOR2_X1 U22461 ( .A(n19335), .B(n19334), .Z(n19338) );
  OAI22_X1 U22462 ( .A1(n19473), .A2(n19442), .B1(n19414), .B2(n19336), .ZN(
        n19337) );
  AOI21_X1 U22463 ( .B1(n19338), .B2(n19416), .A(n19337), .ZN(n19339) );
  OAI211_X1 U22464 ( .C1(n21272), .C2(n19420), .A(n19340), .B(n19339), .ZN(
        P2_U2842) );
  OAI22_X1 U22465 ( .A1(n19341), .A2(n19447), .B1(n19429), .B2(n21145), .ZN(
        n19342) );
  INV_X1 U22466 ( .A(n19342), .ZN(n19343) );
  OAI211_X1 U22467 ( .C1(n20217), .C2(n19440), .A(n19343), .B(n19272), .ZN(
        n19344) );
  AOI21_X1 U22468 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19454), .A(
        n19344), .ZN(n19350) );
  XOR2_X1 U22469 ( .A(n19346), .B(n19345), .Z(n19348) );
  AOI22_X1 U22470 ( .A1(n19348), .A2(n19416), .B1(n19449), .B2(n19347), .ZN(
        n19349) );
  OAI211_X1 U22471 ( .C1(n19475), .C2(n19442), .A(n19350), .B(n19349), .ZN(
        P2_U2843) );
  INV_X1 U22472 ( .A(n19351), .ZN(n19352) );
  AOI22_X1 U22473 ( .A1(n19352), .A2(n19422), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19444), .ZN(n19353) );
  OAI211_X1 U22474 ( .C1(n20215), .C2(n19440), .A(n19353), .B(n19272), .ZN(
        n19354) );
  AOI21_X1 U22475 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19454), .A(
        n19354), .ZN(n19361) );
  NAND2_X1 U22476 ( .A1(n10049), .A2(n19355), .ZN(n19356) );
  XNOR2_X1 U22477 ( .A(n19357), .B(n19356), .ZN(n19359) );
  AOI22_X1 U22478 ( .A1(n19359), .A2(n19416), .B1(n19449), .B2(n19358), .ZN(
        n19360) );
  OAI211_X1 U22479 ( .C1(n19442), .C2(n19480), .A(n19361), .B(n19360), .ZN(
        P2_U2845) );
  OAI22_X1 U22480 ( .A1(n19362), .A2(n19447), .B1(n19429), .B2(n11454), .ZN(
        n19363) );
  AOI211_X1 U22481 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19431), .A(n19643), .B(
        n19363), .ZN(n19371) );
  NOR2_X1 U22482 ( .A1(n19410), .A2(n19364), .ZN(n19365) );
  XNOR2_X1 U22483 ( .A(n19366), .B(n19365), .ZN(n19369) );
  OAI22_X1 U22484 ( .A1(n19483), .A2(n19442), .B1(n19414), .B2(n19367), .ZN(
        n19368) );
  AOI21_X1 U22485 ( .B1(n19369), .B2(n19416), .A(n19368), .ZN(n19370) );
  OAI211_X1 U22486 ( .C1(n19372), .C2(n19420), .A(n19371), .B(n19370), .ZN(
        P2_U2846) );
  NAND2_X1 U22487 ( .A1(n10049), .A2(n19373), .ZN(n19374) );
  XOR2_X1 U22488 ( .A(n19375), .B(n19374), .Z(n19383) );
  AOI22_X1 U22489 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19454), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19444), .ZN(n19376) );
  OAI21_X1 U22490 ( .B1(n19377), .B2(n19447), .A(n19376), .ZN(n19378) );
  AOI211_X1 U22491 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19431), .A(n19643), .B(
        n19378), .ZN(n19382) );
  AOI22_X1 U22492 ( .A1(n19380), .A2(n19449), .B1(n19379), .B2(n19484), .ZN(
        n19381) );
  OAI211_X1 U22493 ( .C1(n19450), .C2(n19383), .A(n19382), .B(n19381), .ZN(
        P2_U2847) );
  NOR2_X1 U22494 ( .A1(n19410), .A2(n19384), .ZN(n19385) );
  XOR2_X1 U22495 ( .A(n19386), .B(n19385), .Z(n19394) );
  AOI22_X1 U22496 ( .A1(n19387), .A2(n19422), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19444), .ZN(n19389) );
  OAI211_X1 U22497 ( .C1(n20211), .C2(n19440), .A(n19389), .B(n19388), .ZN(
        n19392) );
  OAI22_X1 U22498 ( .A1(n19487), .A2(n19442), .B1(n19414), .B2(n19390), .ZN(
        n19391) );
  AOI211_X1 U22499 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19454), .A(
        n19392), .B(n19391), .ZN(n19393) );
  OAI21_X1 U22500 ( .B1(n19450), .B2(n19394), .A(n19393), .ZN(P2_U2848) );
  OAI21_X1 U22501 ( .B1(n20209), .B2(n19440), .A(n19272), .ZN(n19398) );
  INV_X1 U22502 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19395) );
  OAI22_X1 U22503 ( .A1(n19396), .A2(n19447), .B1(n19429), .B2(n19395), .ZN(
        n19397) );
  AOI211_X1 U22504 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19454), .A(
        n19398), .B(n19397), .ZN(n19405) );
  NAND2_X1 U22505 ( .A1(n10049), .A2(n19399), .ZN(n19400) );
  XNOR2_X1 U22506 ( .A(n19401), .B(n19400), .ZN(n19403) );
  AOI22_X1 U22507 ( .A1(n19403), .A2(n19416), .B1(n19449), .B2(n19402), .ZN(
        n19404) );
  OAI211_X1 U22508 ( .C1(n19442), .C2(n19490), .A(n19405), .B(n19404), .ZN(
        P2_U2849) );
  OAI22_X1 U22509 ( .A1(n19407), .A2(n19447), .B1(n19429), .B2(n19406), .ZN(
        n19408) );
  AOI211_X1 U22510 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19431), .A(n19643), .B(
        n19408), .ZN(n19419) );
  NOR2_X1 U22511 ( .A1(n19410), .A2(n19409), .ZN(n19411) );
  XNOR2_X1 U22512 ( .A(n19412), .B(n19411), .ZN(n19417) );
  OAI22_X1 U22513 ( .A1(n19500), .A2(n19442), .B1(n19414), .B2(n19413), .ZN(
        n19415) );
  AOI21_X1 U22514 ( .B1(n19417), .B2(n19416), .A(n19415), .ZN(n19418) );
  OAI211_X1 U22515 ( .C1(n19421), .C2(n19420), .A(n19419), .B(n19418), .ZN(
        P2_U2850) );
  AOI22_X1 U22516 ( .A1(n19423), .A2(n19422), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19454), .ZN(n19438) );
  NAND2_X1 U22517 ( .A1(n19424), .A2(n14329), .ZN(n19427) );
  INV_X1 U22518 ( .A(n19425), .ZN(n19426) );
  NAND2_X1 U22519 ( .A1(n19427), .A2(n19426), .ZN(n19502) );
  OAI22_X1 U22520 ( .A1(n19429), .A2(n19428), .B1(n19442), .B2(n19502), .ZN(
        n19430) );
  AOI211_X1 U22521 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19431), .A(n19643), .B(
        n19430), .ZN(n19437) );
  INV_X1 U22522 ( .A(n19503), .ZN(n19497) );
  AOI22_X1 U22523 ( .A1(n19497), .A2(n19452), .B1(n19449), .B2(n19648), .ZN(
        n19436) );
  AND2_X1 U22524 ( .A1(n10049), .A2(n19432), .ZN(n19434) );
  AOI21_X1 U22525 ( .B1(n19612), .B2(n19434), .A(n19450), .ZN(n19433) );
  OAI21_X1 U22526 ( .B1(n19612), .B2(n19434), .A(n19433), .ZN(n19435) );
  NAND4_X1 U22527 ( .A1(n19438), .A2(n19437), .A3(n19436), .A4(n19435), .ZN(
        P2_U2851) );
  OAI22_X1 U22528 ( .A1(n19442), .A2(n19441), .B1(n19440), .B2(n19439), .ZN(
        n19443) );
  AOI21_X1 U22529 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19444), .A(n19443), .ZN(
        n19445) );
  OAI21_X1 U22530 ( .B1(n19447), .B2(n19446), .A(n19445), .ZN(n19448) );
  AOI21_X1 U22531 ( .B1(n13096), .B2(n19449), .A(n19448), .ZN(n19457) );
  AOI22_X1 U22532 ( .A1(n19453), .A2(n19452), .B1(n19451), .B2(n19416), .ZN(
        n19456) );
  NAND2_X1 U22533 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19454), .ZN(
        n19455) );
  NAND3_X1 U22534 ( .A1(n19457), .A2(n19456), .A3(n19455), .ZN(P2_U2855) );
  AOI22_X1 U22535 ( .A1(n19459), .A2(n19458), .B1(n19522), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19466) );
  AOI22_X1 U22536 ( .A1(n19461), .A2(BUF1_REG_16__SCAN_IN), .B1(n19460), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19465) );
  AOI22_X1 U22537 ( .A1(n19463), .A2(n19505), .B1(n19462), .B2(n19523), .ZN(
        n19464) );
  NAND3_X1 U22538 ( .A1(n19466), .A2(n19465), .A3(n19464), .ZN(P2_U2903) );
  OAI222_X1 U22539 ( .A1(n19468), .A2(n19501), .B1(n13701), .B2(n19489), .C1(
        n19467), .C2(n19531), .ZN(P2_U2904) );
  INV_X1 U22540 ( .A(n19469), .ZN(n19471) );
  AOI22_X1 U22541 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19522), .B1(n19605), 
        .B2(n19491), .ZN(n19470) );
  OAI21_X1 U22542 ( .B1(n19501), .B2(n19471), .A(n19470), .ZN(P2_U2905) );
  INV_X1 U22543 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19575) );
  OAI222_X1 U22544 ( .A1(n19473), .A2(n19501), .B1(n19575), .B2(n19489), .C1(
        n19531), .C2(n19472), .ZN(P2_U2906) );
  INV_X1 U22545 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19577) );
  OAI222_X1 U22546 ( .A1(n19475), .A2(n19501), .B1(n19577), .B2(n19489), .C1(
        n19531), .C2(n19474), .ZN(P2_U2907) );
  INV_X1 U22547 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n21294) );
  OAI222_X1 U22548 ( .A1(n19477), .A2(n19501), .B1(n21294), .B2(n19489), .C1(
        n19531), .C2(n19476), .ZN(P2_U2908) );
  AOI22_X1 U22549 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19522), .B1(n19478), 
        .B2(n19491), .ZN(n19479) );
  OAI21_X1 U22550 ( .B1(n19501), .B2(n19480), .A(n19479), .ZN(P2_U2909) );
  AOI22_X1 U22551 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19522), .B1(n19481), .B2(
        n19491), .ZN(n19482) );
  OAI21_X1 U22552 ( .B1(n19501), .B2(n19483), .A(n19482), .ZN(P2_U2910) );
  INV_X1 U22553 ( .A(n19484), .ZN(n19486) );
  INV_X1 U22554 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19584) );
  OAI222_X1 U22555 ( .A1(n19486), .A2(n19501), .B1(n19584), .B2(n19489), .C1(
        n19531), .C2(n19485), .ZN(P2_U2911) );
  INV_X1 U22556 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19586) );
  OAI222_X1 U22557 ( .A1(n19487), .A2(n19501), .B1(n19586), .B2(n19489), .C1(
        n19531), .C2(n19698), .ZN(P2_U2912) );
  INV_X1 U22558 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19589) );
  OAI222_X1 U22559 ( .A1(n19490), .A2(n19501), .B1(n19589), .B2(n19489), .C1(
        n19531), .C2(n19488), .ZN(P2_U2913) );
  AOI22_X1 U22560 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19522), .B1(n19492), .B2(
        n19491), .ZN(n19499) );
  INV_X1 U22561 ( .A(n20286), .ZN(n19493) );
  XNOR2_X1 U22562 ( .A(n20284), .B(n20286), .ZN(n19525) );
  NOR2_X1 U22563 ( .A1(n19525), .A2(n19526), .ZN(n19524) );
  AOI21_X1 U22564 ( .B1(n20281), .B2(n19493), .A(n19524), .ZN(n19517) );
  XNOR2_X1 U22565 ( .A(n20271), .B(n19668), .ZN(n19518) );
  NOR2_X1 U22566 ( .A1(n19517), .A2(n19518), .ZN(n19516) );
  AOI21_X1 U22567 ( .B1(n19668), .B2(n20271), .A(n19516), .ZN(n19512) );
  XNOR2_X1 U22568 ( .A(n20264), .B(n19494), .ZN(n19511) );
  NOR2_X1 U22569 ( .A1(n19512), .A2(n19511), .ZN(n19510) );
  INV_X1 U22570 ( .A(n19494), .ZN(n20268) );
  NOR2_X1 U22571 ( .A1(n19495), .A2(n20268), .ZN(n19496) );
  OAI21_X1 U22572 ( .B1(n19510), .B2(n19496), .A(n19502), .ZN(n19504) );
  NAND3_X1 U22573 ( .A1(n19504), .A2(n19497), .A3(n19505), .ZN(n19498) );
  OAI211_X1 U22574 ( .C1(n19501), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P2_U2914) );
  INV_X1 U22575 ( .A(n19502), .ZN(n19644) );
  AOI22_X1 U22576 ( .A1(n19523), .A2(n19644), .B1(n19522), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19508) );
  XNOR2_X1 U22577 ( .A(n19504), .B(n19503), .ZN(n19506) );
  NAND2_X1 U22578 ( .A1(n19506), .A2(n19505), .ZN(n19507) );
  OAI211_X1 U22579 ( .C1(n19509), .C2(n19531), .A(n19508), .B(n19507), .ZN(
        P2_U2915) );
  AOI22_X1 U22580 ( .A1(n20268), .A2(n19523), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19522), .ZN(n19515) );
  AOI21_X1 U22581 ( .B1(n19512), .B2(n19511), .A(n19510), .ZN(n19513) );
  OR2_X1 U22582 ( .A1(n19513), .A2(n19527), .ZN(n19514) );
  OAI211_X1 U22583 ( .C1(n19687), .C2(n19531), .A(n19515), .B(n19514), .ZN(
        P2_U2916) );
  INV_X1 U22584 ( .A(n19668), .ZN(n20272) );
  AOI22_X1 U22585 ( .A1(n20272), .A2(n19523), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19522), .ZN(n19521) );
  AOI21_X1 U22586 ( .B1(n19518), .B2(n19517), .A(n19516), .ZN(n19519) );
  OR2_X1 U22587 ( .A1(n19519), .A2(n19527), .ZN(n19520) );
  OAI211_X1 U22588 ( .C1(n19683), .C2(n19531), .A(n19521), .B(n19520), .ZN(
        P2_U2917) );
  AOI22_X1 U22589 ( .A1(n19523), .A2(n20286), .B1(n19522), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19530) );
  AOI21_X1 U22590 ( .B1(n19526), .B2(n19525), .A(n19524), .ZN(n19528) );
  OR2_X1 U22591 ( .A1(n19528), .A2(n19527), .ZN(n19529) );
  OAI211_X1 U22592 ( .C1(n19532), .C2(n19531), .A(n19530), .B(n19529), .ZN(
        P2_U2918) );
  OR2_X1 U22593 ( .A1(n10951), .A2(n19533), .ZN(n19535) );
  OAI21_X1 U22594 ( .B1(n19536), .B2(n19535), .A(n19534), .ZN(n19537) );
  NOR2_X1 U22595 ( .A1(n19558), .A2(n19538), .ZN(P2_U2920) );
  NOR2_X1 U22596 ( .A1(n19602), .A2(n19539), .ZN(n19556) );
  INV_X2 U22597 ( .A(n19540), .ZN(n19598) );
  AOI22_X1 U22598 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19556), .B1(n19598), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19541) );
  OAI21_X1 U22599 ( .B1(n19558), .B2(n19542), .A(n19541), .ZN(P2_U2921) );
  INV_X2 U22600 ( .A(n19558), .ZN(n19587) );
  AOI22_X1 U22601 ( .A1(n19598), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19543) );
  OAI21_X1 U22602 ( .B1(n19544), .B2(n19569), .A(n19543), .ZN(P2_U2922) );
  AOI22_X1 U22603 ( .A1(n19598), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19545) );
  OAI21_X1 U22604 ( .B1(n19546), .B2(n19569), .A(n19545), .ZN(P2_U2923) );
  AOI22_X1 U22605 ( .A1(n19598), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19547) );
  OAI21_X1 U22606 ( .B1(n19548), .B2(n19569), .A(n19547), .ZN(P2_U2924) );
  AOI22_X1 U22607 ( .A1(n19598), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19549) );
  OAI21_X1 U22608 ( .B1(n21071), .B2(n19569), .A(n19549), .ZN(P2_U2925) );
  AOI22_X1 U22609 ( .A1(n19598), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19550) );
  OAI21_X1 U22610 ( .B1(n19551), .B2(n19569), .A(n19550), .ZN(P2_U2926) );
  AOI22_X1 U22611 ( .A1(n19598), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19552) );
  OAI21_X1 U22612 ( .B1(n19553), .B2(n19569), .A(n19552), .ZN(P2_U2927) );
  AOI22_X1 U22613 ( .A1(n19598), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19554) );
  OAI21_X1 U22614 ( .B1(n19555), .B2(n19569), .A(n19554), .ZN(P2_U2928) );
  AOI22_X1 U22615 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n19556), .B1(n19598), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n19557) );
  OAI21_X1 U22616 ( .B1(n21122), .B2(n19558), .A(n19557), .ZN(P2_U2929) );
  INV_X1 U22617 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n21168) );
  AOI22_X1 U22618 ( .A1(n19598), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19559) );
  OAI21_X1 U22619 ( .B1(n21168), .B2(n19569), .A(n19559), .ZN(P2_U2930) );
  INV_X1 U22620 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19561) );
  AOI22_X1 U22621 ( .A1(n19598), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19560) );
  OAI21_X1 U22622 ( .B1(n19561), .B2(n19569), .A(n19560), .ZN(P2_U2931) );
  INV_X1 U22623 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19563) );
  AOI22_X1 U22624 ( .A1(n19598), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19562) );
  OAI21_X1 U22625 ( .B1(n19563), .B2(n19569), .A(n19562), .ZN(P2_U2932) );
  INV_X1 U22626 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19565) );
  AOI22_X1 U22627 ( .A1(n19598), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19564) );
  OAI21_X1 U22628 ( .B1(n19565), .B2(n19569), .A(n19564), .ZN(P2_U2933) );
  INV_X1 U22629 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19567) );
  AOI22_X1 U22630 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n19598), .B1(n19587), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19566) );
  OAI21_X1 U22631 ( .B1(n19567), .B2(n19569), .A(n19566), .ZN(P2_U2934) );
  INV_X1 U22632 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19570) );
  AOI22_X1 U22633 ( .A1(n19598), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19568) );
  OAI21_X1 U22634 ( .B1(n19570), .B2(n19569), .A(n19568), .ZN(P2_U2935) );
  AOI22_X1 U22635 ( .A1(n19598), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19571) );
  OAI21_X1 U22636 ( .B1(n13701), .B2(n19602), .A(n19571), .ZN(P2_U2936) );
  INV_X1 U22637 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U22638 ( .A1(n19598), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19572) );
  OAI21_X1 U22639 ( .B1(n19573), .B2(n19602), .A(n19572), .ZN(P2_U2937) );
  AOI22_X1 U22640 ( .A1(n19598), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19574) );
  OAI21_X1 U22641 ( .B1(n19575), .B2(n19602), .A(n19574), .ZN(P2_U2938) );
  AOI22_X1 U22642 ( .A1(n19598), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19576) );
  OAI21_X1 U22643 ( .B1(n19577), .B2(n19602), .A(n19576), .ZN(P2_U2939) );
  AOI22_X1 U22644 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n19587), .B1(n19598), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19578) );
  OAI21_X1 U22645 ( .B1(n21294), .B2(n19602), .A(n19578), .ZN(P2_U2940) );
  AOI22_X1 U22646 ( .A1(P2_LWORD_REG_10__SCAN_IN), .A2(n19598), .B1(n19587), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19579) );
  OAI21_X1 U22647 ( .B1(n19580), .B2(n19602), .A(n19579), .ZN(P2_U2941) );
  AOI22_X1 U22648 ( .A1(n19598), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19581) );
  OAI21_X1 U22649 ( .B1(n19582), .B2(n19602), .A(n19581), .ZN(P2_U2942) );
  AOI22_X1 U22650 ( .A1(n19598), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19583) );
  OAI21_X1 U22651 ( .B1(n19584), .B2(n19602), .A(n19583), .ZN(P2_U2943) );
  AOI22_X1 U22652 ( .A1(n19598), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19585) );
  OAI21_X1 U22653 ( .B1(n19586), .B2(n19602), .A(n19585), .ZN(P2_U2944) );
  AOI22_X1 U22654 ( .A1(n19598), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19588) );
  OAI21_X1 U22655 ( .B1(n19589), .B2(n19602), .A(n19588), .ZN(P2_U2945) );
  INV_X1 U22656 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19591) );
  AOI22_X1 U22657 ( .A1(n19598), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19590) );
  OAI21_X1 U22658 ( .B1(n19591), .B2(n19602), .A(n19590), .ZN(P2_U2946) );
  INV_X1 U22659 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19593) );
  AOI22_X1 U22660 ( .A1(n19598), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19592) );
  OAI21_X1 U22661 ( .B1(n19593), .B2(n19602), .A(n19592), .ZN(P2_U2947) );
  INV_X1 U22662 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19595) );
  AOI22_X1 U22663 ( .A1(n19598), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19594) );
  OAI21_X1 U22664 ( .B1(n19595), .B2(n19602), .A(n19594), .ZN(P2_U2948) );
  INV_X1 U22665 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19597) );
  AOI22_X1 U22666 ( .A1(n19598), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19596) );
  OAI21_X1 U22667 ( .B1(n19597), .B2(n19602), .A(n19596), .ZN(P2_U2949) );
  INV_X1 U22668 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19600) );
  AOI22_X1 U22669 ( .A1(n19598), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19587), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19599) );
  OAI21_X1 U22670 ( .B1(n19600), .B2(n19602), .A(n19599), .ZN(P2_U2950) );
  INV_X1 U22671 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19603) );
  AOI22_X1 U22672 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n19587), .B1(n19598), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n19601) );
  OAI21_X1 U22673 ( .B1(n19603), .B2(n19602), .A(n19601), .ZN(P2_U2951) );
  AOI22_X1 U22674 ( .A1(n19609), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19604), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19607) );
  NAND2_X1 U22675 ( .A1(n19606), .A2(n19605), .ZN(n19610) );
  NAND2_X1 U22676 ( .A1(n19607), .A2(n19610), .ZN(P2_U2966) );
  AOI22_X1 U22677 ( .A1(n19609), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19608), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19611) );
  NAND2_X1 U22678 ( .A1(n19611), .A2(n19610), .ZN(P2_U2981) );
  AOI22_X1 U22679 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19643), .B1(n19613), 
        .B2(n19612), .ZN(n19624) );
  XOR2_X1 U22680 ( .A(n19614), .B(n19615), .Z(n19653) );
  INV_X1 U22681 ( .A(n19653), .ZN(n19620) );
  XNOR2_X1 U22682 ( .A(n19616), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19617) );
  XNOR2_X1 U22683 ( .A(n19618), .B(n19617), .ZN(n19651) );
  OAI22_X1 U22684 ( .A1(n19620), .A2(n19619), .B1(n19651), .B2(n19636), .ZN(
        n19621) );
  AOI21_X1 U22685 ( .B1(n19622), .B2(n19648), .A(n19621), .ZN(n19623) );
  OAI211_X1 U22686 ( .C1(n19625), .C2(n19642), .A(n19624), .B(n19623), .ZN(
        P2_U3010) );
  INV_X1 U22687 ( .A(n19626), .ZN(n19627) );
  XNOR2_X1 U22688 ( .A(n19628), .B(n19627), .ZN(n19664) );
  NOR2_X1 U22689 ( .A1(n19629), .A2(n14135), .ZN(n19639) );
  AOI21_X1 U22690 ( .B1(n19632), .B2(n19631), .A(n19630), .ZN(n19659) );
  INV_X1 U22691 ( .A(n19659), .ZN(n19637) );
  INV_X1 U22692 ( .A(n19633), .ZN(n19635) );
  OAI22_X1 U22693 ( .A1(n19637), .A2(n19636), .B1(n19635), .B2(n19634), .ZN(
        n19638) );
  AOI211_X1 U22694 ( .C1(n19664), .C2(n12997), .A(n19639), .B(n19638), .ZN(
        n19640) );
  NAND2_X1 U22695 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19643), .ZN(n19661) );
  OAI211_X1 U22696 ( .C1(n19642), .C2(n19641), .A(n19640), .B(n19661), .ZN(
        P2_U3012) );
  AOI22_X1 U22697 ( .A1(n19645), .A2(n19644), .B1(n19643), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n19655) );
  NOR2_X1 U22698 ( .A1(n10787), .A2(n19646), .ZN(n19647) );
  AOI21_X1 U22699 ( .B1(n19648), .B2(n19669), .A(n19647), .ZN(n19649) );
  OAI21_X1 U22700 ( .B1(n19651), .B2(n19650), .A(n19649), .ZN(n19652) );
  AOI21_X1 U22701 ( .B1(n19653), .B2(n19663), .A(n19652), .ZN(n19654) );
  OAI211_X1 U22702 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n19656), .A(
        n19655), .B(n19654), .ZN(P2_U3042) );
  AOI22_X1 U22703 ( .A1(n19660), .A2(n19659), .B1(n19658), .B2(n19657), .ZN(
        n19676) );
  AND2_X1 U22704 ( .A1(n19662), .A2(n19661), .ZN(n19666) );
  NAND2_X1 U22705 ( .A1(n19664), .A2(n19663), .ZN(n19665) );
  OAI211_X1 U22706 ( .C1(n19668), .C2(n19667), .A(n19666), .B(n19665), .ZN(
        n19674) );
  AND2_X1 U22707 ( .A1(n19669), .A2(n9750), .ZN(n19673) );
  NOR2_X1 U22708 ( .A1(n19671), .A2(n19670), .ZN(n19672) );
  NOR3_X1 U22709 ( .A1(n19674), .A2(n19673), .A3(n19672), .ZN(n19675) );
  OAI211_X1 U22710 ( .C1(n19677), .C2(n10577), .A(n19676), .B(n19675), .ZN(
        P2_U3044) );
  INV_X1 U22711 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19681) );
  INV_X1 U22712 ( .A(n19678), .ZN(n20119) );
  AOI22_X1 U22713 ( .A1(n20080), .A2(n20173), .B1(n19697), .B2(n20119), .ZN(
        n19680) );
  AOI22_X1 U22714 ( .A1(n14145), .A2(n19703), .B1(n19731), .B2(n20127), .ZN(
        n19679) );
  OAI211_X1 U22715 ( .C1(n19707), .C2(n19681), .A(n19680), .B(n19679), .ZN(
        P2_U3048) );
  AOI22_X1 U22716 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19693), .ZN(n20141) );
  AOI22_X1 U22717 ( .A1(n20092), .A2(n20173), .B1(n19697), .B2(n20136), .ZN(
        n19685) );
  NOR2_X2 U22718 ( .A1(n19683), .A2(n19874), .ZN(n20137) );
  AOI22_X1 U22719 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19693), .ZN(n20055) );
  AOI22_X1 U22720 ( .A1(n20137), .A2(n19703), .B1(n19731), .B2(n20138), .ZN(
        n19684) );
  OAI211_X1 U22721 ( .C1(n19707), .C2(n13108), .A(n19685), .B(n19684), .ZN(
        P2_U3050) );
  AOI22_X1 U22722 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19693), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19694), .ZN(n20147) );
  AOI22_X1 U22723 ( .A1(n20095), .A2(n20173), .B1(n19697), .B2(n20142), .ZN(
        n19689) );
  NOR2_X2 U22724 ( .A1(n19687), .A2(n19874), .ZN(n20143) );
  AOI22_X1 U22725 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19693), .ZN(n20025) );
  INV_X1 U22726 ( .A(n20025), .ZN(n20144) );
  AOI22_X1 U22727 ( .A1(n20143), .A2(n19703), .B1(n19731), .B2(n20144), .ZN(
        n19688) );
  OAI211_X1 U22728 ( .C1(n19707), .C2(n13093), .A(n19689), .B(n19688), .ZN(
        P2_U3051) );
  AOI22_X1 U22729 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19693), .ZN(n20159) );
  INV_X1 U22730 ( .A(n20159), .ZN(n20102) );
  NOR2_X2 U22731 ( .A1(n11455), .A2(n19695), .ZN(n20154) );
  AOI22_X1 U22732 ( .A1(n20102), .A2(n20173), .B1(n19697), .B2(n20154), .ZN(
        n19692) );
  NOR2_X2 U22733 ( .A1(n19690), .A2(n19874), .ZN(n20155) );
  AOI22_X1 U22734 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19693), .ZN(n19973) );
  AOI22_X1 U22735 ( .A1(n20155), .A2(n19703), .B1(n19731), .B2(n20156), .ZN(
        n19691) );
  OAI211_X1 U22736 ( .C1(n19707), .C2(n13908), .A(n19692), .B(n19691), .ZN(
        P2_U3053) );
  AOI22_X2 U22737 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19694), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19693), .ZN(n20178) );
  INV_X1 U22738 ( .A(n20178), .ZN(n20110) );
  NOR2_X2 U22739 ( .A1(n19696), .A2(n19695), .ZN(n20168) );
  AOI22_X1 U22740 ( .A1(n20110), .A2(n20173), .B1(n19697), .B2(n20168), .ZN(
        n19705) );
  NOR2_X2 U22741 ( .A1(n19698), .A2(n19874), .ZN(n20170) );
  OAI22_X2 U22742 ( .A1(n19702), .A2(n19701), .B1(n19700), .B2(n19699), .ZN(
        n20172) );
  AOI22_X1 U22743 ( .A1(n20170), .A2(n19703), .B1(n19731), .B2(n20172), .ZN(
        n19704) );
  OAI211_X1 U22744 ( .C1(n19707), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P2_U3055) );
  INV_X1 U22745 ( .A(n19931), .ZN(n19708) );
  INV_X1 U22746 ( .A(n10797), .ZN(n19709) );
  NOR2_X1 U22747 ( .A1(n20039), .A2(n19771), .ZN(n19734) );
  NOR3_X1 U22748 ( .A1(n19709), .A2(n19734), .A3(n13514), .ZN(n19712) );
  INV_X1 U22749 ( .A(n19713), .ZN(n19710) );
  AOI21_X1 U22750 ( .B1(n19936), .B2(n19710), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19711) );
  NOR2_X1 U22751 ( .A1(n19712), .A2(n19711), .ZN(n19735) );
  AOI22_X1 U22752 ( .A1(n19735), .A2(n14145), .B1(n20119), .B2(n19734), .ZN(
        n19717) );
  INV_X1 U22753 ( .A(n20258), .ZN(n19873) );
  NAND2_X1 U22754 ( .A1(n19873), .A2(n19931), .ZN(n19714) );
  AOI21_X1 U22755 ( .B1(n19714), .B2(n19713), .A(n19712), .ZN(n19715) );
  OAI211_X1 U22756 ( .C1(n19734), .C2(n19936), .A(n19715), .B(n20125), .ZN(
        n19736) );
  AOI22_X1 U22757 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20080), .ZN(n19716) );
  OAI211_X1 U22758 ( .C1(n19881), .C2(n19770), .A(n19717), .B(n19716), .ZN(
        P2_U3056) );
  INV_X1 U22759 ( .A(n19718), .ZN(n20131) );
  AOI22_X1 U22760 ( .A1(n19735), .A2(n14194), .B1(n20131), .B2(n19734), .ZN(
        n19720) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20132), .ZN(n19719) );
  OAI211_X1 U22762 ( .C1(n20135), .C2(n19770), .A(n19720), .B(n19719), .ZN(
        P2_U3057) );
  AOI22_X1 U22763 ( .A1(n19735), .A2(n20137), .B1(n20136), .B2(n19734), .ZN(
        n19722) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20092), .ZN(n19721) );
  OAI211_X1 U22765 ( .C1(n20055), .C2(n19770), .A(n19722), .B(n19721), .ZN(
        P2_U3058) );
  AOI22_X1 U22766 ( .A1(n19735), .A2(n20143), .B1(n20142), .B2(n19734), .ZN(
        n19724) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20095), .ZN(n19723) );
  OAI211_X1 U22768 ( .C1(n20025), .C2(n19770), .A(n19724), .B(n19723), .ZN(
        P2_U3059) );
  AOI22_X1 U22769 ( .A1(n19735), .A2(n20149), .B1(n20148), .B2(n19734), .ZN(
        n19727) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20098), .ZN(n19726) );
  OAI211_X1 U22771 ( .C1(n19951), .C2(n19770), .A(n19727), .B(n19726), .ZN(
        P2_U3060) );
  AOI22_X1 U22772 ( .A1(n19735), .A2(n20155), .B1(n20154), .B2(n19734), .ZN(
        n19729) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20102), .ZN(n19728) );
  OAI211_X1 U22774 ( .C1(n19973), .C2(n19770), .A(n19729), .B(n19728), .ZN(
        P2_U3061) );
  AOI22_X1 U22775 ( .A1(n19735), .A2(n20161), .B1(n20160), .B2(n19734), .ZN(
        n19733) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19736), .B1(
        n19731), .B2(n20162), .ZN(n19732) );
  OAI211_X1 U22777 ( .C1(n20167), .C2(n19770), .A(n19733), .B(n19732), .ZN(
        P2_U3062) );
  AOI22_X1 U22778 ( .A1(n19735), .A2(n20170), .B1(n20168), .B2(n19734), .ZN(
        n19738) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19736), .B1(
        n19762), .B2(n20172), .ZN(n19737) );
  OAI211_X1 U22780 ( .C1(n20178), .C2(n19739), .A(n19738), .B(n19737), .ZN(
        P2_U3063) );
  NOR2_X1 U22781 ( .A1(n20077), .A2(n19771), .ZN(n19765) );
  OAI21_X1 U22782 ( .B1(n19740), .B2(n19765), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19743) );
  INV_X1 U22783 ( .A(n19771), .ZN(n19741) );
  NAND2_X1 U22784 ( .A1(n19742), .A2(n19741), .ZN(n19746) );
  NAND2_X1 U22785 ( .A1(n19743), .A2(n19746), .ZN(n19766) );
  AOI22_X1 U22786 ( .A1(n19766), .A2(n14145), .B1(n20119), .B2(n19765), .ZN(
        n19751) );
  AOI21_X1 U22787 ( .B1(n10801), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19749) );
  OAI21_X1 U22788 ( .B1(n19792), .B2(n19762), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19747) );
  NAND3_X1 U22789 ( .A1(n19747), .A2(n20259), .A3(n19746), .ZN(n19748) );
  OAI211_X1 U22790 ( .C1(n19765), .C2(n19749), .A(n19748), .B(n20125), .ZN(
        n19767) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19767), .B1(
        n19792), .B2(n20127), .ZN(n19750) );
  OAI211_X1 U22792 ( .C1(n20130), .C2(n19770), .A(n19751), .B(n19750), .ZN(
        P2_U3064) );
  AOI22_X1 U22793 ( .A1(n19766), .A2(n14194), .B1(n20131), .B2(n19765), .ZN(
        n19753) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19767), .B1(
        n19762), .B2(n20132), .ZN(n19752) );
  OAI211_X1 U22795 ( .C1(n20135), .C2(n19800), .A(n19753), .B(n19752), .ZN(
        P2_U3065) );
  AOI22_X1 U22796 ( .A1(n19766), .A2(n20137), .B1(n20136), .B2(n19765), .ZN(
        n19755) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19767), .B1(
        n19792), .B2(n20138), .ZN(n19754) );
  OAI211_X1 U22798 ( .C1(n20141), .C2(n19770), .A(n19755), .B(n19754), .ZN(
        P2_U3066) );
  AOI22_X1 U22799 ( .A1(n19766), .A2(n20143), .B1(n20142), .B2(n19765), .ZN(
        n19757) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19767), .B1(
        n19762), .B2(n20095), .ZN(n19756) );
  OAI211_X1 U22801 ( .C1(n20025), .C2(n19800), .A(n19757), .B(n19756), .ZN(
        P2_U3067) );
  AOI22_X1 U22802 ( .A1(n19766), .A2(n20149), .B1(n20148), .B2(n19765), .ZN(
        n19759) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19767), .B1(
        n19792), .B2(n20150), .ZN(n19758) );
  OAI211_X1 U22804 ( .C1(n20153), .C2(n19770), .A(n19759), .B(n19758), .ZN(
        P2_U3068) );
  AOI22_X1 U22805 ( .A1(n19766), .A2(n20155), .B1(n20154), .B2(n19765), .ZN(
        n19761) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19767), .B1(
        n19762), .B2(n20102), .ZN(n19760) );
  OAI211_X1 U22807 ( .C1(n19973), .C2(n19800), .A(n19761), .B(n19760), .ZN(
        P2_U3069) );
  AOI22_X1 U22808 ( .A1(n19766), .A2(n20161), .B1(n20160), .B2(n19765), .ZN(
        n19764) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19767), .B1(
        n19762), .B2(n20162), .ZN(n19763) );
  OAI211_X1 U22810 ( .C1(n20167), .C2(n19800), .A(n19764), .B(n19763), .ZN(
        P2_U3070) );
  AOI22_X1 U22811 ( .A1(n19766), .A2(n20170), .B1(n20168), .B2(n19765), .ZN(
        n19769) );
  AOI22_X1 U22812 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19767), .B1(
        n19792), .B2(n20172), .ZN(n19768) );
  OAI211_X1 U22813 ( .C1(n20178), .C2(n19770), .A(n19769), .B(n19768), .ZN(
        P2_U3071) );
  INV_X1 U22814 ( .A(n19801), .ZN(n19817) );
  NOR2_X1 U22815 ( .A1(n19870), .A2(n19771), .ZN(n19795) );
  AOI22_X1 U22816 ( .A1(n20080), .A2(n19792), .B1(n20119), .B2(n19795), .ZN(
        n19781) );
  OAI21_X1 U22817 ( .B1(n20258), .B2(n20260), .A(n20259), .ZN(n19779) );
  NOR2_X1 U22818 ( .A1(n20288), .A2(n19771), .ZN(n19775) );
  INV_X1 U22819 ( .A(n19795), .ZN(n19772) );
  OAI211_X1 U22820 ( .C1(n19773), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19772), 
        .B(n20261), .ZN(n19774) );
  OAI211_X1 U22821 ( .C1(n19779), .C2(n19775), .A(n20125), .B(n19774), .ZN(
        n19797) );
  INV_X1 U22822 ( .A(n19775), .ZN(n19778) );
  OAI21_X1 U22823 ( .B1(n19776), .B2(n19795), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19777) );
  OAI21_X1 U22824 ( .B1(n19779), .B2(n19778), .A(n19777), .ZN(n19796) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19797), .B1(
        n14145), .B2(n19796), .ZN(n19780) );
  OAI211_X1 U22826 ( .C1(n19881), .C2(n19817), .A(n19781), .B(n19780), .ZN(
        P2_U3072) );
  AOI22_X1 U22827 ( .A1(n20132), .A2(n19792), .B1(n20131), .B2(n19795), .ZN(
        n19783) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19797), .B1(
        n14194), .B2(n19796), .ZN(n19782) );
  OAI211_X1 U22829 ( .C1(n20135), .C2(n19817), .A(n19783), .B(n19782), .ZN(
        P2_U3073) );
  AOI22_X1 U22830 ( .A1(n20092), .A2(n19792), .B1(n19795), .B2(n20136), .ZN(
        n19785) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19797), .B1(
        n20137), .B2(n19796), .ZN(n19784) );
  OAI211_X1 U22832 ( .C1(n20055), .C2(n19817), .A(n19785), .B(n19784), .ZN(
        P2_U3074) );
  AOI22_X1 U22833 ( .A1(n20144), .A2(n19801), .B1(n19795), .B2(n20142), .ZN(
        n19787) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19797), .B1(
        n20143), .B2(n19796), .ZN(n19786) );
  OAI211_X1 U22835 ( .C1(n20147), .C2(n19800), .A(n19787), .B(n19786), .ZN(
        P2_U3075) );
  AOI22_X1 U22836 ( .A1(n20098), .A2(n19792), .B1(n20148), .B2(n19795), .ZN(
        n19789) );
  AOI22_X1 U22837 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19797), .B1(
        n20149), .B2(n19796), .ZN(n19788) );
  OAI211_X1 U22838 ( .C1(n19951), .C2(n19817), .A(n19789), .B(n19788), .ZN(
        P2_U3076) );
  AOI22_X1 U22839 ( .A1(n20156), .A2(n19801), .B1(n19795), .B2(n20154), .ZN(
        n19791) );
  AOI22_X1 U22840 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19797), .B1(
        n20155), .B2(n19796), .ZN(n19790) );
  OAI211_X1 U22841 ( .C1(n20159), .C2(n19800), .A(n19791), .B(n19790), .ZN(
        P2_U3077) );
  AOI22_X1 U22842 ( .A1(n20162), .A2(n19792), .B1(n20160), .B2(n19795), .ZN(
        n19794) );
  AOI22_X1 U22843 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19797), .B1(
        n20161), .B2(n19796), .ZN(n19793) );
  OAI211_X1 U22844 ( .C1(n20167), .C2(n19817), .A(n19794), .B(n19793), .ZN(
        P2_U3078) );
  AOI22_X1 U22845 ( .A1(n20172), .A2(n19801), .B1(n19795), .B2(n20168), .ZN(
        n19799) );
  AOI22_X1 U22846 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19797), .B1(
        n20170), .B2(n19796), .ZN(n19798) );
  OAI211_X1 U22847 ( .C1(n20178), .C2(n19800), .A(n19799), .B(n19798), .ZN(
        P2_U3079) );
  AOI22_X1 U22848 ( .A1(n19813), .A2(n20137), .B1(n20136), .B2(n19812), .ZN(
        n19803) );
  AOI22_X1 U22849 ( .A1(n19830), .A2(n20138), .B1(n19801), .B2(n20092), .ZN(
        n19802) );
  OAI211_X1 U22850 ( .C1(n19805), .C2(n19804), .A(n19803), .B(n19802), .ZN(
        P2_U3082) );
  AOI22_X1 U22851 ( .A1(n19813), .A2(n20143), .B1(n20142), .B2(n19812), .ZN(
        n19807) );
  AOI22_X1 U22852 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19814), .B1(
        n19830), .B2(n20144), .ZN(n19806) );
  OAI211_X1 U22853 ( .C1(n20147), .C2(n19817), .A(n19807), .B(n19806), .ZN(
        P2_U3083) );
  AOI22_X1 U22854 ( .A1(n19813), .A2(n20149), .B1(n20148), .B2(n19812), .ZN(
        n19809) );
  AOI22_X1 U22855 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19814), .B1(
        n19830), .B2(n20150), .ZN(n19808) );
  OAI211_X1 U22856 ( .C1(n20153), .C2(n19817), .A(n19809), .B(n19808), .ZN(
        P2_U3084) );
  AOI22_X1 U22857 ( .A1(n19813), .A2(n20155), .B1(n20154), .B2(n19812), .ZN(
        n19811) );
  AOI22_X1 U22858 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19814), .B1(
        n19830), .B2(n20156), .ZN(n19810) );
  OAI211_X1 U22859 ( .C1(n20159), .C2(n19817), .A(n19811), .B(n19810), .ZN(
        P2_U3085) );
  AOI22_X1 U22860 ( .A1(n19813), .A2(n20170), .B1(n20168), .B2(n19812), .ZN(
        n19816) );
  AOI22_X1 U22861 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19814), .B1(
        n19830), .B2(n20172), .ZN(n19815) );
  OAI211_X1 U22862 ( .C1(n20178), .C2(n19817), .A(n19816), .B(n19815), .ZN(
        P2_U3087) );
  AOI22_X1 U22863 ( .A1(n20132), .A2(n19830), .B1(n20131), .B2(n19839), .ZN(
        n19819) );
  AOI22_X1 U22864 ( .A1(n14194), .A2(n19831), .B1(n19857), .B2(n20089), .ZN(
        n19818) );
  OAI211_X1 U22865 ( .C1(n19834), .C2(n10676), .A(n19819), .B(n19818), .ZN(
        P2_U3089) );
  AOI22_X1 U22866 ( .A1(n20138), .A2(n19857), .B1(n19839), .B2(n20136), .ZN(
        n19821) );
  AOI22_X1 U22867 ( .A1(n20137), .A2(n19831), .B1(n19830), .B2(n20092), .ZN(
        n19820) );
  OAI211_X1 U22868 ( .C1(n19834), .C2(n10696), .A(n19821), .B(n19820), .ZN(
        P2_U3090) );
  AOI22_X1 U22869 ( .A1(n20144), .A2(n19857), .B1(n19839), .B2(n20142), .ZN(
        n19823) );
  AOI22_X1 U22870 ( .A1(n20143), .A2(n19831), .B1(n19830), .B2(n20095), .ZN(
        n19822) );
  OAI211_X1 U22871 ( .C1(n19834), .C2(n10730), .A(n19823), .B(n19822), .ZN(
        P2_U3091) );
  AOI22_X1 U22872 ( .A1(n20098), .A2(n19830), .B1(n20148), .B2(n19839), .ZN(
        n19825) );
  AOI22_X1 U22873 ( .A1(n20149), .A2(n19831), .B1(n19857), .B2(n20150), .ZN(
        n19824) );
  OAI211_X1 U22874 ( .C1(n19834), .C2(n10762), .A(n19825), .B(n19824), .ZN(
        P2_U3092) );
  AOI22_X1 U22875 ( .A1(n20156), .A2(n19857), .B1(n19839), .B2(n20154), .ZN(
        n19827) );
  AOI22_X1 U22876 ( .A1(n20155), .A2(n19831), .B1(n19830), .B2(n20102), .ZN(
        n19826) );
  OAI211_X1 U22877 ( .C1(n19834), .C2(n10816), .A(n19827), .B(n19826), .ZN(
        P2_U3093) );
  AOI22_X1 U22878 ( .A1(n20162), .A2(n19830), .B1(n20160), .B2(n19839), .ZN(
        n19829) );
  AOI22_X1 U22879 ( .A1(n20161), .A2(n19831), .B1(n19857), .B2(n20105), .ZN(
        n19828) );
  OAI211_X1 U22880 ( .C1(n19834), .C2(n10853), .A(n19829), .B(n19828), .ZN(
        P2_U3094) );
  AOI22_X1 U22881 ( .A1(n20172), .A2(n19857), .B1(n19839), .B2(n20168), .ZN(
        n19833) );
  AOI22_X1 U22882 ( .A1(n20170), .A2(n19831), .B1(n19830), .B2(n20110), .ZN(
        n19832) );
  OAI211_X1 U22883 ( .C1(n19834), .C2(n10886), .A(n19833), .B(n19832), .ZN(
        P2_U3095) );
  NOR2_X1 U22884 ( .A1(n20077), .A2(n19869), .ZN(n19860) );
  OAI21_X1 U22885 ( .B1(n19836), .B2(n19860), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19837) );
  OAI21_X1 U22886 ( .B1(n19869), .B2(n19838), .A(n19837), .ZN(n19861) );
  AOI22_X1 U22887 ( .A1(n19861), .A2(n14145), .B1(n20119), .B2(n19860), .ZN(
        n19846) );
  AOI221_X1 U22888 ( .B1(n19857), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19892), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19839), .ZN(n19840) );
  INV_X1 U22889 ( .A(n19860), .ZN(n19841) );
  OAI21_X1 U22890 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19840), .A(n19841), 
        .ZN(n19844) );
  NAND3_X1 U22891 ( .A1(n19842), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19841), 
        .ZN(n19843) );
  NAND3_X1 U22892 ( .A1(n19844), .A2(n20125), .A3(n19843), .ZN(n19862) );
  AOI22_X1 U22893 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20080), .ZN(n19845) );
  OAI211_X1 U22894 ( .C1(n19881), .C2(n19899), .A(n19846), .B(n19845), .ZN(
        P2_U3096) );
  AOI22_X1 U22895 ( .A1(n19861), .A2(n14194), .B1(n20131), .B2(n19860), .ZN(
        n19848) );
  AOI22_X1 U22896 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20132), .ZN(n19847) );
  OAI211_X1 U22897 ( .C1(n20135), .C2(n19899), .A(n19848), .B(n19847), .ZN(
        P2_U3097) );
  AOI22_X1 U22898 ( .A1(n19861), .A2(n20137), .B1(n20136), .B2(n19860), .ZN(
        n19850) );
  AOI22_X1 U22899 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20092), .ZN(n19849) );
  OAI211_X1 U22900 ( .C1(n20055), .C2(n19899), .A(n19850), .B(n19849), .ZN(
        P2_U3098) );
  AOI22_X1 U22901 ( .A1(n19861), .A2(n20143), .B1(n20142), .B2(n19860), .ZN(
        n19852) );
  AOI22_X1 U22902 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20095), .ZN(n19851) );
  OAI211_X1 U22903 ( .C1(n20025), .C2(n19899), .A(n19852), .B(n19851), .ZN(
        P2_U3099) );
  AOI22_X1 U22904 ( .A1(n19861), .A2(n20149), .B1(n20148), .B2(n19860), .ZN(
        n19854) );
  AOI22_X1 U22905 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20098), .ZN(n19853) );
  OAI211_X1 U22906 ( .C1(n19951), .C2(n19899), .A(n19854), .B(n19853), .ZN(
        P2_U3100) );
  AOI22_X1 U22907 ( .A1(n19861), .A2(n20155), .B1(n20154), .B2(n19860), .ZN(
        n19856) );
  AOI22_X1 U22908 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20102), .ZN(n19855) );
  OAI211_X1 U22909 ( .C1(n19973), .C2(n19899), .A(n19856), .B(n19855), .ZN(
        P2_U3101) );
  AOI22_X1 U22910 ( .A1(n19861), .A2(n20161), .B1(n20160), .B2(n19860), .ZN(
        n19859) );
  AOI22_X1 U22911 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19862), .B1(
        n19857), .B2(n20162), .ZN(n19858) );
  OAI211_X1 U22912 ( .C1(n20167), .C2(n19899), .A(n19859), .B(n19858), .ZN(
        P2_U3102) );
  AOI22_X1 U22913 ( .A1(n19861), .A2(n20170), .B1(n20168), .B2(n19860), .ZN(
        n19864) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19862), .B1(
        n19892), .B2(n20172), .ZN(n19863) );
  OAI211_X1 U22915 ( .C1(n20178), .C2(n19865), .A(n19864), .B(n19863), .ZN(
        P2_U3103) );
  NAND2_X1 U22916 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19867), .ZN(
        n19876) );
  OR2_X1 U22917 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19876), .ZN(n19872) );
  INV_X1 U22918 ( .A(n19868), .ZN(n19871) );
  NOR2_X1 U22919 ( .A1(n19870), .A2(n19869), .ZN(n19904) );
  NOR3_X1 U22920 ( .A1(n19871), .A2(n19904), .A3(n13514), .ZN(n19875) );
  AOI21_X1 U22921 ( .B1(n13514), .B2(n19872), .A(n19875), .ZN(n19895) );
  AOI22_X1 U22922 ( .A1(n19895), .A2(n14145), .B1(n20119), .B2(n19904), .ZN(
        n19880) );
  NAND2_X1 U22923 ( .A1(n19873), .A2(n20071), .ZN(n19877) );
  AOI211_X1 U22924 ( .C1(n19877), .C2(n19876), .A(n19875), .B(n19874), .ZN(
        n19878) );
  OAI21_X1 U22925 ( .B1(n19904), .B2(n19936), .A(n19878), .ZN(n19896) );
  AOI22_X1 U22926 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19896), .B1(
        n19892), .B2(n20080), .ZN(n19879) );
  OAI211_X1 U22927 ( .C1(n19881), .C2(n19930), .A(n19880), .B(n19879), .ZN(
        P2_U3104) );
  AOI22_X1 U22928 ( .A1(n19895), .A2(n14194), .B1(n20131), .B2(n19904), .ZN(
        n19883) );
  AOI22_X1 U22929 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19896), .B1(
        n19892), .B2(n20132), .ZN(n19882) );
  OAI211_X1 U22930 ( .C1(n20135), .C2(n19930), .A(n19883), .B(n19882), .ZN(
        P2_U3105) );
  AOI22_X1 U22931 ( .A1(n19895), .A2(n20137), .B1(n19904), .B2(n20136), .ZN(
        n19885) );
  AOI22_X1 U22932 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19896), .B1(
        n19892), .B2(n20092), .ZN(n19884) );
  OAI211_X1 U22933 ( .C1(n20055), .C2(n19930), .A(n19885), .B(n19884), .ZN(
        P2_U3106) );
  AOI22_X1 U22934 ( .A1(n19895), .A2(n20143), .B1(n19904), .B2(n20142), .ZN(
        n19887) );
  AOI22_X1 U22935 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19896), .B1(
        n19892), .B2(n20095), .ZN(n19886) );
  OAI211_X1 U22936 ( .C1(n20025), .C2(n19930), .A(n19887), .B(n19886), .ZN(
        P2_U3107) );
  AOI22_X1 U22937 ( .A1(n19895), .A2(n20149), .B1(n20148), .B2(n19904), .ZN(
        n19889) );
  AOI22_X1 U22938 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19896), .B1(
        n19892), .B2(n20098), .ZN(n19888) );
  OAI211_X1 U22939 ( .C1(n19951), .C2(n19930), .A(n19889), .B(n19888), .ZN(
        P2_U3108) );
  AOI22_X1 U22940 ( .A1(n19895), .A2(n20155), .B1(n19904), .B2(n20154), .ZN(
        n19891) );
  AOI22_X1 U22941 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19896), .B1(
        n19922), .B2(n20156), .ZN(n19890) );
  OAI211_X1 U22942 ( .C1(n20159), .C2(n19899), .A(n19891), .B(n19890), .ZN(
        P2_U3109) );
  AOI22_X1 U22943 ( .A1(n19895), .A2(n20161), .B1(n20160), .B2(n19904), .ZN(
        n19894) );
  AOI22_X1 U22944 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19896), .B1(
        n19892), .B2(n20162), .ZN(n19893) );
  OAI211_X1 U22945 ( .C1(n20167), .C2(n19930), .A(n19894), .B(n19893), .ZN(
        P2_U3110) );
  AOI22_X1 U22946 ( .A1(n19895), .A2(n20170), .B1(n19904), .B2(n20168), .ZN(
        n19898) );
  AOI22_X1 U22947 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19896), .B1(
        n19922), .B2(n20172), .ZN(n19897) );
  OAI211_X1 U22948 ( .C1(n20178), .C2(n19899), .A(n19898), .B(n19897), .ZN(
        P2_U3111) );
  NAND2_X1 U22949 ( .A1(n19900), .A2(n20288), .ZN(n19939) );
  NOR2_X1 U22950 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19939), .ZN(
        n19925) );
  AOI22_X1 U22951 ( .A1(n20127), .A2(n19954), .B1(n20119), .B2(n19925), .ZN(
        n19911) );
  OAI21_X1 U22952 ( .B1(n19954), .B2(n19922), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19901) );
  NAND2_X1 U22953 ( .A1(n19901), .A2(n20259), .ZN(n19909) );
  NOR2_X1 U22954 ( .A1(n19904), .A2(n19909), .ZN(n19902) );
  AOI211_X1 U22955 ( .C1(n19905), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19902), .ZN(n19903) );
  OAI21_X1 U22956 ( .B1(n19903), .B2(n19925), .A(n20125), .ZN(n19927) );
  NOR2_X1 U22957 ( .A1(n19904), .A2(n19925), .ZN(n19908) );
  INV_X1 U22958 ( .A(n19905), .ZN(n19906) );
  OAI21_X1 U22959 ( .B1(n19906), .B2(n19925), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19907) );
  AOI22_X1 U22960 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19927), .B1(
        n14145), .B2(n19926), .ZN(n19910) );
  OAI211_X1 U22961 ( .C1(n20130), .C2(n19930), .A(n19911), .B(n19910), .ZN(
        P2_U3112) );
  AOI22_X1 U22962 ( .A1(n20132), .A2(n19922), .B1(n20131), .B2(n19925), .ZN(
        n19913) );
  AOI22_X1 U22963 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n14194), .ZN(n19912) );
  OAI211_X1 U22964 ( .C1(n20135), .C2(n19962), .A(n19913), .B(n19912), .ZN(
        P2_U3113) );
  AOI22_X1 U22965 ( .A1(n20138), .A2(n19954), .B1(n19925), .B2(n20136), .ZN(
        n19915) );
  AOI22_X1 U22966 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n20137), .ZN(n19914) );
  OAI211_X1 U22967 ( .C1(n20141), .C2(n19930), .A(n19915), .B(n19914), .ZN(
        P2_U3114) );
  AOI22_X1 U22968 ( .A1(n20095), .A2(n19922), .B1(n20142), .B2(n19925), .ZN(
        n19917) );
  AOI22_X1 U22969 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n20143), .ZN(n19916) );
  OAI211_X1 U22970 ( .C1(n20025), .C2(n19962), .A(n19917), .B(n19916), .ZN(
        P2_U3115) );
  AOI22_X1 U22971 ( .A1(n20150), .A2(n19954), .B1(n20148), .B2(n19925), .ZN(
        n19919) );
  AOI22_X1 U22972 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n20149), .ZN(n19918) );
  OAI211_X1 U22973 ( .C1(n20153), .C2(n19930), .A(n19919), .B(n19918), .ZN(
        P2_U3116) );
  AOI22_X1 U22974 ( .A1(n20102), .A2(n19922), .B1(n20154), .B2(n19925), .ZN(
        n19921) );
  AOI22_X1 U22975 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n20155), .ZN(n19920) );
  OAI211_X1 U22976 ( .C1(n19973), .C2(n19962), .A(n19921), .B(n19920), .ZN(
        P2_U3117) );
  AOI22_X1 U22977 ( .A1(n20162), .A2(n19922), .B1(n20160), .B2(n19925), .ZN(
        n19924) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n20161), .ZN(n19923) );
  OAI211_X1 U22979 ( .C1(n20167), .C2(n19962), .A(n19924), .B(n19923), .ZN(
        P2_U3118) );
  AOI22_X1 U22980 ( .A1(n20172), .A2(n19954), .B1(n20168), .B2(n19925), .ZN(
        n19929) );
  AOI22_X1 U22981 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19927), .B1(
        n19926), .B2(n20170), .ZN(n19928) );
  OAI211_X1 U22982 ( .C1(n20178), .C2(n19930), .A(n19929), .B(n19928), .ZN(
        P2_U3119) );
  AOI22_X1 U22983 ( .A1(n20127), .A2(n19974), .B1(n20119), .B2(n19957), .ZN(
        n19942) );
  INV_X1 U22984 ( .A(n20121), .ZN(n19932) );
  AOI21_X1 U22985 ( .B1(n19932), .B2(n19931), .A(n20261), .ZN(n19937) );
  INV_X1 U22986 ( .A(n19933), .ZN(n19934) );
  NOR2_X1 U22987 ( .A1(n19934), .A2(n19957), .ZN(n19938) );
  AOI22_X1 U22988 ( .A1(n19937), .A2(n19939), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19938), .ZN(n19935) );
  OAI211_X1 U22989 ( .C1(n19957), .C2(n19936), .A(n19935), .B(n20125), .ZN(
        n19959) );
  INV_X1 U22990 ( .A(n19937), .ZN(n19940) );
  AOI22_X1 U22991 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19959), .B1(
        n14145), .B2(n19958), .ZN(n19941) );
  OAI211_X1 U22992 ( .C1(n20130), .C2(n19962), .A(n19942), .B(n19941), .ZN(
        P2_U3120) );
  AOI22_X1 U22993 ( .A1(n20132), .A2(n19954), .B1(n20131), .B2(n19957), .ZN(
        n19944) );
  AOI22_X1 U22994 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19959), .B1(
        n14194), .B2(n19958), .ZN(n19943) );
  OAI211_X1 U22995 ( .C1(n20135), .C2(n19982), .A(n19944), .B(n19943), .ZN(
        P2_U3121) );
  AOI22_X1 U22996 ( .A1(n20138), .A2(n19974), .B1(n20136), .B2(n19957), .ZN(
        n19946) );
  AOI22_X1 U22997 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19959), .B1(
        n20137), .B2(n19958), .ZN(n19945) );
  OAI211_X1 U22998 ( .C1(n20141), .C2(n19962), .A(n19946), .B(n19945), .ZN(
        P2_U3122) );
  AOI22_X1 U22999 ( .A1(n20095), .A2(n19954), .B1(n20142), .B2(n19957), .ZN(
        n19948) );
  AOI22_X1 U23000 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19959), .B1(
        n20143), .B2(n19958), .ZN(n19947) );
  OAI211_X1 U23001 ( .C1(n20025), .C2(n19982), .A(n19948), .B(n19947), .ZN(
        P2_U3123) );
  AOI22_X1 U23002 ( .A1(n20098), .A2(n19954), .B1(n20148), .B2(n19957), .ZN(
        n19950) );
  AOI22_X1 U23003 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19959), .B1(
        n20149), .B2(n19958), .ZN(n19949) );
  OAI211_X1 U23004 ( .C1(n19951), .C2(n19982), .A(n19950), .B(n19949), .ZN(
        P2_U3124) );
  AOI22_X1 U23005 ( .A1(n20156), .A2(n19974), .B1(n20154), .B2(n19957), .ZN(
        n19953) );
  AOI22_X1 U23006 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19959), .B1(
        n20155), .B2(n19958), .ZN(n19952) );
  OAI211_X1 U23007 ( .C1(n20159), .C2(n19962), .A(n19953), .B(n19952), .ZN(
        P2_U3125) );
  AOI22_X1 U23008 ( .A1(n20162), .A2(n19954), .B1(n20160), .B2(n19957), .ZN(
        n19956) );
  AOI22_X1 U23009 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19959), .B1(
        n20161), .B2(n19958), .ZN(n19955) );
  OAI211_X1 U23010 ( .C1(n20167), .C2(n19982), .A(n19956), .B(n19955), .ZN(
        P2_U3126) );
  AOI22_X1 U23011 ( .A1(n20172), .A2(n19974), .B1(n20168), .B2(n19957), .ZN(
        n19961) );
  AOI22_X1 U23012 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19959), .B1(
        n20170), .B2(n19958), .ZN(n19960) );
  OAI211_X1 U23013 ( .C1(n20178), .C2(n19962), .A(n19961), .B(n19960), .ZN(
        P2_U3127) );
  AOI22_X1 U23014 ( .A1(n19978), .A2(n14194), .B1(n20131), .B2(n19977), .ZN(
        n19964) );
  AOI22_X1 U23015 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19979), .B1(
        n19974), .B2(n20132), .ZN(n19963) );
  OAI211_X1 U23016 ( .C1(n20135), .C2(n20001), .A(n19964), .B(n19963), .ZN(
        P2_U3129) );
  AOI22_X1 U23017 ( .A1(n19978), .A2(n20137), .B1(n20136), .B2(n19977), .ZN(
        n19966) );
  AOI22_X1 U23018 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19979), .B1(
        n19992), .B2(n20138), .ZN(n19965) );
  OAI211_X1 U23019 ( .C1(n20141), .C2(n19982), .A(n19966), .B(n19965), .ZN(
        P2_U3130) );
  AOI22_X1 U23020 ( .A1(n19978), .A2(n20143), .B1(n20142), .B2(n19977), .ZN(
        n19968) );
  AOI22_X1 U23021 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19979), .B1(
        n19974), .B2(n20095), .ZN(n19967) );
  OAI211_X1 U23022 ( .C1(n20025), .C2(n20001), .A(n19968), .B(n19967), .ZN(
        P2_U3131) );
  AOI22_X1 U23023 ( .A1(n19978), .A2(n20149), .B1(n20148), .B2(n19977), .ZN(
        n19970) );
  AOI22_X1 U23024 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19979), .B1(
        n19992), .B2(n20150), .ZN(n19969) );
  OAI211_X1 U23025 ( .C1(n20153), .C2(n19982), .A(n19970), .B(n19969), .ZN(
        P2_U3132) );
  AOI22_X1 U23026 ( .A1(n19978), .A2(n20155), .B1(n20154), .B2(n19977), .ZN(
        n19972) );
  AOI22_X1 U23027 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19979), .B1(
        n19974), .B2(n20102), .ZN(n19971) );
  OAI211_X1 U23028 ( .C1(n19973), .C2(n20001), .A(n19972), .B(n19971), .ZN(
        P2_U3133) );
  AOI22_X1 U23029 ( .A1(n19978), .A2(n20161), .B1(n20160), .B2(n19977), .ZN(
        n19976) );
  AOI22_X1 U23030 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19979), .B1(
        n19974), .B2(n20162), .ZN(n19975) );
  OAI211_X1 U23031 ( .C1(n20167), .C2(n20001), .A(n19976), .B(n19975), .ZN(
        P2_U3134) );
  AOI22_X1 U23032 ( .A1(n19978), .A2(n20170), .B1(n20168), .B2(n19977), .ZN(
        n19981) );
  AOI22_X1 U23033 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19979), .B1(
        n19992), .B2(n20172), .ZN(n19980) );
  OAI211_X1 U23034 ( .C1(n20178), .C2(n19982), .A(n19981), .B(n19980), .ZN(
        P2_U3135) );
  AOI22_X1 U23035 ( .A1(n19997), .A2(n20137), .B1(n19996), .B2(n20136), .ZN(
        n19984) );
  AOI22_X1 U23036 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19998), .B1(
        n20030), .B2(n20138), .ZN(n19983) );
  OAI211_X1 U23037 ( .C1(n20141), .C2(n20001), .A(n19984), .B(n19983), .ZN(
        P2_U3138) );
  AOI22_X1 U23038 ( .A1(n19997), .A2(n20143), .B1(n19996), .B2(n20142), .ZN(
        n19986) );
  AOI22_X1 U23039 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19998), .B1(
        n20030), .B2(n20144), .ZN(n19985) );
  OAI211_X1 U23040 ( .C1(n20147), .C2(n20001), .A(n19986), .B(n19985), .ZN(
        P2_U3139) );
  INV_X1 U23041 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U23042 ( .A1(n19997), .A2(n20149), .B1(n20148), .B2(n19996), .ZN(
        n19988) );
  AOI22_X1 U23043 ( .A1(n20030), .A2(n20150), .B1(n19992), .B2(n20098), .ZN(
        n19987) );
  OAI211_X1 U23044 ( .C1(n19995), .C2(n19989), .A(n19988), .B(n19987), .ZN(
        P2_U3140) );
  AOI22_X1 U23045 ( .A1(n19997), .A2(n20155), .B1(n19996), .B2(n20154), .ZN(
        n19991) );
  AOI22_X1 U23046 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19998), .B1(
        n20030), .B2(n20156), .ZN(n19990) );
  OAI211_X1 U23047 ( .C1(n20159), .C2(n20001), .A(n19991), .B(n19990), .ZN(
        P2_U3141) );
  AOI22_X1 U23048 ( .A1(n19997), .A2(n20161), .B1(n20160), .B2(n19996), .ZN(
        n19994) );
  AOI22_X1 U23049 ( .A1(n19992), .A2(n20162), .B1(n20030), .B2(n20105), .ZN(
        n19993) );
  OAI211_X1 U23050 ( .C1(n19995), .C2(n10836), .A(n19994), .B(n19993), .ZN(
        P2_U3142) );
  AOI22_X1 U23051 ( .A1(n19997), .A2(n20170), .B1(n19996), .B2(n20168), .ZN(
        n20000) );
  AOI22_X1 U23052 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19998), .B1(
        n20030), .B2(n20172), .ZN(n19999) );
  OAI211_X1 U23053 ( .C1(n20178), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P2_U3143) );
  AOI21_X1 U23054 ( .B1(n20038), .B2(n20070), .A(n21288), .ZN(n20003) );
  AOI21_X1 U23055 ( .B1(n20009), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20003), .ZN(n20007) );
  NAND2_X1 U23056 ( .A1(n13089), .A2(n20288), .ZN(n20043) );
  NOR2_X1 U23057 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20043), .ZN(
        n20033) );
  NOR2_X1 U23058 ( .A1(n20259), .A2(n20033), .ZN(n20004) );
  OAI21_X1 U23059 ( .B1(n20010), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20004), 
        .ZN(n20005) );
  NAND2_X1 U23060 ( .A1(n20005), .A2(n20125), .ZN(n20006) );
  INV_X1 U23061 ( .A(n20035), .ZN(n20018) );
  INV_X1 U23062 ( .A(n20008), .ZN(n20014) );
  INV_X1 U23063 ( .A(n20009), .ZN(n20013) );
  INV_X1 U23064 ( .A(n20010), .ZN(n20011) );
  OAI21_X1 U23065 ( .B1(n20011), .B2(n20033), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20012) );
  OAI21_X1 U23066 ( .B1(n20014), .B2(n20013), .A(n20012), .ZN(n20034) );
  AOI22_X1 U23067 ( .A1(n20034), .A2(n14145), .B1(n20119), .B2(n20033), .ZN(
        n20016) );
  AOI22_X1 U23068 ( .A1(n20062), .A2(n20127), .B1(n20030), .B2(n20080), .ZN(
        n20015) );
  OAI211_X1 U23069 ( .C1(n20018), .C2(n20017), .A(n20016), .B(n20015), .ZN(
        P2_U3144) );
  AOI22_X1 U23070 ( .A1(n20034), .A2(n14194), .B1(n20131), .B2(n20033), .ZN(
        n20020) );
  AOI22_X1 U23071 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20035), .B1(
        n20030), .B2(n20132), .ZN(n20019) );
  OAI211_X1 U23072 ( .C1(n20135), .C2(n20070), .A(n20020), .B(n20019), .ZN(
        P2_U3145) );
  AOI22_X1 U23073 ( .A1(n20034), .A2(n20137), .B1(n20136), .B2(n20033), .ZN(
        n20022) );
  AOI22_X1 U23074 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20035), .B1(
        n20030), .B2(n20092), .ZN(n20021) );
  OAI211_X1 U23075 ( .C1(n20055), .C2(n20070), .A(n20022), .B(n20021), .ZN(
        P2_U3146) );
  AOI22_X1 U23076 ( .A1(n20034), .A2(n20143), .B1(n20142), .B2(n20033), .ZN(
        n20024) );
  AOI22_X1 U23077 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20035), .B1(
        n20030), .B2(n20095), .ZN(n20023) );
  OAI211_X1 U23078 ( .C1(n20025), .C2(n20070), .A(n20024), .B(n20023), .ZN(
        P2_U3147) );
  AOI22_X1 U23079 ( .A1(n20034), .A2(n20149), .B1(n20148), .B2(n20033), .ZN(
        n20027) );
  AOI22_X1 U23080 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20035), .B1(
        n20062), .B2(n20150), .ZN(n20026) );
  OAI211_X1 U23081 ( .C1(n20153), .C2(n20038), .A(n20027), .B(n20026), .ZN(
        P2_U3148) );
  AOI22_X1 U23082 ( .A1(n20034), .A2(n20155), .B1(n20154), .B2(n20033), .ZN(
        n20029) );
  AOI22_X1 U23083 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20035), .B1(
        n20062), .B2(n20156), .ZN(n20028) );
  OAI211_X1 U23084 ( .C1(n20159), .C2(n20038), .A(n20029), .B(n20028), .ZN(
        P2_U3149) );
  AOI22_X1 U23085 ( .A1(n20034), .A2(n20161), .B1(n20160), .B2(n20033), .ZN(
        n20032) );
  AOI22_X1 U23086 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20035), .B1(
        n20030), .B2(n20162), .ZN(n20031) );
  OAI211_X1 U23087 ( .C1(n20167), .C2(n20070), .A(n20032), .B(n20031), .ZN(
        P2_U3150) );
  AOI22_X1 U23088 ( .A1(n20034), .A2(n20170), .B1(n20168), .B2(n20033), .ZN(
        n20037) );
  AOI22_X1 U23089 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20035), .B1(
        n20062), .B2(n20172), .ZN(n20036) );
  OAI211_X1 U23090 ( .C1(n20178), .C2(n20038), .A(n20037), .B(n20036), .ZN(
        P2_U3151) );
  INV_X1 U23091 ( .A(n20042), .ZN(n20040) );
  NOR2_X1 U23092 ( .A1(n20120), .A2(n20039), .ZN(n20065) );
  OAI21_X1 U23093 ( .B1(n20040), .B2(n20065), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20041) );
  OAI21_X1 U23094 ( .B1(n20043), .B2(n20261), .A(n20041), .ZN(n20066) );
  AOI22_X1 U23095 ( .A1(n20066), .A2(n14145), .B1(n20119), .B2(n20065), .ZN(
        n20050) );
  AOI21_X1 U23096 ( .B1(n20042), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20045) );
  OAI21_X1 U23097 ( .B1(n20121), .B2(n20046), .A(n20043), .ZN(n20044) );
  OAI211_X1 U23098 ( .C1(n20065), .C2(n20045), .A(n20044), .B(n20125), .ZN(
        n20067) );
  INV_X1 U23099 ( .A(n20046), .ZN(n20047) );
  AOI22_X1 U23100 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20067), .B1(
        n20109), .B2(n20127), .ZN(n20049) );
  OAI211_X1 U23101 ( .C1(n20130), .C2(n20070), .A(n20050), .B(n20049), .ZN(
        P2_U3152) );
  AOI22_X1 U23102 ( .A1(n20066), .A2(n14194), .B1(n20131), .B2(n20065), .ZN(
        n20052) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20067), .B1(
        n20062), .B2(n20132), .ZN(n20051) );
  OAI211_X1 U23104 ( .C1(n20135), .C2(n20073), .A(n20052), .B(n20051), .ZN(
        P2_U3153) );
  AOI22_X1 U23105 ( .A1(n20066), .A2(n20137), .B1(n20136), .B2(n20065), .ZN(
        n20054) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20067), .B1(
        n20062), .B2(n20092), .ZN(n20053) );
  OAI211_X1 U23107 ( .C1(n20055), .C2(n20073), .A(n20054), .B(n20053), .ZN(
        P2_U3154) );
  AOI22_X1 U23108 ( .A1(n20066), .A2(n20143), .B1(n20142), .B2(n20065), .ZN(
        n20057) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20067), .B1(
        n20109), .B2(n20144), .ZN(n20056) );
  OAI211_X1 U23110 ( .C1(n20147), .C2(n20070), .A(n20057), .B(n20056), .ZN(
        P2_U3155) );
  AOI22_X1 U23111 ( .A1(n20066), .A2(n20149), .B1(n20148), .B2(n20065), .ZN(
        n20059) );
  AOI22_X1 U23112 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20067), .B1(
        n20109), .B2(n20150), .ZN(n20058) );
  OAI211_X1 U23113 ( .C1(n20153), .C2(n20070), .A(n20059), .B(n20058), .ZN(
        P2_U3156) );
  AOI22_X1 U23114 ( .A1(n20066), .A2(n20155), .B1(n20154), .B2(n20065), .ZN(
        n20061) );
  AOI22_X1 U23115 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20067), .B1(
        n20109), .B2(n20156), .ZN(n20060) );
  OAI211_X1 U23116 ( .C1(n20159), .C2(n20070), .A(n20061), .B(n20060), .ZN(
        P2_U3157) );
  AOI22_X1 U23117 ( .A1(n20066), .A2(n20161), .B1(n20160), .B2(n20065), .ZN(
        n20064) );
  AOI22_X1 U23118 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20067), .B1(
        n20062), .B2(n20162), .ZN(n20063) );
  OAI211_X1 U23119 ( .C1(n20167), .C2(n20073), .A(n20064), .B(n20063), .ZN(
        P2_U3158) );
  AOI22_X1 U23120 ( .A1(n20066), .A2(n20170), .B1(n20168), .B2(n20065), .ZN(
        n20069) );
  AOI22_X1 U23121 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20067), .B1(
        n20109), .B2(n20172), .ZN(n20068) );
  OAI211_X1 U23122 ( .C1(n20178), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P2_U3159) );
  AOI21_X1 U23123 ( .B1(n20073), .B2(n20177), .A(n21288), .ZN(n20074) );
  NOR2_X1 U23124 ( .A1(n20074), .A2(n20261), .ZN(n20081) );
  NAND2_X1 U23125 ( .A1(n20075), .A2(n13089), .ZN(n20084) );
  AOI21_X1 U23126 ( .B1(n20076), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20078) );
  NOR2_X1 U23127 ( .A1(n20120), .A2(n20077), .ZN(n20108) );
  OAI21_X1 U23128 ( .B1(n20078), .B2(n20108), .A(n20125), .ZN(n20079) );
  AOI22_X1 U23129 ( .A1(n20080), .A2(n20109), .B1(n20119), .B2(n20108), .ZN(
        n20087) );
  INV_X1 U23130 ( .A(n20081), .ZN(n20085) );
  OAI21_X1 U23131 ( .B1(n20082), .B2(n20108), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20083) );
  AOI22_X1 U23132 ( .A1(n14145), .A2(n20111), .B1(n20163), .B2(n20127), .ZN(
        n20086) );
  OAI211_X1 U23133 ( .C1(n20115), .C2(n20088), .A(n20087), .B(n20086), .ZN(
        P2_U3160) );
  AOI22_X1 U23134 ( .A1(n20132), .A2(n20109), .B1(n20131), .B2(n20108), .ZN(
        n20091) );
  AOI22_X1 U23135 ( .A1(n14194), .A2(n20111), .B1(n20163), .B2(n20089), .ZN(
        n20090) );
  OAI211_X1 U23136 ( .C1(n20115), .C2(n11056), .A(n20091), .B(n20090), .ZN(
        P2_U3161) );
  AOI22_X1 U23137 ( .A1(n20092), .A2(n20109), .B1(n20136), .B2(n20108), .ZN(
        n20094) );
  AOI22_X1 U23138 ( .A1(n20137), .A2(n20111), .B1(n20163), .B2(n20138), .ZN(
        n20093) );
  OAI211_X1 U23139 ( .C1(n20115), .C2(n11072), .A(n20094), .B(n20093), .ZN(
        P2_U3162) );
  AOI22_X1 U23140 ( .A1(n20095), .A2(n20109), .B1(n20142), .B2(n20108), .ZN(
        n20097) );
  AOI22_X1 U23141 ( .A1(n20143), .A2(n20111), .B1(n20163), .B2(n20144), .ZN(
        n20096) );
  OAI211_X1 U23142 ( .C1(n20115), .C2(n11106), .A(n20097), .B(n20096), .ZN(
        P2_U3163) );
  INV_X1 U23143 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20101) );
  AOI22_X1 U23144 ( .A1(n20098), .A2(n20109), .B1(n20148), .B2(n20108), .ZN(
        n20100) );
  AOI22_X1 U23145 ( .A1(n20149), .A2(n20111), .B1(n20163), .B2(n20150), .ZN(
        n20099) );
  OAI211_X1 U23146 ( .C1(n20115), .C2(n20101), .A(n20100), .B(n20099), .ZN(
        P2_U3164) );
  AOI22_X1 U23147 ( .A1(n20102), .A2(n20109), .B1(n20154), .B2(n20108), .ZN(
        n20104) );
  AOI22_X1 U23148 ( .A1(n20155), .A2(n20111), .B1(n20163), .B2(n20156), .ZN(
        n20103) );
  OAI211_X1 U23149 ( .C1(n20115), .C2(n11143), .A(n20104), .B(n20103), .ZN(
        P2_U3165) );
  AOI22_X1 U23150 ( .A1(n20162), .A2(n20109), .B1(n20160), .B2(n20108), .ZN(
        n20107) );
  AOI22_X1 U23151 ( .A1(n20161), .A2(n20111), .B1(n20163), .B2(n20105), .ZN(
        n20106) );
  OAI211_X1 U23152 ( .C1(n20115), .C2(n11161), .A(n20107), .B(n20106), .ZN(
        P2_U3166) );
  AOI22_X1 U23153 ( .A1(n20110), .A2(n20109), .B1(n20168), .B2(n20108), .ZN(
        n20113) );
  AOI22_X1 U23154 ( .A1(n20170), .A2(n20111), .B1(n20163), .B2(n20172), .ZN(
        n20112) );
  OAI211_X1 U23155 ( .C1(n20115), .C2(n20114), .A(n20113), .B(n20112), .ZN(
        P2_U3167) );
  NAND2_X1 U23156 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n13089), .ZN(
        n20118) );
  INV_X1 U23157 ( .A(n20123), .ZN(n20116) );
  INV_X1 U23158 ( .A(n20122), .ZN(n20169) );
  OAI21_X1 U23159 ( .B1(n20116), .B2(n20169), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20117) );
  OAI21_X1 U23160 ( .B1(n20118), .B2(n20261), .A(n20117), .ZN(n20171) );
  AOI22_X1 U23161 ( .A1(n20171), .A2(n14145), .B1(n20169), .B2(n20119), .ZN(
        n20129) );
  OAI22_X1 U23162 ( .A1(n20121), .A2(n20257), .B1(n20120), .B2(n20288), .ZN(
        n20126) );
  OAI211_X1 U23163 ( .C1(n20123), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20122), 
        .B(n20261), .ZN(n20124) );
  NAND3_X1 U23164 ( .A1(n20126), .A2(n20125), .A3(n20124), .ZN(n20174) );
  AOI22_X1 U23165 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20127), .ZN(n20128) );
  OAI211_X1 U23166 ( .C1(n20130), .C2(n20177), .A(n20129), .B(n20128), .ZN(
        P2_U3168) );
  AOI22_X1 U23167 ( .A1(n20171), .A2(n14194), .B1(n20169), .B2(n20131), .ZN(
        n20134) );
  AOI22_X1 U23168 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20174), .B1(
        n20163), .B2(n20132), .ZN(n20133) );
  OAI211_X1 U23169 ( .C1(n20135), .C2(n20166), .A(n20134), .B(n20133), .ZN(
        P2_U3169) );
  AOI22_X1 U23170 ( .A1(n20171), .A2(n20137), .B1(n20169), .B2(n20136), .ZN(
        n20140) );
  AOI22_X1 U23171 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20138), .ZN(n20139) );
  OAI211_X1 U23172 ( .C1(n20141), .C2(n20177), .A(n20140), .B(n20139), .ZN(
        P2_U3170) );
  AOI22_X1 U23173 ( .A1(n20171), .A2(n20143), .B1(n20169), .B2(n20142), .ZN(
        n20146) );
  AOI22_X1 U23174 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20144), .ZN(n20145) );
  OAI211_X1 U23175 ( .C1(n20147), .C2(n20177), .A(n20146), .B(n20145), .ZN(
        P2_U3171) );
  AOI22_X1 U23176 ( .A1(n20171), .A2(n20149), .B1(n20169), .B2(n20148), .ZN(
        n20152) );
  AOI22_X1 U23177 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20150), .ZN(n20151) );
  OAI211_X1 U23178 ( .C1(n20153), .C2(n20177), .A(n20152), .B(n20151), .ZN(
        P2_U3172) );
  AOI22_X1 U23179 ( .A1(n20171), .A2(n20155), .B1(n20169), .B2(n20154), .ZN(
        n20158) );
  AOI22_X1 U23180 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20156), .ZN(n20157) );
  OAI211_X1 U23181 ( .C1(n20159), .C2(n20177), .A(n20158), .B(n20157), .ZN(
        P2_U3173) );
  AOI22_X1 U23182 ( .A1(n20171), .A2(n20161), .B1(n20169), .B2(n20160), .ZN(
        n20165) );
  AOI22_X1 U23183 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20174), .B1(
        n20163), .B2(n20162), .ZN(n20164) );
  OAI211_X1 U23184 ( .C1(n20167), .C2(n20166), .A(n20165), .B(n20164), .ZN(
        P2_U3174) );
  AOI22_X1 U23185 ( .A1(n20171), .A2(n20170), .B1(n20169), .B2(n20168), .ZN(
        n20176) );
  AOI22_X1 U23186 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20172), .ZN(n20175) );
  OAI211_X1 U23187 ( .C1(n20178), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        P2_U3175) );
  NOR2_X1 U23188 ( .A1(n21090), .A2(n20256), .ZN(P2_U3179) );
  AND2_X1 U23189 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20179), .ZN(
        P2_U3180) );
  AND2_X1 U23190 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20179), .ZN(
        P2_U3181) );
  AND2_X1 U23191 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20179), .ZN(
        P2_U3182) );
  AND2_X1 U23192 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20179), .ZN(
        P2_U3183) );
  AND2_X1 U23193 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20179), .ZN(
        P2_U3184) );
  AND2_X1 U23194 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20179), .ZN(
        P2_U3185) );
  AND2_X1 U23195 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20179), .ZN(
        P2_U3186) );
  AND2_X1 U23196 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20179), .ZN(
        P2_U3187) );
  INV_X1 U23197 ( .A(P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n21142) );
  NOR2_X1 U23198 ( .A1(n21142), .A2(n20256), .ZN(P2_U3188) );
  AND2_X1 U23199 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20179), .ZN(
        P2_U3189) );
  AND2_X1 U23200 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20179), .ZN(
        P2_U3190) );
  AND2_X1 U23201 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20179), .ZN(
        P2_U3191) );
  AND2_X1 U23202 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20179), .ZN(
        P2_U3192) );
  AND2_X1 U23203 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20179), .ZN(
        P2_U3193) );
  AND2_X1 U23204 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20179), .ZN(
        P2_U3194) );
  AND2_X1 U23205 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20179), .ZN(
        P2_U3195) );
  AND2_X1 U23206 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20179), .ZN(
        P2_U3196) );
  AND2_X1 U23207 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20179), .ZN(
        P2_U3197) );
  AND2_X1 U23208 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20179), .ZN(
        P2_U3198) );
  AND2_X1 U23209 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20179), .ZN(
        P2_U3199) );
  AND2_X1 U23210 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20179), .ZN(
        P2_U3200) );
  AND2_X1 U23211 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20179), .ZN(P2_U3201) );
  AND2_X1 U23212 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20179), .ZN(P2_U3202) );
  AND2_X1 U23213 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20179), .ZN(P2_U3203) );
  AND2_X1 U23214 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20179), .ZN(P2_U3204) );
  AND2_X1 U23215 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20179), .ZN(P2_U3205) );
  AND2_X1 U23216 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20179), .ZN(P2_U3206) );
  AND2_X1 U23217 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20179), .ZN(P2_U3207) );
  NOR2_X1 U23218 ( .A1(n20180), .A2(n20256), .ZN(P2_U3208) );
  AOI21_X1 U23219 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n20981), .A(n20181), .ZN(n20185) );
  INV_X1 U23220 ( .A(NA), .ZN(n20993) );
  OAI21_X1 U23221 ( .B1(n20993), .B2(n20190), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20199) );
  NOR2_X1 U23222 ( .A1(n20183), .A2(n20182), .ZN(n20187) );
  INV_X1 U23223 ( .A(n20187), .ZN(n20197) );
  NAND3_X1 U23224 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20197), .ZN(n20184) );
  AOI22_X1 U23225 ( .A1(n20185), .A2(n20315), .B1(n20199), .B2(n20184), .ZN(
        n20186) );
  INV_X1 U23226 ( .A(n20186), .ZN(P2_U3209) );
  NOR2_X1 U23227 ( .A1(n20188), .A2(n20187), .ZN(n20192) );
  NOR2_X1 U23228 ( .A1(HOLD), .A2(n20189), .ZN(n20198) );
  OAI211_X1 U23229 ( .C1(n20198), .C2(n20200), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n20190), .ZN(n20191) );
  OAI211_X1 U23230 ( .C1(n20193), .C2(n20981), .A(n20192), .B(n20191), .ZN(
        P2_U3210) );
  OAI22_X1 U23231 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20194), .B1(NA), 
        .B2(n20197), .ZN(n20195) );
  OAI211_X1 U23232 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20195), .ZN(n20196) );
  OAI221_X1 U23233 ( .B1(n20199), .B2(n20198), .C1(n20199), .C2(n20197), .A(
        n20196), .ZN(P2_U3211) );
  OAI222_X1 U23234 ( .A1(n20247), .A2(n20202), .B1(n20201), .B2(n20314), .C1(
        n20204), .C2(n20249), .ZN(P2_U3212) );
  OAI222_X1 U23235 ( .A1(n20247), .A2(n20204), .B1(n20203), .B2(n20314), .C1(
        n20205), .C2(n20249), .ZN(P2_U3213) );
  INV_X1 U23236 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20206) );
  OAI222_X1 U23237 ( .A1(n20247), .A2(n20205), .B1(n21237), .B2(n20314), .C1(
        n20206), .C2(n20249), .ZN(P2_U3214) );
  OAI222_X1 U23238 ( .A1(n20249), .A2(n15768), .B1(n20207), .B2(n20314), .C1(
        n20206), .C2(n20247), .ZN(P2_U3215) );
  OAI222_X1 U23239 ( .A1(n20249), .A2(n20209), .B1(n20208), .B2(n20314), .C1(
        n15768), .C2(n20247), .ZN(P2_U3216) );
  OAI222_X1 U23240 ( .A1(n20249), .A2(n20211), .B1(n20210), .B2(n20314), .C1(
        n20209), .C2(n20247), .ZN(P2_U3217) );
  INV_X1 U23241 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20212) );
  OAI222_X1 U23242 ( .A1(n20249), .A2(n20212), .B1(n21080), .B2(n20314), .C1(
        n20211), .C2(n20247), .ZN(P2_U3218) );
  OAI222_X1 U23243 ( .A1(n20249), .A2(n15748), .B1(n20213), .B2(n20314), .C1(
        n20212), .C2(n20247), .ZN(P2_U3219) );
  OAI222_X1 U23244 ( .A1(n20249), .A2(n20215), .B1(n20214), .B2(n20314), .C1(
        n15748), .C2(n20247), .ZN(P2_U3220) );
  OAI222_X1 U23245 ( .A1(n20249), .A2(n21297), .B1(n20216), .B2(n20314), .C1(
        n20215), .C2(n20247), .ZN(P2_U3221) );
  OAI222_X1 U23246 ( .A1(n20249), .A2(n20217), .B1(n21227), .B2(n20314), .C1(
        n21297), .C2(n20247), .ZN(P2_U3222) );
  INV_X1 U23247 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20219) );
  OAI222_X1 U23248 ( .A1(n20249), .A2(n20219), .B1(n20218), .B2(n20314), .C1(
        n20217), .C2(n20247), .ZN(P2_U3223) );
  OAI222_X1 U23249 ( .A1(n20249), .A2(n11265), .B1(n20220), .B2(n20314), .C1(
        n20219), .C2(n20247), .ZN(P2_U3224) );
  OAI222_X1 U23250 ( .A1(n20249), .A2(n20222), .B1(n20221), .B2(n20314), .C1(
        n11265), .C2(n20247), .ZN(P2_U3225) );
  INV_X1 U23251 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20224) );
  OAI222_X1 U23252 ( .A1(n20249), .A2(n20224), .B1(n20223), .B2(n20314), .C1(
        n20222), .C2(n20247), .ZN(P2_U3226) );
  OAI222_X1 U23253 ( .A1(n20249), .A2(n20226), .B1(n20225), .B2(n20314), .C1(
        n20224), .C2(n20247), .ZN(P2_U3227) );
  OAI222_X1 U23254 ( .A1(n20249), .A2(n20227), .B1(n21202), .B2(n20314), .C1(
        n20226), .C2(n20247), .ZN(P2_U3228) );
  OAI222_X1 U23255 ( .A1(n20249), .A2(n20229), .B1(n20228), .B2(n20314), .C1(
        n20227), .C2(n20247), .ZN(P2_U3229) );
  OAI222_X1 U23256 ( .A1(n20249), .A2(n20230), .B1(n21280), .B2(n20314), .C1(
        n20229), .C2(n20247), .ZN(P2_U3230) );
  OAI222_X1 U23257 ( .A1(n20249), .A2(n20232), .B1(n20231), .B2(n20314), .C1(
        n20230), .C2(n20247), .ZN(P2_U3231) );
  OAI222_X1 U23258 ( .A1(n20249), .A2(n21096), .B1(n20233), .B2(n20314), .C1(
        n20232), .C2(n20247), .ZN(P2_U3232) );
  OAI222_X1 U23259 ( .A1(n20249), .A2(n21139), .B1(n20234), .B2(n20314), .C1(
        n21096), .C2(n20247), .ZN(P2_U3233) );
  OAI222_X1 U23260 ( .A1(n20249), .A2(n20236), .B1(n20235), .B2(n20314), .C1(
        n21139), .C2(n20247), .ZN(P2_U3234) );
  OAI222_X1 U23261 ( .A1(n20249), .A2(n20238), .B1(n20237), .B2(n20314), .C1(
        n20236), .C2(n20247), .ZN(P2_U3235) );
  OAI222_X1 U23262 ( .A1(n20249), .A2(n20240), .B1(n20239), .B2(n20314), .C1(
        n20238), .C2(n20247), .ZN(P2_U3236) );
  OAI222_X1 U23263 ( .A1(n20249), .A2(n20243), .B1(n20241), .B2(n20314), .C1(
        n20240), .C2(n20247), .ZN(P2_U3237) );
  OAI222_X1 U23264 ( .A1(n20247), .A2(n20243), .B1(n20242), .B2(n20314), .C1(
        n11601), .C2(n20249), .ZN(P2_U3238) );
  INV_X1 U23265 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20245) );
  OAI222_X1 U23266 ( .A1(n20249), .A2(n20245), .B1(n20244), .B2(n20314), .C1(
        n11601), .C2(n20247), .ZN(P2_U3239) );
  OAI222_X1 U23267 ( .A1(n20249), .A2(n13083), .B1(n20246), .B2(n20314), .C1(
        n20245), .C2(n20247), .ZN(P2_U3240) );
  OAI222_X1 U23268 ( .A1(n20249), .A2(n21234), .B1(n20248), .B2(n20314), .C1(
        n13083), .C2(n20247), .ZN(P2_U3241) );
  OAI22_X1 U23269 ( .A1(n20315), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20314), .ZN(n20250) );
  INV_X1 U23270 ( .A(n20250), .ZN(P2_U3585) );
  MUX2_X1 U23271 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20315), .Z(P2_U3586) );
  OAI22_X1 U23272 ( .A1(n20315), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20314), .ZN(n20251) );
  INV_X1 U23273 ( .A(n20251), .ZN(P2_U3587) );
  OAI22_X1 U23274 ( .A1(n20315), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20314), .ZN(n20252) );
  INV_X1 U23275 ( .A(n20252), .ZN(P2_U3588) );
  OAI21_X1 U23276 ( .B1(n20256), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20254), 
        .ZN(n20253) );
  INV_X1 U23277 ( .A(n20253), .ZN(P2_U3591) );
  OAI21_X1 U23278 ( .B1(n20256), .B2(n20255), .A(n20254), .ZN(P2_U3592) );
  INV_X1 U23279 ( .A(n20296), .ZN(n20299) );
  NOR3_X1 U23280 ( .A1(n20258), .A2(n20261), .A3(n20257), .ZN(n20267) );
  NAND2_X1 U23281 ( .A1(n20259), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20283) );
  NOR2_X1 U23282 ( .A1(n20260), .A2(n20283), .ZN(n20275) );
  INV_X1 U23283 ( .A(n20275), .ZN(n20265) );
  AOI21_X1 U23284 ( .B1(n20284), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20261), 
        .ZN(n20263) );
  NOR2_X1 U23285 ( .A1(n20263), .A2(n20262), .ZN(n20270) );
  AOI21_X1 U23286 ( .B1(n20265), .B2(n20270), .A(n20264), .ZN(n20266) );
  AOI211_X1 U23287 ( .C1(n20268), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20267), 
        .B(n20266), .ZN(n20269) );
  AOI22_X1 U23288 ( .A1(n20299), .A2(n21171), .B1(n20269), .B2(n20296), .ZN(
        P2_U3602) );
  INV_X1 U23289 ( .A(n20270), .ZN(n20274) );
  INV_X1 U23290 ( .A(n20271), .ZN(n20273) );
  AOI22_X1 U23291 ( .A1(n20274), .A2(n20273), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20272), .ZN(n20277) );
  NOR2_X1 U23292 ( .A1(n20299), .A2(n20275), .ZN(n20276) );
  AOI22_X1 U23293 ( .A1(n20278), .A2(n20299), .B1(n20277), .B2(n20276), .ZN(
        P2_U3603) );
  INV_X1 U23294 ( .A(n20279), .ZN(n20291) );
  AND2_X1 U23295 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20280) );
  OR3_X1 U23296 ( .A1(n20281), .A2(n20291), .A3(n20280), .ZN(n20282) );
  OAI21_X1 U23297 ( .B1(n20284), .B2(n20283), .A(n20282), .ZN(n20285) );
  AOI21_X1 U23298 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20286), .A(n20285), 
        .ZN(n20287) );
  AOI22_X1 U23299 ( .A1(n20299), .A2(n20288), .B1(n20287), .B2(n20296), .ZN(
        P2_U3604) );
  INV_X1 U23300 ( .A(n20289), .ZN(n20290) );
  OAI21_X1 U23301 ( .B1(n20292), .B2(n20291), .A(n20290), .ZN(n20293) );
  AOI21_X1 U23302 ( .B1(n20295), .B2(n20294), .A(n20293), .ZN(n20297) );
  AOI22_X1 U23303 ( .A1(n20299), .A2(n20298), .B1(n20297), .B2(n20296), .ZN(
        P2_U3605) );
  INV_X1 U23304 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20300) );
  AOI22_X1 U23305 ( .A1(n20314), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20300), 
        .B2(n20315), .ZN(P2_U3608) );
  INV_X1 U23306 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20313) );
  INV_X1 U23307 ( .A(n20301), .ZN(n20312) );
  INV_X1 U23308 ( .A(n20302), .ZN(n20307) );
  AOI21_X1 U23309 ( .B1(n20305), .B2(n20304), .A(n20303), .ZN(n20306) );
  AOI21_X1 U23310 ( .B1(n20308), .B2(n20307), .A(n20306), .ZN(n20311) );
  NOR2_X1 U23311 ( .A1(n20312), .A2(n20309), .ZN(n20310) );
  AOI22_X1 U23312 ( .A1(n20313), .A2(n20312), .B1(n20311), .B2(n20310), .ZN(
        P2_U3609) );
  OAI22_X1 U23313 ( .A1(n20315), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20314), .ZN(n20316) );
  INV_X1 U23314 ( .A(n20316), .ZN(P2_U3611) );
  INV_X1 U23315 ( .A(n20317), .ZN(n20989) );
  NOR2_X1 U23316 ( .A1(n20989), .A2(n20992), .ZN(n20319) );
  INV_X1 U23317 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20318) );
  NAND2_X2 U23318 ( .A1(n20992), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21056) );
  AOI21_X1 U23319 ( .B1(n20319), .B2(n20318), .A(n21058), .ZN(P1_U2802) );
  NOR2_X1 U23320 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20984) );
  OAI21_X1 U23321 ( .B1(n20984), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21056), .ZN(
        n20320) );
  OAI21_X1 U23322 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21056), .A(n20320), 
        .ZN(P1_U2804) );
  OAI21_X1 U23323 ( .B1(n20992), .B2(n20989), .A(n21056), .ZN(n20979) );
  INV_X1 U23324 ( .A(n20979), .ZN(n21048) );
  OAI21_X1 U23325 ( .B1(BS16), .B2(n20984), .A(n21048), .ZN(n21046) );
  OAI21_X1 U23326 ( .B1(n21048), .B2(n20683), .A(n21046), .ZN(P1_U2805) );
  INV_X1 U23327 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20322) );
  OAI21_X1 U23328 ( .B1(n20323), .B2(n20322), .A(n20321), .ZN(P1_U2806) );
  NOR4_X1 U23329 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20327) );
  NOR4_X1 U23330 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20326) );
  NOR4_X1 U23331 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20325) );
  NOR4_X1 U23332 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20324) );
  NAND4_X1 U23333 ( .A1(n20327), .A2(n20326), .A3(n20325), .A4(n20324), .ZN(
        n20333) );
  NOR4_X1 U23334 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20331) );
  AOI211_X1 U23335 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_28__SCAN_IN), .B(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20330) );
  NOR4_X1 U23336 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20329) );
  NOR4_X1 U23337 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20328) );
  NAND4_X1 U23338 ( .A1(n20331), .A2(n20330), .A3(n20329), .A4(n20328), .ZN(
        n20332) );
  NOR2_X1 U23339 ( .A1(n20333), .A2(n20332), .ZN(n21055) );
  INV_X1 U23340 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20335) );
  NOR3_X1 U23341 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20336) );
  OAI21_X1 U23342 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20336), .A(n21055), .ZN(
        n20334) );
  OAI21_X1 U23343 ( .B1(n21055), .B2(n20335), .A(n20334), .ZN(P1_U2807) );
  INV_X1 U23344 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21047) );
  AOI21_X1 U23345 ( .B1(n20337), .B2(n21047), .A(n20336), .ZN(n20339) );
  INV_X1 U23346 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20338) );
  INV_X1 U23347 ( .A(n21055), .ZN(n21052) );
  AOI22_X1 U23348 ( .A1(n21055), .A2(n20339), .B1(n20338), .B2(n21052), .ZN(
        P1_U2808) );
  NAND2_X1 U23349 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20340), .ZN(n20351) );
  AOI22_X1 U23350 ( .A1(n20342), .A2(n20341), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n20353), .ZN(n20343) );
  OAI211_X1 U23351 ( .C1(n20389), .C2(n20344), .A(n20343), .B(n20379), .ZN(
        n20345) );
  AOI21_X1 U23352 ( .B1(n20377), .B2(n20346), .A(n20345), .ZN(n20350) );
  AOI22_X1 U23353 ( .A1(n20348), .A2(n20368), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20347), .ZN(n20349) );
  OAI211_X1 U23354 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20351), .A(n20350), .B(
        n20349), .ZN(P1_U2831) );
  AOI22_X1 U23355 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20353), .B1(n20377), .B2(
        n20352), .ZN(n20354) );
  OAI21_X1 U23356 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20357), .A(n20354), .ZN(
        n20355) );
  AOI211_X1 U23357 ( .C1(n21395), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21393), .B(n20355), .ZN(n20360) );
  AND2_X1 U23358 ( .A1(n20357), .A2(n20356), .ZN(n20367) );
  AOI22_X1 U23359 ( .A1(n20358), .A2(n20368), .B1(n20367), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n20359) );
  OAI211_X1 U23360 ( .C1(n20361), .C2(n21398), .A(n20360), .B(n20359), .ZN(
        P1_U2833) );
  AOI22_X1 U23361 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20378), .B1(n20363), .B2(
        n20362), .ZN(n20364) );
  OAI21_X1 U23362 ( .B1(n21390), .B2(n20365), .A(n20364), .ZN(n20366) );
  AOI211_X1 U23363 ( .C1(n21395), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21393), .B(n20366), .ZN(n20371) );
  AOI22_X1 U23364 ( .A1(n20369), .A2(n20368), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20367), .ZN(n20370) );
  OAI211_X1 U23365 ( .C1(n20372), .C2(n21398), .A(n20371), .B(n20370), .ZN(
        P1_U2834) );
  NOR2_X1 U23366 ( .A1(n20374), .A2(n20373), .ZN(n20384) );
  NAND2_X1 U23367 ( .A1(n20375), .A2(n20374), .ZN(n20397) );
  NAND2_X1 U23368 ( .A1(n20376), .A2(n20397), .ZN(n20392) );
  AOI22_X1 U23369 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20378), .B1(n20377), .B2(
        n20403), .ZN(n20380) );
  OAI211_X1 U23370 ( .C1(n20389), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        n20382) );
  AOI221_X1 U23371 ( .B1(n20384), .B2(n20383), .C1(n20392), .C2(
        P1_REIP_REG_5__SCAN_IN), .A(n20382), .ZN(n20386) );
  NAND2_X1 U23372 ( .A1(n20406), .A2(n20400), .ZN(n20385) );
  OAI211_X1 U23373 ( .C1(n21398), .C2(n20387), .A(n20386), .B(n20385), .ZN(
        P1_U2835) );
  INV_X1 U23374 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20390) );
  OAI22_X1 U23375 ( .A1(n20390), .A2(n20389), .B1(n20388), .B2(n21391), .ZN(
        n20391) );
  AOI211_X1 U23376 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n20392), .A(n21393), .B(
        n20391), .ZN(n20402) );
  OAI22_X1 U23377 ( .A1(n20395), .A2(n20394), .B1(n21390), .B2(n20393), .ZN(
        n20399) );
  NAND3_X1 U23378 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20396) );
  NOR2_X1 U23379 ( .A1(n20397), .A2(n20396), .ZN(n20398) );
  AOI211_X1 U23380 ( .C1(n20476), .C2(n20400), .A(n20399), .B(n20398), .ZN(
        n20401) );
  OAI211_X1 U23381 ( .C1(n20481), .C2(n21398), .A(n20402), .B(n20401), .ZN(
        P1_U2836) );
  INV_X1 U23382 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21226) );
  AOI22_X1 U23383 ( .A1(n20406), .A2(n20405), .B1(n20404), .B2(n20403), .ZN(
        n20407) );
  OAI21_X1 U23384 ( .B1(n20408), .B2(n21226), .A(n20407), .ZN(P1_U2867) );
  INV_X1 U23385 ( .A(n20409), .ZN(n20410) );
  AOI22_X1 U23386 ( .A1(n20410), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n21067), .ZN(n20411) );
  OAI21_X1 U23387 ( .B1(n20413), .B2(n20412), .A(n20411), .ZN(P1_U2906) );
  AOI22_X1 U23388 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20437), .B1(
        P1_LWORD_REG_15__SCAN_IN), .B2(n20432), .ZN(n20415) );
  OAI21_X1 U23389 ( .B1(n13771), .B2(n20440), .A(n20415), .ZN(P1_U2921) );
  INV_X1 U23390 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20417) );
  AOI22_X1 U23391 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20416) );
  OAI21_X1 U23392 ( .B1(n20417), .B2(n20440), .A(n20416), .ZN(P1_U2922) );
  INV_X1 U23393 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20419) );
  AOI22_X1 U23394 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20418) );
  OAI21_X1 U23395 ( .B1(n20419), .B2(n20440), .A(n20418), .ZN(P1_U2923) );
  INV_X1 U23396 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U23397 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20420) );
  OAI21_X1 U23398 ( .B1(n20421), .B2(n20440), .A(n20420), .ZN(P1_U2924) );
  AOI22_X1 U23399 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20422) );
  OAI21_X1 U23400 ( .B1(n14986), .B2(n20440), .A(n20422), .ZN(P1_U2925) );
  INV_X1 U23401 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20424) );
  AOI22_X1 U23402 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20423) );
  OAI21_X1 U23403 ( .B1(n20424), .B2(n20440), .A(n20423), .ZN(P1_U2926) );
  INV_X1 U23404 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20426) );
  AOI22_X1 U23405 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20425) );
  OAI21_X1 U23406 ( .B1(n20426), .B2(n20440), .A(n20425), .ZN(P1_U2927) );
  AOI22_X1 U23407 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20427) );
  OAI21_X1 U23408 ( .B1(n14394), .B2(n20440), .A(n20427), .ZN(P1_U2928) );
  AOI22_X1 U23409 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20428) );
  OAI21_X1 U23410 ( .B1(n12544), .B2(n20440), .A(n20428), .ZN(P1_U2929) );
  AOI22_X1 U23411 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20429) );
  OAI21_X1 U23412 ( .B1(n20430), .B2(n20440), .A(n20429), .ZN(P1_U2930) );
  AOI22_X1 U23413 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20437), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20432), .ZN(n20431) );
  OAI21_X1 U23414 ( .B1(n14236), .B2(n20440), .A(n20431), .ZN(P1_U2931) );
  AOI22_X1 U23415 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20437), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20432), .ZN(n20433) );
  OAI21_X1 U23416 ( .B1(n20434), .B2(n20440), .A(n20433), .ZN(P1_U2932) );
  AOI22_X1 U23417 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20435) );
  OAI21_X1 U23418 ( .B1(n12511), .B2(n20440), .A(n20435), .ZN(P1_U2933) );
  AOI22_X1 U23419 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20436) );
  OAI21_X1 U23420 ( .B1(n12484), .B2(n20440), .A(n20436), .ZN(P1_U2934) );
  AOI22_X1 U23421 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20438) );
  OAI21_X1 U23422 ( .B1(n12491), .B2(n20440), .A(n20438), .ZN(P1_U2935) );
  AOI22_X1 U23423 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21067), .B1(n20437), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20439) );
  OAI21_X1 U23424 ( .B1(n20441), .B2(n20440), .A(n20439), .ZN(P1_U2936) );
  AOI22_X1 U23425 ( .A1(n20465), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20470), .ZN(n20443) );
  NAND2_X1 U23426 ( .A1(n20455), .A2(n20442), .ZN(n20457) );
  NAND2_X1 U23427 ( .A1(n20443), .A2(n20457), .ZN(P1_U2945) );
  AOI22_X1 U23428 ( .A1(n20465), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20445) );
  NAND2_X1 U23429 ( .A1(n20455), .A2(n20444), .ZN(n20459) );
  NAND2_X1 U23430 ( .A1(n20445), .A2(n20459), .ZN(P1_U2946) );
  AOI22_X1 U23431 ( .A1(n20465), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20447) );
  NAND2_X1 U23432 ( .A1(n20455), .A2(n20446), .ZN(n20461) );
  NAND2_X1 U23433 ( .A1(n20447), .A2(n20461), .ZN(P1_U2947) );
  AOI22_X1 U23434 ( .A1(n20465), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20449) );
  NAND2_X1 U23435 ( .A1(n20455), .A2(n20448), .ZN(n20463) );
  NAND2_X1 U23436 ( .A1(n20449), .A2(n20463), .ZN(P1_U2948) );
  AOI22_X1 U23437 ( .A1(n20465), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20451) );
  NAND2_X1 U23438 ( .A1(n20455), .A2(n20450), .ZN(n20466) );
  NAND2_X1 U23439 ( .A1(n20451), .A2(n20466), .ZN(P1_U2949) );
  AOI22_X1 U23440 ( .A1(n20465), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20453) );
  NAND2_X1 U23441 ( .A1(n20455), .A2(n20452), .ZN(n20468) );
  NAND2_X1 U23442 ( .A1(n20453), .A2(n20468), .ZN(P1_U2950) );
  AOI22_X1 U23443 ( .A1(n20465), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20470), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20456) );
  NAND2_X1 U23444 ( .A1(n20455), .A2(n20454), .ZN(n20471) );
  NAND2_X1 U23445 ( .A1(n20456), .A2(n20471), .ZN(P1_U2951) );
  AOI22_X1 U23446 ( .A1(n20465), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20458) );
  NAND2_X1 U23447 ( .A1(n20458), .A2(n20457), .ZN(P1_U2960) );
  AOI22_X1 U23448 ( .A1(n20465), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20470), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20460) );
  NAND2_X1 U23449 ( .A1(n20460), .A2(n20459), .ZN(P1_U2961) );
  AOI22_X1 U23450 ( .A1(n20465), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20470), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20462) );
  NAND2_X1 U23451 ( .A1(n20462), .A2(n20461), .ZN(P1_U2962) );
  AOI22_X1 U23452 ( .A1(n20465), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20470), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20464) );
  NAND2_X1 U23453 ( .A1(n20464), .A2(n20463), .ZN(P1_U2963) );
  AOI22_X1 U23454 ( .A1(n20465), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20470), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20467) );
  NAND2_X1 U23455 ( .A1(n20467), .A2(n20466), .ZN(P1_U2964) );
  AOI22_X1 U23456 ( .A1(n20465), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20470), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20469) );
  NAND2_X1 U23457 ( .A1(n20469), .A2(n20468), .ZN(P1_U2965) );
  AOI22_X1 U23458 ( .A1(n20465), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20470), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20472) );
  NAND2_X1 U23459 ( .A1(n20472), .A2(n20471), .ZN(P1_U2966) );
  AOI22_X1 U23460 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20480) );
  INV_X1 U23461 ( .A(n20475), .ZN(n20478) );
  AOI22_X1 U23462 ( .A1(n20478), .A2(n12479), .B1(n20477), .B2(n20476), .ZN(
        n20479) );
  OAI211_X1 U23463 ( .C1(n20482), .C2(n20481), .A(n20480), .B(n20479), .ZN(
        P1_U2995) );
  INV_X1 U23464 ( .A(n20483), .ZN(n20484) );
  AOI21_X1 U23465 ( .B1(n20486), .B2(n20485), .A(n20484), .ZN(n20491) );
  INV_X1 U23466 ( .A(n20487), .ZN(n20489) );
  AOI22_X1 U23467 ( .A1(n20489), .A2(n20507), .B1(n20488), .B2(n12159), .ZN(
        n20490) );
  OAI211_X1 U23468 ( .C1(n20492), .C2(n12159), .A(n20491), .B(n20490), .ZN(
        P1_U3028) );
  NAND2_X1 U23469 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20493), .ZN(
        n20512) );
  OAI21_X1 U23470 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20495), .A(
        n20494), .ZN(n20496) );
  INV_X1 U23471 ( .A(n20496), .ZN(n20510) );
  INV_X1 U23472 ( .A(n20497), .ZN(n20508) );
  NOR2_X1 U23473 ( .A1(n13613), .A2(n20498), .ZN(n20500) );
  AOI21_X1 U23474 ( .B1(n20500), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20499), .ZN(n20501) );
  NOR2_X1 U23475 ( .A1(n20502), .A2(n20501), .ZN(n20506) );
  INV_X1 U23476 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21001) );
  OAI22_X1 U23477 ( .A1(n20504), .A2(n20503), .B1(n21001), .B2(n12460), .ZN(
        n20505) );
  AOI211_X1 U23478 ( .C1(n20508), .C2(n20507), .A(n20506), .B(n20505), .ZN(
        n20509) );
  OAI221_X1 U23479 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20512), .C1(
        n20511), .C2(n20510), .A(n20509), .ZN(P1_U3029) );
  NOR2_X1 U23480 ( .A1(n20514), .A2(n20513), .ZN(P1_U3032) );
  NAND2_X1 U23481 ( .A1(n20517), .A2(n20911), .ZN(n20518) );
  NOR2_X1 U23482 ( .A1(n20915), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20863) );
  INV_X1 U23483 ( .A(n20863), .ZN(n20576) );
  OAI21_X1 U23484 ( .B1(n20570), .B2(n20518), .A(n20576), .ZN(n20525) );
  OR2_X1 U23485 ( .A1(n9749), .A2(n20519), .ZN(n20617) );
  NOR2_X1 U23486 ( .A1(n20617), .A2(n20865), .ZN(n20521) );
  INV_X1 U23487 ( .A(n20741), .ZN(n20520) );
  NOR2_X1 U23488 ( .A1(n20520), .A2(n20742), .ZN(n20654) );
  NOR3_X1 U23489 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20553) );
  INV_X1 U23490 ( .A(n20553), .ZN(n20550) );
  NOR2_X1 U23491 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20550), .ZN(
        n20541) );
  AOI22_X1 U23492 ( .A1(n20542), .A2(n9852), .B1(n20918), .B2(n20541), .ZN(
        n20528) );
  INV_X1 U23493 ( .A(n20521), .ZN(n20524) );
  NAND2_X1 U23494 ( .A1(n20522), .A2(n20656), .ZN(n20747) );
  OAI22_X1 U23495 ( .A1(n20913), .A2(n20654), .B1(n20817), .B2(n20541), .ZN(
        n20523) );
  AOI211_X1 U23496 ( .C1(n20525), .C2(n20524), .A(n20747), .B(n20523), .ZN(
        n20526) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20919), .ZN(n20527) );
  OAI211_X1 U23498 ( .C1(n20546), .C2(n20879), .A(n20528), .B(n20527), .ZN(
        P1_U3033) );
  AOI22_X1 U23499 ( .A1(n20542), .A2(n9858), .B1(n20924), .B2(n20541), .ZN(
        n20530) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20925), .ZN(n20529) );
  OAI211_X1 U23501 ( .C1(n20546), .C2(n20882), .A(n20530), .B(n20529), .ZN(
        P1_U3034) );
  AOI22_X1 U23502 ( .A1(n20542), .A2(n9854), .B1(n20931), .B2(n20541), .ZN(
        n20532) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20932), .ZN(n20531) );
  OAI211_X1 U23504 ( .C1(n20546), .C2(n20885), .A(n20532), .B(n20531), .ZN(
        P1_U3035) );
  AOI22_X1 U23505 ( .A1(n20542), .A2(n20940), .B1(n20938), .B2(n20541), .ZN(
        n20534) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20939), .ZN(n20533) );
  OAI211_X1 U23507 ( .C1(n20546), .C2(n20888), .A(n20534), .B(n20533), .ZN(
        P1_U3036) );
  AOI22_X1 U23508 ( .A1(n20542), .A2(n20947), .B1(n20945), .B2(n20541), .ZN(
        n20536) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20946), .ZN(n20535) );
  OAI211_X1 U23510 ( .C1(n20546), .C2(n20891), .A(n20536), .B(n20535), .ZN(
        P1_U3037) );
  AOI22_X1 U23511 ( .A1(n20542), .A2(n20954), .B1(n20952), .B2(n20541), .ZN(
        n20538) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20953), .ZN(n20537) );
  OAI211_X1 U23513 ( .C1(n20546), .C2(n20894), .A(n20538), .B(n20537), .ZN(
        P1_U3038) );
  AOI22_X1 U23514 ( .A1(n20542), .A2(n9860), .B1(n20959), .B2(n20541), .ZN(
        n20540) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20960), .ZN(n20539) );
  OAI211_X1 U23516 ( .C1(n20546), .C2(n20897), .A(n20540), .B(n20539), .ZN(
        P1_U3039) );
  AOI22_X1 U23517 ( .A1(n20542), .A2(n9856), .B1(n20968), .B2(n20541), .ZN(
        n20545) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20543), .B1(
        n20570), .B2(n20969), .ZN(n20544) );
  OAI211_X1 U23519 ( .C1(n20546), .C2(n20903), .A(n20545), .B(n20544), .ZN(
        P1_U3040) );
  NOR2_X1 U23520 ( .A1(n20905), .A2(n20550), .ZN(n20569) );
  INV_X1 U23521 ( .A(n20617), .ZN(n20549) );
  INV_X1 U23522 ( .A(n20548), .ZN(n20906) );
  AOI21_X1 U23523 ( .B1(n20549), .B2(n20906), .A(n20569), .ZN(n20551) );
  OAI22_X1 U23524 ( .A1(n20551), .A2(n20915), .B1(n20550), .B2(n20913), .ZN(
        n20568) );
  AOI22_X1 U23525 ( .A1(n20918), .A2(n20569), .B1(n20568), .B2(n20917), .ZN(
        n20555) );
  OAI211_X1 U23526 ( .C1(n20615), .C2(n20779), .A(n20911), .B(n20551), .ZN(
        n20552) );
  OAI211_X1 U23527 ( .C1(n20911), .C2(n20553), .A(n20781), .B(n20552), .ZN(
        n20571) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n9852), .ZN(n20554) );
  OAI211_X1 U23529 ( .C1(n20751), .C2(n20607), .A(n20555), .B(n20554), .ZN(
        P1_U3041) );
  AOI22_X1 U23530 ( .A1(n20924), .A2(n20569), .B1(n20568), .B2(n20923), .ZN(
        n20557) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n9858), .ZN(n20556) );
  OAI211_X1 U23532 ( .C1(n20754), .C2(n20607), .A(n20557), .B(n20556), .ZN(
        P1_U3042) );
  AOI22_X1 U23533 ( .A1(n20931), .A2(n20569), .B1(n20568), .B2(n20930), .ZN(
        n20559) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n9854), .ZN(n20558) );
  OAI211_X1 U23535 ( .C1(n20757), .C2(n20607), .A(n20559), .B(n20558), .ZN(
        P1_U3043) );
  AOI22_X1 U23536 ( .A1(n20938), .A2(n20569), .B1(n20568), .B2(n20937), .ZN(
        n20561) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20940), .ZN(n20560) );
  OAI211_X1 U23538 ( .C1(n20760), .C2(n20607), .A(n20561), .B(n20560), .ZN(
        P1_U3044) );
  AOI22_X1 U23539 ( .A1(n20945), .A2(n20569), .B1(n20568), .B2(n20944), .ZN(
        n20563) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20947), .ZN(n20562) );
  OAI211_X1 U23541 ( .C1(n20763), .C2(n20607), .A(n20563), .B(n20562), .ZN(
        P1_U3045) );
  AOI22_X1 U23542 ( .A1(n20952), .A2(n20569), .B1(n20568), .B2(n20951), .ZN(
        n20565) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20954), .ZN(n20564) );
  OAI211_X1 U23544 ( .C1(n20766), .C2(n20607), .A(n20565), .B(n20564), .ZN(
        P1_U3046) );
  AOI22_X1 U23545 ( .A1(n20959), .A2(n20569), .B1(n20568), .B2(n20958), .ZN(
        n20567) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n9860), .ZN(n20566) );
  OAI211_X1 U23547 ( .C1(n20769), .C2(n20607), .A(n20567), .B(n20566), .ZN(
        P1_U3047) );
  AOI22_X1 U23548 ( .A1(n20968), .A2(n20569), .B1(n20568), .B2(n20966), .ZN(
        n20573) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n9856), .ZN(n20572) );
  OAI211_X1 U23550 ( .C1(n20776), .C2(n20607), .A(n20573), .B(n20572), .ZN(
        P1_U3048) );
  INV_X1 U23551 ( .A(n20645), .ZN(n20575) );
  NAND3_X1 U23552 ( .A1(n20575), .A2(n20911), .A3(n20607), .ZN(n20577) );
  NAND2_X1 U23553 ( .A1(n20577), .A2(n20576), .ZN(n20581) );
  OR2_X1 U23554 ( .A1(n20617), .A2(n14172), .ZN(n20580) );
  INV_X1 U23555 ( .A(n20580), .ZN(n20578) );
  NAND3_X1 U23556 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20740), .A3(
        n20653), .ZN(n20626) );
  NOR2_X1 U23557 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20626), .ZN(
        n20585) );
  INV_X1 U23558 ( .A(n20585), .ZN(n20606) );
  OAI22_X1 U23559 ( .A1(n20607), .A2(n9851), .B1(n20812), .B2(n20606), .ZN(
        n20579) );
  INV_X1 U23560 ( .A(n20579), .ZN(n20587) );
  NAND2_X1 U23561 ( .A1(n20581), .A2(n20580), .ZN(n20584) );
  NOR2_X1 U23562 ( .A1(n10262), .A2(n20582), .ZN(n20712) );
  NOR2_X1 U23563 ( .A1(n20712), .A2(n20747), .ZN(n20583) );
  AOI22_X1 U23564 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n20919), .B2(n20645), .ZN(n20586) );
  OAI211_X1 U23565 ( .C1(n20612), .C2(n20879), .A(n20587), .B(n20586), .ZN(
        P1_U3049) );
  OAI22_X1 U23566 ( .A1(n20607), .A2(n9857), .B1(n20824), .B2(n20606), .ZN(
        n20588) );
  INV_X1 U23567 ( .A(n20588), .ZN(n20590) );
  AOI22_X1 U23568 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n20925), .B2(n20645), .ZN(n20589) );
  OAI211_X1 U23569 ( .C1(n20612), .C2(n20882), .A(n20590), .B(n20589), .ZN(
        P1_U3050) );
  OAI22_X1 U23570 ( .A1(n20607), .A2(n9853), .B1(n20828), .B2(n20606), .ZN(
        n20591) );
  INV_X1 U23571 ( .A(n20591), .ZN(n20593) );
  AOI22_X1 U23572 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n20932), .B2(n20645), .ZN(n20592) );
  OAI211_X1 U23573 ( .C1(n20612), .C2(n20885), .A(n20593), .B(n20592), .ZN(
        P1_U3051) );
  OAI22_X1 U23574 ( .A1(n20607), .A2(n20833), .B1(n20832), .B2(n20606), .ZN(
        n20594) );
  INV_X1 U23575 ( .A(n20594), .ZN(n20596) );
  AOI22_X1 U23576 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n20939), .B2(n20645), .ZN(n20595) );
  OAI211_X1 U23577 ( .C1(n20612), .C2(n20888), .A(n20596), .B(n20595), .ZN(
        P1_U3052) );
  OAI22_X1 U23578 ( .A1(n20607), .A2(n20838), .B1(n20837), .B2(n20606), .ZN(
        n20597) );
  INV_X1 U23579 ( .A(n20597), .ZN(n20599) );
  AOI22_X1 U23580 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n20946), .B2(n20645), .ZN(n20598) );
  OAI211_X1 U23581 ( .C1(n20612), .C2(n20891), .A(n20599), .B(n20598), .ZN(
        P1_U3053) );
  OAI22_X1 U23582 ( .A1(n20607), .A2(n20843), .B1(n20842), .B2(n20606), .ZN(
        n20600) );
  INV_X1 U23583 ( .A(n20600), .ZN(n20602) );
  AOI22_X1 U23584 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n20953), .B2(n20645), .ZN(n20601) );
  OAI211_X1 U23585 ( .C1(n20612), .C2(n20894), .A(n20602), .B(n20601), .ZN(
        P1_U3054) );
  OAI22_X1 U23586 ( .A1(n20607), .A2(n9859), .B1(n20847), .B2(n20606), .ZN(
        n20603) );
  INV_X1 U23587 ( .A(n20603), .ZN(n20605) );
  AOI22_X1 U23588 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n20960), .B2(n20645), .ZN(n20604) );
  OAI211_X1 U23589 ( .C1(n20612), .C2(n20897), .A(n20605), .B(n20604), .ZN(
        P1_U3055) );
  OAI22_X1 U23590 ( .A1(n20607), .A2(n9855), .B1(n20852), .B2(n20606), .ZN(
        n20608) );
  INV_X1 U23591 ( .A(n20608), .ZN(n20611) );
  AOI22_X1 U23592 ( .A1(n20609), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9850), .B2(n20645), .ZN(n20610) );
  OAI211_X1 U23593 ( .C1(n20612), .C2(n20903), .A(n20611), .B(n20610), .ZN(
        P1_U3056) );
  INV_X1 U23594 ( .A(n20613), .ZN(n20614) );
  AOI21_X1 U23595 ( .B1(n20615), .B2(n20911), .A(n20614), .ZN(n20629) );
  OR2_X1 U23596 ( .A1(n20617), .A2(n20616), .ZN(n20620) );
  INV_X1 U23597 ( .A(n20618), .ZN(n20619) );
  NAND2_X1 U23598 ( .A1(n20619), .A2(n20740), .ZN(n20624) );
  OAI22_X1 U23599 ( .A1(n20913), .A2(n20626), .B1(n20629), .B2(n20625), .ZN(
        n20621) );
  INV_X1 U23600 ( .A(n20624), .ZN(n20644) );
  AOI22_X1 U23601 ( .A1(n20677), .A2(n20919), .B1(n20918), .B2(n20644), .ZN(
        n20631) );
  INV_X1 U23602 ( .A(n20625), .ZN(n20628) );
  AOI21_X1 U23603 ( .B1(n20915), .B2(n20626), .A(n20910), .ZN(n20627) );
  OAI21_X1 U23604 ( .B1(n20629), .B2(n20628), .A(n20627), .ZN(n20646) );
  AOI22_X1 U23605 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9852), .B2(n20645), .ZN(n20630) );
  OAI211_X1 U23606 ( .C1(n20649), .C2(n20879), .A(n20631), .B(n20630), .ZN(
        P1_U3057) );
  AOI22_X1 U23607 ( .A1(n20645), .A2(n9858), .B1(n20924), .B2(n20644), .ZN(
        n20633) );
  AOI22_X1 U23608 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n20925), .B2(n20677), .ZN(n20632) );
  OAI211_X1 U23609 ( .C1(n20649), .C2(n20882), .A(n20633), .B(n20632), .ZN(
        P1_U3058) );
  AOI22_X1 U23610 ( .A1(n20677), .A2(n20932), .B1(n20931), .B2(n20644), .ZN(
        n20635) );
  AOI22_X1 U23611 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9854), .B2(n20645), .ZN(n20634) );
  OAI211_X1 U23612 ( .C1(n20649), .C2(n20885), .A(n20635), .B(n20634), .ZN(
        P1_U3059) );
  AOI22_X1 U23613 ( .A1(n20677), .A2(n20939), .B1(n20938), .B2(n20644), .ZN(
        n20637) );
  AOI22_X1 U23614 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n20940), .B2(n20645), .ZN(n20636) );
  OAI211_X1 U23615 ( .C1(n20649), .C2(n20888), .A(n20637), .B(n20636), .ZN(
        P1_U3060) );
  AOI22_X1 U23616 ( .A1(n20645), .A2(n20947), .B1(n20945), .B2(n20644), .ZN(
        n20639) );
  AOI22_X1 U23617 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n20946), .B2(n20677), .ZN(n20638) );
  OAI211_X1 U23618 ( .C1(n20649), .C2(n20891), .A(n20639), .B(n20638), .ZN(
        P1_U3061) );
  AOI22_X1 U23619 ( .A1(n20645), .A2(n20954), .B1(n20952), .B2(n20644), .ZN(
        n20641) );
  AOI22_X1 U23620 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n20953), .B2(n20677), .ZN(n20640) );
  OAI211_X1 U23621 ( .C1(n20649), .C2(n20894), .A(n20641), .B(n20640), .ZN(
        P1_U3062) );
  AOI22_X1 U23622 ( .A1(n20645), .A2(n9860), .B1(n20959), .B2(n20644), .ZN(
        n20643) );
  AOI22_X1 U23623 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n20960), .B2(n20677), .ZN(n20642) );
  OAI211_X1 U23624 ( .C1(n20649), .C2(n20897), .A(n20643), .B(n20642), .ZN(
        P1_U3063) );
  AOI22_X1 U23625 ( .A1(n20645), .A2(n9856), .B1(n20968), .B2(n20644), .ZN(
        n20648) );
  AOI22_X1 U23626 ( .A1(n20646), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9850), .B2(n20677), .ZN(n20647) );
  OAI211_X1 U23627 ( .C1(n20649), .C2(n20903), .A(n20648), .B(n20647), .ZN(
        P1_U3064) );
  NOR2_X1 U23628 ( .A1(n9897), .A2(n20650), .ZN(n20651) );
  NOR3_X1 U23629 ( .A1(n20653), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20686) );
  INV_X1 U23630 ( .A(n20686), .ZN(n20681) );
  NOR2_X1 U23631 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20681), .ZN(
        n20676) );
  NAND2_X1 U23632 ( .A1(n20709), .A2(n14172), .ZN(n20658) );
  INV_X1 U23633 ( .A(n20654), .ZN(n20655) );
  OAI22_X1 U23634 ( .A1(n20658), .A2(n20915), .B1(n20656), .B2(n20655), .ZN(
        n20675) );
  AOI22_X1 U23635 ( .A1(n20918), .A2(n20676), .B1(n20917), .B2(n20675), .ZN(
        n20662) );
  INV_X1 U23636 ( .A(n20707), .ZN(n20657) );
  OAI21_X1 U23637 ( .B1(n20677), .B2(n20657), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20659) );
  AOI21_X1 U23638 ( .B1(n20659), .B2(n20658), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20660) );
  AOI22_X1 U23639 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9852), .B2(n20677), .ZN(n20661) );
  OAI211_X1 U23640 ( .C1(n20751), .C2(n20707), .A(n20662), .B(n20661), .ZN(
        P1_U3065) );
  AOI22_X1 U23641 ( .A1(n20924), .A2(n20676), .B1(n20923), .B2(n20675), .ZN(
        n20664) );
  AOI22_X1 U23642 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9858), .B2(n20677), .ZN(n20663) );
  OAI211_X1 U23643 ( .C1(n20754), .C2(n20707), .A(n20664), .B(n20663), .ZN(
        P1_U3066) );
  AOI22_X1 U23644 ( .A1(n20931), .A2(n20676), .B1(n20930), .B2(n20675), .ZN(
        n20666) );
  AOI22_X1 U23645 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9854), .B2(n20677), .ZN(n20665) );
  OAI211_X1 U23646 ( .C1(n20757), .C2(n20707), .A(n20666), .B(n20665), .ZN(
        P1_U3067) );
  AOI22_X1 U23647 ( .A1(n20938), .A2(n20676), .B1(n20937), .B2(n20675), .ZN(
        n20668) );
  AOI22_X1 U23648 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n20940), .B2(n20677), .ZN(n20667) );
  OAI211_X1 U23649 ( .C1(n20760), .C2(n20707), .A(n20668), .B(n20667), .ZN(
        P1_U3068) );
  AOI22_X1 U23650 ( .A1(n20945), .A2(n20676), .B1(n20944), .B2(n20675), .ZN(
        n20670) );
  AOI22_X1 U23651 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n20947), .B2(n20677), .ZN(n20669) );
  OAI211_X1 U23652 ( .C1(n20763), .C2(n20707), .A(n20670), .B(n20669), .ZN(
        P1_U3069) );
  AOI22_X1 U23653 ( .A1(n20952), .A2(n20676), .B1(n20951), .B2(n20675), .ZN(
        n20672) );
  AOI22_X1 U23654 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n20954), .B2(n20677), .ZN(n20671) );
  OAI211_X1 U23655 ( .C1(n20766), .C2(n20707), .A(n20672), .B(n20671), .ZN(
        P1_U3070) );
  AOI22_X1 U23656 ( .A1(n20959), .A2(n20676), .B1(n20958), .B2(n20675), .ZN(
        n20674) );
  AOI22_X1 U23657 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9860), .B2(n20677), .ZN(n20673) );
  OAI211_X1 U23658 ( .C1(n20769), .C2(n20707), .A(n20674), .B(n20673), .ZN(
        P1_U3071) );
  AOI22_X1 U23659 ( .A1(n20968), .A2(n20676), .B1(n20966), .B2(n20675), .ZN(
        n20680) );
  AOI22_X1 U23660 ( .A1(n20678), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9856), .B2(n20677), .ZN(n20679) );
  OAI211_X1 U23661 ( .C1(n20776), .C2(n20707), .A(n20680), .B(n20679), .ZN(
        P1_U3072) );
  NOR2_X1 U23662 ( .A1(n20905), .A2(n20681), .ZN(n20703) );
  AOI21_X1 U23663 ( .B1(n20709), .B2(n20906), .A(n20703), .ZN(n20682) );
  OAI22_X1 U23664 ( .A1(n20682), .A2(n20915), .B1(n20681), .B2(n20913), .ZN(
        n20702) );
  AOI22_X1 U23665 ( .A1(n20918), .A2(n20703), .B1(n20917), .B2(n20702), .ZN(
        n20689) );
  INV_X1 U23666 ( .A(n20687), .ZN(n20684) );
  NOR3_X1 U23667 ( .A1(n20684), .A2(n20915), .A3(n20683), .ZN(n20685) );
  OAI21_X1 U23668 ( .B1(n20686), .B2(n20685), .A(n20781), .ZN(n20704) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20919), .ZN(n20688) );
  OAI211_X1 U23670 ( .C1(n9851), .C2(n20707), .A(n20689), .B(n20688), .ZN(
        P1_U3073) );
  AOI22_X1 U23671 ( .A1(n20924), .A2(n20703), .B1(n20923), .B2(n20702), .ZN(
        n20691) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20925), .ZN(n20690) );
  OAI211_X1 U23673 ( .C1(n9857), .C2(n20707), .A(n20691), .B(n20690), .ZN(
        P1_U3074) );
  AOI22_X1 U23674 ( .A1(n20931), .A2(n20703), .B1(n20930), .B2(n20702), .ZN(
        n20693) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20932), .ZN(n20692) );
  OAI211_X1 U23676 ( .C1(n9853), .C2(n20707), .A(n20693), .B(n20692), .ZN(
        P1_U3075) );
  AOI22_X1 U23677 ( .A1(n20938), .A2(n20703), .B1(n20937), .B2(n20702), .ZN(
        n20695) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20939), .ZN(n20694) );
  OAI211_X1 U23679 ( .C1(n20833), .C2(n20707), .A(n20695), .B(n20694), .ZN(
        P1_U3076) );
  AOI22_X1 U23680 ( .A1(n20945), .A2(n20703), .B1(n20944), .B2(n20702), .ZN(
        n20697) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20946), .ZN(n20696) );
  OAI211_X1 U23682 ( .C1(n20838), .C2(n20707), .A(n20697), .B(n20696), .ZN(
        P1_U3077) );
  AOI22_X1 U23683 ( .A1(n20952), .A2(n20703), .B1(n20951), .B2(n20702), .ZN(
        n20699) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20953), .ZN(n20698) );
  OAI211_X1 U23685 ( .C1(n20843), .C2(n20707), .A(n20699), .B(n20698), .ZN(
        P1_U3078) );
  AOI22_X1 U23686 ( .A1(n20959), .A2(n20703), .B1(n20958), .B2(n20702), .ZN(
        n20701) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n20960), .ZN(n20700) );
  OAI211_X1 U23688 ( .C1(n9859), .C2(n20707), .A(n20701), .B(n20700), .ZN(
        P1_U3079) );
  AOI22_X1 U23689 ( .A1(n20968), .A2(n20703), .B1(n20966), .B2(n20702), .ZN(
        n20706) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20704), .B1(
        n20732), .B2(n9850), .ZN(n20705) );
  OAI211_X1 U23691 ( .C1(n9855), .C2(n20707), .A(n20706), .B(n20705), .ZN(
        P1_U3080) );
  NOR3_X1 U23692 ( .A1(n20732), .A2(n20733), .A3(n20915), .ZN(n20708) );
  NOR2_X1 U23693 ( .A1(n20708), .A2(n20863), .ZN(n20716) );
  INV_X1 U23694 ( .A(n20716), .ZN(n20710) );
  AND2_X1 U23695 ( .A1(n20709), .A2(n20865), .ZN(n20715) );
  NOR2_X1 U23696 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20711), .ZN(
        n20731) );
  AOI22_X1 U23697 ( .A1(n20732), .A2(n9852), .B1(n20918), .B2(n20731), .ZN(
        n20718) );
  INV_X1 U23698 ( .A(n20731), .ZN(n20713) );
  AOI21_X1 U23699 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20713), .A(n20712), 
        .ZN(n20714) );
  OAI211_X1 U23700 ( .C1(n20716), .C2(n20715), .A(n20874), .B(n20714), .ZN(
        n20734) );
  AOI22_X1 U23701 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20919), .B2(n20733), .ZN(n20717) );
  OAI211_X1 U23702 ( .C1(n20737), .C2(n20879), .A(n20718), .B(n20717), .ZN(
        P1_U3081) );
  AOI22_X1 U23703 ( .A1(n20732), .A2(n9858), .B1(n20924), .B2(n20731), .ZN(
        n20720) );
  AOI22_X1 U23704 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20925), .B2(n20733), .ZN(n20719) );
  OAI211_X1 U23705 ( .C1(n20737), .C2(n20882), .A(n20720), .B(n20719), .ZN(
        P1_U3082) );
  AOI22_X1 U23706 ( .A1(n20732), .A2(n9854), .B1(n20931), .B2(n20731), .ZN(
        n20722) );
  AOI22_X1 U23707 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n20932), .B2(n20733), .ZN(n20721) );
  OAI211_X1 U23708 ( .C1(n20737), .C2(n20885), .A(n20722), .B(n20721), .ZN(
        P1_U3083) );
  AOI22_X1 U23709 ( .A1(n20732), .A2(n20940), .B1(n20938), .B2(n20731), .ZN(
        n20724) );
  AOI22_X1 U23710 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20939), .B2(n20733), .ZN(n20723) );
  OAI211_X1 U23711 ( .C1(n20737), .C2(n20888), .A(n20724), .B(n20723), .ZN(
        P1_U3084) );
  AOI22_X1 U23712 ( .A1(n20732), .A2(n20947), .B1(n20945), .B2(n20731), .ZN(
        n20726) );
  AOI22_X1 U23713 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20946), .B2(n20733), .ZN(n20725) );
  OAI211_X1 U23714 ( .C1(n20737), .C2(n20891), .A(n20726), .B(n20725), .ZN(
        P1_U3085) );
  AOI22_X1 U23715 ( .A1(n20732), .A2(n20954), .B1(n20952), .B2(n20731), .ZN(
        n20728) );
  AOI22_X1 U23716 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n20953), .B2(n20733), .ZN(n20727) );
  OAI211_X1 U23717 ( .C1(n20737), .C2(n20894), .A(n20728), .B(n20727), .ZN(
        P1_U3086) );
  AOI22_X1 U23718 ( .A1(n20732), .A2(n9860), .B1(n20959), .B2(n20731), .ZN(
        n20730) );
  AOI22_X1 U23719 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n20960), .B2(n20733), .ZN(n20729) );
  OAI211_X1 U23720 ( .C1(n20737), .C2(n20897), .A(n20730), .B(n20729), .ZN(
        P1_U3087) );
  AOI22_X1 U23721 ( .A1(n20732), .A2(n9856), .B1(n20968), .B2(n20731), .ZN(
        n20736) );
  AOI22_X1 U23722 ( .A1(n20734), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9850), .B2(n20733), .ZN(n20735) );
  OAI211_X1 U23723 ( .C1(n20737), .C2(n20903), .A(n20736), .B(n20735), .ZN(
        P1_U3088) );
  INV_X1 U23724 ( .A(n20738), .ZN(n20861) );
  NOR3_X1 U23725 ( .A1(n20740), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20782) );
  INV_X1 U23726 ( .A(n20782), .ZN(n20777) );
  NOR2_X1 U23727 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20777), .ZN(
        n20771) );
  AOI21_X1 U23728 ( .B1(n20807), .B2(n14172), .A(n20771), .ZN(n20745) );
  NAND2_X1 U23729 ( .A1(n20742), .A2(n20741), .ZN(n20872) );
  INV_X1 U23730 ( .A(n20808), .ZN(n20743) );
  OAI22_X1 U23731 ( .A1(n20745), .A2(n20915), .B1(n20872), .B2(n20743), .ZN(
        n20770) );
  AOI22_X1 U23732 ( .A1(n20918), .A2(n20771), .B1(n20770), .B2(n20917), .ZN(
        n20750) );
  INV_X1 U23733 ( .A(n20804), .ZN(n20744) );
  OAI21_X1 U23734 ( .B1(n20744), .B2(n20772), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20746) );
  NAND2_X1 U23735 ( .A1(n20746), .A2(n20745), .ZN(n20748) );
  INV_X1 U23736 ( .A(n20747), .ZN(n20814) );
  AOI22_X1 U23737 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9852), .B2(n20772), .ZN(n20749) );
  OAI211_X1 U23738 ( .C1(n20751), .C2(n20804), .A(n20750), .B(n20749), .ZN(
        P1_U3097) );
  AOI22_X1 U23739 ( .A1(n20924), .A2(n20771), .B1(n20770), .B2(n20923), .ZN(
        n20753) );
  AOI22_X1 U23740 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9858), .B2(n20772), .ZN(n20752) );
  OAI211_X1 U23741 ( .C1(n20754), .C2(n20804), .A(n20753), .B(n20752), .ZN(
        P1_U3098) );
  AOI22_X1 U23742 ( .A1(n20931), .A2(n20771), .B1(n20770), .B2(n20930), .ZN(
        n20756) );
  AOI22_X1 U23743 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9854), .B2(n20772), .ZN(n20755) );
  OAI211_X1 U23744 ( .C1(n20757), .C2(n20804), .A(n20756), .B(n20755), .ZN(
        P1_U3099) );
  AOI22_X1 U23745 ( .A1(n20938), .A2(n20771), .B1(n20770), .B2(n20937), .ZN(
        n20759) );
  AOI22_X1 U23746 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20940), .B2(n20772), .ZN(n20758) );
  OAI211_X1 U23747 ( .C1(n20760), .C2(n20804), .A(n20759), .B(n20758), .ZN(
        P1_U3100) );
  AOI22_X1 U23748 ( .A1(n20945), .A2(n20771), .B1(n20770), .B2(n20944), .ZN(
        n20762) );
  AOI22_X1 U23749 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20947), .B2(n20772), .ZN(n20761) );
  OAI211_X1 U23750 ( .C1(n20763), .C2(n20804), .A(n20762), .B(n20761), .ZN(
        P1_U3101) );
  AOI22_X1 U23751 ( .A1(n20952), .A2(n20771), .B1(n20770), .B2(n20951), .ZN(
        n20765) );
  AOI22_X1 U23752 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20954), .B2(n20772), .ZN(n20764) );
  OAI211_X1 U23753 ( .C1(n20766), .C2(n20804), .A(n20765), .B(n20764), .ZN(
        P1_U3102) );
  AOI22_X1 U23754 ( .A1(n20959), .A2(n20771), .B1(n20770), .B2(n20958), .ZN(
        n20768) );
  AOI22_X1 U23755 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9860), .B2(n20772), .ZN(n20767) );
  OAI211_X1 U23756 ( .C1(n20769), .C2(n20804), .A(n20768), .B(n20767), .ZN(
        P1_U3103) );
  AOI22_X1 U23757 ( .A1(n20968), .A2(n20771), .B1(n20770), .B2(n20966), .ZN(
        n20775) );
  AOI22_X1 U23758 ( .A1(n20773), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9856), .B2(n20772), .ZN(n20774) );
  OAI211_X1 U23759 ( .C1(n20776), .C2(n20804), .A(n20775), .B(n20774), .ZN(
        P1_U3104) );
  NOR2_X1 U23760 ( .A1(n20905), .A2(n20777), .ZN(n20800) );
  AOI21_X1 U23761 ( .B1(n20807), .B2(n20906), .A(n20800), .ZN(n20778) );
  OAI22_X1 U23762 ( .A1(n20778), .A2(n20915), .B1(n20777), .B2(n20913), .ZN(
        n20799) );
  AOI22_X1 U23763 ( .A1(n20918), .A2(n20800), .B1(n20799), .B2(n20917), .ZN(
        n20786) );
  OAI211_X1 U23764 ( .C1(n20784), .C2(n20779), .A(n20911), .B(n20778), .ZN(
        n20780) );
  OAI211_X1 U23765 ( .C1(n20911), .C2(n20782), .A(n20781), .B(n20780), .ZN(
        n20801) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20919), .ZN(n20785) );
  OAI211_X1 U23767 ( .C1(n9851), .C2(n20804), .A(n20786), .B(n20785), .ZN(
        P1_U3105) );
  AOI22_X1 U23768 ( .A1(n20924), .A2(n20800), .B1(n20799), .B2(n20923), .ZN(
        n20788) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20925), .ZN(n20787) );
  OAI211_X1 U23770 ( .C1(n9857), .C2(n20804), .A(n20788), .B(n20787), .ZN(
        P1_U3106) );
  AOI22_X1 U23771 ( .A1(n20931), .A2(n20800), .B1(n20799), .B2(n20930), .ZN(
        n20790) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20932), .ZN(n20789) );
  OAI211_X1 U23773 ( .C1(n9853), .C2(n20804), .A(n20790), .B(n20789), .ZN(
        P1_U3107) );
  AOI22_X1 U23774 ( .A1(n20938), .A2(n20800), .B1(n20799), .B2(n20937), .ZN(
        n20792) );
  AOI22_X1 U23775 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20939), .ZN(n20791) );
  OAI211_X1 U23776 ( .C1(n20833), .C2(n20804), .A(n20792), .B(n20791), .ZN(
        P1_U3108) );
  AOI22_X1 U23777 ( .A1(n20945), .A2(n20800), .B1(n20799), .B2(n20944), .ZN(
        n20794) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20946), .ZN(n20793) );
  OAI211_X1 U23779 ( .C1(n20838), .C2(n20804), .A(n20794), .B(n20793), .ZN(
        P1_U3109) );
  AOI22_X1 U23780 ( .A1(n20952), .A2(n20800), .B1(n20799), .B2(n20951), .ZN(
        n20796) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20953), .ZN(n20795) );
  OAI211_X1 U23782 ( .C1(n20843), .C2(n20804), .A(n20796), .B(n20795), .ZN(
        P1_U3110) );
  AOI22_X1 U23783 ( .A1(n20959), .A2(n20800), .B1(n20799), .B2(n20958), .ZN(
        n20798) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20960), .ZN(n20797) );
  OAI211_X1 U23785 ( .C1(n9859), .C2(n20804), .A(n20798), .B(n20797), .ZN(
        P1_U3111) );
  AOI22_X1 U23786 ( .A1(n20968), .A2(n20800), .B1(n20799), .B2(n20966), .ZN(
        n20803) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20801), .B1(
        n20805), .B2(n20969), .ZN(n20802) );
  OAI211_X1 U23788 ( .C1(n9855), .C2(n20804), .A(n20803), .B(n20802), .ZN(
        P1_U3112) );
  NOR3_X1 U23789 ( .A1(n20805), .A2(n20855), .A3(n20915), .ZN(n20806) );
  NOR2_X1 U23790 ( .A1(n20806), .A2(n20863), .ZN(n20821) );
  INV_X1 U23791 ( .A(n20821), .ZN(n20810) );
  AND2_X1 U23792 ( .A1(n20807), .A2(n20865), .ZN(n20820) );
  NOR2_X1 U23793 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20811), .ZN(
        n20816) );
  INV_X1 U23794 ( .A(n20816), .ZN(n20851) );
  OAI22_X1 U23795 ( .A1(n20853), .A2(n9851), .B1(n20812), .B2(n20851), .ZN(
        n20813) );
  INV_X1 U23796 ( .A(n20813), .ZN(n20823) );
  OAI211_X1 U23797 ( .C1(n20817), .C2(n20816), .A(n20815), .B(n20814), .ZN(
        n20818) );
  INV_X1 U23798 ( .A(n20818), .ZN(n20819) );
  AOI22_X1 U23799 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n20919), .B2(n20855), .ZN(n20822) );
  OAI211_X1 U23800 ( .C1(n20859), .C2(n20879), .A(n20823), .B(n20822), .ZN(
        P1_U3113) );
  OAI22_X1 U23801 ( .A1(n20853), .A2(n9857), .B1(n20824), .B2(n20851), .ZN(
        n20825) );
  INV_X1 U23802 ( .A(n20825), .ZN(n20827) );
  AOI22_X1 U23803 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n20925), .B2(n20855), .ZN(n20826) );
  OAI211_X1 U23804 ( .C1(n20859), .C2(n20882), .A(n20827), .B(n20826), .ZN(
        P1_U3114) );
  OAI22_X1 U23805 ( .A1(n20853), .A2(n9853), .B1(n20828), .B2(n20851), .ZN(
        n20829) );
  INV_X1 U23806 ( .A(n20829), .ZN(n20831) );
  AOI22_X1 U23807 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n20932), .B2(n20855), .ZN(n20830) );
  OAI211_X1 U23808 ( .C1(n20859), .C2(n20885), .A(n20831), .B(n20830), .ZN(
        P1_U3115) );
  OAI22_X1 U23809 ( .A1(n20853), .A2(n20833), .B1(n20832), .B2(n20851), .ZN(
        n20834) );
  INV_X1 U23810 ( .A(n20834), .ZN(n20836) );
  AOI22_X1 U23811 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20939), .B2(n20855), .ZN(n20835) );
  OAI211_X1 U23812 ( .C1(n20859), .C2(n20888), .A(n20836), .B(n20835), .ZN(
        P1_U3116) );
  OAI22_X1 U23813 ( .A1(n20853), .A2(n20838), .B1(n20837), .B2(n20851), .ZN(
        n20839) );
  INV_X1 U23814 ( .A(n20839), .ZN(n20841) );
  AOI22_X1 U23815 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n20946), .B2(n20855), .ZN(n20840) );
  OAI211_X1 U23816 ( .C1(n20859), .C2(n20891), .A(n20841), .B(n20840), .ZN(
        P1_U3117) );
  OAI22_X1 U23817 ( .A1(n20853), .A2(n20843), .B1(n20842), .B2(n20851), .ZN(
        n20844) );
  INV_X1 U23818 ( .A(n20844), .ZN(n20846) );
  AOI22_X1 U23819 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n20953), .B2(n20855), .ZN(n20845) );
  OAI211_X1 U23820 ( .C1(n20859), .C2(n20894), .A(n20846), .B(n20845), .ZN(
        P1_U3118) );
  OAI22_X1 U23821 ( .A1(n20853), .A2(n9859), .B1(n20847), .B2(n20851), .ZN(
        n20848) );
  INV_X1 U23822 ( .A(n20848), .ZN(n20850) );
  AOI22_X1 U23823 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n20960), .B2(n20855), .ZN(n20849) );
  OAI211_X1 U23824 ( .C1(n20859), .C2(n20897), .A(n20850), .B(n20849), .ZN(
        P1_U3119) );
  OAI22_X1 U23825 ( .A1(n20853), .A2(n9855), .B1(n20852), .B2(n20851), .ZN(
        n20854) );
  INV_X1 U23826 ( .A(n20854), .ZN(n20858) );
  AOI22_X1 U23827 ( .A1(n20856), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9850), .B2(n20855), .ZN(n20857) );
  OAI211_X1 U23828 ( .C1(n20859), .C2(n20903), .A(n20858), .B(n20857), .ZN(
        P1_U3120) );
  NOR3_X1 U23829 ( .A1(n20899), .A2(n20972), .A3(n20915), .ZN(n20864) );
  NOR2_X1 U23830 ( .A1(n20864), .A2(n20863), .ZN(n20876) );
  INV_X1 U23831 ( .A(n20876), .ZN(n20869) );
  NOR2_X1 U23832 ( .A1(n20866), .A2(n20865), .ZN(n20875) );
  INV_X1 U23833 ( .A(n20872), .ZN(n20867) );
  NAND3_X1 U23834 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20870), .ZN(n20914) );
  NOR2_X1 U23835 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20914), .ZN(
        n20898) );
  AOI22_X1 U23836 ( .A1(n20972), .A2(n20919), .B1(n20918), .B2(n20898), .ZN(
        n20878) );
  INV_X1 U23837 ( .A(n20898), .ZN(n20871) );
  AOI22_X1 U23838 ( .A1(n20872), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20871), .ZN(n20873) );
  OAI211_X1 U23839 ( .C1(n20876), .C2(n20875), .A(n20874), .B(n20873), .ZN(
        n20900) );
  AOI22_X1 U23840 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9852), .B2(n20899), .ZN(n20877) );
  OAI211_X1 U23841 ( .C1(n20904), .C2(n20879), .A(n20878), .B(n20877), .ZN(
        P1_U3129) );
  AOI22_X1 U23842 ( .A1(n20972), .A2(n20925), .B1(n20924), .B2(n20898), .ZN(
        n20881) );
  AOI22_X1 U23843 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9858), .B2(n20899), .ZN(n20880) );
  OAI211_X1 U23844 ( .C1(n20904), .C2(n20882), .A(n20881), .B(n20880), .ZN(
        P1_U3130) );
  AOI22_X1 U23845 ( .A1(n20972), .A2(n20932), .B1(n20931), .B2(n20898), .ZN(
        n20884) );
  AOI22_X1 U23846 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9854), .B2(n20899), .ZN(n20883) );
  OAI211_X1 U23847 ( .C1(n20904), .C2(n20885), .A(n20884), .B(n20883), .ZN(
        P1_U3131) );
  AOI22_X1 U23848 ( .A1(n20972), .A2(n20939), .B1(n20938), .B2(n20898), .ZN(
        n20887) );
  AOI22_X1 U23849 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20940), .B2(n20899), .ZN(n20886) );
  OAI211_X1 U23850 ( .C1(n20904), .C2(n20888), .A(n20887), .B(n20886), .ZN(
        P1_U3132) );
  AOI22_X1 U23851 ( .A1(n20972), .A2(n20946), .B1(n20945), .B2(n20898), .ZN(
        n20890) );
  AOI22_X1 U23852 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20947), .B2(n20899), .ZN(n20889) );
  OAI211_X1 U23853 ( .C1(n20904), .C2(n20891), .A(n20890), .B(n20889), .ZN(
        P1_U3133) );
  AOI22_X1 U23854 ( .A1(n20972), .A2(n20953), .B1(n20952), .B2(n20898), .ZN(
        n20893) );
  AOI22_X1 U23855 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20954), .B2(n20899), .ZN(n20892) );
  OAI211_X1 U23856 ( .C1(n20904), .C2(n20894), .A(n20893), .B(n20892), .ZN(
        P1_U3134) );
  AOI22_X1 U23857 ( .A1(n20972), .A2(n20960), .B1(n20959), .B2(n20898), .ZN(
        n20896) );
  AOI22_X1 U23858 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9860), .B2(n20899), .ZN(n20895) );
  OAI211_X1 U23859 ( .C1(n20904), .C2(n20897), .A(n20896), .B(n20895), .ZN(
        P1_U3135) );
  AOI22_X1 U23860 ( .A1(n20972), .A2(n9850), .B1(n20968), .B2(n20898), .ZN(
        n20902) );
  AOI22_X1 U23861 ( .A1(n20900), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9856), .B2(n20899), .ZN(n20901) );
  OAI211_X1 U23862 ( .C1(n20904), .C2(n20903), .A(n20902), .B(n20901), .ZN(
        P1_U3136) );
  NOR2_X1 U23863 ( .A1(n20905), .A2(n20914), .ZN(n20967) );
  AOI21_X1 U23864 ( .B1(n20907), .B2(n20906), .A(n20967), .ZN(n20916) );
  INV_X1 U23865 ( .A(n20916), .ZN(n20908) );
  NOR2_X1 U23866 ( .A1(n20909), .A2(n20908), .ZN(n20912) );
  INV_X1 U23867 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n21273) );
  OAI22_X1 U23868 ( .A1(n20916), .A2(n20915), .B1(n20914), .B2(n20913), .ZN(
        n20965) );
  AOI22_X1 U23869 ( .A1(n20918), .A2(n20967), .B1(n20917), .B2(n20965), .ZN(
        n20922) );
  AOI22_X1 U23870 ( .A1(n20972), .A2(n9852), .B1(n20970), .B2(n20919), .ZN(
        n20921) );
  OAI211_X1 U23871 ( .C1(n20976), .C2(n21273), .A(n20922), .B(n20921), .ZN(
        P1_U3137) );
  INV_X1 U23872 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20929) );
  AOI22_X1 U23873 ( .A1(n20924), .A2(n20967), .B1(n20923), .B2(n20965), .ZN(
        n20928) );
  AOI22_X1 U23874 ( .A1(n20972), .A2(n9858), .B1(n20970), .B2(n20925), .ZN(
        n20927) );
  OAI211_X1 U23875 ( .C1(n20976), .C2(n20929), .A(n20928), .B(n20927), .ZN(
        P1_U3138) );
  INV_X1 U23876 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U23877 ( .A1(n20931), .A2(n20967), .B1(n20930), .B2(n20965), .ZN(
        n20935) );
  AOI22_X1 U23878 ( .A1(n20972), .A2(n9854), .B1(n20970), .B2(n20932), .ZN(
        n20934) );
  OAI211_X1 U23879 ( .C1(n20976), .C2(n20936), .A(n20935), .B(n20934), .ZN(
        P1_U3139) );
  INV_X1 U23880 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20943) );
  AOI22_X1 U23881 ( .A1(n20938), .A2(n20967), .B1(n20937), .B2(n20965), .ZN(
        n20942) );
  AOI22_X1 U23882 ( .A1(n20972), .A2(n20940), .B1(n20970), .B2(n20939), .ZN(
        n20941) );
  OAI211_X1 U23883 ( .C1(n20976), .C2(n20943), .A(n20942), .B(n20941), .ZN(
        P1_U3140) );
  INV_X1 U23884 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20950) );
  AOI22_X1 U23885 ( .A1(n20945), .A2(n20967), .B1(n20944), .B2(n20965), .ZN(
        n20949) );
  AOI22_X1 U23886 ( .A1(n20972), .A2(n20947), .B1(n20970), .B2(n20946), .ZN(
        n20948) );
  OAI211_X1 U23887 ( .C1(n20976), .C2(n20950), .A(n20949), .B(n20948), .ZN(
        P1_U3141) );
  INV_X1 U23888 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20957) );
  AOI22_X1 U23889 ( .A1(n20952), .A2(n20967), .B1(n20951), .B2(n20965), .ZN(
        n20956) );
  AOI22_X1 U23890 ( .A1(n20972), .A2(n20954), .B1(n20970), .B2(n20953), .ZN(
        n20955) );
  OAI211_X1 U23891 ( .C1(n20976), .C2(n20957), .A(n20956), .B(n20955), .ZN(
        P1_U3142) );
  INV_X1 U23892 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n20964) );
  AOI22_X1 U23893 ( .A1(n20959), .A2(n20967), .B1(n20958), .B2(n20965), .ZN(
        n20963) );
  AOI22_X1 U23894 ( .A1(n20972), .A2(n9860), .B1(n20970), .B2(n20960), .ZN(
        n20962) );
  OAI211_X1 U23895 ( .C1(n20976), .C2(n20964), .A(n20963), .B(n20962), .ZN(
        P1_U3143) );
  INV_X1 U23896 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U23897 ( .A1(n20968), .A2(n20967), .B1(n20966), .B2(n20965), .ZN(
        n20974) );
  AOI22_X1 U23898 ( .A1(n20972), .A2(n9856), .B1(n20970), .B2(n9850), .ZN(
        n20973) );
  OAI211_X1 U23899 ( .C1(n20976), .C2(n20975), .A(n20974), .B(n20973), .ZN(
        P1_U3144) );
  NOR2_X1 U23900 ( .A1(n9919), .A2(n21247), .ZN(n20978) );
  OAI21_X1 U23901 ( .B1(n20978), .B2(n20913), .A(n20977), .ZN(P1_U3163) );
  AND2_X1 U23902 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20979), .ZN(
        P1_U3164) );
  AND2_X1 U23903 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20980), .ZN(
        P1_U3165) );
  AND2_X1 U23904 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20980), .ZN(
        P1_U3166) );
  AND2_X1 U23905 ( .A1(n20980), .A2(P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(
        P1_U3167) );
  AND2_X1 U23906 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20980), .ZN(
        P1_U3168) );
  AND2_X1 U23907 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20980), .ZN(
        P1_U3169) );
  AND2_X1 U23908 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20980), .ZN(
        P1_U3170) );
  AND2_X1 U23909 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20979), .ZN(
        P1_U3171) );
  AND2_X1 U23910 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20980), .ZN(
        P1_U3172) );
  AND2_X1 U23911 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20979), .ZN(
        P1_U3173) );
  AND2_X1 U23912 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20979), .ZN(
        P1_U3174) );
  AND2_X1 U23913 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20979), .ZN(
        P1_U3175) );
  AND2_X1 U23914 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20979), .ZN(
        P1_U3176) );
  AND2_X1 U23915 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20979), .ZN(
        P1_U3177) );
  AND2_X1 U23916 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20980), .ZN(
        P1_U3178) );
  AND2_X1 U23917 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20980), .ZN(
        P1_U3179) );
  AND2_X1 U23918 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20980), .ZN(
        P1_U3180) );
  AND2_X1 U23919 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20980), .ZN(
        P1_U3181) );
  AND2_X1 U23920 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20979), .ZN(
        P1_U3182) );
  AND2_X1 U23921 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20979), .ZN(
        P1_U3183) );
  AND2_X1 U23922 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20979), .ZN(
        P1_U3184) );
  AND2_X1 U23923 ( .A1(n20980), .A2(P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P1_U3185) );
  AND2_X1 U23924 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20979), .ZN(P1_U3186) );
  AND2_X1 U23925 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20979), .ZN(P1_U3187) );
  AND2_X1 U23926 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20980), .ZN(P1_U3188) );
  AND2_X1 U23927 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20979), .ZN(P1_U3189) );
  AND2_X1 U23928 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20980), .ZN(P1_U3190) );
  AND2_X1 U23929 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20979), .ZN(P1_U3191) );
  AND2_X1 U23930 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20980), .ZN(P1_U3192) );
  AND2_X1 U23931 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20980), .ZN(P1_U3193) );
  AOI21_X1 U23932 ( .B1(n20982), .B2(n20998), .A(n20981), .ZN(n20983) );
  AOI211_X1 U23933 ( .C1(NA), .C2(n20992), .A(n20983), .B(n20991), .ZN(n20987)
         );
  AOI21_X1 U23934 ( .B1(n20989), .B2(n20985), .A(n20984), .ZN(n20986) );
  OAI21_X1 U23935 ( .B1(n21058), .B2(n20987), .A(n20986), .ZN(P1_U3194) );
  AOI21_X1 U23936 ( .B1(n20988), .B2(n20993), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20997) );
  AOI221_X1 U23937 ( .B1(NA), .B2(n20989), .C1(n21066), .C2(n20989), .A(n20992), .ZN(n20990) );
  OAI211_X1 U23938 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20991), .A(HOLD), .B(
        n20990), .ZN(n20995) );
  OAI211_X1 U23939 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20993), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20992), .ZN(n20994) );
  OAI211_X1 U23940 ( .C1(n20997), .C2(n20996), .A(n20995), .B(n20994), .ZN(
        P1_U3196) );
  OR2_X1 U23941 ( .A1(n21056), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21034) );
  OR2_X1 U23942 ( .A1(n20998), .A2(n21056), .ZN(n21031) );
  INV_X1 U23943 ( .A(n21031), .ZN(n21039) );
  AOI222_X1 U23944 ( .A1(n21038), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21039), .ZN(n20999) );
  INV_X1 U23945 ( .A(n20999), .ZN(P1_U3197) );
  AOI22_X1 U23946 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n21038), .ZN(n21000) );
  OAI21_X1 U23947 ( .B1(n21001), .B2(n21031), .A(n21000), .ZN(P1_U3198) );
  AOI222_X1 U23948 ( .A1(n21038), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21039), .ZN(n21002) );
  INV_X1 U23949 ( .A(n21002), .ZN(P1_U3199) );
  AOI222_X1 U23950 ( .A1(n21038), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21039), .ZN(n21003) );
  INV_X1 U23951 ( .A(n21003), .ZN(P1_U3200) );
  AOI222_X1 U23952 ( .A1(n21039), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21038), .ZN(n21004) );
  INV_X1 U23953 ( .A(n21004), .ZN(P1_U3201) );
  AOI222_X1 U23954 ( .A1(n21039), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21038), .ZN(n21005) );
  INV_X1 U23955 ( .A(n21005), .ZN(P1_U3202) );
  AOI22_X1 U23956 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21038), .ZN(n21006) );
  OAI21_X1 U23957 ( .B1(n21007), .B2(n21031), .A(n21006), .ZN(P1_U3203) );
  AOI22_X1 U23958 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21039), .ZN(n21008) );
  OAI21_X1 U23959 ( .B1(n21009), .B2(n21034), .A(n21008), .ZN(P1_U3204) );
  AOI222_X1 U23960 ( .A1(n21038), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n21039), .ZN(n21010) );
  INV_X1 U23961 ( .A(n21010), .ZN(P1_U3205) );
  AOI222_X1 U23962 ( .A1(n21038), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21039), .ZN(n21011) );
  INV_X1 U23963 ( .A(n21011), .ZN(P1_U3206) );
  AOI222_X1 U23964 ( .A1(n21039), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21038), .ZN(n21012) );
  INV_X1 U23965 ( .A(n21012), .ZN(P1_U3207) );
  AOI222_X1 U23966 ( .A1(n21039), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21038), .ZN(n21013) );
  INV_X1 U23967 ( .A(n21013), .ZN(P1_U3208) );
  INV_X1 U23968 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21152) );
  OAI222_X1 U23969 ( .A1(n21031), .A2(n21387), .B1(n21152), .B2(n21058), .C1(
        n21385), .C2(n21034), .ZN(P1_U3209) );
  AOI222_X1 U23970 ( .A1(n21038), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21039), .ZN(n21014) );
  INV_X1 U23971 ( .A(n21014), .ZN(P1_U3210) );
  AOI22_X1 U23972 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21038), .ZN(n21015) );
  OAI21_X1 U23973 ( .B1(n21016), .B2(n21031), .A(n21015), .ZN(P1_U3211) );
  AOI22_X1 U23974 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21039), .ZN(n21017) );
  OAI21_X1 U23975 ( .B1(n21018), .B2(n21034), .A(n21017), .ZN(P1_U3212) );
  AOI222_X1 U23976 ( .A1(n21038), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21039), .ZN(n21019) );
  INV_X1 U23977 ( .A(n21019), .ZN(P1_U3213) );
  AOI22_X1 U23978 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21038), .ZN(n21020) );
  OAI21_X1 U23979 ( .B1(n16238), .B2(n21031), .A(n21020), .ZN(P1_U3214) );
  AOI22_X1 U23980 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21039), .ZN(n21021) );
  OAI21_X1 U23981 ( .B1(n21022), .B2(n21034), .A(n21021), .ZN(P1_U3215) );
  AOI222_X1 U23982 ( .A1(n21038), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n21039), .ZN(n21023) );
  INV_X1 U23983 ( .A(n21023), .ZN(P1_U3216) );
  AOI222_X1 U23984 ( .A1(n21038), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21039), .ZN(n21024) );
  INV_X1 U23985 ( .A(n21024), .ZN(P1_U3217) );
  AOI222_X1 U23986 ( .A1(n21039), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21038), .ZN(n21025) );
  INV_X1 U23987 ( .A(n21025), .ZN(P1_U3218) );
  AOI222_X1 U23988 ( .A1(n21038), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21039), .ZN(n21026) );
  INV_X1 U23989 ( .A(n21026), .ZN(P1_U3219) );
  AOI22_X1 U23990 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21038), .ZN(n21027) );
  OAI21_X1 U23991 ( .B1(n21028), .B2(n21031), .A(n21027), .ZN(P1_U3220) );
  AOI22_X1 U23992 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(n21056), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21039), .ZN(n21029) );
  OAI21_X1 U23993 ( .B1(n21032), .B2(n21034), .A(n21029), .ZN(P1_U3221) );
  AOI22_X1 U23994 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n21038), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21056), .ZN(n21030) );
  OAI21_X1 U23995 ( .B1(n21032), .B2(n21031), .A(n21030), .ZN(P1_U3222) );
  AOI22_X1 U23996 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n21039), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21056), .ZN(n21033) );
  OAI21_X1 U23997 ( .B1(n21035), .B2(n21034), .A(n21033), .ZN(P1_U3223) );
  AOI222_X1 U23998 ( .A1(n21039), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21038), .ZN(n21036) );
  INV_X1 U23999 ( .A(n21036), .ZN(P1_U3224) );
  AOI222_X1 U24000 ( .A1(n21039), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n21038), .ZN(n21037) );
  INV_X1 U24001 ( .A(n21037), .ZN(P1_U3225) );
  AOI222_X1 U24002 ( .A1(n21039), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21056), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21038), .ZN(n21040) );
  INV_X1 U24003 ( .A(n21040), .ZN(P1_U3226) );
  OAI22_X1 U24004 ( .A1(n21056), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21058), .ZN(n21041) );
  INV_X1 U24005 ( .A(n21041), .ZN(P1_U3458) );
  OAI22_X1 U24006 ( .A1(n21056), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21058), .ZN(n21042) );
  INV_X1 U24007 ( .A(n21042), .ZN(P1_U3459) );
  OAI22_X1 U24008 ( .A1(n21056), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21058), .ZN(n21043) );
  INV_X1 U24009 ( .A(n21043), .ZN(P1_U3460) );
  OAI22_X1 U24010 ( .A1(n21056), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21058), .ZN(n21044) );
  INV_X1 U24011 ( .A(n21044), .ZN(P1_U3461) );
  OAI21_X1 U24012 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21048), .A(n21046), 
        .ZN(n21045) );
  INV_X1 U24013 ( .A(n21045), .ZN(P1_U3464) );
  OAI21_X1 U24014 ( .B1(n21048), .B2(n21047), .A(n21046), .ZN(P1_U3465) );
  AOI211_X1 U24015 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21049) );
  AOI21_X1 U24016 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21049), .ZN(n21051) );
  INV_X1 U24017 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21050) );
  AOI22_X1 U24018 ( .A1(n21055), .A2(n21051), .B1(n21050), .B2(n21052), .ZN(
        P1_U3481) );
  NOR2_X1 U24019 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21054) );
  INV_X1 U24020 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21053) );
  AOI22_X1 U24021 ( .A1(n21055), .A2(n21054), .B1(n21053), .B2(n21052), .ZN(
        P1_U3482) );
  AOI22_X1 U24022 ( .A1(n21058), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21057), 
        .B2(n21056), .ZN(P1_U3483) );
  OAI211_X1 U24023 ( .C1(n21059), .C2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .B(n21066), .ZN(n21060) );
  OAI21_X1 U24024 ( .B1(n21061), .B2(n21060), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n21063) );
  NAND2_X1 U24025 ( .A1(n21063), .A2(n21062), .ZN(n21069) );
  AOI211_X1 U24026 ( .C1(n21067), .C2(n21066), .A(n21065), .B(n21064), .ZN(
        n21068) );
  MUX2_X1 U24027 ( .A(n21069), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21068), 
        .Z(P1_U3485) );
  MUX2_X1 U24028 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21056), .Z(P1_U3486) );
  AOI22_X1 U24029 ( .A1(n21072), .A2(keyinput120), .B1(n21071), .B2(
        keyinput111), .ZN(n21070) );
  OAI221_X1 U24030 ( .B1(n21072), .B2(keyinput120), .C1(n21071), .C2(
        keyinput111), .A(n21070), .ZN(n21084) );
  INV_X1 U24031 ( .A(keyinput28), .ZN(n21074) );
  AOI22_X1 U24032 ( .A1(n21075), .A2(keyinput109), .B1(BUF2_REG_5__SCAN_IN), 
        .B2(n21074), .ZN(n21073) );
  OAI221_X1 U24033 ( .B1(n21075), .B2(keyinput109), .C1(n21074), .C2(
        BUF2_REG_5__SCAN_IN), .A(n21073), .ZN(n21083) );
  AOI22_X1 U24034 ( .A1(n21077), .A2(keyinput117), .B1(n11451), .B2(keyinput97), .ZN(n21076) );
  OAI221_X1 U24035 ( .B1(n21077), .B2(keyinput117), .C1(n11451), .C2(
        keyinput97), .A(n21076), .ZN(n21082) );
  INV_X1 U24036 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U24037 ( .A1(n21080), .A2(keyinput124), .B1(keyinput71), .B2(n21079), .ZN(n21078) );
  OAI221_X1 U24038 ( .B1(n21080), .B2(keyinput124), .C1(n21079), .C2(
        keyinput71), .A(n21078), .ZN(n21081) );
  NOR4_X1 U24039 ( .A1(n21084), .A2(n21083), .A3(n21082), .A4(n21081), .ZN(
        n21384) );
  OAI22_X1 U24040 ( .A1(n21087), .A2(keyinput45), .B1(n21086), .B2(keyinput72), 
        .ZN(n21085) );
  AOI221_X1 U24041 ( .B1(n21087), .B2(keyinput45), .C1(keyinput72), .C2(n21086), .A(n21085), .ZN(n21100) );
  INV_X1 U24042 ( .A(keyinput86), .ZN(n21089) );
  OAI22_X1 U24043 ( .A1(keyinput108), .A2(n21090), .B1(n21089), .B2(
        P1_DATAO_REG_4__SCAN_IN), .ZN(n21088) );
  AOI221_X1 U24044 ( .B1(n21090), .B2(keyinput108), .C1(n21089), .C2(
        P1_DATAO_REG_4__SCAN_IN), .A(n21088), .ZN(n21099) );
  INV_X1 U24045 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21093) );
  INV_X1 U24046 ( .A(keyinput96), .ZN(n21092) );
  OAI22_X1 U24047 ( .A1(n21093), .A2(keyinput103), .B1(n21092), .B2(
        P3_ADDRESS_REG_28__SCAN_IN), .ZN(n21091) );
  AOI221_X1 U24048 ( .B1(n21093), .B2(keyinput103), .C1(
        P3_ADDRESS_REG_28__SCAN_IN), .C2(n21092), .A(n21091), .ZN(n21098) );
  INV_X1 U24049 ( .A(keyinput3), .ZN(n21095) );
  OAI22_X1 U24050 ( .A1(n21096), .A2(keyinput59), .B1(n21095), .B2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21094) );
  AOI221_X1 U24051 ( .B1(n21096), .B2(keyinput59), .C1(
        P2_DATAWIDTH_REG_2__SCAN_IN), .C2(n21095), .A(n21094), .ZN(n21097) );
  NAND4_X1 U24052 ( .A1(n21100), .A2(n21099), .A3(n21098), .A4(n21097), .ZN(
        n21133) );
  INV_X1 U24053 ( .A(keyinput64), .ZN(n21102) );
  OAI22_X1 U24054 ( .A1(n12866), .A2(keyinput105), .B1(n21102), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n21101) );
  AOI221_X1 U24055 ( .B1(n12866), .B2(keyinput105), .C1(P3_REIP_REG_6__SCAN_IN), .C2(n21102), .A(n21101), .ZN(n21115) );
  INV_X1 U24056 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21105) );
  OAI22_X1 U24057 ( .A1(n21105), .A2(keyinput73), .B1(n21104), .B2(keyinput43), 
        .ZN(n21103) );
  AOI221_X1 U24058 ( .B1(n21105), .B2(keyinput73), .C1(keyinput43), .C2(n21104), .A(n21103), .ZN(n21114) );
  INV_X1 U24059 ( .A(keyinput101), .ZN(n21107) );
  OAI22_X1 U24060 ( .A1(n21108), .A2(keyinput84), .B1(n21107), .B2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21106) );
  AOI221_X1 U24061 ( .B1(n21108), .B2(keyinput84), .C1(
        P2_DATAWIDTH_REG_8__SCAN_IN), .C2(n21107), .A(n21106), .ZN(n21113) );
  OAI22_X1 U24062 ( .A1(keyinput114), .A2(n21111), .B1(n21110), .B2(keyinput56), .ZN(n21109) );
  AOI221_X1 U24063 ( .B1(n21111), .B2(keyinput114), .C1(n21110), .C2(
        keyinput56), .A(n21109), .ZN(n21112) );
  NAND4_X1 U24064 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21132) );
  INV_X1 U24065 ( .A(keyinput49), .ZN(n21117) );
  OAI22_X1 U24066 ( .A1(n21118), .A2(keyinput88), .B1(n21117), .B2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21116) );
  AOI221_X1 U24067 ( .B1(n21118), .B2(keyinput88), .C1(
        P1_DATAWIDTH_REG_10__SCAN_IN), .C2(n21117), .A(n21116), .ZN(n21130) );
  INV_X1 U24068 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n21120) );
  OAI22_X1 U24069 ( .A1(n21120), .A2(keyinput30), .B1(n11731), .B2(keyinput20), 
        .ZN(n21119) );
  AOI221_X1 U24070 ( .B1(n21120), .B2(keyinput30), .C1(keyinput20), .C2(n11731), .A(n21119), .ZN(n21129) );
  OAI22_X1 U24071 ( .A1(keyinput6), .A2(n21123), .B1(n21122), .B2(keyinput95), 
        .ZN(n21121) );
  AOI221_X1 U24072 ( .B1(n21123), .B2(keyinput6), .C1(n21122), .C2(keyinput95), 
        .A(n21121), .ZN(n21128) );
  INV_X1 U24073 ( .A(keyinput5), .ZN(n21125) );
  OAI22_X1 U24074 ( .A1(n21126), .A2(keyinput19), .B1(n21125), .B2(
        P3_REIP_REG_15__SCAN_IN), .ZN(n21124) );
  AOI221_X1 U24075 ( .B1(n21126), .B2(keyinput19), .C1(P3_REIP_REG_15__SCAN_IN), .C2(n21125), .A(n21124), .ZN(n21127) );
  NAND4_X1 U24076 ( .A1(n21130), .A2(n21129), .A3(n21128), .A4(n21127), .ZN(
        n21131) );
  NOR3_X1 U24077 ( .A1(n21133), .A2(n21132), .A3(n21131), .ZN(n21383) );
  INV_X1 U24078 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21136) );
  INV_X1 U24079 ( .A(keyinput126), .ZN(n21135) );
  OAI22_X1 U24080 ( .A1(n21136), .A2(keyinput67), .B1(n21135), .B2(
        P3_DATAO_REG_24__SCAN_IN), .ZN(n21134) );
  AOI221_X1 U24081 ( .B1(n21136), .B2(keyinput67), .C1(
        P3_DATAO_REG_24__SCAN_IN), .C2(n21135), .A(n21134), .ZN(n21149) );
  INV_X1 U24082 ( .A(keyinput18), .ZN(n21138) );
  OAI22_X1 U24083 ( .A1(n21139), .A2(keyinput121), .B1(n21138), .B2(
        P3_EBX_REG_15__SCAN_IN), .ZN(n21137) );
  AOI221_X1 U24084 ( .B1(n21139), .B2(keyinput121), .C1(P3_EBX_REG_15__SCAN_IN), .C2(n21138), .A(n21137), .ZN(n21148) );
  OAI22_X1 U24085 ( .A1(keyinput57), .A2(n21142), .B1(n21141), .B2(keyinput115), .ZN(n21140) );
  AOI221_X1 U24086 ( .B1(n21142), .B2(keyinput57), .C1(n21141), .C2(
        keyinput115), .A(n21140), .ZN(n21147) );
  INV_X1 U24087 ( .A(keyinput80), .ZN(n21144) );
  OAI22_X1 U24088 ( .A1(n21145), .A2(keyinput79), .B1(n21144), .B2(
        P2_DATAO_REG_0__SCAN_IN), .ZN(n21143) );
  AOI221_X1 U24089 ( .B1(n21145), .B2(keyinput79), .C1(P2_DATAO_REG_0__SCAN_IN), .C2(n21144), .A(n21143), .ZN(n21146) );
  NAND4_X1 U24090 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21328) );
  AOI22_X1 U24091 ( .A1(n21152), .A2(keyinput100), .B1(n21151), .B2(keyinput9), 
        .ZN(n21150) );
  OAI221_X1 U24092 ( .B1(n21152), .B2(keyinput100), .C1(n21151), .C2(keyinput9), .A(n21150), .ZN(n21165) );
  INV_X1 U24093 ( .A(keyinput125), .ZN(n21154) );
  AOI22_X1 U24094 ( .A1(n21155), .A2(keyinput77), .B1(P3_DATAO_REG_23__SCAN_IN), .B2(n21154), .ZN(n21153) );
  OAI221_X1 U24095 ( .B1(n21155), .B2(keyinput77), .C1(n21154), .C2(
        P3_DATAO_REG_23__SCAN_IN), .A(n21153), .ZN(n21164) );
  INV_X1 U24096 ( .A(DATAI_11_), .ZN(n21158) );
  INV_X1 U24097 ( .A(DATAI_4_), .ZN(n21157) );
  AOI22_X1 U24098 ( .A1(n21158), .A2(keyinput41), .B1(keyinput68), .B2(n21157), 
        .ZN(n21156) );
  OAI221_X1 U24099 ( .B1(n21158), .B2(keyinput41), .C1(n21157), .C2(keyinput68), .A(n21156), .ZN(n21163) );
  INV_X1 U24100 ( .A(keyinput31), .ZN(n21160) );
  AOI22_X1 U24101 ( .A1(n21161), .A2(keyinput107), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n21160), .ZN(n21159) );
  OAI221_X1 U24102 ( .B1(n21161), .B2(keyinput107), .C1(n21160), .C2(
        P1_UWORD_REG_13__SCAN_IN), .A(n21159), .ZN(n21162) );
  NOR4_X1 U24103 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21199) );
  INV_X1 U24104 ( .A(keyinput33), .ZN(n21167) );
  AOI22_X1 U24105 ( .A1(n21168), .A2(keyinput14), .B1(P2_LWORD_REG_10__SCAN_IN), .B2(n21167), .ZN(n21166) );
  OAI221_X1 U24106 ( .B1(n21168), .B2(keyinput14), .C1(n21167), .C2(
        P2_LWORD_REG_10__SCAN_IN), .A(n21166), .ZN(n21181) );
  INV_X1 U24107 ( .A(keyinput10), .ZN(n21170) );
  AOI22_X1 U24108 ( .A1(n21171), .A2(keyinput48), .B1(P1_DATAO_REG_30__SCAN_IN), .B2(n21170), .ZN(n21169) );
  OAI221_X1 U24109 ( .B1(n21171), .B2(keyinput48), .C1(n21170), .C2(
        P1_DATAO_REG_30__SCAN_IN), .A(n21169), .ZN(n21180) );
  INV_X1 U24110 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21173) );
  AOI22_X1 U24111 ( .A1(n21174), .A2(keyinput38), .B1(n21173), .B2(keyinput47), 
        .ZN(n21172) );
  OAI221_X1 U24112 ( .B1(n21174), .B2(keyinput38), .C1(n21173), .C2(keyinput47), .A(n21172), .ZN(n21179) );
  INV_X1 U24113 ( .A(keyinput91), .ZN(n21175) );
  XOR2_X1 U24114 ( .A(P1_LWORD_REG_3__SCAN_IN), .B(n21175), .Z(n21177) );
  XNOR2_X1 U24115 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput98), 
        .ZN(n21176) );
  NAND2_X1 U24116 ( .A1(n21177), .A2(n21176), .ZN(n21178) );
  NOR4_X1 U24117 ( .A1(n21181), .A2(n21180), .A3(n21179), .A4(n21178), .ZN(
        n21198) );
  INV_X1 U24118 ( .A(keyinput66), .ZN(n21183) );
  OAI22_X1 U24119 ( .A1(keyinput53), .A2(n21184), .B1(n21183), .B2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21182) );
  AOI221_X1 U24120 ( .B1(n21184), .B2(keyinput53), .C1(n21183), .C2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A(n21182), .ZN(n21197) );
  AOI22_X1 U24121 ( .A1(n21187), .A2(keyinput35), .B1(keyinput110), .B2(n21186), .ZN(n21185) );
  OAI221_X1 U24122 ( .B1(n21187), .B2(keyinput35), .C1(n21186), .C2(
        keyinput110), .A(n21185), .ZN(n21195) );
  INV_X1 U24123 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21190) );
  INV_X1 U24124 ( .A(keyinput46), .ZN(n21189) );
  AOI22_X1 U24125 ( .A1(n21190), .A2(keyinput123), .B1(
        P3_DATAWIDTH_REG_9__SCAN_IN), .B2(n21189), .ZN(n21188) );
  OAI221_X1 U24126 ( .B1(n21190), .B2(keyinput123), .C1(n21189), .C2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A(n21188), .ZN(n21194) );
  AOI22_X1 U24127 ( .A1(n21192), .A2(keyinput25), .B1(keyinput69), .B2(n12721), 
        .ZN(n21191) );
  OAI221_X1 U24128 ( .B1(n21192), .B2(keyinput25), .C1(n12721), .C2(keyinput69), .A(n21191), .ZN(n21193) );
  NOR3_X1 U24129 ( .A1(n21195), .A2(n21194), .A3(n21193), .ZN(n21196) );
  NAND4_X1 U24130 ( .A1(n21199), .A2(n21198), .A3(n21197), .A4(n21196), .ZN(
        n21327) );
  INV_X1 U24131 ( .A(keyinput102), .ZN(n21201) );
  AOI22_X1 U24132 ( .A1(n21202), .A2(keyinput27), .B1(P2_UWORD_REG_1__SCAN_IN), 
        .B2(n21201), .ZN(n21200) );
  OAI221_X1 U24133 ( .B1(n21202), .B2(keyinput27), .C1(n21201), .C2(
        P2_UWORD_REG_1__SCAN_IN), .A(n21200), .ZN(n21213) );
  INV_X1 U24134 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21204) );
  INV_X1 U24135 ( .A(keyinput17), .ZN(n21352) );
  AOI22_X1 U24136 ( .A1(n21204), .A2(keyinput7), .B1(P1_DATAO_REG_18__SCAN_IN), 
        .B2(n21352), .ZN(n21203) );
  OAI221_X1 U24137 ( .B1(n21204), .B2(keyinput7), .C1(n21352), .C2(
        P1_DATAO_REG_18__SCAN_IN), .A(n21203), .ZN(n21212) );
  AOI22_X1 U24138 ( .A1(n15083), .A2(keyinput116), .B1(n21206), .B2(keyinput89), .ZN(n21205) );
  OAI221_X1 U24139 ( .B1(n15083), .B2(keyinput116), .C1(n21206), .C2(
        keyinput89), .A(n21205), .ZN(n21211) );
  INV_X1 U24140 ( .A(keyinput4), .ZN(n21207) );
  XOR2_X1 U24141 ( .A(P3_FLUSH_REG_SCAN_IN), .B(n21207), .Z(n21209) );
  XNOR2_X1 U24142 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B(keyinput44), .ZN(
        n21208) );
  NAND2_X1 U24143 ( .A1(n21209), .A2(n21208), .ZN(n21210) );
  NOR4_X1 U24144 ( .A1(n21213), .A2(n21212), .A3(n21211), .A4(n21210), .ZN(
        n21262) );
  AOI22_X1 U24145 ( .A1(n21216), .A2(keyinput15), .B1(n21215), .B2(keyinput61), 
        .ZN(n21214) );
  OAI221_X1 U24146 ( .B1(n21216), .B2(keyinput15), .C1(n21215), .C2(keyinput61), .A(n21214), .ZN(n21217) );
  INV_X1 U24147 ( .A(n21217), .ZN(n21221) );
  INV_X1 U24148 ( .A(keyinput82), .ZN(n21218) );
  XOR2_X1 U24149 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n21218), .Z(n21220) );
  XNOR2_X1 U24150 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B(keyinput23), .ZN(
        n21219) );
  NAND3_X1 U24151 ( .A1(n21221), .A2(n21220), .A3(n21219), .ZN(n21230) );
  INV_X1 U24152 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21224) );
  AOI22_X1 U24153 ( .A1(n21224), .A2(keyinput62), .B1(keyinput74), .B2(n21223), 
        .ZN(n21222) );
  OAI221_X1 U24154 ( .B1(n21224), .B2(keyinput62), .C1(n21223), .C2(keyinput74), .A(n21222), .ZN(n21229) );
  AOI22_X1 U24155 ( .A1(n21227), .A2(keyinput83), .B1(keyinput8), .B2(n21226), 
        .ZN(n21225) );
  OAI221_X1 U24156 ( .B1(n21227), .B2(keyinput83), .C1(n21226), .C2(keyinput8), 
        .A(n21225), .ZN(n21228) );
  NOR3_X1 U24157 ( .A1(n21230), .A2(n21229), .A3(n21228), .ZN(n21261) );
  AOI22_X1 U24158 ( .A1(n11568), .A2(keyinput93), .B1(keyinput65), .B2(n14852), 
        .ZN(n21231) );
  OAI221_X1 U24159 ( .B1(n11568), .B2(keyinput93), .C1(n14852), .C2(keyinput65), .A(n21231), .ZN(n21244) );
  INV_X1 U24160 ( .A(keyinput37), .ZN(n21233) );
  AOI22_X1 U24161 ( .A1(n21234), .A2(keyinput75), .B1(P3_EAX_REG_2__SCAN_IN), 
        .B2(n21233), .ZN(n21232) );
  OAI221_X1 U24162 ( .B1(n21234), .B2(keyinput75), .C1(n21233), .C2(
        P3_EAX_REG_2__SCAN_IN), .A(n21232), .ZN(n21243) );
  INV_X1 U24163 ( .A(keyinput13), .ZN(n21236) );
  AOI22_X1 U24164 ( .A1(n21237), .A2(keyinput1), .B1(P3_EBX_REG_25__SCAN_IN), 
        .B2(n21236), .ZN(n21235) );
  OAI221_X1 U24165 ( .B1(n21237), .B2(keyinput1), .C1(n21236), .C2(
        P3_EBX_REG_25__SCAN_IN), .A(n21235), .ZN(n21242) );
  INV_X1 U24166 ( .A(keyinput24), .ZN(n21239) );
  AOI22_X1 U24167 ( .A1(n21240), .A2(keyinput29), .B1(
        P2_DATAWIDTH_REG_15__SCAN_IN), .B2(n21239), .ZN(n21238) );
  OAI221_X1 U24168 ( .B1(n21240), .B2(keyinput29), .C1(n21239), .C2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A(n21238), .ZN(n21241) );
  NOR4_X1 U24169 ( .A1(n21244), .A2(n21243), .A3(n21242), .A4(n21241), .ZN(
        n21260) );
  AOI22_X1 U24170 ( .A1(n21247), .A2(keyinput70), .B1(keyinput87), .B2(n21246), 
        .ZN(n21245) );
  OAI221_X1 U24171 ( .B1(n21247), .B2(keyinput70), .C1(n21246), .C2(keyinput87), .A(n21245), .ZN(n21258) );
  AOI22_X1 U24172 ( .A1(n21249), .A2(keyinput16), .B1(keyinput81), .B2(n9961), 
        .ZN(n21248) );
  OAI221_X1 U24173 ( .B1(n21249), .B2(keyinput16), .C1(n9961), .C2(keyinput81), 
        .A(n21248), .ZN(n21257) );
  INV_X1 U24174 ( .A(keyinput50), .ZN(n21252) );
  INV_X1 U24175 ( .A(keyinput63), .ZN(n21251) );
  AOI22_X1 U24176 ( .A1(n21252), .A2(P3_BE_N_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n21251), .ZN(n21250) );
  OAI221_X1 U24177 ( .B1(n21252), .B2(P3_BE_N_REG_2__SCAN_IN), .C1(n21251), 
        .C2(P3_ADDRESS_REG_9__SCAN_IN), .A(n21250), .ZN(n21256) );
  XNOR2_X1 U24178 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput106), .ZN(
        n21254) );
  XNOR2_X1 U24179 ( .A(keyinput85), .B(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n21253) );
  NAND2_X1 U24180 ( .A1(n21254), .A2(n21253), .ZN(n21255) );
  NOR4_X1 U24181 ( .A1(n21258), .A2(n21257), .A3(n21256), .A4(n21255), .ZN(
        n21259) );
  NAND4_X1 U24182 ( .A1(n21262), .A2(n21261), .A3(n21260), .A4(n21259), .ZN(
        n21326) );
  INV_X1 U24183 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21265) );
  AOI22_X1 U24184 ( .A1(n21265), .A2(keyinput55), .B1(keyinput34), .B2(n21264), 
        .ZN(n21263) );
  OAI221_X1 U24185 ( .B1(n21265), .B2(keyinput55), .C1(n21264), .C2(keyinput34), .A(n21263), .ZN(n21277) );
  INV_X1 U24186 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21268) );
  INV_X1 U24187 ( .A(keyinput58), .ZN(n21267) );
  AOI22_X1 U24188 ( .A1(n21268), .A2(keyinput51), .B1(P3_EBX_REG_9__SCAN_IN), 
        .B2(n21267), .ZN(n21266) );
  OAI221_X1 U24189 ( .B1(n21268), .B2(keyinput51), .C1(n21267), .C2(
        P3_EBX_REG_9__SCAN_IN), .A(n21266), .ZN(n21276) );
  INV_X1 U24190 ( .A(keyinput21), .ZN(n21270) );
  AOI22_X1 U24191 ( .A1(n10077), .A2(keyinput76), .B1(P3_DATAO_REG_8__SCAN_IN), 
        .B2(n21270), .ZN(n21269) );
  OAI221_X1 U24192 ( .B1(n10077), .B2(keyinput76), .C1(n21270), .C2(
        P3_DATAO_REG_8__SCAN_IN), .A(n21269), .ZN(n21275) );
  AOI22_X1 U24193 ( .A1(n21273), .A2(keyinput122), .B1(n21272), .B2(
        keyinput104), .ZN(n21271) );
  OAI221_X1 U24194 ( .B1(n21273), .B2(keyinput122), .C1(n21272), .C2(
        keyinput104), .A(n21271), .ZN(n21274) );
  NOR4_X1 U24195 ( .A1(n21277), .A2(n21276), .A3(n21275), .A4(n21274), .ZN(
        n21324) );
  AOI22_X1 U24196 ( .A1(n21280), .A2(keyinput36), .B1(keyinput90), .B2(n21279), 
        .ZN(n21278) );
  OAI221_X1 U24197 ( .B1(n21280), .B2(keyinput36), .C1(n21279), .C2(keyinput90), .A(n21278), .ZN(n21292) );
  INV_X1 U24198 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n21282) );
  AOI22_X1 U24199 ( .A1(n21282), .A2(keyinput2), .B1(keyinput94), .B2(n9948), 
        .ZN(n21281) );
  OAI221_X1 U24200 ( .B1(n21282), .B2(keyinput2), .C1(n9948), .C2(keyinput94), 
        .A(n21281), .ZN(n21291) );
  INV_X1 U24201 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21285) );
  AOI22_X1 U24202 ( .A1(n21285), .A2(keyinput22), .B1(n21284), .B2(keyinput0), 
        .ZN(n21283) );
  OAI221_X1 U24203 ( .B1(n21285), .B2(keyinput22), .C1(n21284), .C2(keyinput0), 
        .A(n21283), .ZN(n21290) );
  AOI22_X1 U24204 ( .A1(n21288), .A2(keyinput78), .B1(keyinput54), .B2(n21287), 
        .ZN(n21286) );
  OAI221_X1 U24205 ( .B1(n21288), .B2(keyinput78), .C1(n21287), .C2(keyinput54), .A(n21286), .ZN(n21289) );
  NOR4_X1 U24206 ( .A1(n21292), .A2(n21291), .A3(n21290), .A4(n21289), .ZN(
        n21323) );
  XOR2_X1 U24207 ( .A(keyinput112), .B(P3_DATAO_REG_29__SCAN_IN), .Z(n21307)
         );
  AOI22_X1 U24208 ( .A1(n21295), .A2(keyinput52), .B1(n21294), .B2(keyinput60), 
        .ZN(n21293) );
  OAI221_X1 U24209 ( .B1(n21295), .B2(keyinput52), .C1(n21294), .C2(keyinput60), .A(n21293), .ZN(n21306) );
  AOI22_X1 U24210 ( .A1(n11072), .A2(keyinput42), .B1(keyinput39), .B2(n21297), 
        .ZN(n21296) );
  OAI221_X1 U24211 ( .B1(n11072), .B2(keyinput42), .C1(n21297), .C2(keyinput39), .A(n21296), .ZN(n21305) );
  INV_X1 U24212 ( .A(keyinput32), .ZN(n21302) );
  INV_X1 U24213 ( .A(keyinput127), .ZN(n21299) );
  OAI22_X1 U24214 ( .A1(keyinput92), .A2(n21300), .B1(n21299), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n21298) );
  AOI221_X1 U24215 ( .B1(n21300), .B2(keyinput92), .C1(n21299), .C2(
        P1_DATAO_REG_15__SCAN_IN), .A(n21298), .ZN(n21301) );
  OAI221_X1 U24216 ( .B1(keyinput32), .B2(n21303), .C1(n21302), .C2(
        P3_REIP_REG_2__SCAN_IN), .A(n21301), .ZN(n21304) );
  NOR4_X1 U24217 ( .A1(n21307), .A2(n21306), .A3(n21305), .A4(n21304), .ZN(
        n21322) );
  INV_X1 U24218 ( .A(keyinput118), .ZN(n21309) );
  AOI22_X1 U24219 ( .A1(n21310), .A2(keyinput119), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n21309), .ZN(n21308) );
  OAI221_X1 U24220 ( .B1(n21310), .B2(keyinput119), .C1(n21309), .C2(
        P2_DATAO_REG_11__SCAN_IN), .A(n21308), .ZN(n21320) );
  INV_X1 U24221 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n21312) );
  AOI22_X1 U24222 ( .A1(n10710), .A2(keyinput113), .B1(keyinput40), .B2(n21312), .ZN(n21311) );
  OAI221_X1 U24223 ( .B1(n10710), .B2(keyinput113), .C1(n21312), .C2(
        keyinput40), .A(n21311), .ZN(n21319) );
  AOI22_X1 U24224 ( .A1(n21314), .A2(keyinput99), .B1(n14836), .B2(keyinput11), 
        .ZN(n21313) );
  OAI221_X1 U24225 ( .B1(n21314), .B2(keyinput99), .C1(n14836), .C2(keyinput11), .A(n21313), .ZN(n21318) );
  XNOR2_X1 U24226 ( .A(P2_STATE2_REG_2__SCAN_IN), .B(keyinput26), .ZN(n21316)
         );
  XNOR2_X1 U24227 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput12), 
        .ZN(n21315) );
  NAND2_X1 U24228 ( .A1(n21316), .A2(n21315), .ZN(n21317) );
  NOR4_X1 U24229 ( .A1(n21320), .A2(n21319), .A3(n21318), .A4(n21317), .ZN(
        n21321) );
  NAND4_X1 U24230 ( .A1(n21324), .A2(n21323), .A3(n21322), .A4(n21321), .ZN(
        n21325) );
  NOR4_X1 U24231 ( .A1(n21328), .A2(n21327), .A3(n21326), .A4(n21325), .ZN(
        n21382) );
  NAND2_X1 U24232 ( .A1(keyinput42), .A2(keyinput52), .ZN(n21329) );
  NOR3_X1 U24233 ( .A1(keyinput60), .A2(keyinput39), .A3(n21329), .ZN(n21330)
         );
  NAND3_X1 U24234 ( .A1(keyinput127), .A2(keyinput32), .A3(n21330), .ZN(n21342) );
  NAND2_X1 U24235 ( .A1(keyinput78), .A2(keyinput90), .ZN(n21331) );
  NOR3_X1 U24236 ( .A1(keyinput36), .A2(keyinput54), .A3(n21331), .ZN(n21340)
         );
  NOR4_X1 U24237 ( .A1(keyinput2), .A2(keyinput94), .A3(keyinput22), .A4(
        keyinput0), .ZN(n21339) );
  NAND4_X1 U24238 ( .A1(keyinput122), .A2(keyinput104), .A3(keyinput76), .A4(
        keyinput21), .ZN(n21337) );
  INV_X1 U24239 ( .A(keyinput34), .ZN(n21332) );
  NAND4_X1 U24240 ( .A1(keyinput58), .A2(keyinput51), .A3(keyinput55), .A4(
        n21332), .ZN(n21336) );
  NAND4_X1 U24241 ( .A1(keyinput113), .A2(keyinput40), .A3(keyinput118), .A4(
        keyinput119), .ZN(n21335) );
  NOR3_X1 U24242 ( .A1(keyinput99), .A2(keyinput12), .A3(keyinput11), .ZN(
        n21333) );
  NAND2_X1 U24243 ( .A1(keyinput26), .A2(n21333), .ZN(n21334) );
  NOR4_X1 U24244 ( .A1(n21337), .A2(n21336), .A3(n21335), .A4(n21334), .ZN(
        n21338) );
  NAND3_X1 U24245 ( .A1(n21340), .A2(n21339), .A3(n21338), .ZN(n21341) );
  NOR4_X1 U24246 ( .A1(keyinput92), .A2(keyinput112), .A3(n21342), .A4(n21341), 
        .ZN(n21380) );
  NAND4_X1 U24247 ( .A1(keyinput14), .A2(keyinput3), .A3(keyinput107), .A4(
        keyinput98), .ZN(n21346) );
  NAND4_X1 U24248 ( .A1(keyinput84), .A2(keyinput108), .A3(keyinput47), .A4(
        keyinput59), .ZN(n21345) );
  NAND4_X1 U24249 ( .A1(keyinput71), .A2(keyinput67), .A3(keyinput91), .A4(
        keyinput86), .ZN(n21344) );
  NAND4_X1 U24250 ( .A1(keyinput123), .A2(keyinput103), .A3(keyinput115), .A4(
        keyinput66), .ZN(n21343) );
  NOR4_X1 U24251 ( .A1(n21346), .A2(n21345), .A3(n21344), .A4(n21343), .ZN(
        n21379) );
  NAND4_X1 U24252 ( .A1(keyinput57), .A2(keyinput49), .A3(keyinput69), .A4(
        keyinput77), .ZN(n21351) );
  NOR3_X1 U24253 ( .A1(keyinput114), .A2(keyinput95), .A3(keyinput79), .ZN(
        n21347) );
  NAND2_X1 U24254 ( .A1(keyinput9), .A2(n21347), .ZN(n21350) );
  NAND4_X1 U24255 ( .A1(keyinput20), .A2(keyinput28), .A3(keyinput56), .A4(
        keyinput88), .ZN(n21349) );
  NAND4_X1 U24256 ( .A1(keyinput101), .A2(keyinput97), .A3(keyinput121), .A4(
        keyinput64), .ZN(n21348) );
  NOR4_X1 U24257 ( .A1(n21351), .A2(n21350), .A3(n21349), .A4(n21348), .ZN(
        n21378) );
  NAND4_X1 U24258 ( .A1(keyinput27), .A2(keyinput102), .A3(keyinput7), .A4(
        n21352), .ZN(n21357) );
  NAND4_X1 U24259 ( .A1(keyinput116), .A2(keyinput89), .A3(keyinput4), .A4(
        keyinput44), .ZN(n21356) );
  NOR2_X1 U24260 ( .A1(keyinput70), .A2(keyinput81), .ZN(n21353) );
  NAND3_X1 U24261 ( .A1(keyinput87), .A2(keyinput16), .A3(n21353), .ZN(n21355)
         );
  NAND4_X1 U24262 ( .A1(keyinput85), .A2(keyinput106), .A3(keyinput50), .A4(
        keyinput63), .ZN(n21354) );
  OR4_X1 U24263 ( .A1(n21357), .A2(n21356), .A3(n21355), .A4(n21354), .ZN(
        n21376) );
  NAND3_X1 U24264 ( .A1(keyinput23), .A2(keyinput15), .A3(keyinput61), .ZN(
        n21358) );
  NOR2_X1 U24265 ( .A1(keyinput82), .A2(n21358), .ZN(n21364) );
  NOR4_X1 U24266 ( .A1(keyinput83), .A2(keyinput8), .A3(keyinput62), .A4(
        keyinput74), .ZN(n21363) );
  NAND2_X1 U24267 ( .A1(keyinput13), .A2(keyinput29), .ZN(n21359) );
  NOR3_X1 U24268 ( .A1(keyinput24), .A2(keyinput1), .A3(n21359), .ZN(n21362)
         );
  INV_X1 U24269 ( .A(keyinput75), .ZN(n21360) );
  NOR4_X1 U24270 ( .A1(keyinput37), .A2(keyinput93), .A3(keyinput65), .A4(
        n21360), .ZN(n21361) );
  NAND4_X1 U24271 ( .A1(n21364), .A2(n21363), .A3(n21362), .A4(n21361), .ZN(
        n21375) );
  NOR4_X1 U24272 ( .A1(keyinput46), .A2(keyinput35), .A3(keyinput38), .A4(
        keyinput10), .ZN(n21368) );
  NOR4_X1 U24273 ( .A1(keyinput72), .A2(keyinput80), .A3(keyinput100), .A4(
        keyinput43), .ZN(n21367) );
  NOR4_X1 U24274 ( .A1(keyinput18), .A2(keyinput111), .A3(keyinput110), .A4(
        keyinput126), .ZN(n21366) );
  NOR4_X1 U24275 ( .A1(keyinput6), .A2(keyinput31), .A3(keyinput30), .A4(
        keyinput19), .ZN(n21365) );
  NAND4_X1 U24276 ( .A1(n21368), .A2(n21367), .A3(n21366), .A4(n21365), .ZN(
        n21374) );
  NOR4_X1 U24277 ( .A1(keyinput45), .A2(keyinput53), .A3(keyinput73), .A4(
        keyinput105), .ZN(n21372) );
  NOR4_X1 U24278 ( .A1(keyinput5), .A2(keyinput25), .A3(keyinput33), .A4(
        keyinput41), .ZN(n21371) );
  NOR4_X1 U24279 ( .A1(keyinput124), .A2(keyinput96), .A3(keyinput48), .A4(
        keyinput68), .ZN(n21370) );
  NOR4_X1 U24280 ( .A1(keyinput109), .A2(keyinput117), .A3(keyinput125), .A4(
        keyinput120), .ZN(n21369) );
  NAND4_X1 U24281 ( .A1(n21372), .A2(n21371), .A3(n21370), .A4(n21369), .ZN(
        n21373) );
  NOR4_X1 U24282 ( .A1(n21376), .A2(n21375), .A3(n21374), .A4(n21373), .ZN(
        n21377) );
  NAND4_X1 U24283 ( .A1(n21380), .A2(n21379), .A3(n21378), .A4(n21377), .ZN(
        n21381) );
  NAND4_X1 U24284 ( .A1(n21384), .A2(n21383), .A3(n21382), .A4(n21381), .ZN(
        n21406) );
  OAI21_X1 U24285 ( .B1(n21387), .B2(n21386), .A(n21385), .ZN(n21401) );
  INV_X1 U24286 ( .A(n21388), .ZN(n21397) );
  OAI22_X1 U24287 ( .A1(n21392), .A2(n21391), .B1(n21390), .B2(n21389), .ZN(
        n21394) );
  AOI211_X1 U24288 ( .C1(n21395), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21394), .B(n21393), .ZN(n21396) );
  OAI21_X1 U24289 ( .B1(n21398), .B2(n21397), .A(n21396), .ZN(n21399) );
  AOI21_X1 U24290 ( .B1(n21401), .B2(n21400), .A(n21399), .ZN(n21402) );
  OAI21_X1 U24291 ( .B1(n21404), .B2(n21403), .A(n21402), .ZN(n21405) );
  XNOR2_X1 U24292 ( .A(n21406), .B(n21405), .ZN(P1_U2826) );
  AND2_X1 U15135 ( .A1(n13644), .A2(n11849), .ZN(n11924) );
  INV_X1 U11306 ( .A(n11656), .ZN(n10310) );
  AOI221_X2 U11247 ( .B1(n20912), .B2(n20911), .C1(n20914), .C2(n20915), .A(
        n20910), .ZN(n20976) );
  NOR2_X4 U13677 ( .A1(n10658), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13288) );
  BUF_X2 U11183 ( .A(n11645), .Z(n9718) );
  CLKBUF_X1 U11190 ( .A(n12032), .Z(n12933) );
  OR2_X1 U11224 ( .A1(n11524), .A2(n10155), .ZN(n10154) );
  CLKBUF_X1 U11237 ( .A(n12057), .Z(n12077) );
  CLKBUF_X1 U11257 ( .A(n15112), .Z(n16348) );
  NAND2_X1 U11265 ( .A1(n12020), .A2(n12019), .ZN(n12137) );
  CLKBUF_X1 U11270 ( .A(n11645), .Z(n9719) );
  CLKBUF_X2 U11280 ( .A(n11966), .Z(n13962) );
  CLKBUF_X1 U11284 ( .A(n14783), .Z(n14799) );
  NAND2_X1 U11546 ( .A1(n13693), .A2(n13114), .ZN(n13777) );
  CLKBUF_X1 U11659 ( .A(n10601), .Z(n10603) );
  CLKBUF_X1 U12151 ( .A(n10493), .Z(n19696) );
  CLKBUF_X1 U12201 ( .A(n18197), .Z(n9733) );
  CLKBUF_X1 U12421 ( .A(n12497), .Z(n12498) );
  CLKBUF_X1 U12423 ( .A(n15033), .Z(n15065) );
  CLKBUF_X1 U12479 ( .A(n15096), .Z(n15106) );
  CLKBUF_X1 U12521 ( .A(n13099), .Z(n16001) );
  NOR2_X1 U12755 ( .A1(n10372), .A2(n10371), .ZN(n18552) );
  AND2_X2 U12903 ( .A1(n12198), .A2(n12135), .ZN(n21407) );
endmodule

