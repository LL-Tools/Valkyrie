

module b15_C_AntiSAT_k_256_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380;

  NAND2_X1 U3642 ( .A1(n4351), .A2(n4350), .ZN(n6822) );
  XNOR2_X1 U3643 ( .A(n4514), .B(n4513), .ZN(n6450) );
  NAND2_X1 U3644 ( .A1(n4512), .A2(n4511), .ZN(n4514) );
  BUF_X1 U3645 ( .A(n4304), .Z(n4534) );
  CLKBUF_X2 U3647 ( .A(n3441), .Z(n3722) );
  INV_X1 U3648 ( .A(n4594), .ZN(n3624) );
  CLKBUF_X2 U3649 ( .A(n3430), .Z(n3554) );
  CLKBUF_X2 U3650 ( .A(n3414), .Z(n3635) );
  NAND2_X2 U3651 ( .A1(n3525), .A2(n4806), .ZN(n6204) );
  NAND4_X1 U3652 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3439)
         );
  AND4_X1 U3653 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3348)
         );
  AND4_X1 U3654 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3329)
         );
  AND4_X1 U3655 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3328)
         );
  AND2_X1 U3656 ( .A1(n3320), .A2(n3322), .ZN(n3441) );
  NAND2_X1 U3657 ( .A1(n4952), .A2(n6830), .ZN(n3453) );
  AND2_X2 U3658 ( .A1(n3321), .A2(n3314), .ZN(n4148) );
  AND2_X1 U3659 ( .A1(n3305), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3320)
         );
  AND2_X2 U3660 ( .A1(n4735), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3314)
         );
  NOR2_X2 U3661 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3322) );
  INV_X1 U3662 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3304) );
  CLKBUF_X1 U3663 ( .A(n6990), .Z(n3194) );
  NOR2_X1 U3664 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6877), .ZN(n6990) );
  CLKBUF_X1 U3665 ( .A(n5260), .Z(n3195) );
  AND2_X1 U3666 ( .A1(n5877), .A2(n4573), .ZN(n3196) );
  NAND2_X2 U3667 ( .A1(n3702), .A2(n4889), .ZN(n3197) );
  AND2_X1 U3668 ( .A1(n3540), .A2(n3615), .ZN(n3198) );
  NAND2_X1 U3670 ( .A1(n3702), .A2(n4889), .ZN(n3738) );
  INV_X2 U3671 ( .A(n3703), .ZN(n3702) );
  NAND3_X1 U3672 ( .A1(n3505), .A2(n3504), .A3(n3295), .ZN(n3617) );
  INV_X1 U3673 ( .A(n3510), .ZN(n3525) );
  INV_X1 U3674 ( .A(n4368), .ZN(n4466) );
  NOR2_X2 U3675 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4736) );
  INV_X1 U3678 ( .A(n6357), .ZN(n6343) );
  OR2_X1 U3679 ( .A1(n4816), .A2(n6825), .ZN(n6468) );
  NAND4_X1 U3680 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3468)
         );
  BUF_X1 U3681 ( .A(n3468), .Z(n3201) );
  AND2_X2 U3682 ( .A1(n5127), .A2(n3225), .ZN(n5461) );
  NAND2_X2 U3683 ( .A1(n5852), .A2(n4572), .ZN(n5877) );
  NAND2_X2 U3684 ( .A1(n5920), .A2(n4570), .ZN(n5852) );
  BUF_X4 U3686 ( .A(n3439), .Z(n3522) );
  INV_X2 U3688 ( .A(n3494), .ZN(n3515) );
  NAND4_X4 U3689 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3494)
         );
  NAND2_X2 U3690 ( .A1(n3470), .A2(n3469), .ZN(n3516) );
  AOI21_X1 U3692 ( .B1(n4556), .B2(n3286), .A(n3216), .ZN(n3285) );
  NAND2_X1 U3695 ( .A1(n6380), .A2(n3499), .ZN(n6152) );
  INV_X1 U3696 ( .A(n4360), .ZN(n4394) );
  INV_X4 U3698 ( .A(n4385), .ZN(n4470) );
  INV_X2 U3699 ( .A(n3511), .ZN(n4804) );
  INV_X1 U3700 ( .A(n3499), .ZN(n5811) );
  AND4_X2 U3701 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3511)
         );
  BUF_X2 U3702 ( .A(n3429), .Z(n4156) );
  BUF_X2 U3703 ( .A(n3442), .Z(n3774) );
  AOI22_X1 U3704 ( .A1(n5856), .A2(n5864), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5855), .ZN(n5857) );
  NAND2_X1 U3705 ( .A1(n5927), .A2(n3288), .ZN(n5886) );
  NOR2_X1 U3706 ( .A1(n3242), .A2(n5543), .ZN(n3241) );
  INV_X1 U3707 ( .A(n4560), .ZN(n3242) );
  NOR2_X1 U3708 ( .A1(n3287), .A2(n3284), .ZN(n3283) );
  AND2_X1 U3709 ( .A1(n6433), .A2(n4559), .ZN(n4560) );
  NAND2_X1 U3710 ( .A1(n4561), .A2(n6485), .ZN(n4556) );
  NOR2_X1 U3712 ( .A1(n5125), .A2(n3224), .ZN(n3278) );
  INV_X1 U3713 ( .A(n5126), .ZN(n3279) );
  AOI21_X1 U3714 ( .B1(n4535), .B2(n3953), .A(n3802), .ZN(n5125) );
  XNOR2_X1 U3715 ( .A(n4545), .B(n3797), .ZN(n4535) );
  NOR2_X1 U3716 ( .A1(n5104), .A2(n5266), .ZN(n6809) );
  AND2_X1 U3717 ( .A1(n3677), .A2(n4874), .ZN(n4839) );
  OAI21_X1 U3718 ( .B1(n4978), .B2(n3877), .A(n3712), .ZN(n4841) );
  AND2_X1 U3719 ( .A1(n4767), .A2(n4766), .ZN(n4769) );
  CLKBUF_X1 U3720 ( .A(n4890), .Z(n6073) );
  NAND2_X1 U3721 ( .A1(n3701), .A2(n3700), .ZN(n4889) );
  AND2_X1 U3722 ( .A1(n3666), .A2(n3612), .ZN(n3646) );
  NOR3_X1 U3723 ( .A1(n5796), .A2(n3210), .A3(n3228), .ZN(n5780) );
  NAND2_X2 U3724 ( .A1(n3657), .A2(n3656), .ZN(n4891) );
  NAND2_X1 U3725 ( .A1(n6833), .A2(n6861), .ZN(n3651) );
  NAND2_X1 U3726 ( .A1(n4294), .A2(n3521), .ZN(n3584) );
  NAND2_X1 U3727 ( .A1(n3302), .A2(n3512), .ZN(n4294) );
  NAND2_X1 U3728 ( .A1(n3235), .A2(n3526), .ZN(n3234) );
  INV_X1 U3729 ( .A(n4694), .ZN(n3526) );
  NAND2_X1 U3730 ( .A1(n3685), .A2(n3684), .ZN(n4349) );
  INV_X1 U3731 ( .A(n3685), .ZN(n3643) );
  AND2_X1 U3732 ( .A1(n3214), .A2(n4904), .ZN(n3235) );
  NAND2_X1 U3733 ( .A1(n4310), .A2(n4929), .ZN(n4335) );
  AND2_X2 U3734 ( .A1(n3201), .A2(n4904), .ZN(n4770) );
  AND2_X1 U3735 ( .A1(n3510), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4310) );
  AND2_X2 U3736 ( .A1(n4806), .A2(n3510), .ZN(n4774) );
  NOR2_X2 U3737 ( .A1(n3499), .A2(n3658), .ZN(n4623) );
  NAND4_X2 U3738 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3514)
         );
  AND4_X1 U3739 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3491)
         );
  AND3_X1 U3740 ( .A1(n3461), .A2(n3460), .A3(n3459), .ZN(n3462) );
  AOI21_X1 U3741 ( .B1(n4602), .B2(INSTQUEUE_REG_10__3__SCAN_IN), .A(n3457), 
        .ZN(n3463) );
  AND4_X1 U3742 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3464)
         );
  AND4_X1 U3743 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(n3435)
         );
  AND4_X1 U3744 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3489)
         );
  AND4_X1 U3745 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3436)
         );
  NAND4_X2 U3746 ( .A1(n3392), .A2(n3391), .A3(n3390), .A4(n3389), .ZN(n3499)
         );
  AND4_X1 U3747 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3437)
         );
  AND4_X1 U3748 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3347)
         );
  AND4_X1 U3749 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3349)
         );
  AND4_X1 U3750 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3368)
         );
  AND4_X1 U3751 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  AND4_X1 U3752 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3370)
         );
  AND4_X1 U3753 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3350)
         );
  AND4_X1 U3754 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n3465)
         );
  AND4_X1 U3755 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  AND4_X1 U3756 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3391)
         );
  AND4_X1 U3757 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3392)
         );
  AND4_X1 U3758 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3490)
         );
  AND4_X1 U3759 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3371)
         );
  AND4_X1 U3760 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3369)
         );
  BUF_X2 U3761 ( .A(n3372), .Z(n4273) );
  AND4_X1 U3762 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3438)
         );
  AND4_X1 U3763 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3410)
         );
  AND4_X1 U3764 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3411)
         );
  AND4_X1 U3765 ( .A1(n3217), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3330)
         );
  AND4_X1 U3766 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3327)
         );
  AND4_X1 U3767 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3412)
         );
  NOR2_X1 U3768 ( .A1(n3458), .A2(n3298), .ZN(n3461) );
  CLKBUF_X3 U3769 ( .A(n4265), .Z(n4602) );
  BUF_X2 U3770 ( .A(n3483), .Z(n3542) );
  BUF_X2 U3771 ( .A(n3447), .Z(n4605) );
  BUF_X2 U3772 ( .A(n3447), .Z(n4246) );
  BUF_X2 U3773 ( .A(n3553), .Z(n3723) );
  BUF_X2 U3774 ( .A(n4148), .Z(n4245) );
  AND2_X2 U3775 ( .A1(n3321), .A2(n4736), .ZN(n3419) );
  AND2_X2 U3776 ( .A1(n3314), .A2(n3322), .ZN(n3483) );
  AND2_X2 U3777 ( .A1(n3321), .A2(n4950), .ZN(n3414) );
  BUF_X2 U3778 ( .A(n3424), .Z(n4604) );
  AND2_X2 U3779 ( .A1(n3314), .A2(n3319), .ZN(n3447) );
  AND2_X2 U3780 ( .A1(n3320), .A2(n3321), .ZN(n3413) );
  AND2_X2 U3781 ( .A1(n4949), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3321)
         );
  INV_X1 U3782 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3305) );
  INV_X1 U3783 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6830) );
  INV_X2 U3784 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n3658) );
  AND2_X2 U3785 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4950) );
  AND2_X2 U3786 ( .A1(n3703), .A2(n3650), .ZN(n6580) );
  OAI21_X1 U3787 ( .B1(n5920), .B2(n3290), .A(n3289), .ZN(n3293) );
  AOI21_X1 U3788 ( .B1(n3503), .B2(n3514), .A(n5811), .ZN(n3500) );
  NAND2_X1 U3789 ( .A1(n3281), .A2(n4481), .ZN(n4505) );
  AOI22_X2 U3790 ( .A1(n6458), .A2(n4504), .B1(n4503), .B2(n6564), .ZN(n4939)
         );
  AOI21_X2 U3791 ( .B1(n6580), .B2(n4534), .A(n4486), .ZN(n6458) );
  NAND2_X2 U3792 ( .A1(n3282), .A2(n3285), .ZN(n5534) );
  INV_X1 U3793 ( .A(n3554), .ZN(n3202) );
  NAND2_X4 U3795 ( .A1(n3678), .A2(n3623), .ZN(n4755) );
  XNOR2_X1 U3796 ( .A(n3678), .B(n6654), .ZN(n4892) );
  OAI21_X2 U3797 ( .B1(n5580), .B2(n5581), .A(n5582), .ZN(n5945) );
  AND2_X1 U3798 ( .A1(n3320), .A2(n3322), .ZN(n3205) );
  NAND2_X1 U3799 ( .A1(n3525), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3685) );
  INV_X2 U3800 ( .A(n3200), .ZN(n4806) );
  NOR2_X1 U3801 ( .A1(n5710), .A2(n5723), .ZN(n3276) );
  OR2_X1 U3802 ( .A1(n3561), .A2(n3560), .ZN(n4494) );
  NAND2_X1 U3803 ( .A1(n3511), .A2(n3514), .ZN(n4495) );
  INV_X1 U3804 ( .A(n3514), .ZN(n4352) );
  INV_X1 U3805 ( .A(n5785), .ZN(n3270) );
  INV_X1 U3806 ( .A(n3758), .ZN(n4621) );
  NAND2_X1 U3807 ( .A1(n5877), .A2(n4573), .ZN(n4575) );
  INV_X1 U3808 ( .A(n5878), .ZN(n4573) );
  NOR2_X1 U3809 ( .A1(n5377), .A2(n3255), .ZN(n3254) );
  INV_X1 U3810 ( .A(n5254), .ZN(n3255) );
  INV_X1 U3811 ( .A(n4335), .ZN(n4305) );
  OR2_X1 U3812 ( .A1(n4929), .A2(n6861), .ZN(n3684) );
  OR2_X1 U3813 ( .A1(n4335), .A2(n4288), .ZN(n3295) );
  INV_X1 U3814 ( .A(n4774), .ZN(n6984) );
  AND2_X1 U3815 ( .A1(n3276), .A2(n3275), .ZN(n3274) );
  INV_X1 U3816 ( .A(n4285), .ZN(n3275) );
  OR2_X1 U3817 ( .A1(n6822), .A2(n6865), .ZN(n4816) );
  AND2_X1 U3818 ( .A1(n3209), .A2(n4566), .ZN(n3288) );
  NOR2_X1 U3819 ( .A1(n5920), .A2(n5919), .ZN(n5918) );
  NAND2_X1 U3820 ( .A1(n3244), .A2(n5541), .ZN(n6166) );
  NAND2_X1 U3821 ( .A1(n3243), .A2(n3241), .ZN(n3244) );
  AND2_X1 U3822 ( .A1(n6952), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4357) );
  INV_X1 U3823 ( .A(n4953), .ZN(n3309) );
  AND2_X2 U3824 ( .A1(n3304), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3319)
         );
  OR2_X1 U3825 ( .A1(n3578), .A2(n3577), .ZN(n4539) );
  OR2_X1 U3826 ( .A1(n3453), .A2(n5490), .ZN(n3478) );
  AND2_X1 U3827 ( .A1(n4025), .A2(n3273), .ZN(n3272) );
  INV_X1 U3828 ( .A(n5736), .ZN(n3273) );
  INV_X1 U3829 ( .A(n5733), .ZN(n3271) );
  INV_X1 U3830 ( .A(n4618), .ZN(n4282) );
  AND2_X1 U3831 ( .A1(n6831), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4618) );
  NOR2_X1 U3832 ( .A1(n5762), .A2(n3264), .ZN(n3263) );
  INV_X1 U3833 ( .A(n4687), .ZN(n3264) );
  AOI21_X1 U3834 ( .B1(n5919), .B2(n3292), .A(n3296), .ZN(n3291) );
  INV_X1 U3835 ( .A(n3301), .ZN(n3292) );
  NOR2_X1 U3836 ( .A1(n4548), .A2(n4547), .ZN(n4549) );
  OR2_X1 U3837 ( .A1(n6196), .A2(n6065), .ZN(n3251) );
  NAND2_X1 U3838 ( .A1(n3530), .A2(n3529), .ZN(n4295) );
  AND3_X1 U3839 ( .A1(n3351), .A2(n4352), .A3(n3511), .ZN(n3529) );
  INV_X1 U3840 ( .A(n4287), .ZN(n3524) );
  XNOR2_X1 U3841 ( .A(n3609), .B(n3610), .ZN(n3662) );
  NAND2_X1 U3842 ( .A1(n3508), .A2(n3507), .ZN(n3583) );
  AND4_X1 U3843 ( .A1(n3513), .A2(n6868), .A3(n3520), .A4(n3519), .ZN(n3521)
         );
  NAND2_X1 U3844 ( .A1(n3583), .A2(n3584), .ZN(n3614) );
  OR2_X1 U3845 ( .A1(n4978), .A2(n6580), .ZN(n5268) );
  AND2_X1 U3846 ( .A1(n3619), .A2(n6740), .ZN(n5010) );
  INV_X1 U3847 ( .A(n5151), .ZN(n5054) );
  NAND4_X2 U3848 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3435), .ZN(n3510)
         );
  INV_X1 U3849 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6844) );
  INV_X1 U3850 ( .A(n6825), .ZN(n3238) );
  AND2_X1 U3851 ( .A1(n4663), .A2(n4662), .ZN(n6820) );
  AND2_X1 U3852 ( .A1(n4654), .A2(n4655), .ZN(n6819) );
  AND3_X1 U3853 ( .A1(n3502), .A2(n3500), .A3(n3501), .ZN(n4654) );
  NAND2_X1 U3854 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6333), .ZN(n5294) );
  INV_X1 U3855 ( .A(n6269), .ZN(n3253) );
  AND2_X1 U3856 ( .A1(n3267), .A2(n3266), .ZN(n3265) );
  INV_X1 U3857 ( .A(n4683), .ZN(n3266) );
  AOI21_X1 U3858 ( .B1(n6580), .B2(n3953), .A(n4622), .ZN(n4875) );
  NAND2_X1 U3859 ( .A1(n4360), .A2(n4385), .ZN(n5658) );
  OAI21_X1 U3860 ( .B1(n5620), .B2(n4470), .A(n3303), .ZN(n5654) );
  OR2_X1 U3861 ( .A1(n4467), .A2(n4469), .ZN(n5620) );
  NOR2_X1 U3862 ( .A1(n5757), .A2(n5725), .ZN(n5727) );
  NAND2_X1 U3863 ( .A1(n5851), .A2(n3300), .ZN(n5865) );
  AND2_X1 U3864 ( .A1(n5780), .A2(n5773), .ZN(n5775) );
  AND2_X1 U3865 ( .A1(n4443), .A2(n4442), .ZN(n5779) );
  INV_X1 U3866 ( .A(n6029), .ZN(n4435) );
  OR2_X1 U3867 ( .A1(n3204), .A2(n4567), .ZN(n4568) );
  OR2_X1 U3868 ( .A1(n3221), .A2(n5739), .ZN(n5796) );
  INV_X1 U3869 ( .A(n4554), .ZN(n3286) );
  NAND2_X1 U3870 ( .A1(n3260), .A2(n3261), .ZN(n4879) );
  AND2_X1 U3871 ( .A1(n4909), .A2(n3499), .ZN(n5684) );
  INV_X1 U3872 ( .A(n4770), .ZN(n5657) );
  CLKBUF_X1 U3873 ( .A(n4694), .Z(n4695) );
  NAND2_X1 U3874 ( .A1(n4818), .A2(n4817), .ZN(n4831) );
  OR2_X1 U3875 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  OAI21_X2 U3876 ( .B1(n4891), .B2(n4547), .A(n4489), .ZN(n6467) );
  OR2_X1 U3877 ( .A1(n4478), .A2(n3684), .ZN(n3642) );
  INV_X1 U3878 ( .A(n4891), .ZN(n5266) );
  BUF_X1 U3879 ( .A(n3494), .Z(n4909) );
  AND2_X1 U3880 ( .A1(n6580), .A2(n4889), .ZN(n4976) );
  NAND2_X1 U3881 ( .A1(n4349), .A2(n4656), .ZN(n4350) );
  NAND2_X1 U3882 ( .A1(n4348), .A2(n4347), .ZN(n4351) );
  CLKBUF_X1 U3883 ( .A(n4892), .Z(n4893) );
  XNOR2_X1 U3884 ( .A(n4365), .B(n4788), .ZN(n6363) );
  AND2_X1 U3885 ( .A1(n4358), .A2(n6867), .ZN(n6380) );
  AND2_X1 U3886 ( .A1(n6394), .A2(n5685), .ZN(n6387) );
  INV_X1 U3887 ( .A(n6394), .ZN(n6386) );
  NOR2_X1 U3888 ( .A1(n4286), .A2(n4644), .ZN(n5849) );
  INV_X1 U3889 ( .A(n6474), .ZN(n6456) );
  INV_X1 U3890 ( .A(n3452), .ZN(n3543) );
  INV_X1 U3891 ( .A(n4265), .ZN(n3768) );
  NAND2_X1 U3892 ( .A1(n4353), .A2(n4826), .ZN(n3498) );
  OR2_X1 U3893 ( .A1(n3755), .A2(n3754), .ZN(n4525) );
  OR2_X1 U3894 ( .A1(n3780), .A2(n3779), .ZN(n4537) );
  OR2_X1 U3895 ( .A1(n3729), .A2(n3728), .ZN(n4526) );
  AND2_X1 U3896 ( .A1(n3522), .A2(n3468), .ZN(n4304) );
  NAND2_X1 U3897 ( .A1(n3214), .A2(n3351), .ZN(n3492) );
  OR2_X1 U3898 ( .A1(n3453), .A2(n5511), .ZN(n3418) );
  OR2_X1 U3899 ( .A1(n3699), .A2(n3698), .ZN(n4508) );
  NAND2_X1 U3900 ( .A1(n4305), .A2(n4534), .ZN(n4338) );
  NOR2_X1 U3901 ( .A1(n5771), .A2(n3268), .ZN(n3267) );
  INV_X1 U3902 ( .A(n5778), .ZN(n3268) );
  NAND2_X1 U3903 ( .A1(n3980), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4002)
         );
  INV_X1 U3904 ( .A(n5253), .ZN(n3280) );
  INV_X1 U3905 ( .A(n5360), .ZN(n3284) );
  INV_X1 U3906 ( .A(n4556), .ZN(n3287) );
  NAND2_X1 U3907 ( .A1(n4770), .A2(n4385), .ZN(n4461) );
  INV_X1 U3908 ( .A(n4842), .ZN(n3259) );
  OR2_X1 U3909 ( .A1(n3602), .A2(n3601), .ZN(n4493) );
  OR2_X1 U3910 ( .A1(n3641), .A2(n3640), .ZN(n4483) );
  AND3_X1 U3911 ( .A1(n3582), .A2(n3581), .A3(n3580), .ZN(n3610) );
  AOI21_X1 U3912 ( .B1(n3617), .B2(n4954), .A(n3537), .ZN(n3539) );
  OR2_X1 U3913 ( .A1(n3503), .A2(n3961), .ZN(n4581) );
  INV_X1 U3914 ( .A(n6073), .ZN(n5047) );
  OR2_X1 U3915 ( .A1(n3453), .A2(n5502), .ZN(n3454) );
  AND2_X1 U3916 ( .A1(n3553), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3458) );
  OAI21_X1 U3917 ( .B1(n6985), .B2(n4984), .A(n6953), .ZN(n4897) );
  INV_X1 U3918 ( .A(n4338), .ZN(n4346) );
  AND2_X1 U3919 ( .A1(n4345), .A2(n4344), .ZN(n4656) );
  OR2_X1 U3920 ( .A1(n4343), .A2(n4342), .ZN(n4345) );
  AND2_X1 U3921 ( .A1(n7293), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4342)
         );
  INV_X1 U3922 ( .A(n5899), .ZN(n6112) );
  NAND2_X1 U3923 ( .A1(n3260), .A2(n3257), .ZN(n4994) );
  AND2_X1 U3924 ( .A1(n3261), .A2(n3258), .ZN(n3257) );
  AND2_X1 U3925 ( .A1(n3259), .A2(n6318), .ZN(n3258) );
  OR2_X1 U3926 ( .A1(n6817), .A2(n6207), .ZN(n4728) );
  AND2_X1 U3927 ( .A1(n3860), .A2(n3859), .ZN(n5528) );
  AND2_X1 U3928 ( .A1(n4214), .A2(n4213), .ZN(n5753) );
  OR2_X1 U3929 ( .A1(n6089), .A2(n3758), .ZN(n4214) );
  OR2_X1 U3930 ( .A1(n4144), .A2(n7223), .ZN(n4190) );
  NOR2_X1 U3931 ( .A1(n4089), .A2(n4088), .ZN(n4110) );
  NAND2_X1 U3932 ( .A1(n5913), .A2(n3211), .ZN(n3269) );
  NAND2_X1 U3933 ( .A1(n4046), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4089)
         );
  NOR2_X1 U3934 ( .A1(n4002), .A2(n5740), .ZN(n4003) );
  AND2_X1 U3935 ( .A1(n4003), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4045)
         );
  CLKBUF_X1 U3936 ( .A(n5733), .Z(n5807) );
  OR2_X1 U3937 ( .A1(n3941), .A2(n5571), .ZN(n3960) );
  AND2_X1 U3938 ( .A1(n3886), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3883)
         );
  NAND2_X1 U3939 ( .A1(n3883), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3941)
         );
  NAND2_X1 U3940 ( .A1(n3861), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3842)
         );
  NOR2_X1 U3941 ( .A1(n3841), .A2(n3840), .ZN(n3861) );
  NAND2_X1 U3942 ( .A1(n3279), .A2(n3277), .ZN(n5371) );
  NOR2_X1 U3943 ( .A1(n5125), .A2(n3280), .ZN(n3277) );
  AND2_X1 U3944 ( .A1(n3798), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3821)
         );
  NOR2_X1 U3945 ( .A1(n3785), .A2(n5092), .ZN(n3786) );
  AOI21_X1 U3946 ( .B1(n4524), .B2(n3953), .A(n3790), .ZN(n5096) );
  AND2_X1 U3947 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3705), .ZN(n3732)
         );
  NAND2_X1 U3948 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3706) );
  MUX2_X1 U3949 ( .A(n4789), .B(n4621), .S(n4790), .Z(n4767) );
  NAND2_X1 U3950 ( .A1(n5775), .A2(n3229), .ZN(n5757) );
  INV_X1 U3951 ( .A(n5755), .ZN(n3262) );
  NAND2_X1 U3952 ( .A1(n5775), .A2(n3263), .ZN(n5765) );
  OR2_X1 U3953 ( .A1(n6007), .A2(n5628), .ZN(n5988) );
  NAND2_X1 U3954 ( .A1(n3204), .A2(n4571), .ZN(n4572) );
  NAND2_X1 U3955 ( .A1(n5775), .A2(n4687), .ZN(n5763) );
  INV_X1 U3956 ( .A(n3293), .ZN(n5906) );
  INV_X1 U3957 ( .A(n3291), .ZN(n3290) );
  AOI21_X1 U3958 ( .B1(n3291), .B2(n3301), .A(n3223), .ZN(n3289) );
  AND2_X1 U3959 ( .A1(n4431), .A2(n5787), .ZN(n6029) );
  AND2_X1 U3960 ( .A1(n4430), .A2(n4429), .ZN(n5791) );
  OR2_X1 U3961 ( .A1(n3252), .A2(n3250), .ZN(n3249) );
  INV_X1 U3962 ( .A(n5808), .ZN(n3250) );
  INV_X1 U3963 ( .A(n5569), .ZN(n3252) );
  NOR3_X1 U3964 ( .A1(n6195), .A2(n3251), .A3(n3252), .ZN(n6064) );
  CLKBUF_X1 U3965 ( .A(n5927), .Z(n5928) );
  AND2_X1 U3966 ( .A1(n4831), .A2(n4824), .ZN(n5588) );
  NAND2_X1 U3967 ( .A1(n5461), .A2(n5462), .ZN(n6195) );
  NOR2_X1 U3968 ( .A1(n6195), .A2(n6196), .ZN(n6194) );
  NAND2_X1 U3969 ( .A1(n5534), .A2(n3208), .ZN(n3243) );
  NOR2_X1 U3970 ( .A1(n5550), .A2(n5552), .ZN(n5597) );
  NAND2_X1 U3971 ( .A1(n5127), .A2(n5254), .ZN(n5376) );
  NAND2_X1 U3972 ( .A1(n6443), .A2(n6442), .ZN(n3233) );
  INV_X1 U3973 ( .A(n6550), .ZN(n6527) );
  NOR2_X1 U3974 ( .A1(n4367), .A2(n3256), .ZN(n6319) );
  NAND2_X1 U3975 ( .A1(n3261), .A2(n3259), .ZN(n3256) );
  NOR2_X1 U3976 ( .A1(n5605), .A2(n5588), .ZN(n5599) );
  OR2_X1 U3977 ( .A1(n5588), .A2(n5611), .ZN(n5607) );
  INV_X1 U3978 ( .A(n5585), .ZN(n5605) );
  CLKBUF_X1 U3979 ( .A(n4730), .Z(n6350) );
  AOI21_X1 U3980 ( .B1(n3199), .B2(n4955), .A(n3620), .ZN(n3621) );
  NAND2_X1 U3981 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  INV_X1 U3982 ( .A(n3584), .ZN(n3585) );
  INV_X1 U3983 ( .A(n6835), .ZN(n4965) );
  NOR2_X1 U3984 ( .A1(n5268), .A2(n6073), .ZN(n5274) );
  INV_X1 U3985 ( .A(n5268), .ZN(n6745) );
  NAND2_X1 U3986 ( .A1(n4976), .A2(n5047), .ZN(n5104) );
  AND2_X1 U3987 ( .A1(n6943), .A2(n4897), .ZN(n4930) );
  AND2_X1 U3988 ( .A1(n4976), .A2(n6649), .ZN(n5207) );
  OR2_X1 U3989 ( .A1(n4721), .A2(n4584), .ZN(n6825) );
  OAI21_X1 U3990 ( .B1(n6205), .B2(n6820), .A(n3236), .ZN(n6206) );
  NAND2_X1 U3991 ( .A1(n6818), .A2(n3237), .ZN(n6821) );
  AOI21_X1 U3992 ( .B1(n5697), .B2(REIP_REG_31__SCAN_IN), .A(n5696), .ZN(n3247) );
  AND2_X1 U3993 ( .A1(n6137), .A2(n4679), .ZN(n6103) );
  AND2_X1 U3994 ( .A1(n6234), .A2(n4676), .ZN(n6125) );
  NOR2_X1 U3995 ( .A1(n7268), .A2(n5568), .ZN(n6244) );
  INV_X1 U3996 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U3997 ( .A1(n5127), .A2(n3207), .ZN(n6268) );
  NOR2_X1 U3998 ( .A1(n6334), .A2(n4673), .ZN(n6289) );
  NOR2_X2 U3999 ( .A1(n4686), .A2(n4685), .ZN(n6315) );
  AND2_X1 U4000 ( .A1(n4770), .A2(n4690), .ZN(n6322) );
  AND2_X1 U4001 ( .A1(n4689), .A2(n5692), .ZN(n4690) );
  NAND2_X1 U4002 ( .A1(n6333), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6354) );
  INV_X1 U4003 ( .A(n6322), .ZN(n6362) );
  AND2_X1 U4004 ( .A1(n4671), .A2(n5352), .ZN(n6346) );
  AND2_X1 U4005 ( .A1(n4686), .A2(n4680), .ZN(n6357) );
  INV_X1 U4006 ( .A(n6354), .ZN(n6332) );
  NOR2_X1 U4007 ( .A1(n4367), .A2(n4366), .ZN(n4878) );
  INV_X1 U4008 ( .A(n6380), .ZN(n5802) );
  NAND2_X1 U4009 ( .A1(n4887), .A2(n4799), .ZN(n6394) );
  INV_X1 U4010 ( .A(n6390), .ZN(n5577) );
  INV_X1 U4011 ( .A(n4886), .ZN(n6430) );
  XNOR2_X1 U4012 ( .A(n4629), .B(n5695), .ZN(n4686) );
  OR2_X1 U4013 ( .A1(n4628), .A2(n4645), .ZN(n4629) );
  NAND2_X1 U4014 ( .A1(n3213), .A2(n5711), .ZN(n5858) );
  AND2_X1 U4015 ( .A1(n5784), .A2(n5795), .ZN(n6381) );
  NAND2_X1 U4016 ( .A1(n5534), .A2(n5535), .ZN(n6434) );
  INV_X1 U4017 ( .A(n6468), .ZN(n6460) );
  INV_X2 U4018 ( .A(n6470), .ZN(n6461) );
  NAND2_X1 U4019 ( .A1(n6468), .A2(n4630), .ZN(n6474) );
  XNOR2_X1 U4020 ( .A(n5660), .B(n5659), .ZN(n5748) );
  XNOR2_X1 U4021 ( .A(n4580), .B(n4579), .ZN(n5669) );
  NOR2_X1 U4022 ( .A1(n5988), .A2(n5990), .ZN(n5983) );
  INV_X1 U4023 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7174) );
  AOI22_X1 U4024 ( .A1(n5888), .A2(n5889), .B1(n5641), .B2(n5640), .ZN(n5642)
         );
  NOR2_X1 U4025 ( .A1(n4555), .A2(n5637), .ZN(n5641) );
  NOR2_X1 U4026 ( .A1(n5918), .A2(n3301), .ZN(n5912) );
  NAND2_X1 U4027 ( .A1(n4831), .A2(n4829), .ZN(n6551) );
  INV_X1 U4028 ( .A(n6478), .ZN(n6571) );
  INV_X1 U4029 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U4030 ( .A1(n3655), .A2(n3654), .ZN(n3656) );
  NAND2_X1 U4031 ( .A1(n3653), .A2(n3652), .ZN(n3657) );
  INV_X1 U4032 ( .A(n6350), .ZN(n6074) );
  NAND2_X1 U4033 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  AND2_X1 U4034 ( .A1(n6073), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6744) );
  INV_X1 U4035 ( .A(n6753), .ZN(n6658) );
  INV_X1 U4036 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7293) );
  INV_X1 U4037 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U4038 ( .A1(n7315), .A2(n6952), .ZN(n6962) );
  INV_X1 U4039 ( .A(n6622), .ZN(n5088) );
  NOR2_X2 U4040 ( .A1(n5386), .A2(n5266), .ZN(n6621) );
  NOR2_X1 U4041 ( .A1(n5386), .A2(n4891), .ZN(n6644) );
  NAND2_X1 U4042 ( .A1(n6745), .A2(n6649), .ZN(n7370) );
  INV_X1 U4043 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5511) );
  INV_X1 U4044 ( .A(n6741), .ZN(n6698) );
  INV_X1 U4045 ( .A(n6761), .ZN(n6711) );
  INV_X1 U4046 ( .A(n6768), .ZN(n6715) );
  INV_X1 U4047 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5502) );
  INV_X1 U4048 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5494) );
  INV_X1 U4049 ( .A(n7368), .ZN(n6723) );
  INV_X1 U4050 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5498) );
  INV_X1 U4051 ( .A(n6782), .ZN(n6727) );
  INV_X1 U4052 ( .A(n6789), .ZN(n6800) );
  INV_X1 U4053 ( .A(n6794), .ZN(n6808) );
  INV_X1 U4054 ( .A(n5483), .ZN(n5525) );
  AND3_X1 U4055 ( .A1(n5479), .A2(n6753), .A3(n5486), .ZN(n5481) );
  INV_X1 U4056 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6861) );
  INV_X1 U4057 ( .A(n6867), .ZN(n6865) );
  OR2_X1 U4058 ( .A1(n6822), .A2(n7315), .ZN(n6953) );
  INV_X1 U4059 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7315) );
  INV_X1 U4060 ( .A(n6874), .ZN(n6946) );
  INV_X1 U4061 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6877) );
  CLKBUF_X1 U4062 ( .A(n6974), .Z(n6936) );
  NAND2_X1 U4063 ( .A1(n3248), .A2(n3245), .ZN(U2796) );
  OR2_X1 U4064 ( .A1(n5748), .A2(n6362), .ZN(n3248) );
  INV_X1 U4065 ( .A(n3246), .ZN(n3245) );
  OAI211_X1 U4066 ( .C1(n5700), .C2(n5699), .A(n5698), .B(n3247), .ZN(n3246)
         );
  AOI21_X1 U4067 ( .B1(n4475), .B2(n4474), .A(n4473), .ZN(n4476) );
  NOR2_X1 U4068 ( .A1(n6380), .A2(n5701), .ZN(n4473) );
  AND2_X1 U4069 ( .A1(n3271), .A2(n3211), .ZN(n3206) );
  NAND2_X1 U4070 ( .A1(n5777), .A2(n5778), .ZN(n5770) );
  AND2_X1 U4071 ( .A1(n3254), .A2(n5459), .ZN(n3207) );
  AND2_X1 U4072 ( .A1(n3219), .A2(n5535), .ZN(n3208) );
  AND2_X1 U4073 ( .A1(n3218), .A2(n4565), .ZN(n3209) );
  NAND2_X1 U4074 ( .A1(n4437), .A2(n4436), .ZN(n3210) );
  AND2_X1 U4075 ( .A1(n3272), .A2(n3270), .ZN(n3211) );
  OR3_X1 U4076 ( .A1(n5796), .A2(n3210), .A3(n3227), .ZN(n3212) );
  NAND2_X1 U4077 ( .A1(n4545), .A2(n4549), .ZN(n4561) );
  INV_X1 U4078 ( .A(n3414), .ZN(n3440) );
  AND2_X1 U4079 ( .A1(n5777), .A2(n3265), .ZN(n4681) );
  NOR2_X1 U4080 ( .A1(n5733), .A2(n3269), .ZN(n5902) );
  NAND2_X1 U4081 ( .A1(n4236), .A2(n4235), .ZN(n5709) );
  AND2_X1 U4082 ( .A1(n5927), .A2(n3209), .ZN(n5924) );
  AND2_X1 U4083 ( .A1(n4681), .A2(n5760), .ZN(n5752) );
  NAND2_X1 U4084 ( .A1(n4236), .A2(n3276), .ZN(n3213) );
  AND2_X1 U4085 ( .A1(n5902), .A2(n5903), .ZN(n5777) );
  OR2_X1 U4086 ( .A1(n3201), .A2(n4653), .ZN(n3214) );
  INV_X1 U4087 ( .A(n4826), .ZN(n4929) );
  AND4_X2 U4088 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n4826)
         );
  AND2_X1 U4089 ( .A1(n4826), .A2(n3499), .ZN(n3215) );
  AND2_X1 U4090 ( .A1(n3467), .A2(n4732), .ZN(n3513) );
  NOR2_X1 U4091 ( .A1(n3203), .A2(n6485), .ZN(n3216) );
  INV_X1 U4092 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U4093 ( .A1(n5777), .A2(n3267), .ZN(n4682) );
  OR2_X1 U4094 ( .A1(n3453), .A2(n5498), .ZN(n3217) );
  NAND2_X1 U4095 ( .A1(n3271), .A2(n3272), .ZN(n5784) );
  NAND2_X1 U4096 ( .A1(n3203), .A2(n7164), .ZN(n3218) );
  NAND2_X1 U4097 ( .A1(n3204), .A2(n4558), .ZN(n3219) );
  AND2_X1 U4098 ( .A1(n5927), .A2(n4565), .ZN(n3220) );
  NAND2_X1 U4099 ( .A1(n3197), .A2(n3704), .ZN(n4978) );
  OR3_X1 U4100 ( .A1(n6195), .A2(n3251), .A3(n3249), .ZN(n3221) );
  AND2_X1 U4101 ( .A1(n3233), .A2(n3232), .ZN(n3222) );
  NAND2_X1 U4102 ( .A1(n5727), .A2(n5712), .ZN(n4467) );
  NAND2_X1 U4103 ( .A1(n5359), .A2(n4554), .ZN(n5471) );
  NAND2_X1 U4104 ( .A1(n3243), .A2(n4560), .ZN(n5540) );
  AND2_X1 U4105 ( .A1(n4555), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4106 ( .A1(n5361), .A2(n5360), .ZN(n5359) );
  OR3_X1 U4107 ( .A1(n3882), .A2(n3280), .A3(n5372), .ZN(n3224) );
  NOR2_X1 U4108 ( .A1(n5126), .A2(n5125), .ZN(n5252) );
  NAND2_X1 U4109 ( .A1(n4353), .A2(n3215), .ZN(n4287) );
  NOR2_X1 U4110 ( .A1(n5733), .A2(n5736), .ZN(n5734) );
  INV_X1 U4111 ( .A(n5723), .ZN(n4235) );
  AND2_X1 U4112 ( .A1(n4067), .A2(n4066), .ZN(n5913) );
  OAI21_X1 U4113 ( .B1(n4368), .B2(EBX_REG_1__SCAN_IN), .A(n4362), .ZN(n4365)
         );
  AND2_X1 U4114 ( .A1(n3207), .A2(n3253), .ZN(n3225) );
  AND2_X1 U4116 ( .A1(n4877), .A2(n4365), .ZN(n3261) );
  INV_X1 U4117 ( .A(n4367), .ZN(n3260) );
  NOR2_X1 U4118 ( .A1(n4994), .A2(n4995), .ZN(n4996) );
  AND2_X1 U4119 ( .A1(n5127), .A2(n3254), .ZN(n3226) );
  OR2_X1 U4120 ( .A1(n5791), .A2(n6020), .ZN(n3227) );
  NOR2_X1 U4121 ( .A1(n5128), .A2(n5129), .ZN(n5127) );
  OR2_X1 U4122 ( .A1(n3227), .A2(n5779), .ZN(n3228) );
  AND2_X1 U4123 ( .A1(n3263), .A2(n3262), .ZN(n3229) );
  OR3_X1 U4124 ( .A1(n5796), .A2(n3210), .A3(n5791), .ZN(n3230) );
  OR3_X1 U4125 ( .A1(n6195), .A2(n3252), .A3(n6196), .ZN(n3231) );
  INV_X1 U4126 ( .A(n3236), .ZN(n3239) );
  NAND2_X1 U4127 ( .A1(n3526), .A2(n4904), .ZN(n3236) );
  INV_X1 U4128 ( .A(n4623), .ZN(n4616) );
  NAND2_X1 U4129 ( .A1(n3233), .A2(n4533), .ZN(n5262) );
  OR2_X1 U4130 ( .A1(n6443), .A2(n6442), .ZN(n3232) );
  NAND3_X1 U4131 ( .A1(n4819), .A2(n4715), .A3(n3234), .ZN(n3531) );
  NOR2_X1 U4132 ( .A1(n3238), .A2(n3239), .ZN(n3237) );
  NAND2_X1 U4133 ( .A1(n3240), .A2(n3239), .ZN(n4778) );
  INV_X1 U4134 ( .A(n4816), .ZN(n3240) );
  NAND2_X1 U4135 ( .A1(n6166), .A2(n6167), .ZN(n4564) );
  AND2_X2 U4136 ( .A1(n5886), .A2(n4568), .ZN(n5920) );
  OR2_X2 U4137 ( .A1(n5945), .A2(n5947), .ZN(n5927) );
  NOR2_X2 U4138 ( .A1(n5865), .A2(n5972), .ZN(n5844) );
  AND2_X2 U4139 ( .A1(n4575), .A2(n4574), .ZN(n5851) );
  NOR2_X1 U4140 ( .A1(n5796), .A2(n5791), .ZN(n6031) );
  AND2_X2 U4141 ( .A1(n4236), .A2(n3274), .ZN(n4644) );
  AND2_X2 U4142 ( .A1(n3279), .A2(n3278), .ZN(n6168) );
  NAND3_X1 U4143 ( .A1(n3279), .A2(n3278), .A3(n3922), .ZN(n6171) );
  NAND3_X1 U4144 ( .A1(n3197), .A2(n3704), .A3(n4534), .ZN(n3281) );
  NAND4_X1 U4145 ( .A1(n3502), .A2(n3500), .A3(n3501), .A4(n4806), .ZN(n3527)
         );
  NAND2_X1 U4146 ( .A1(n5361), .A2(n3283), .ZN(n3282) );
  NAND2_X2 U4147 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4953) );
  AND2_X2 U4148 ( .A1(n4736), .A2(n3309), .ZN(n3372) );
  OR2_X1 U4149 ( .A1(n5654), .A2(n4472), .ZN(n5962) );
  NAND2_X1 U4150 ( .A1(n4304), .A2(n4826), .ZN(n3509) );
  OR2_X1 U4151 ( .A1(n5748), .A2(n6551), .ZN(n5668) );
  INV_X1 U4152 ( .A(n5877), .ZN(n5879) );
  AOI22_X1 U4153 ( .A1(n5844), .A2(n4578), .B1(n3196), .B2(n4577), .ZN(n4580)
         );
  INV_X1 U4154 ( .A(n3583), .ZN(n3586) );
  NAND2_X1 U4155 ( .A1(n3527), .A2(n3643), .ZN(n3504) );
  NAND2_X2 U4156 ( .A1(n3351), .A2(n3494), .ZN(n4353) );
  NAND2_X1 U4157 ( .A1(n5091), .A2(n5090), .ZN(n5089) );
  XNOR2_X1 U4158 ( .A(n4642), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5636)
         );
  NAND2_X1 U4159 ( .A1(n4641), .A2(n4640), .ZN(n4642) );
  INV_X1 U4160 ( .A(n3413), .ZN(n3572) );
  AND2_X1 U4161 ( .A1(n5668), .A2(n5667), .ZN(n3294) );
  OR2_X1 U4162 ( .A1(n4634), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U4163 ( .A1(n6380), .A2(n5811), .ZN(n6371) );
  INV_X1 U4164 ( .A(n6371), .ZN(n4474) );
  INV_X1 U4165 ( .A(n6152), .ZN(n4359) );
  AND2_X1 U4166 ( .A1(n6170), .A2(n5460), .ZN(n3922) );
  INV_X1 U4167 ( .A(n5372), .ZN(n5373) );
  AND2_X1 U4168 ( .A1(n3203), .A2(n5910), .ZN(n3296) );
  OR3_X1 U4169 ( .A1(n5959), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5664), 
        .ZN(n3297) );
  AND2_X1 U4170 ( .A1(n3372), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3298) );
  OR2_X1 U4171 ( .A1(n3537), .A2(n4954), .ZN(n3299) );
  AND2_X1 U4172 ( .A1(n3204), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3300)
         );
  INV_X1 U4173 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6272) );
  AND2_X1 U4174 ( .A1(n4555), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3301)
         );
  NAND2_X1 U4175 ( .A1(n3204), .A2(n5997), .ZN(n4574) );
  INV_X1 U4176 ( .A(n6204), .ZN(n3530) );
  AND2_X1 U4177 ( .A1(n3509), .A2(n3527), .ZN(n3302) );
  OR2_X1 U4178 ( .A1(n4467), .A2(n4468), .ZN(n3303) );
  INV_X1 U4179 ( .A(n5962), .ZN(n4475) );
  AND2_X2 U4180 ( .A1(n3322), .A2(n4950), .ZN(n3424) );
  INV_X1 U4181 ( .A(n3542), .ZN(n4594) );
  INV_X1 U4182 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4949) );
  INV_X1 U4183 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4242) );
  INV_X1 U4184 ( .A(n3503), .ZN(n4288) );
  INV_X1 U4185 ( .A(n4483), .ZN(n4478) );
  NAND2_X1 U4186 ( .A1(n3452), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3475)
         );
  AND2_X1 U4187 ( .A1(n5388), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4308)
         );
  OR2_X1 U4188 ( .A1(n3453), .A2(n5524), .ZN(n3342) );
  NAND2_X1 U4189 ( .A1(n4435), .A2(n4385), .ZN(n4436) );
  INV_X1 U4190 ( .A(n5460), .ZN(n3904) );
  NAND2_X1 U4191 ( .A1(n4288), .A2(n4826), .ZN(n3470) );
  OR2_X1 U4192 ( .A1(n3204), .A2(n4558), .ZN(n4559) );
  NAND2_X1 U4193 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  NOR2_X1 U4194 ( .A1(n4495), .A2(n3522), .ZN(n3523) );
  OR2_X1 U4195 ( .A1(n3453), .A2(n5507), .ZN(n3380) );
  OR2_X1 U4196 ( .A1(n4237), .A2(n5867), .ZN(n4239) );
  INV_X1 U4197 ( .A(n5794), .ZN(n4025) );
  NAND2_X1 U4198 ( .A1(n3782), .A2(n3781), .ZN(n3794) );
  NAND2_X1 U4199 ( .A1(n3731), .A2(n3730), .ZN(n3739) );
  AND4_X1 U4200 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3409)
         );
  NAND2_X1 U4201 ( .A1(n3665), .A2(n3664), .ZN(n3667) );
  OR3_X1 U4202 ( .A1(n4343), .A2(n7293), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n4662) );
  NOR2_X1 U4203 ( .A1(n4731), .A2(n4298), .ZN(n4823) );
  AND2_X1 U4204 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5352), .ZN(n5692) );
  AND4_X1 U4205 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  OR2_X1 U4206 ( .A1(n4239), .A2(n4238), .ZN(n4585) );
  AND2_X1 U4207 ( .A1(n4045), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4046)
         );
  INV_X1 U4208 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3840) );
  XNOR2_X1 U4209 ( .A(n3793), .B(n3794), .ZN(n4524) );
  AND2_X1 U4210 ( .A1(n3658), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4622) );
  AND2_X1 U4211 ( .A1(n3203), .A2(n7224), .ZN(n5581) );
  INV_X1 U4212 ( .A(n4534), .ZN(n4547) );
  NOR2_X1 U4213 ( .A1(n4581), .A2(n4804), .ZN(n6831) );
  NAND2_X1 U4214 ( .A1(n3683), .A2(n3682), .ZN(n6654) );
  AND2_X1 U4215 ( .A1(n6652), .A2(n6753), .ZN(n6660) );
  INV_X1 U4216 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6838) );
  NOR2_X1 U4217 ( .A1(n4190), .A2(n5880), .ZN(n4191) );
  INV_X1 U4218 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6248) );
  OR2_X1 U4219 ( .A1(n4673), .A2(n6351), .ZN(n6277) );
  NAND2_X1 U4220 ( .A1(n4811), .A2(n4668), .ZN(n6334) );
  OR2_X1 U4221 ( .A1(n5528), .A2(n5456), .ZN(n3882) );
  INV_X1 U4222 ( .A(n4624), .ZN(n4625) );
  NOR2_X1 U4223 ( .A1(n3960), .A2(n6248), .ZN(n3980) );
  NOR2_X1 U4224 ( .A1(n6272), .A2(n3842), .ZN(n3886) );
  NAND2_X1 U4225 ( .A1(n3821), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3841)
         );
  NAND2_X1 U4226 ( .A1(n5843), .A2(n5958), .ZN(n4640) );
  NAND2_X1 U4227 ( .A1(n3203), .A2(n5638), .ZN(n5639) );
  OR2_X1 U4228 ( .A1(n3204), .A2(n7224), .ZN(n5582) );
  NOR2_X1 U4229 ( .A1(n5607), .A2(n5605), .ZN(n6518) );
  INV_X1 U4230 ( .A(n5136), .ZN(n5203) );
  AND2_X1 U4231 ( .A1(n4978), .A2(n5003), .ZN(n5135) );
  NAND2_X1 U4232 ( .A1(n6650), .A2(n5047), .ZN(n5386) );
  NAND2_X1 U4233 ( .A1(n4976), .A2(n5416), .ZN(n5519) );
  NAND2_X1 U4234 ( .A1(n4778), .A2(n4698), .ZN(n6979) );
  OR2_X1 U4235 ( .A1(n6081), .A2(n5673), .ZN(n5717) );
  NAND2_X1 U4236 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4237)
         );
  NOR4_X1 U4237 ( .A1(n6256), .A2(n6913), .A3(n5940), .A4(n6912), .ZN(n6234)
         );
  NOR2_X1 U4238 ( .A1(n5467), .A2(n6257), .ZN(n6264) );
  INV_X1 U4239 ( .A(n6312), .ZN(n6323) );
  OR2_X1 U4240 ( .A1(n6315), .A2(n5295), .ZN(n6348) );
  AND2_X1 U4241 ( .A1(n4364), .A2(n4363), .ZN(n4788) );
  AND2_X1 U4242 ( .A1(n6394), .A2(n5684), .ZN(n6384) );
  AND2_X1 U4243 ( .A1(n6394), .A2(n4801), .ZN(n6390) );
  INV_X1 U4244 ( .A(n6422), .ZN(n6415) );
  INV_X1 U4245 ( .A(n4887), .ZN(n4858) );
  INV_X1 U4246 ( .A(n4778), .ZN(n4777) );
  AND2_X1 U4247 ( .A1(n3786), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3798)
         );
  NAND2_X1 U4248 ( .A1(n3732), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3785)
         );
  INV_X1 U4249 ( .A(n6466), .ZN(n6438) );
  INV_X1 U4250 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4579) );
  OR2_X1 U4251 ( .A1(n5996), .A2(n5613), .ZN(n5971) );
  NAND2_X1 U4252 ( .A1(n5904), .A2(n5639), .ZN(n5895) );
  OR2_X1 U4253 ( .A1(n6962), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U4254 ( .A1(n4831), .A2(n4825), .ZN(n6558) );
  NOR2_X1 U4255 ( .A1(n5599), .A2(n5362), .ZN(n6550) );
  INV_X1 U4256 ( .A(n6551), .ZN(n6569) );
  NAND2_X1 U4257 ( .A1(n6861), .A2(n4897), .ZN(n5151) );
  AND2_X1 U4258 ( .A1(n5135), .A2(n4891), .ZN(n5248) );
  AND2_X1 U4259 ( .A1(n5135), .A2(n5266), .ZN(n5136) );
  INV_X1 U4260 ( .A(n6626), .ZN(n6646) );
  AND2_X1 U4261 ( .A1(n6580), .A2(n4979), .ZN(n6650) );
  AND2_X1 U4262 ( .A1(n5274), .A2(n4891), .ZN(n6735) );
  INV_X1 U4263 ( .A(n5315), .ZN(n5347) );
  OAI211_X1 U4264 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n3658), .A(n5314), .B(n5313), .ZN(n5344) );
  AND2_X1 U4265 ( .A1(n6073), .A2(n4891), .ZN(n5416) );
  INV_X1 U4266 ( .A(n7370), .ZN(n5181) );
  AND2_X1 U4267 ( .A1(n6073), .A2(n5266), .ZN(n6649) );
  INV_X1 U4268 ( .A(n6775), .ZN(n6719) );
  NOR2_X1 U4269 ( .A1(n5104), .A2(n4891), .ZN(n5521) );
  INV_X1 U4270 ( .A(n5519), .ZN(n5477) );
  AND2_X1 U4271 ( .A1(n4357), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6867) );
  INV_X1 U4272 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6213) );
  INV_X1 U4273 ( .A(n3194), .ZN(n6974) );
  INV_X1 U4274 ( .A(n6244), .ZN(n6256) );
  INV_X1 U4275 ( .A(n6315), .ZN(n6302) );
  INV_X1 U4276 ( .A(n6346), .ZN(n6331) );
  OR2_X1 U4277 ( .A1(n5530), .A2(n6168), .ZN(n6372) );
  OR2_X1 U4278 ( .A1(n4816), .A2(n4697), .ZN(n6422) );
  INV_X1 U4279 ( .A(n6429), .ZN(n4884) );
  NAND2_X1 U4280 ( .A1(n4777), .A2(n4776), .ZN(n4887) );
  NAND2_X1 U4281 ( .A1(n6474), .A2(n4633), .ZN(n6466) );
  AND2_X1 U4282 ( .A1(n5603), .A2(n5602), .ZN(n6186) );
  NAND2_X1 U4283 ( .A1(n4831), .A2(n4822), .ZN(n6478) );
  INV_X1 U4284 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6850) );
  AND2_X1 U4285 ( .A1(n5213), .A2(n5212), .ZN(n5251) );
  INV_X1 U4286 ( .A(n5009), .ZN(n5046) );
  NAND2_X1 U4287 ( .A1(n5005), .A2(n4978), .ZN(n6613) );
  NAND2_X1 U4288 ( .A1(n5049), .A2(n4978), .ZN(n6625) );
  INV_X1 U4289 ( .A(n6644), .ZN(n5415) );
  AND3_X1 U4290 ( .A1(n5422), .A2(n5421), .A3(n6850), .ZN(n6626) );
  NAND2_X1 U4291 ( .A1(n6650), .A2(n5416), .ZN(n6685) );
  NAND2_X1 U4292 ( .A1(n6650), .A2(n6649), .ZN(n6739) );
  NAND2_X1 U4293 ( .A1(n5274), .A2(n5266), .ZN(n5315) );
  NAND2_X1 U4294 ( .A1(n6745), .A2(n5416), .ZN(n7377) );
  INV_X1 U4295 ( .A(n6811), .ZN(n5184) );
  INV_X1 U4296 ( .A(n5521), .ZN(n5124) );
  INV_X1 U4297 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5515) );
  INV_X1 U4298 ( .A(n5207), .ZN(n5246) );
  AND2_X1 U4299 ( .A1(n6858), .A2(n6857), .ZN(n6874) );
  INV_X1 U4300 ( .A(n6942), .ZN(n6939) );
  INV_X1 U4301 ( .A(n6932), .ZN(n6931) );
  NAND2_X1 U4302 ( .A1(n4477), .A2(n4476), .ZN(U2830) );
  AND2_X4 U4304 ( .A1(n3319), .A2(n3320), .ZN(n4265) );
  NAND2_X1 U4305 ( .A1(n4265), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3308)
         );
  NAND2_X1 U4306 ( .A1(n3483), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3307) );
  AND2_X2 U4307 ( .A1(n3309), .A2(n4950), .ZN(n3452) );
  NAND2_X1 U4308 ( .A1(n3452), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3306)
         );
  AND2_X2 U4309 ( .A1(n3319), .A2(n4950), .ZN(n3553) );
  NAND2_X1 U4310 ( .A1(n3553), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3313)
         );
  NAND2_X1 U4311 ( .A1(n3430), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3312)
         );
  NAND2_X1 U4312 ( .A1(n3372), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4313 ( .A1(n3205), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4314 ( .A1(n4148), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4315 ( .A1(n3447), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4316 ( .A1(n3414), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4317 ( .A1(n3424), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3315) );
  AND2_X2 U4318 ( .A1(n3319), .A2(n4736), .ZN(n3429) );
  NAND2_X1 U4319 ( .A1(n3429), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4320 ( .A1(n3413), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4321 ( .A1(n3419), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3324) );
  AND2_X2 U4322 ( .A1(n3322), .A2(n4736), .ZN(n3442) );
  NAND2_X1 U4323 ( .A1(n3442), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3323) );
  INV_X1 U4324 ( .A(n3439), .ZN(n3351) );
  NAND2_X1 U4325 ( .A1(n4148), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4326 ( .A1(n3414), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4327 ( .A1(n3441), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4328 ( .A1(n3442), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3331) );
  NAND2_X1 U4329 ( .A1(n3419), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4330 ( .A1(n3429), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4331 ( .A1(n3447), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3336) );
  NAND2_X1 U4332 ( .A1(n3424), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3335) );
  INV_X1 U4333 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U4334 ( .A1(n4265), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3341)
         );
  NAND2_X1 U4335 ( .A1(n3483), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4336 ( .A1(n3452), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3339)
         );
  NAND2_X1 U4337 ( .A1(n3413), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4338 ( .A1(n3553), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3345)
         );
  NAND2_X1 U4339 ( .A1(n3430), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3344)
         );
  NAND2_X1 U4340 ( .A1(n3372), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3343)
         );
  NAND2_X1 U4341 ( .A1(n4148), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4342 ( .A1(n3414), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4343 ( .A1(n3441), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4344 ( .A1(n3442), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U4345 ( .A1(n3419), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4346 ( .A1(n3429), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4347 ( .A1(n3447), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4348 ( .A1(n3424), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3356) );
  OR2_X1 U4349 ( .A1(n3453), .A2(n5494), .ZN(n3363) );
  NAND2_X1 U4350 ( .A1(n4265), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3362)
         );
  NAND2_X1 U4351 ( .A1(n3483), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4352 ( .A1(n3452), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3360)
         );
  NAND2_X1 U4353 ( .A1(n3413), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4354 ( .A1(n3553), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3366)
         );
  NAND2_X1 U4355 ( .A1(n3430), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3365)
         );
  NAND2_X1 U4356 ( .A1(n3372), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4357 ( .A1(n3413), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4358 ( .A1(n3553), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3375)
         );
  NAND2_X1 U4359 ( .A1(n3430), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3374)
         );
  NAND2_X1 U4360 ( .A1(n3372), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3373)
         );
  INV_X1 U4361 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U4362 ( .A1(n4265), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3379)
         );
  NAND2_X1 U4363 ( .A1(n3483), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U4364 ( .A1(n3452), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3377)
         );
  NAND2_X1 U4365 ( .A1(n3414), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4366 ( .A1(n4148), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4367 ( .A1(n3441), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4368 ( .A1(n3442), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4369 ( .A1(n3419), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3388) );
  NAND2_X1 U4370 ( .A1(n3429), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4371 ( .A1(n3447), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U4372 ( .A1(n3424), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4373 ( .A1(n4148), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U4374 ( .A1(n3414), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4375 ( .A1(n3441), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4376 ( .A1(n3442), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4377 ( .A1(n3419), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3400) );
  NAND2_X1 U4378 ( .A1(n3429), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4379 ( .A1(n3447), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4380 ( .A1(n3424), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3397) );
  OR2_X1 U4381 ( .A1(n3453), .A2(n5515), .ZN(n3404) );
  NAND2_X1 U4382 ( .A1(n4265), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3403)
         );
  NAND2_X1 U4383 ( .A1(n3483), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4384 ( .A1(n3452), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3401)
         );
  NAND2_X1 U4385 ( .A1(n3413), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4386 ( .A1(n3553), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3407)
         );
  NAND2_X1 U4387 ( .A1(n3430), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3406)
         );
  NAND2_X1 U4388 ( .A1(n3372), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3405)
         );
  NAND2_X1 U4389 ( .A1(n3413), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3417) );
  NAND2_X1 U4390 ( .A1(n4265), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3416)
         );
  NAND2_X1 U4391 ( .A1(n3414), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4392 ( .A1(n3419), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4393 ( .A1(n4148), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4394 ( .A1(n3441), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3421) );
  NAND2_X1 U4395 ( .A1(n3542), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4396 ( .A1(n3553), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3428)
         );
  NAND2_X1 U4397 ( .A1(n4605), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U4398 ( .A1(n3442), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4399 ( .A1(n3424), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4400 ( .A1(n4156), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3434) );
  NAND2_X1 U4401 ( .A1(n3430), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3433)
         );
  NAND2_X1 U4402 ( .A1(n3452), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3432)
         );
  NAND2_X1 U4403 ( .A1(n3372), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3431)
         );
  NAND2_X1 U4404 ( .A1(n4287), .A2(n4774), .ZN(n3467) );
  INV_X1 U4405 ( .A(n3509), .ZN(n3466) );
  NAND2_X1 U4406 ( .A1(n4148), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3446) );
  NAND2_X1 U4407 ( .A1(n3414), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3445) );
  NAND2_X1 U4408 ( .A1(n3205), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U4409 ( .A1(n3442), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U4410 ( .A1(n3419), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3451) );
  NAND2_X1 U4411 ( .A1(n4156), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3450) );
  NAND2_X1 U4412 ( .A1(n4605), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U4413 ( .A1(n3424), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4414 ( .A1(n3483), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U4415 ( .A1(n3452), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3455)
         );
  NAND3_X1 U4416 ( .A1(n3456), .A2(n3455), .A3(n3454), .ZN(n3457) );
  NAND2_X1 U4417 ( .A1(n3430), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3460)
         );
  NAND2_X1 U4418 ( .A1(n3413), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U4419 ( .A1(n3466), .A2(n3514), .ZN(n4732) );
  XNOR2_X1 U4420 ( .A(n6877), .B(STATE_REG_2__SCAN_IN), .ZN(n4653) );
  NAND2_X2 U4421 ( .A1(n3515), .A2(n3522), .ZN(n3503) );
  AND2_X1 U4422 ( .A1(n4353), .A2(n3499), .ZN(n3469) );
  NAND2_X1 U4423 ( .A1(n3419), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U4424 ( .A1(n4156), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4425 ( .A1(n3372), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3472)
         );
  NAND2_X1 U4426 ( .A1(n3442), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3471) );
  INV_X1 U4427 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U4428 ( .A1(n4265), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3477)
         );
  NAND2_X1 U4429 ( .A1(n3414), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3476) );
  NAND2_X1 U4430 ( .A1(n3553), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3482)
         );
  NAND2_X1 U4431 ( .A1(n4605), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4432 ( .A1(n3441), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4433 ( .A1(n3430), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3479)
         );
  NAND2_X1 U4434 ( .A1(n3413), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U4435 ( .A1(n4148), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3486) );
  NAND2_X1 U4436 ( .A1(n3483), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3485) );
  NAND2_X1 U4437 ( .A1(n3424), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3484) );
  NOR2_X2 U4438 ( .A1(n3516), .A2(n4495), .ZN(n4583) );
  NAND3_X1 U4439 ( .A1(n3513), .A2(n3492), .A3(n4583), .ZN(n3493) );
  NAND2_X1 U4440 ( .A1(n3493), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U4441 ( .A1(n3498), .A2(n3515), .ZN(n3497) );
  NAND2_X1 U4442 ( .A1(n4353), .A2(n3511), .ZN(n3495) );
  NAND2_X1 U4443 ( .A1(n3495), .A2(n3494), .ZN(n3496) );
  NAND2_X1 U4444 ( .A1(n3497), .A2(n3496), .ZN(n3502) );
  NAND2_X1 U4445 ( .A1(n3498), .A2(n4804), .ZN(n3501) );
  NAND2_X1 U4446 ( .A1(n3617), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3508) );
  INV_X1 U4447 ( .A(n4357), .ZN(n3533) );
  INV_X1 U4448 ( .A(n4634), .ZN(n3532) );
  MUX2_X1 U4449 ( .A(n3533), .B(n3532), .S(n5388), .Z(n3506) );
  INV_X1 U4450 ( .A(n3506), .ZN(n3507) );
  NAND2_X1 U4451 ( .A1(n4904), .A2(n3511), .ZN(n3512) );
  NOR2_X1 U4452 ( .A1(n6962), .A2(n6861), .ZN(n6868) );
  NAND2_X1 U4453 ( .A1(n4352), .A2(n3515), .ZN(n3520) );
  NAND2_X1 U4454 ( .A1(n3503), .A2(n4929), .ZN(n3517) );
  NAND2_X1 U4455 ( .A1(n3517), .A2(n3514), .ZN(n3518) );
  OAI21_X1 U4456 ( .B1(n3516), .B2(n3518), .A(n6204), .ZN(n3519) );
  INV_X1 U4457 ( .A(n3614), .ZN(n3541) );
  NAND2_X1 U4458 ( .A1(n3524), .A2(n3523), .ZN(n4694) );
  INV_X1 U4459 ( .A(n3527), .ZN(n3528) );
  AND3_X1 U4460 ( .A1(n4826), .A2(n3525), .A3(n3522), .ZN(n4655) );
  NAND2_X1 U4461 ( .A1(n3528), .A2(n4655), .ZN(n4715) );
  INV_X1 U4462 ( .A(n4295), .ZN(n4827) );
  NAND2_X1 U4463 ( .A1(n4827), .A2(n5684), .ZN(n4819) );
  NAND2_X1 U4464 ( .A1(n3531), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3538) );
  INV_X1 U4465 ( .A(n3538), .ZN(n3536) );
  XNOR2_X1 U4466 ( .A(n5388), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5484)
         );
  NAND2_X1 U4467 ( .A1(n3532), .A2(n5484), .ZN(n3535) );
  NAND2_X1 U4468 ( .A1(n3533), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U4469 ( .A1(n3535), .A2(n3534), .ZN(n3537) );
  NAND2_X1 U4470 ( .A1(n3536), .A2(n3299), .ZN(n3540) );
  NAND2_X1 U4471 ( .A1(n3539), .A2(n3538), .ZN(n3615) );
  NAND2_X1 U4472 ( .A1(n3540), .A2(n3615), .ZN(n3613) );
  XNOR2_X1 U4473 ( .A(n3541), .B(n3613), .ZN(n4730) );
  NAND2_X1 U4474 ( .A1(n4730), .A2(n6861), .ZN(n3563) );
  INV_X1 U4475 ( .A(n3684), .ZN(n3579) );
  AOI22_X1 U4476 ( .A1(n4605), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3552) );
  INV_X1 U4477 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4478 ( .A1(n3624), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3545) );
  NAND2_X1 U4479 ( .A1(n4589), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3544) );
  OAI211_X1 U4480 ( .C1(n3546), .C2(n3768), .A(n3545), .B(n3544), .ZN(n3547)
         );
  INV_X1 U4481 ( .A(n3547), .ZN(n3551) );
  AOI22_X1 U4482 ( .A1(n3774), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3550) );
  BUF_X1 U4483 ( .A(n3453), .Z(n3629) );
  INV_X1 U4484 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3548) );
  OR2_X1 U4485 ( .A1(n3629), .A2(n3548), .ZN(n3549) );
  NAND4_X1 U4486 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3561)
         );
  INV_X2 U4487 ( .A(n3572), .ZN(n4603) );
  INV_X1 U4488 ( .A(n3419), .ZN(n4596) );
  INV_X2 U4489 ( .A(n4596), .ZN(n4196) );
  AOI22_X1 U4490 ( .A1(n4603), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4491 ( .A1(n3723), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4492 ( .A1(n4245), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3557) );
  INV_X1 U4493 ( .A(n3372), .ZN(n4597) );
  AOI22_X1 U4494 ( .A1(n4590), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4495 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3560)
         );
  NAND2_X1 U4496 ( .A1(n3579), .A2(n4494), .ZN(n3562) );
  NAND2_X1 U4497 ( .A1(n4305), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3582) );
  INV_X1 U4498 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U4499 ( .A1(n3635), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3565) );
  NAND2_X1 U4500 ( .A1(n3372), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3564)
         );
  OAI211_X1 U4501 ( .C1(n4598), .C2(n3768), .A(n3565), .B(n3564), .ZN(n3566)
         );
  INV_X1 U4502 ( .A(n3566), .ZN(n3571) );
  AOI22_X1 U4503 ( .A1(n4196), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4504 ( .A1(n3774), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3569) );
  INV_X1 U4505 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3567) );
  OR2_X1 U4506 ( .A1(n3629), .A2(n3567), .ZN(n3568) );
  NAND4_X1 U4507 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3578)
         );
  AOI22_X1 U4508 ( .A1(n4605), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4509 ( .A1(n4603), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4510 ( .A1(n4245), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3624), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4511 ( .A1(n3723), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4512 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3577)
         );
  INV_X1 U4513 ( .A(n4539), .ZN(n4550) );
  NAND2_X1 U4514 ( .A1(n3579), .A2(n4550), .ZN(n3581) );
  NAND2_X1 U4515 ( .A1(n3643), .A2(n4494), .ZN(n3580) );
  AND2_X2 U4516 ( .A1(n3587), .A2(n3614), .ZN(n6833) );
  NAND2_X1 U4517 ( .A1(n4826), .A2(n4539), .ZN(n3607) );
  NAND2_X1 U4518 ( .A1(n4550), .A2(n4826), .ZN(n3603) );
  INV_X1 U4519 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4520 ( .A1(n4603), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4521 ( .A1(n3624), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3588) );
  OAI211_X1 U4522 ( .C1(n3768), .C2(n3590), .A(n3589), .B(n3588), .ZN(n3591)
         );
  INV_X1 U4523 ( .A(n3591), .ZN(n3596) );
  AOI22_X1 U4524 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3635), .B1(n3722), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4525 ( .A1(n4196), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3594) );
  INV_X1 U4526 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3592) );
  OR2_X1 U4527 ( .A1(n3629), .A2(n3592), .ZN(n3593) );
  NAND4_X1 U4528 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3602)
         );
  AOI22_X1 U4529 ( .A1(n4605), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4530 ( .A1(n3723), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4531 ( .A1(n4245), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4532 ( .A1(n3372), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3597) );
  NAND4_X1 U4533 ( .A1(n3600), .A2(n3599), .A3(n3598), .A4(n3597), .ZN(n3601)
         );
  MUX2_X1 U4534 ( .A(n3607), .B(n3603), .S(n4493), .Z(n3604) );
  INV_X1 U4535 ( .A(n3604), .ZN(n3605) );
  NAND2_X1 U4536 ( .A1(n3605), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4537 ( .A1(n3651), .A2(n3652), .ZN(n3608) );
  INV_X1 U4538 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5234) );
  AOI21_X1 U4539 ( .B1(n3525), .B2(n4493), .A(n6861), .ZN(n3606) );
  OAI211_X1 U4540 ( .C1(n4335), .C2(n5234), .A(n3606), .B(n3607), .ZN(n3654)
         );
  NOR2_X1 U4541 ( .A1(n3607), .A2(n6861), .ZN(n4546) );
  AOI21_X1 U4542 ( .B1(n3608), .B2(n3654), .A(n4546), .ZN(n3663) );
  NAND2_X1 U4543 ( .A1(n3662), .A2(n3663), .ZN(n3666) );
  INV_X1 U4544 ( .A(n3609), .ZN(n3611) );
  NAND2_X1 U4545 ( .A1(n3198), .A2(n3614), .ZN(n3616) );
  NAND2_X1 U4546 ( .A1(n3616), .A2(n3615), .ZN(n3622) );
  NAND2_X1 U4547 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3618) );
  NAND2_X1 U4548 ( .A1(n3618), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3619) );
  NOR2_X1 U4549 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6838), .ZN(n5310)
         );
  NAND2_X1 U4550 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5310), .ZN(n6740) );
  OAI22_X1 U4551 ( .A1(n4634), .A2(n5010), .B1(n4357), .B2(n6844), .ZN(n3620)
         );
  NAND2_X1 U4552 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  AOI22_X1 U4553 ( .A1(n4590), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3634) );
  INV_X1 U4554 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3627) );
  NAND2_X1 U4555 ( .A1(n3624), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3626) );
  INV_X1 U4556 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n7263) );
  NAND2_X1 U4557 ( .A1(n4589), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3625) );
  OAI211_X1 U4558 ( .C1(n3627), .C2(n3768), .A(n3626), .B(n3625), .ZN(n3628)
         );
  INV_X1 U4559 ( .A(n3628), .ZN(n3633) );
  AOI22_X1 U4560 ( .A1(n4605), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3632) );
  INV_X1 U4561 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3630) );
  OR2_X1 U4562 ( .A1(n3629), .A2(n3630), .ZN(n3631) );
  NAND4_X1 U4563 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3641)
         );
  AOI22_X1 U4564 ( .A1(n4245), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4565 ( .A1(n4603), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4566 ( .A1(n3722), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4567 ( .A1(n3723), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3636) );
  NAND4_X1 U4568 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3640)
         );
  OAI21_X2 U4569 ( .B1(n4755), .B2(STATE2_REG_0__SCAN_IN), .A(n3642), .ZN(
        n3645) );
  AOI22_X1 U4570 ( .A1(n4305), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3643), 
        .B2(n4483), .ZN(n3644) );
  XNOR2_X2 U4571 ( .A(n3645), .B(n3644), .ZN(n3647) );
  NAND2_X2 U4572 ( .A1(n3646), .A2(n3647), .ZN(n3703) );
  INV_X1 U4573 ( .A(n3646), .ZN(n3649) );
  INV_X1 U4574 ( .A(n3647), .ZN(n3648) );
  NOR2_X2 U4575 ( .A1(n4909), .A2(n3658), .ZN(n3953) );
  NAND2_X1 U4576 ( .A1(n3651), .A2(n3654), .ZN(n3653) );
  INV_X1 U4577 ( .A(n3652), .ZN(n3655) );
  AOI21_X1 U4578 ( .B1(n4891), .B2(n3515), .A(n3658), .ZN(n4789) );
  NAND2_X1 U4579 ( .A1(n3658), .A2(n6213), .ZN(n3758) );
  NAND2_X1 U4580 ( .A1(n5684), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4581 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3660)
         );
  NAND2_X1 U4582 ( .A1(n4623), .A2(EAX_REG_0__SCAN_IN), .ZN(n3659) );
  OAI211_X1 U4583 ( .C1(n3735), .C2(n6830), .A(n3660), .B(n3659), .ZN(n3661)
         );
  AOI21_X1 U4584 ( .B1(n6833), .B2(n3953), .A(n3661), .ZN(n4790) );
  INV_X1 U4585 ( .A(n3662), .ZN(n3665) );
  INV_X1 U4586 ( .A(n3663), .ZN(n3664) );
  NAND2_X1 U4587 ( .A1(n3667), .A2(n3666), .ZN(n4890) );
  NAND2_X1 U4588 ( .A1(n4890), .A2(n3953), .ZN(n3670) );
  INV_X1 U4589 ( .A(n3735), .ZN(n3711) );
  INV_X1 U4590 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6356) );
  OAI22_X1 U4591 ( .A1(n4616), .A2(n6418), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6356), .ZN(n3668) );
  AOI21_X1 U4592 ( .B1(n4954), .B2(n3711), .A(n3668), .ZN(n3669) );
  NAND2_X1 U4593 ( .A1(n3670), .A2(n3669), .ZN(n4766) );
  OAI21_X1 U4594 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3706), .ZN(n6465) );
  AOI22_X1 U4595 ( .A1(n4621), .A2(n6465), .B1(n4622), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4596 ( .A1(n4623), .A2(EAX_REG_2__SCAN_IN), .ZN(n3671) );
  OAI211_X1 U4597 ( .C1(n3735), .C2(n3304), .A(n3672), .B(n3671), .ZN(n3674)
         );
  NAND2_X1 U4598 ( .A1(n4769), .A2(n3674), .ZN(n3673) );
  NAND2_X1 U4599 ( .A1(n4875), .A2(n3673), .ZN(n3677) );
  INV_X1 U4600 ( .A(n4769), .ZN(n3676) );
  INV_X1 U4601 ( .A(n3674), .ZN(n3675) );
  NAND2_X1 U4602 ( .A1(n3676), .A2(n3675), .ZN(n4874) );
  NAND2_X1 U4603 ( .A1(n3199), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3683) );
  NAND3_X1 U4604 ( .A1(n6850), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6661) );
  INV_X1 U4605 ( .A(n6661), .ZN(n3679) );
  NAND2_X1 U4606 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3679), .ZN(n6684) );
  NAND2_X1 U4607 ( .A1(n6850), .A2(n6684), .ZN(n3680) );
  NAND3_X1 U4608 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5476) );
  INV_X1 U4609 ( .A(n5476), .ZN(n4899) );
  NAND2_X1 U4610 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4899), .ZN(n4933) );
  NAND2_X1 U4611 ( .A1(n3680), .A2(n4933), .ZN(n5150) );
  OAI22_X1 U4612 ( .A1(n4634), .A2(n5150), .B1(n4357), .B2(n6850), .ZN(n3681)
         );
  INV_X1 U4613 ( .A(n3681), .ZN(n3682) );
  NAND2_X1 U4614 ( .A1(n4892), .A2(n6861), .ZN(n3701) );
  INV_X1 U4615 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U4616 ( .A1(n3635), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3687) );
  INV_X2 U4617 ( .A(n3543), .ZN(n4589) );
  NAND2_X1 U4618 ( .A1(n4589), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3686) );
  OAI211_X1 U4619 ( .C1(n3688), .C2(n3768), .A(n3687), .B(n3686), .ZN(n3689)
         );
  INV_X1 U4620 ( .A(n3689), .ZN(n3693) );
  AOI22_X1 U4621 ( .A1(n4605), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4622 ( .A1(n3723), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3691) );
  OR2_X1 U4623 ( .A1(n3629), .A2(n7138), .ZN(n3690) );
  NAND4_X1 U4624 ( .A1(n3693), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3699)
         );
  AOI22_X1 U4625 ( .A1(n4590), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4626 ( .A1(n3722), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4627 ( .A1(n3624), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4628 ( .A1(n4603), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3694) );
  NAND4_X1 U4629 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3698)
         );
  AOI22_X1 U4630 ( .A1(n4349), .A2(n4508), .B1(n4305), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3700) );
  INV_X1 U4631 ( .A(n4889), .ZN(n4979) );
  NAND2_X1 U4632 ( .A1(n4979), .A2(n3703), .ZN(n3704) );
  INV_X1 U4633 ( .A(n3953), .ZN(n3877) );
  INV_X1 U4634 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7183) );
  INV_X1 U4635 ( .A(n3706), .ZN(n3705) );
  INV_X1 U4636 ( .A(n3732), .ZN(n3708) );
  INV_X1 U4637 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U4638 ( .A1(n5449), .A2(n3706), .ZN(n3707) );
  NAND2_X1 U4639 ( .A1(n3708), .A2(n3707), .ZN(n5450) );
  AOI22_X1 U4640 ( .A1(n5450), .A2(n4621), .B1(n4622), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3709) );
  OAI21_X1 U4641 ( .B1(n4616), .B2(n7183), .A(n3709), .ZN(n3710) );
  AOI21_X1 U4642 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n3711), .A(n3710), 
        .ZN(n3712) );
  NAND2_X1 U4643 ( .A1(n4839), .A2(n4841), .ZN(n4840) );
  AOI22_X1 U4644 ( .A1(n4590), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3721) );
  INV_X1 U4645 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4646 ( .A1(n3624), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3714) );
  NAND2_X1 U4647 ( .A1(n4589), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3713) );
  OAI211_X1 U4648 ( .C1(n3715), .C2(n3768), .A(n3714), .B(n3713), .ZN(n3716)
         );
  INV_X1 U4649 ( .A(n3716), .ZN(n3720) );
  AOI22_X1 U4650 ( .A1(n4605), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3719) );
  INV_X1 U4651 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3717) );
  OR2_X1 U4652 ( .A1(n3629), .A2(n3717), .ZN(n3718) );
  NAND4_X1 U4653 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3729)
         );
  AOI22_X1 U4654 ( .A1(n4245), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4655 ( .A1(n4603), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4656 ( .A1(n3722), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4657 ( .A1(n3723), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3724) );
  NAND4_X1 U4658 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3728)
         );
  NAND2_X1 U4659 ( .A1(n4349), .A2(n4526), .ZN(n3731) );
  NAND2_X1 U4660 ( .A1(n4305), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3730) );
  XNOR2_X1 U4661 ( .A(n3738), .B(n3739), .ZN(n4507) );
  OAI21_X1 U4662 ( .B1(n3732), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3785), 
        .ZN(n6455) );
  INV_X1 U4663 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U4664 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3734)
         );
  NAND2_X1 U4665 ( .A1(n4623), .A2(EAX_REG_4__SCAN_IN), .ZN(n3733) );
  OAI211_X1 U4666 ( .C1(n3735), .C2(n4743), .A(n3734), .B(n3733), .ZN(n3736)
         );
  MUX2_X1 U4667 ( .A(n6455), .B(n3736), .S(n3758), .Z(n3737) );
  AOI21_X1 U4668 ( .B1(n4507), .B2(n3953), .A(n3737), .ZN(n5000) );
  NOR2_X2 U4669 ( .A1(n4840), .A2(n5000), .ZN(n4991) );
  INV_X1 U4670 ( .A(n3197), .ZN(n3740) );
  NAND2_X1 U4671 ( .A1(n3740), .A2(n3739), .ZN(n3762) );
  INV_X1 U4672 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3743) );
  NAND2_X1 U4673 ( .A1(n3722), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U4674 ( .A1(n3774), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3741) );
  OAI211_X1 U4675 ( .C1(n3572), .C2(n3743), .A(n3742), .B(n3741), .ZN(n3744)
         );
  INV_X1 U4676 ( .A(n3744), .ZN(n3749) );
  AOI22_X1 U4677 ( .A1(n3723), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4678 ( .A1(n4245), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3747) );
  INV_X1 U4679 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3745) );
  OR2_X1 U4680 ( .A1(n3629), .A2(n3745), .ZN(n3746) );
  NAND4_X1 U4681 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3755)
         );
  AOI22_X1 U4682 ( .A1(n4246), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4683 ( .A1(n4196), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4684 ( .A1(n3624), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4685 ( .A1(n4602), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4686 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3754)
         );
  NAND2_X1 U4687 ( .A1(n4349), .A2(n4525), .ZN(n3757) );
  NAND2_X1 U4688 ( .A1(n4305), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U4689 ( .A1(n3757), .A2(n3756), .ZN(n3763) );
  XNOR2_X1 U4690 ( .A(n3762), .B(n3763), .ZN(n4516) );
  NAND2_X1 U4691 ( .A1(n4516), .A2(n3953), .ZN(n3761) );
  XNOR2_X1 U4692 ( .A(n3785), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5303) );
  INV_X1 U4693 ( .A(n4622), .ZN(n4163) );
  INV_X1 U4694 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5092) );
  OAI22_X1 U4695 ( .A1(n5303), .A2(n3758), .B1(n4163), .B2(n5092), .ZN(n3759)
         );
  AOI21_X1 U4696 ( .B1(n4623), .B2(EAX_REG_5__SCAN_IN), .A(n3759), .ZN(n3760)
         );
  NAND2_X1 U4697 ( .A1(n3761), .A2(n3760), .ZN(n4990) );
  NAND2_X1 U4698 ( .A1(n4991), .A2(n4990), .ZN(n4989) );
  INV_X1 U4699 ( .A(n4989), .ZN(n3792) );
  INV_X1 U4700 ( .A(n3762), .ZN(n3764) );
  NAND2_X1 U4701 ( .A1(n3764), .A2(n3763), .ZN(n3793) );
  AOI22_X1 U4702 ( .A1(n4590), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3773) );
  INV_X1 U4703 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3767) );
  NAND2_X1 U4704 ( .A1(n3624), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4705 ( .A1(n4589), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3765) );
  OAI211_X1 U4706 ( .C1(n3768), .C2(n3767), .A(n3766), .B(n3765), .ZN(n3769)
         );
  INV_X1 U4707 ( .A(n3769), .ZN(n3772) );
  AOI22_X1 U4708 ( .A1(n4246), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3771) );
  INV_X1 U4709 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n7266) );
  OR2_X1 U4710 ( .A1(n3629), .A2(n7266), .ZN(n3770) );
  NAND4_X1 U4711 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3780)
         );
  AOI22_X1 U4712 ( .A1(n4245), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4713 ( .A1(n4603), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4714 ( .A1(n3722), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4715 ( .A1(n3723), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4716 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NAND2_X1 U4717 ( .A1(n4349), .A2(n4537), .ZN(n3782) );
  NAND2_X1 U4718 ( .A1(n4305), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3781) );
  INV_X1 U4719 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6411) );
  INV_X1 U4720 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3783) );
  OAI22_X1 U4721 ( .A1(n4616), .A2(n6411), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3783), .ZN(n3784) );
  NAND2_X1 U4722 ( .A1(n3784), .A2(n3758), .ZN(n3789) );
  NOR2_X1 U4723 ( .A1(n3786), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3787)
         );
  OR2_X1 U4724 ( .A1(n3798), .A2(n3787), .ZN(n6447) );
  NAND2_X1 U4725 ( .A1(n6447), .A2(n4621), .ZN(n3788) );
  NAND2_X1 U4726 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  INV_X1 U4727 ( .A(n5096), .ZN(n3791) );
  NAND2_X1 U4728 ( .A1(n3792), .A2(n3791), .ZN(n5126) );
  INV_X1 U4729 ( .A(n3793), .ZN(n3795) );
  NAND2_X1 U4730 ( .A1(n3795), .A2(n3794), .ZN(n4545) );
  INV_X1 U4731 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U4732 ( .A1(n4349), .A2(n4539), .ZN(n3796) );
  OAI21_X1 U4733 ( .B1(n5242), .B2(n4335), .A(n3796), .ZN(n3797) );
  INV_X1 U4734 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4871) );
  NOR2_X1 U4735 ( .A1(n3798), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3799)
         );
  OR2_X1 U4736 ( .A1(n3821), .A2(n3799), .ZN(n5439) );
  INV_X1 U4737 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n7310) );
  NOR2_X1 U4738 ( .A1(n4163), .A2(n7310), .ZN(n3800) );
  AOI21_X1 U4739 ( .B1(n5439), .B2(n4621), .A(n3800), .ZN(n3801) );
  OAI21_X1 U4740 ( .B1(n4616), .B2(n4871), .A(n3801), .ZN(n3802) );
  AOI22_X1 U4741 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4246), .B1(n3722), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4742 ( .A1(n4196), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4743 ( .A1(n3723), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4744 ( .A1(n4245), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4745 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3815)
         );
  NAND2_X1 U4746 ( .A1(n4603), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U4747 ( .A1(n4602), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3808)
         );
  NAND2_X1 U4748 ( .A1(n4590), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3807)
         );
  AND3_X1 U4749 ( .A1(n3809), .A2(n3808), .A3(n3807), .ZN(n3813) );
  AOI22_X1 U4750 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3624), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4751 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3635), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3811) );
  OR2_X1 U4752 ( .A1(n3629), .A2(n5234), .ZN(n3810) );
  NAND4_X1 U4753 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  OAI21_X1 U4754 ( .B1(n3815), .B2(n3814), .A(n3953), .ZN(n3820) );
  NAND2_X1 U4755 ( .A1(n4623), .A2(EAX_REG_8__SCAN_IN), .ZN(n3819) );
  INV_X1 U4756 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3816) );
  XNOR2_X1 U4757 ( .A(n3821), .B(n3816), .ZN(n6305) );
  OR2_X1 U4758 ( .A1(n6305), .A2(n3758), .ZN(n3818) );
  NAND2_X1 U4759 ( .A1(n4622), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3817)
         );
  NAND4_X1 U4760 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n5253)
         );
  XNOR2_X1 U4761 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3841), .ZN(n6291) );
  INV_X1 U4762 ( .A(n6291), .ZN(n3839) );
  AOI22_X1 U4763 ( .A1(n3723), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4764 ( .A1(n4603), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4765 ( .A1(n3635), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4766 ( .A1(n3554), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3822) );
  NAND4_X1 U4767 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3834)
         );
  AOI22_X1 U4768 ( .A1(n4156), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4769 ( .A1(n4602), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3828)
         );
  NAND2_X1 U4770 ( .A1(n3624), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4771 ( .A1(n4589), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3826) );
  AND3_X1 U4772 ( .A1(n3828), .A2(n3827), .A3(n3826), .ZN(n3831) );
  AOI22_X1 U4773 ( .A1(n4196), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3830) );
  INV_X1 U4774 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5219) );
  OR2_X1 U4775 ( .A1(n3629), .A2(n5219), .ZN(n3829) );
  NAND4_X1 U4776 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3833)
         );
  OAI21_X1 U4777 ( .B1(n3834), .B2(n3833), .A(n3953), .ZN(n3837) );
  NAND2_X1 U4778 ( .A1(n4623), .A2(EAX_REG_9__SCAN_IN), .ZN(n3836) );
  NAND2_X1 U4779 ( .A1(n4622), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3835)
         );
  NAND3_X1 U4780 ( .A1(n3837), .A2(n3836), .A3(n3835), .ZN(n3838) );
  AOI21_X1 U4781 ( .B1(n3839), .B2(n4621), .A(n3838), .ZN(n5372) );
  AOI21_X1 U4782 ( .B1(n6272), .B2(n3842), .A(n3886), .ZN(n6437) );
  OR2_X1 U4783 ( .A1(n6437), .A2(n3758), .ZN(n3860) );
  AOI22_X1 U4784 ( .A1(n4603), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4785 ( .A1(n3723), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4786 ( .A1(n3635), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4787 ( .A1(n4245), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4788 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3855)
         );
  AOI22_X1 U4789 ( .A1(n4590), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3853) );
  NAND2_X1 U4790 ( .A1(n4602), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3849)
         );
  NAND2_X1 U4791 ( .A1(n3624), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4792 ( .A1(n4589), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3847) );
  AND3_X1 U4793 ( .A1(n3849), .A2(n3848), .A3(n3847), .ZN(n3852) );
  AOI22_X1 U4794 ( .A1(n4246), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3851) );
  INV_X1 U4795 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5227) );
  OR2_X1 U4796 ( .A1(n3629), .A2(n5227), .ZN(n3850) );
  NAND4_X1 U4797 ( .A1(n3853), .A2(n3852), .A3(n3851), .A4(n3850), .ZN(n3854)
         );
  NOR2_X1 U4798 ( .A1(n3855), .A2(n3854), .ZN(n3856) );
  OAI22_X1 U4799 ( .A1(n3877), .A2(n3856), .B1(n4163), .B2(n6272), .ZN(n3858)
         );
  INV_X1 U4800 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5532) );
  NOR2_X1 U4801 ( .A1(n4616), .A2(n5532), .ZN(n3857) );
  NOR2_X1 U4802 ( .A1(n3858), .A2(n3857), .ZN(n3859) );
  INV_X1 U4803 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6280) );
  XNOR2_X1 U4804 ( .A(n3861), .B(n6280), .ZN(n6285) );
  OR2_X1 U4805 ( .A1(n6285), .A2(n3758), .ZN(n3881) );
  INV_X1 U4806 ( .A(EAX_REG_10__SCAN_IN), .ZN(n3862) );
  OAI22_X1 U4807 ( .A1(n4616), .A2(n3862), .B1(n4163), .B2(n6280), .ZN(n3879)
         );
  INV_X1 U4808 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4009) );
  NAND2_X1 U4809 ( .A1(n3635), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4810 ( .A1(n3722), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3863) );
  OAI211_X1 U4811 ( .C1(n3543), .C2(n4009), .A(n3864), .B(n3863), .ZN(n3865)
         );
  INV_X1 U4812 ( .A(n3865), .ZN(n3869) );
  AOI22_X1 U4813 ( .A1(n4590), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4814 ( .A1(n4196), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3867) );
  OR2_X1 U4815 ( .A1(n3629), .A2(n7263), .ZN(n3866) );
  NAND4_X1 U4816 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3875)
         );
  AOI22_X1 U4817 ( .A1(n3723), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4818 ( .A1(n4602), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4819 ( .A1(n4603), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3624), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4820 ( .A1(n4604), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4821 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3874)
         );
  NOR2_X1 U4822 ( .A1(n3875), .A2(n3874), .ZN(n3876) );
  NOR2_X1 U4823 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  NOR2_X1 U4824 ( .A1(n3879), .A2(n3878), .ZN(n3880) );
  NAND2_X1 U4825 ( .A1(n3881), .A2(n3880), .ZN(n5457) );
  INV_X1 U4826 ( .A(n5457), .ZN(n5456) );
  INV_X1 U4827 ( .A(EAX_REG_13__SCAN_IN), .ZN(n3885) );
  OAI21_X1 U4828 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3883), .A(n3941), 
        .ZN(n6267) );
  AOI22_X1 U4829 ( .A1(n4621), .A2(n6267), .B1(n4622), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3884) );
  OAI21_X1 U4830 ( .B1(n4616), .B2(n3885), .A(n3884), .ZN(n6170) );
  XNOR2_X1 U4831 ( .A(n3886), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5546)
         );
  INV_X1 U4832 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5464) );
  AOI21_X1 U4833 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5464), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3888) );
  INV_X1 U4834 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5526) );
  NOR2_X1 U4835 ( .A1(n4616), .A2(n5526), .ZN(n3887) );
  OAI22_X1 U4836 ( .A1(n5546), .A2(n3758), .B1(n3888), .B2(n3887), .ZN(n3903)
         );
  AOI22_X1 U4837 ( .A1(n4196), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4838 ( .A1(n4246), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4839 ( .A1(n4245), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4840 ( .A1(n4603), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4841 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3901)
         );
  NAND2_X1 U4842 ( .A1(n4602), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3895)
         );
  NAND2_X1 U4843 ( .A1(n3723), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3894)
         );
  NAND2_X1 U4844 ( .A1(n3624), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3893) );
  AND3_X1 U4845 ( .A1(n3895), .A2(n3894), .A3(n3893), .ZN(n3899) );
  AOI22_X1 U4846 ( .A1(n4604), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4847 ( .A1(n3554), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3897) );
  INV_X1 U4848 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5223) );
  OR2_X1 U4849 ( .A1(n3629), .A2(n5223), .ZN(n3896) );
  NAND4_X1 U4850 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3900)
         );
  OAI21_X1 U4851 ( .B1(n3901), .B2(n3900), .A(n3953), .ZN(n3902) );
  NAND2_X1 U4852 ( .A1(n3903), .A2(n3902), .ZN(n5460) );
  NOR2_X1 U4853 ( .A1(n3922), .A2(n3904), .ZN(n6169) );
  NAND2_X1 U4854 ( .A1(n4603), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3907) );
  NAND2_X1 U4855 ( .A1(n4602), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3906)
         );
  NAND2_X1 U4856 ( .A1(n4590), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3905)
         );
  AND3_X1 U4857 ( .A1(n3907), .A2(n3906), .A3(n3905), .ZN(n3911) );
  AOI22_X1 U4858 ( .A1(n4245), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4859 ( .A1(n3722), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3909) );
  INV_X1 U4860 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5250) );
  OR2_X1 U4861 ( .A1(n3629), .A2(n5250), .ZN(n3908) );
  NAND4_X1 U4862 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3917)
         );
  AOI22_X1 U4863 ( .A1(n3635), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4864 ( .A1(n3723), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4865 ( .A1(n4196), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3624), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4866 ( .A1(n4273), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4867 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3916)
         );
  OR2_X1 U4868 ( .A1(n3917), .A2(n3916), .ZN(n3918) );
  NAND2_X1 U4869 ( .A1(n3953), .A2(n3918), .ZN(n6174) );
  INV_X1 U4870 ( .A(n6174), .ZN(n3919) );
  AND2_X1 U4871 ( .A1(n6169), .A2(n3919), .ZN(n3921) );
  AND2_X1 U4872 ( .A1(n3919), .A2(n6170), .ZN(n3920) );
  AOI21_X1 U4873 ( .B1(n6168), .B2(n3921), .A(n3920), .ZN(n6177) );
  NAND2_X1 U4874 ( .A1(n6177), .A2(n6171), .ZN(n5566) );
  INV_X1 U4875 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5579) );
  OAI21_X1 U4876 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6213), .A(n3658), 
        .ZN(n3923) );
  OAI21_X1 U4877 ( .B1(n4616), .B2(n5579), .A(n3923), .ZN(n3925) );
  XNOR2_X1 U4878 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3941), .ZN(n5574)
         );
  INV_X1 U4879 ( .A(n5574), .ZN(n5953) );
  OR2_X1 U4880 ( .A1(n3758), .A2(n5953), .ZN(n3924) );
  NAND2_X1 U4881 ( .A1(n3925), .A2(n3924), .ZN(n3940) );
  AOI22_X1 U4882 ( .A1(n4603), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4883 ( .A1(n4602), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3723), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4884 ( .A1(n4196), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4885 ( .A1(n4246), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4886 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3938)
         );
  AOI22_X1 U4887 ( .A1(n4156), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3936) );
  NAND2_X1 U4888 ( .A1(n3624), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U4889 ( .A1(n4273), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3931)
         );
  NAND2_X1 U4890 ( .A1(n4589), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3930) );
  AND3_X1 U4891 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3935) );
  AOI22_X1 U4892 ( .A1(n4245), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3934) );
  INV_X1 U4893 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5238) );
  OR2_X1 U4894 ( .A1(n3629), .A2(n5238), .ZN(n3933) );
  NAND4_X1 U4895 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3937)
         );
  OAI21_X1 U4896 ( .B1(n3938), .B2(n3937), .A(n3953), .ZN(n3939) );
  NAND2_X1 U4897 ( .A1(n3940), .A2(n3939), .ZN(n5565) );
  NAND2_X1 U4898 ( .A1(n5566), .A2(n5565), .ZN(n5564) );
  XNOR2_X1 U4899 ( .A(n3960), .B(n6248), .ZN(n6252) );
  AOI22_X1 U4900 ( .A1(n4196), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4901 ( .A1(n4603), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4902 ( .A1(n3723), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4903 ( .A1(n4246), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4904 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3955)
         );
  INV_X1 U4905 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4128) );
  NAND2_X1 U4906 ( .A1(n4590), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3947)
         );
  NAND2_X1 U4907 ( .A1(n4265), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3946)
         );
  OAI211_X1 U4908 ( .C1(n3543), .C2(n4128), .A(n3947), .B(n3946), .ZN(n3948)
         );
  INV_X1 U4909 ( .A(n3948), .ZN(n3952) );
  AOI22_X1 U4910 ( .A1(n3624), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4911 ( .A1(n4245), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3950) );
  OR2_X1 U4912 ( .A1(n3629), .A2(n5242), .ZN(n3949) );
  NAND4_X1 U4913 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3954)
         );
  OAI21_X1 U4914 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n3958) );
  NAND2_X1 U4915 ( .A1(n4623), .A2(EAX_REG_15__SCAN_IN), .ZN(n3957) );
  NAND2_X1 U4916 ( .A1(n4622), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3956)
         );
  NAND3_X1 U4917 ( .A1(n3958), .A2(n3957), .A3(n3956), .ZN(n3959) );
  AOI21_X1 U4918 ( .B1(n6252), .B2(n4621), .A(n3959), .ZN(n5840) );
  NOR2_X2 U4919 ( .A1(n5564), .A2(n5840), .ZN(n5805) );
  XOR2_X1 U4920 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3980), .Z(n6239) );
  NAND2_X1 U4921 ( .A1(n4929), .A2(n3499), .ZN(n3961) );
  INV_X1 U4922 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U4923 ( .A1(n4196), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3963) );
  NAND2_X1 U4924 ( .A1(n4602), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3962)
         );
  OAI211_X1 U4925 ( .C1(n3543), .C2(n5035), .A(n3963), .B(n3962), .ZN(n3964)
         );
  INV_X1 U4926 ( .A(n3964), .ZN(n3969) );
  AOI22_X1 U4927 ( .A1(n4246), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4928 ( .A1(n3722), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3967) );
  INV_X1 U4929 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3965) );
  OR2_X1 U4930 ( .A1(n3629), .A2(n3965), .ZN(n3966) );
  NAND4_X1 U4931 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3975)
         );
  AOI22_X1 U4932 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4590), .B1(n3635), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4933 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4603), .B1(n3554), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4934 ( .A1(n3723), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4935 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3542), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4936 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3974)
         );
  OR2_X1 U4937 ( .A1(n3975), .A2(n3974), .ZN(n3978) );
  INV_X1 U4938 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3976) );
  INV_X1 U4939 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5941) );
  OAI22_X1 U4940 ( .A1(n4616), .A2(n3976), .B1(n4163), .B2(n5941), .ZN(n3977)
         );
  AOI21_X1 U4941 ( .B1(n4618), .B2(n3978), .A(n3977), .ZN(n3979) );
  OAI21_X1 U4942 ( .B1(n6239), .B2(n3758), .A(n3979), .ZN(n5804) );
  NAND2_X1 U4943 ( .A1(n5805), .A2(n5804), .ZN(n5733) );
  XNOR2_X1 U4944 ( .A(n4002), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5738)
         );
  NAND2_X1 U4945 ( .A1(n5738), .A2(n4621), .ZN(n4001) );
  NAND2_X1 U4946 ( .A1(n4603), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U4947 ( .A1(n4590), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3982)
         );
  NAND2_X1 U4948 ( .A1(n3554), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3981) );
  AND3_X1 U4949 ( .A1(n3983), .A2(n3982), .A3(n3981), .ZN(n3988) );
  AOI22_X1 U4950 ( .A1(n3723), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4951 ( .A1(n3635), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3624), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3986) );
  INV_X1 U4952 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3984) );
  OR2_X1 U4953 ( .A1(n3629), .A2(n3984), .ZN(n3985) );
  NAND4_X1 U4954 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3994)
         );
  AOI22_X1 U4955 ( .A1(n4245), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4956 ( .A1(n4602), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4957 ( .A1(n4604), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4958 ( .A1(n4196), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U4959 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3993)
         );
  NOR2_X1 U4960 ( .A1(n3994), .A2(n3993), .ZN(n3999) );
  INV_X1 U4961 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3996) );
  NAND2_X1 U4962 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3995)
         );
  OAI211_X1 U4963 ( .C1(n4616), .C2(n3996), .A(n3758), .B(n3995), .ZN(n3997)
         );
  INV_X1 U4964 ( .A(n3997), .ZN(n3998) );
  OAI21_X1 U4965 ( .B1(n4282), .B2(n3999), .A(n3998), .ZN(n4000) );
  NAND2_X1 U4966 ( .A1(n4001), .A2(n4000), .ZN(n5736) );
  INV_X1 U4967 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5740) );
  INV_X1 U4968 ( .A(n4045), .ZN(n4005) );
  OR2_X1 U4969 ( .A1(n4003), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4004)
         );
  NAND2_X1 U4970 ( .A1(n4005), .A2(n4004), .ZN(n6232) );
  NAND2_X1 U4971 ( .A1(n4603), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U4972 ( .A1(n4602), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4007)
         );
  NAND2_X1 U4973 ( .A1(n4590), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4006)
         );
  AND3_X1 U4974 ( .A1(n4008), .A2(n4007), .A3(n4006), .ZN(n4013) );
  AOI22_X1 U4975 ( .A1(n3723), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4976 ( .A1(n4245), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4011) );
  OR2_X1 U4977 ( .A1(n3629), .A2(n4009), .ZN(n4010) );
  NAND4_X1 U4978 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U4979 ( .A1(n3722), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4980 ( .A1(n4196), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4981 ( .A1(n3635), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4982 ( .A1(n3554), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4983 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  NOR2_X1 U4984 ( .A1(n4019), .A2(n4018), .ZN(n4020) );
  NOR2_X1 U4985 ( .A1(n4282), .A2(n4020), .ZN(n4024) );
  INV_X1 U4986 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4022) );
  NAND2_X1 U4987 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4021)
         );
  OAI211_X1 U4988 ( .C1(n4616), .C2(n4022), .A(n3758), .B(n4021), .ZN(n4023)
         );
  OAI22_X1 U4989 ( .A1(n6232), .A2(n3758), .B1(n4024), .B2(n4023), .ZN(n5794)
         );
  INV_X1 U4990 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U4991 ( .A(n4045), .B(n6141), .ZN(n6139) );
  NAND2_X1 U4992 ( .A1(n6139), .A2(n4621), .ZN(n4044) );
  INV_X1 U4993 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U4994 ( .A1(n4246), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4027)
         );
  NAND2_X1 U4995 ( .A1(n4602), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4026)
         );
  OAI211_X1 U4996 ( .C1(n3543), .C2(n5045), .A(n4027), .B(n4026), .ZN(n4028)
         );
  INV_X1 U4997 ( .A(n4028), .ZN(n4033) );
  AOI22_X1 U4998 ( .A1(n3723), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4999 ( .A1(n4590), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4031) );
  INV_X1 U5000 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4029) );
  OR2_X1 U5001 ( .A1(n3629), .A2(n4029), .ZN(n4030) );
  NAND4_X1 U5002 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4039)
         );
  AOI22_X1 U5003 ( .A1(n4245), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5004 ( .A1(n4603), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5005 ( .A1(n4196), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5006 ( .A1(n3624), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U5007 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  NOR2_X1 U5008 ( .A1(n4039), .A2(n4038), .ZN(n4042) );
  OAI21_X1 U5009 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6141), .A(n3758), .ZN(
        n4040) );
  AOI21_X1 U5010 ( .B1(n4623), .B2(EAX_REG_19__SCAN_IN), .A(n4040), .ZN(n4041)
         );
  OAI21_X1 U5011 ( .B1(n4282), .B2(n4042), .A(n4041), .ZN(n4043) );
  NAND2_X1 U5012 ( .A1(n4044), .A2(n4043), .ZN(n5785) );
  OAI21_X1 U5013 ( .B1(n4046), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4089), 
        .ZN(n6131) );
  OR2_X1 U5014 ( .A1(n6131), .A2(n3758), .ZN(n4067) );
  NAND2_X1 U5015 ( .A1(n4602), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4049)
         );
  NAND2_X1 U5016 ( .A1(n4590), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U5017 ( .A1(n3722), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4047) );
  AND3_X1 U5018 ( .A1(n4049), .A2(n4048), .A3(n4047), .ZN(n4054) );
  AOI22_X1 U5019 ( .A1(n3635), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5020 ( .A1(n4246), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4052) );
  INV_X1 U5021 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4050) );
  OR2_X1 U5022 ( .A1(n3629), .A2(n4050), .ZN(n4051) );
  NAND4_X1 U5023 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4060)
         );
  AOI22_X1 U5024 ( .A1(n4603), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5025 ( .A1(n4245), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5026 ( .A1(n3723), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5027 ( .A1(n4273), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U5028 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4059)
         );
  NOR2_X1 U5029 ( .A1(n4060), .A2(n4059), .ZN(n4065) );
  INV_X1 U5030 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5031 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4061)
         );
  OAI211_X1 U5032 ( .C1(n4616), .C2(n4062), .A(n3758), .B(n4061), .ZN(n4063)
         );
  INV_X1 U5033 ( .A(n4063), .ZN(n4064) );
  OAI21_X1 U5034 ( .B1(n4282), .B2(n4065), .A(n4064), .ZN(n4066) );
  XNOR2_X1 U5035 ( .A(n4089), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6121)
         );
  AOI22_X1 U5036 ( .A1(n4590), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4074) );
  NAND2_X1 U5037 ( .A1(n4265), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4070)
         );
  NAND2_X1 U5038 ( .A1(n3542), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4069) );
  NAND2_X1 U5039 ( .A1(n4589), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4068) );
  AND3_X1 U5040 ( .A1(n4070), .A2(n4069), .A3(n4068), .ZN(n4073) );
  AOI22_X1 U5041 ( .A1(n4246), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4072) );
  INV_X1 U5042 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4241) );
  OR2_X1 U5043 ( .A1(n3629), .A2(n4241), .ZN(n4071) );
  NAND4_X1 U5044 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4080)
         );
  AOI22_X1 U5045 ( .A1(n4245), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5046 ( .A1(n4603), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5047 ( .A1(n3722), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5048 ( .A1(n3723), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5049 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  OR2_X1 U5050 ( .A1(n4080), .A2(n4079), .ZN(n4084) );
  INV_X1 U5051 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4082) );
  OAI21_X1 U5052 ( .B1(n6213), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3658), 
        .ZN(n4081) );
  OAI21_X1 U5053 ( .B1(n4616), .B2(n4082), .A(n4081), .ZN(n4083) );
  AOI21_X1 U5054 ( .B1(n4618), .B2(n4084), .A(n4083), .ZN(n4085) );
  AOI21_X1 U5055 ( .B1(n6121), .B2(n4621), .A(n4085), .ZN(n5903) );
  INV_X1 U5056 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6123) );
  INV_X1 U5057 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4086) );
  OAI21_X1 U5058 ( .B1(n4089), .B2(n6123), .A(n4086), .ZN(n4087) );
  INV_X1 U5059 ( .A(n4087), .ZN(n4090) );
  NAND2_X1 U5060 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4088) );
  OR2_X1 U5061 ( .A1(n4090), .A2(n4110), .ZN(n5899) );
  NAND2_X1 U5062 ( .A1(n4265), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4093)
         );
  NAND2_X1 U5063 ( .A1(n3542), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4092) );
  NAND2_X1 U5064 ( .A1(n3554), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4091) );
  AND3_X1 U5065 ( .A1(n4093), .A2(n4092), .A3(n4091), .ZN(n4098) );
  AOI22_X1 U5066 ( .A1(n3635), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5067 ( .A1(n4590), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4096) );
  INV_X1 U5068 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4094) );
  OR2_X1 U5069 ( .A1(n3629), .A2(n4094), .ZN(n4095) );
  NAND4_X1 U5070 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4104)
         );
  AOI22_X1 U5071 ( .A1(n4246), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5072 ( .A1(n3723), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5073 ( .A1(n4245), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5074 ( .A1(n4603), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5075 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4103)
         );
  OR2_X1 U5076 ( .A1(n4104), .A2(n4103), .ZN(n4108) );
  INV_X1 U5077 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4106) );
  NAND2_X1 U5078 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4105)
         );
  OAI211_X1 U5079 ( .C1(n4616), .C2(n4106), .A(n3758), .B(n4105), .ZN(n4107)
         );
  AOI21_X1 U5080 ( .B1(n4618), .B2(n4108), .A(n4107), .ZN(n4109) );
  AOI21_X1 U5081 ( .B1(n6112), .B2(n4621), .A(n4109), .ZN(n5778) );
  NAND2_X1 U5082 ( .A1(n4110), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4144)
         );
  OR2_X1 U5083 ( .A1(n4110), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4111)
         );
  AND2_X1 U5084 ( .A1(n4144), .A2(n4111), .ZN(n6101) );
  NAND2_X1 U5085 ( .A1(n6101), .A2(n4621), .ZN(n4143) );
  AOI22_X1 U5086 ( .A1(n4590), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U5087 ( .A1(n4602), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4114)
         );
  NAND2_X1 U5088 ( .A1(n3542), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4113) );
  NAND2_X1 U5089 ( .A1(n4589), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4112) );
  AND3_X1 U5090 ( .A1(n4114), .A2(n4113), .A3(n4112), .ZN(n4117) );
  AOI22_X1 U5091 ( .A1(n4246), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4116) );
  OR2_X1 U5092 ( .A1(n3629), .A2(n5035), .ZN(n4115) );
  NAND4_X1 U5093 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4124)
         );
  AOI22_X1 U5094 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3635), .B1(n4245), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5095 ( .A1(n4603), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5096 ( .A1(n3722), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5097 ( .A1(n3723), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U5098 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4123)
         );
  OR2_X1 U5099 ( .A1(n4124), .A2(n4123), .ZN(n4147) );
  AOI22_X1 U5100 ( .A1(n4590), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4132) );
  NAND2_X1 U5101 ( .A1(n4602), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4127)
         );
  NAND2_X1 U5102 ( .A1(n3624), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U5103 ( .A1(n4589), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4125) );
  AND3_X1 U5104 ( .A1(n4127), .A2(n4126), .A3(n4125), .ZN(n4131) );
  AOI22_X1 U5105 ( .A1(n4246), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4130) );
  OR2_X1 U5106 ( .A1(n3629), .A2(n4128), .ZN(n4129) );
  NAND4_X1 U5107 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4138)
         );
  AOI22_X1 U5108 ( .A1(n4245), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5109 ( .A1(n4603), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5110 ( .A1(n3722), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5111 ( .A1(n3723), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U5112 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4137)
         );
  OR2_X1 U5113 ( .A1(n4138), .A2(n4137), .ZN(n4146) );
  XNOR2_X1 U5114 ( .A(n4147), .B(n4146), .ZN(n4141) );
  INV_X1 U5115 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n7299) );
  OAI21_X1 U5116 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7299), .A(n3758), .ZN(
        n4139) );
  AOI21_X1 U5117 ( .B1(n4623), .B2(EAX_REG_23__SCAN_IN), .A(n4139), .ZN(n4140)
         );
  OAI21_X1 U5118 ( .B1(n4282), .B2(n4141), .A(n4140), .ZN(n4142) );
  NAND2_X1 U5119 ( .A1(n4143), .A2(n4142), .ZN(n5771) );
  INV_X1 U5120 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n7223) );
  NAND2_X1 U5121 ( .A1(n4144), .A2(n7223), .ZN(n4145) );
  NAND2_X1 U5122 ( .A1(n4190), .A2(n4145), .ZN(n5648) );
  NAND2_X1 U5123 ( .A1(n4147), .A2(n4146), .ZN(n4182) );
  NAND2_X1 U5124 ( .A1(n4148), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4151) );
  NAND2_X1 U5125 ( .A1(n3722), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4150) );
  NAND2_X1 U5126 ( .A1(n3774), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4149) );
  AND3_X1 U5127 ( .A1(n4151), .A2(n4150), .A3(n4149), .ZN(n4155) );
  AOI22_X1 U5128 ( .A1(n4603), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5129 ( .A1(n3723), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4153) );
  INV_X1 U5130 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5023) );
  OR2_X1 U5131 ( .A1(n3629), .A2(n5023), .ZN(n4152) );
  NAND4_X1 U5132 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4162)
         );
  AOI22_X1 U5133 ( .A1(n4196), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5134 ( .A1(n4246), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4156), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5135 ( .A1(n3624), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5136 ( .A1(n4602), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U5137 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4161)
         );
  NOR2_X1 U5138 ( .A1(n4162), .A2(n4161), .ZN(n4183) );
  XNOR2_X1 U5139 ( .A(n4182), .B(n4183), .ZN(n4167) );
  INV_X1 U5140 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4164) );
  OAI22_X1 U5141 ( .A1(n4616), .A2(n4164), .B1(n7223), .B2(n4163), .ZN(n4165)
         );
  INV_X1 U5142 ( .A(n4165), .ZN(n4166) );
  OAI21_X1 U5143 ( .B1(n4282), .B2(n4167), .A(n4166), .ZN(n4168) );
  AOI21_X1 U5144 ( .B1(n5648), .B2(n4621), .A(n4168), .ZN(n4683) );
  XNOR2_X1 U5145 ( .A(n4190), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6091)
         );
  AOI22_X1 U5146 ( .A1(n4590), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4175) );
  NAND2_X1 U5147 ( .A1(n4602), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4171)
         );
  NAND2_X1 U5148 ( .A1(n3624), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U5149 ( .A1(n4589), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4169) );
  AND3_X1 U5150 ( .A1(n4171), .A2(n4170), .A3(n4169), .ZN(n4174) );
  AOI22_X1 U5151 ( .A1(n4246), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4173) );
  INV_X1 U5152 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5019) );
  OR2_X1 U5153 ( .A1(n3629), .A2(n5019), .ZN(n4172) );
  NAND4_X1 U5154 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4181)
         );
  AOI22_X1 U5155 ( .A1(n4245), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5156 ( .A1(n4603), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5157 ( .A1(n3722), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5158 ( .A1(n3723), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4176) );
  NAND4_X1 U5159 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4180)
         );
  OR2_X1 U5160 ( .A1(n4181), .A2(n4180), .ZN(n4206) );
  NOR2_X1 U5161 ( .A1(n4183), .A2(n4182), .ZN(n4207) );
  INV_X1 U5162 ( .A(n4207), .ZN(n4184) );
  XNOR2_X1 U5163 ( .A(n4206), .B(n4184), .ZN(n4188) );
  INV_X1 U5164 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4186) );
  OAI21_X1 U5165 ( .B1(n6213), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n3658), 
        .ZN(n4185) );
  OAI21_X1 U5166 ( .B1(n4616), .B2(n4186), .A(n4185), .ZN(n4187) );
  AOI21_X1 U5167 ( .B1(n4618), .B2(n4188), .A(n4187), .ZN(n4189) );
  AOI21_X1 U5168 ( .B1(n6091), .B2(n4621), .A(n4189), .ZN(n5760) );
  INV_X1 U5169 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5880) );
  OR2_X1 U5170 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4192)
         );
  NAND2_X1 U5171 ( .A1(n4237), .A2(n4192), .ZN(n6089) );
  AOI22_X1 U5172 ( .A1(n4603), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U5173 ( .A1(n3624), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4193) );
  OAI211_X1 U5174 ( .C1(n5045), .C2(n3629), .A(n4194), .B(n4193), .ZN(n4195)
         );
  INV_X1 U5175 ( .A(n4195), .ZN(n4199) );
  AOI22_X1 U5176 ( .A1(n4590), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5177 ( .A1(n4196), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4197) );
  NAND3_X1 U5178 ( .A1(n4199), .A2(n4198), .A3(n4197), .ZN(n4205) );
  AOI22_X1 U5179 ( .A1(n4246), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5180 ( .A1(n3723), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5181 ( .A1(n4602), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5182 ( .A1(n4245), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4200) );
  NAND4_X1 U5183 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4204)
         );
  NOR2_X1 U5184 ( .A1(n4205), .A2(n4204), .ZN(n4216) );
  NAND2_X1 U5185 ( .A1(n4207), .A2(n4206), .ZN(n4215) );
  XNOR2_X1 U5186 ( .A(n4216), .B(n4215), .ZN(n4212) );
  INV_X1 U5187 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4209) );
  NAND2_X1 U5188 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4208)
         );
  OAI211_X1 U5189 ( .C1(n4616), .C2(n4209), .A(n3758), .B(n4208), .ZN(n4210)
         );
  INV_X1 U5190 ( .A(n4210), .ZN(n4211) );
  OAI21_X1 U5191 ( .B1(n4212), .B2(n4282), .A(n4211), .ZN(n4213) );
  NAND2_X1 U5192 ( .A1(n5752), .A2(n5753), .ZN(n5721) );
  INV_X1 U5193 ( .A(n5721), .ZN(n4236) );
  XNOR2_X1 U5194 ( .A(n4237), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5869)
         );
  NAND2_X1 U5195 ( .A1(n5869), .A2(n4621), .ZN(n4234) );
  NOR2_X1 U5196 ( .A1(n4216), .A2(n4215), .ZN(n4257) );
  AOI22_X1 U5197 ( .A1(n4590), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4223) );
  NAND2_X1 U5198 ( .A1(n4602), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4219)
         );
  NAND2_X1 U5199 ( .A1(n3624), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U5200 ( .A1(n4589), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4217) );
  AND3_X1 U5201 ( .A1(n4219), .A2(n4218), .A3(n4217), .ZN(n4222) );
  AOI22_X1 U5202 ( .A1(n4246), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4221) );
  INV_X1 U5203 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5015) );
  OR2_X1 U5204 ( .A1(n3629), .A2(n5015), .ZN(n4220) );
  NAND4_X1 U5205 ( .A1(n4223), .A2(n4222), .A3(n4221), .A4(n4220), .ZN(n4229)
         );
  AOI22_X1 U5206 ( .A1(n4245), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U5207 ( .A1(n4603), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U5208 ( .A1(n3722), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U5209 ( .A1(n3723), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4224) );
  NAND4_X1 U5210 ( .A1(n4227), .A2(n4226), .A3(n4225), .A4(n4224), .ZN(n4228)
         );
  OR2_X1 U5211 ( .A1(n4229), .A2(n4228), .ZN(n4256) );
  XNOR2_X1 U5212 ( .A(n4257), .B(n4256), .ZN(n4232) );
  INV_X1 U5213 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5867) );
  AOI21_X1 U5214 ( .B1(n5867), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4230) );
  AOI21_X1 U5215 ( .B1(n4623), .B2(EAX_REG_27__SCAN_IN), .A(n4230), .ZN(n4231)
         );
  OAI21_X1 U5216 ( .B1(n4232), .B2(n4282), .A(n4231), .ZN(n4233) );
  NAND2_X1 U5217 ( .A1(n4234), .A2(n4233), .ZN(n5723) );
  INV_X1 U5218 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U5219 ( .A1(n4239), .A2(n4238), .ZN(n4240) );
  NAND2_X1 U5220 ( .A1(n4585), .A2(n4240), .ZN(n5860) );
  INV_X1 U5221 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U5222 ( .A1(n3629), .A2(n5031), .ZN(n4244) );
  OAI22_X1 U5223 ( .A1(n3572), .A2(n4242), .B1(n3202), .B2(n4241), .ZN(n4243)
         );
  AOI211_X1 U5224 ( .C1(INSTQUEUE_REG_11__5__SCAN_IN), .C2(n3635), .A(n4244), 
        .B(n4243), .ZN(n4249) );
  AOI22_X1 U5225 ( .A1(n3723), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4248) );
  AOI22_X1 U5226 ( .A1(n4246), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4247) );
  NAND3_X1 U5227 ( .A1(n4249), .A2(n4248), .A3(n4247), .ZN(n4255) );
  AOI22_X1 U5228 ( .A1(n4590), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5229 ( .A1(n3774), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U5230 ( .A1(n3542), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U5231 ( .A1(n4602), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4250) );
  NAND4_X1 U5232 ( .A1(n4253), .A2(n4252), .A3(n4251), .A4(n4250), .ZN(n4254)
         );
  NOR2_X1 U5233 ( .A1(n4255), .A2(n4254), .ZN(n4264) );
  NAND2_X1 U5234 ( .A1(n4257), .A2(n4256), .ZN(n4263) );
  XNOR2_X1 U5235 ( .A(n4264), .B(n4263), .ZN(n4258) );
  NOR2_X1 U5236 ( .A1(n4258), .A2(n4282), .ZN(n4262) );
  INV_X1 U5237 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U5238 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4259)
         );
  OAI211_X1 U5239 ( .C1(n4616), .C2(n4260), .A(n3758), .B(n4259), .ZN(n4261)
         );
  OAI22_X1 U5240 ( .A1(n5860), .A2(n3758), .B1(n4262), .B2(n4261), .ZN(n5710)
         );
  INV_X1 U5241 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5702) );
  XNOR2_X1 U5242 ( .A(n4585), .B(n5702), .ZN(n5847) );
  NOR2_X1 U5243 ( .A1(n4264), .A2(n4263), .ZN(n4588) );
  AOI22_X1 U5244 ( .A1(n4156), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4272) );
  NAND2_X1 U5245 ( .A1(n4265), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4268)
         );
  NAND2_X1 U5246 ( .A1(n3624), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5247 ( .A1(n4589), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4266) );
  AND3_X1 U5248 ( .A1(n4268), .A2(n4267), .A3(n4266), .ZN(n4271) );
  AOI22_X1 U5249 ( .A1(n4246), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4270) );
  INV_X1 U5250 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5027) );
  OR2_X1 U5251 ( .A1(n3629), .A2(n5027), .ZN(n4269) );
  NAND4_X1 U5252 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), .ZN(n4279)
         );
  AOI22_X1 U5253 ( .A1(n4245), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3635), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5254 ( .A1(n4603), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5255 ( .A1(n3722), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5256 ( .A1(n3723), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5257 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4278)
         );
  OR2_X1 U5258 ( .A1(n4279), .A2(n4278), .ZN(n4587) );
  XNOR2_X1 U5259 ( .A(n4588), .B(n4587), .ZN(n4283) );
  AOI21_X1 U5260 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n3658), .A(n4621), 
        .ZN(n4281) );
  NAND2_X1 U5261 ( .A1(n4623), .A2(EAX_REG_29__SCAN_IN), .ZN(n4280) );
  OAI211_X1 U5262 ( .C1(n4283), .C2(n4282), .A(n4281), .B(n4280), .ZN(n4284)
         );
  OAI21_X1 U5263 ( .B1(n5847), .B2(n3758), .A(n4284), .ZN(n4285) );
  AND2_X1 U5264 ( .A1(n3213), .A2(n4285), .ZN(n4286) );
  NAND2_X1 U5265 ( .A1(n4287), .A2(n4904), .ZN(n4289) );
  MUX2_X1 U5266 ( .A(n4289), .B(n6984), .S(n4288), .Z(n4722) );
  NAND2_X2 U5267 ( .A1(n3201), .A2(n3514), .ZN(n4385) );
  NOR2_X1 U5268 ( .A1(n5684), .A2(n3511), .ZN(n4290) );
  AOI21_X1 U5269 ( .B1(n3516), .B2(n4470), .A(n4290), .ZN(n4292) );
  AND2_X1 U5270 ( .A1(n3525), .A2(n3201), .ZN(n5353) );
  AND2_X1 U5271 ( .A1(n5353), .A2(n3511), .ZN(n4720) );
  NAND2_X1 U5272 ( .A1(n4352), .A2(n4904), .ZN(n4360) );
  OAI21_X1 U5273 ( .B1(n4720), .B2(n5658), .A(n4495), .ZN(n4291) );
  AND3_X1 U5274 ( .A1(n4722), .A2(n4292), .A3(n4291), .ZN(n4293) );
  NAND2_X1 U5275 ( .A1(n4294), .A2(n4293), .ZN(n4731) );
  NAND2_X1 U5276 ( .A1(n6831), .A2(n4352), .ZN(n4959) );
  NAND2_X1 U5277 ( .A1(n3525), .A2(n3514), .ZN(n4487) );
  OAI22_X1 U5278 ( .A1(n4295), .A2(n4909), .B1(n3509), .B2(n4487), .ZN(n4296)
         );
  INV_X1 U5279 ( .A(n4296), .ZN(n4297) );
  NAND2_X1 U5280 ( .A1(n4959), .A2(n4297), .ZN(n4298) );
  AND2_X1 U5281 ( .A1(n6831), .A2(n3201), .ZN(n4803) );
  NAND2_X1 U5282 ( .A1(n4823), .A2(n4803), .ZN(n6817) );
  NAND2_X1 U5283 ( .A1(n4806), .A2(n3522), .ZN(n4299) );
  NAND2_X1 U5284 ( .A1(n6204), .A2(n4299), .ZN(n4313) );
  INV_X1 U5285 ( .A(n4313), .ZN(n4324) );
  XNOR2_X1 U5286 ( .A(n4954), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4302)
         );
  NAND2_X1 U5287 ( .A1(n4308), .A2(n4302), .ZN(n4301) );
  NAND2_X1 U5288 ( .A1(n6838), .A2(n4954), .ZN(n4300) );
  NAND2_X1 U5289 ( .A1(n4301), .A2(n4300), .ZN(n4327) );
  XNOR2_X1 U5290 ( .A(n6844), .B(n4955), .ZN(n4325) );
  XNOR2_X1 U5291 ( .A(n4327), .B(n4325), .ZN(n4658) );
  NAND2_X1 U5292 ( .A1(n4349), .A2(n4658), .ZN(n4323) );
  INV_X1 U5293 ( .A(n4302), .ZN(n4303) );
  XNOR2_X1 U5294 ( .A(n4303), .B(n4308), .ZN(n4659) );
  NAND2_X1 U5295 ( .A1(n4349), .A2(n3201), .ZN(n4306) );
  NAND2_X1 U5296 ( .A1(n4306), .A2(n3522), .ZN(n4317) );
  AND2_X1 U5297 ( .A1(n6830), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4307)
         );
  NOR2_X1 U5298 ( .A1(n4308), .A2(n4307), .ZN(n4312) );
  NAND2_X1 U5299 ( .A1(n4349), .A2(n4312), .ZN(n4309) );
  NAND2_X1 U5300 ( .A1(n4338), .A2(n4309), .ZN(n4316) );
  NAND2_X1 U5301 ( .A1(n4826), .A2(n3522), .ZN(n4584) );
  INV_X1 U5302 ( .A(n4310), .ZN(n4311) );
  AOI21_X1 U5303 ( .B1(n4584), .B2(n4312), .A(n4311), .ZN(n4314) );
  OR2_X1 U5304 ( .A1(n4314), .A2(n4313), .ZN(n4315) );
  OAI211_X1 U5305 ( .C1(n4317), .C2(n4659), .A(n4316), .B(n4315), .ZN(n4319)
         );
  NAND3_X1 U5306 ( .A1(n4317), .A2(STATE2_REG_0__SCAN_IN), .A3(n4659), .ZN(
        n4318) );
  OAI211_X1 U5307 ( .C1(n4659), .C2(n4338), .A(n4319), .B(n4318), .ZN(n4321)
         );
  OAI211_X1 U5308 ( .C1(n4658), .C2(n4335), .A(n4323), .B(n4324), .ZN(n4320)
         );
  NAND2_X1 U5309 ( .A1(n4321), .A2(n4320), .ZN(n4322) );
  OAI21_X1 U5310 ( .B1(n4324), .B2(n4323), .A(n4322), .ZN(n4337) );
  INV_X1 U5311 ( .A(n4325), .ZN(n4326) );
  NAND2_X1 U5312 ( .A1(n4327), .A2(n4326), .ZN(n4329) );
  NAND2_X1 U5313 ( .A1(n6844), .A2(n4955), .ZN(n4328) );
  NAND2_X1 U5314 ( .A1(n4329), .A2(n4328), .ZN(n4334) );
  XNOR2_X1 U5315 ( .A(n6850), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4333)
         );
  INV_X1 U5316 ( .A(n4333), .ZN(n4330) );
  NAND2_X1 U5317 ( .A1(n4334), .A2(n4330), .ZN(n4332) );
  NAND2_X1 U5318 ( .A1(n6850), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4331) );
  NAND2_X1 U5319 ( .A1(n4332), .A2(n4331), .ZN(n4343) );
  XNOR2_X1 U5320 ( .A(n4334), .B(n4333), .ZN(n4657) );
  NAND2_X1 U5321 ( .A1(n4662), .A2(n4657), .ZN(n4339) );
  NAND2_X1 U5322 ( .A1(n4335), .A2(n4339), .ZN(n4336) );
  NAND2_X1 U5323 ( .A1(n4337), .A2(n4336), .ZN(n4341) );
  AOI22_X1 U5324 ( .A1(n4346), .A2(n4339), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6861), .ZN(n4340) );
  NAND2_X1 U5325 ( .A1(n4341), .A2(n4340), .ZN(n4348) );
  NAND2_X1 U5326 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4743), .ZN(n4344) );
  NAND2_X1 U5327 ( .A1(n4346), .A2(n4656), .ZN(n4347) );
  INV_X1 U5328 ( .A(n6822), .ZN(n6207) );
  NAND4_X1 U5329 ( .A1(n4826), .A2(n5811), .A3(n4352), .A4(n3511), .ZN(n4795)
         );
  INV_X1 U5330 ( .A(n4795), .ZN(n4355) );
  INV_X1 U5331 ( .A(n4353), .ZN(n4354) );
  NAND3_X1 U5332 ( .A1(n4355), .A2(n4354), .A3(n4770), .ZN(n4356) );
  NAND2_X1 U5333 ( .A1(n4728), .A2(n4356), .ZN(n4358) );
  NAND2_X1 U5334 ( .A1(n5849), .A2(n4359), .ZN(n4477) );
  INV_X1 U5335 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U5336 ( .A1(n4770), .A2(n4771), .ZN(n4361) );
  OAI211_X1 U5337 ( .C1(n4394), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4361), 
        .B(n4385), .ZN(n4362) );
  NAND2_X1 U5338 ( .A1(n4360), .A2(EBX_REG_0__SCAN_IN), .ZN(n4364) );
  INV_X1 U5339 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U5340 ( .A1(n4385), .A2(n4791), .ZN(n4363) );
  NOR2_X1 U5341 ( .A1(n6363), .A2(n5657), .ZN(n4367) );
  INV_X1 U5342 ( .A(n4365), .ZN(n4366) );
  INV_X1 U5343 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5344 ( .A1(n4466), .A2(n4369), .ZN(n4373) );
  INV_X1 U5345 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U5346 ( .A1(n4360), .A2(n6564), .ZN(n4371) );
  NAND2_X1 U5347 ( .A1(n4770), .A2(n4369), .ZN(n4370) );
  NAND3_X1 U5348 ( .A1(n4371), .A2(n4385), .A3(n4370), .ZN(n4372) );
  NAND2_X1 U5349 ( .A1(n4373), .A2(n4372), .ZN(n4877) );
  INV_X1 U5350 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4482) );
  INV_X1 U5351 ( .A(EBX_REG_3__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U5352 ( .A1(n4770), .A2(n7254), .ZN(n4374) );
  OAI211_X1 U5353 ( .C1(n4470), .C2(n4482), .A(n4360), .B(n4374), .ZN(n4375)
         );
  OAI21_X1 U5354 ( .B1(EBX_REG_3__SCAN_IN), .B2(n4461), .A(n4375), .ZN(n4842)
         );
  INV_X1 U5355 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U5356 ( .A1(n4770), .A2(n6379), .ZN(n4376) );
  OAI211_X1 U5357 ( .C1(n4394), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4376), 
        .B(n4385), .ZN(n4377) );
  OAI21_X1 U5358 ( .B1(n4368), .B2(EBX_REG_4__SCAN_IN), .A(n4377), .ZN(n6318)
         );
  OR2_X1 U5359 ( .A1(n4461), .A2(EBX_REG_5__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5360 ( .A1(n4470), .A2(EBX_REG_5__SCAN_IN), .ZN(n4379) );
  OR2_X1 U5361 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4378)
         );
  NAND3_X1 U5362 ( .A1(n4380), .A2(n4379), .A3(n4378), .ZN(n4995) );
  INV_X1 U5363 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U5364 ( .A1(n4770), .A2(n6377), .ZN(n4381) );
  OAI211_X1 U5365 ( .C1(n4394), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4381), 
        .B(n4385), .ZN(n4382) );
  OAI21_X1 U5366 ( .B1(n4368), .B2(EBX_REG_6__SCAN_IN), .A(n4382), .ZN(n6311)
         );
  NAND2_X1 U5367 ( .A1(n4996), .A2(n6311), .ZN(n5128) );
  NOR2_X1 U5368 ( .A1(n4461), .A2(EBX_REG_7__SCAN_IN), .ZN(n4383) );
  AOI21_X1 U5369 ( .B1(n4470), .B2(EBX_REG_7__SCAN_IN), .A(n4383), .ZN(n4384)
         );
  OAI21_X1 U5370 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5658), .A(n4384), 
        .ZN(n5129) );
  INV_X1 U5371 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U5372 ( .A1(n4466), .A2(n4386), .ZN(n4390) );
  INV_X1 U5373 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U5374 ( .A1(n4360), .A2(n5366), .ZN(n4388) );
  NAND2_X1 U5375 ( .A1(n4770), .A2(n4386), .ZN(n4387) );
  NAND3_X1 U5376 ( .A1(n4388), .A2(n4385), .A3(n4387), .ZN(n4389) );
  NAND2_X1 U5377 ( .A1(n4390), .A2(n4389), .ZN(n5254) );
  NAND2_X1 U5378 ( .A1(EBX_REG_9__SCAN_IN), .A2(n4470), .ZN(n4393) );
  INV_X1 U5379 ( .A(n5658), .ZN(n4391) );
  INV_X1 U5380 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U5381 ( .A1(n4391), .A2(n6485), .ZN(n4392) );
  OAI211_X1 U5382 ( .C1(EBX_REG_9__SCAN_IN), .C2(n4461), .A(n4393), .B(n4392), 
        .ZN(n5377) );
  INV_X1 U5383 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5384 ( .A1(n4466), .A2(n4396), .ZN(n4400) );
  NAND2_X1 U5385 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5386 ( .A1(n4360), .A2(n4395), .ZN(n4398) );
  NAND2_X1 U5387 ( .A1(n4770), .A2(n4396), .ZN(n4397) );
  NAND2_X1 U5388 ( .A1(n4398), .A2(n4397), .ZN(n4399) );
  NAND2_X1 U5389 ( .A1(n4400), .A2(n4399), .ZN(n5459) );
  OR2_X1 U5390 ( .A1(n4461), .A2(EBX_REG_11__SCAN_IN), .ZN(n4404) );
  INV_X1 U5391 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U5392 ( .A1(n4770), .A2(n6375), .ZN(n4402) );
  NAND2_X1 U5393 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4401) );
  NAND3_X1 U5394 ( .A1(n4402), .A2(n4360), .A3(n4401), .ZN(n4403) );
  NAND2_X1 U5395 ( .A1(n4404), .A2(n4403), .ZN(n6269) );
  INV_X1 U5396 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5397 ( .A1(n4466), .A2(n4406), .ZN(n4410) );
  NAND2_X1 U5398 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U5399 ( .A1(n4360), .A2(n4405), .ZN(n4408) );
  NAND2_X1 U5400 ( .A1(n4770), .A2(n4406), .ZN(n4407) );
  NAND2_X1 U5401 ( .A1(n4408), .A2(n4407), .ZN(n4409) );
  NAND2_X1 U5402 ( .A1(n4410), .A2(n4409), .ZN(n5462) );
  OR2_X1 U5403 ( .A1(n4461), .A2(EBX_REG_13__SCAN_IN), .ZN(n4414) );
  INV_X1 U5404 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U5405 ( .A1(n4770), .A2(n6369), .ZN(n4412) );
  NAND2_X1 U5406 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4411) );
  NAND3_X1 U5407 ( .A1(n4412), .A2(n4360), .A3(n4411), .ZN(n4413) );
  NAND2_X1 U5408 ( .A1(n4414), .A2(n4413), .ZN(n6196) );
  INV_X1 U5409 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n7224) );
  OAI21_X1 U5410 ( .B1(n4470), .B2(n7224), .A(n4360), .ZN(n4415) );
  OAI21_X1 U5411 ( .B1(EBX_REG_14__SCAN_IN), .B2(n5657), .A(n4415), .ZN(n4416)
         );
  OAI21_X1 U5412 ( .B1(n4368), .B2(EBX_REG_14__SCAN_IN), .A(n4416), .ZN(n5569)
         );
  INV_X1 U5413 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7218) );
  INV_X1 U5414 ( .A(EBX_REG_15__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U5415 ( .A1(n4770), .A2(n7109), .ZN(n4417) );
  OAI211_X1 U5416 ( .C1(n4470), .C2(n7218), .A(n4417), .B(n4360), .ZN(n4418)
         );
  OAI21_X1 U5417 ( .B1(EBX_REG_15__SCAN_IN), .B2(n4461), .A(n4418), .ZN(n6065)
         );
  INV_X1 U5418 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U5419 ( .A1(n4466), .A2(n5810), .ZN(n4423) );
  NAND2_X1 U5420 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4419) );
  NAND2_X1 U5421 ( .A1(n4360), .A2(n4419), .ZN(n4421) );
  NAND2_X1 U5422 ( .A1(n4770), .A2(n5810), .ZN(n4420) );
  NAND2_X1 U5423 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  NAND2_X1 U5424 ( .A1(n4423), .A2(n4422), .ZN(n5808) );
  NAND2_X1 U5425 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4424) );
  OAI211_X1 U5426 ( .C1(n5657), .C2(EBX_REG_17__SCAN_IN), .A(n4360), .B(n4424), 
        .ZN(n4425) );
  OAI21_X1 U5427 ( .B1(n4461), .B2(EBX_REG_17__SCAN_IN), .A(n4425), .ZN(n5739)
         );
  INV_X1 U5428 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U5429 ( .A1(n4466), .A2(n4426), .ZN(n4430) );
  INV_X1 U5430 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U5431 ( .A1(n4360), .A2(n7237), .ZN(n4428) );
  NAND2_X1 U5432 ( .A1(n4770), .A2(n4426), .ZN(n4427) );
  NAND3_X1 U5433 ( .A1(n4428), .A2(n4385), .A3(n4427), .ZN(n4429) );
  OR2_X1 U5434 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4431)
         );
  INV_X1 U5435 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U5436 ( .A1(n4770), .A2(n5800), .ZN(n5787) );
  OR2_X1 U5437 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4434)
         );
  INV_X1 U5438 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U5439 ( .A1(n4770), .A2(n4432), .ZN(n4433) );
  NAND2_X1 U5440 ( .A1(n4434), .A2(n4433), .ZN(n6032) );
  AOI22_X1 U5441 ( .A1(n6029), .A2(n6032), .B1(n4470), .B2(EBX_REG_20__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U5442 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4438) );
  OAI211_X1 U5443 ( .C1(n5657), .C2(EBX_REG_21__SCAN_IN), .A(n4360), .B(n4438), 
        .ZN(n4439) );
  OAI21_X1 U5444 ( .B1(n4461), .B2(EBX_REG_21__SCAN_IN), .A(n4439), .ZN(n6020)
         );
  INV_X1 U5445 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U5446 ( .A1(n4466), .A2(n6110), .ZN(n4443) );
  INV_X1 U5447 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U5448 ( .A1(n4360), .A2(n7269), .ZN(n4441) );
  NAND2_X1 U5449 ( .A1(n4770), .A2(n6110), .ZN(n4440) );
  NAND3_X1 U5450 ( .A1(n4441), .A2(n4385), .A3(n4440), .ZN(n4442) );
  INV_X1 U5451 ( .A(n4461), .ZN(n4444) );
  INV_X1 U5452 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U5453 ( .A1(n4444), .A2(n6109), .ZN(n4447) );
  NAND2_X1 U5454 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4445) );
  OAI211_X1 U5455 ( .C1(n5657), .C2(EBX_REG_23__SCAN_IN), .A(n4360), .B(n4445), 
        .ZN(n4446) );
  AND2_X1 U5456 ( .A1(n4447), .A2(n4446), .ZN(n5773) );
  INV_X1 U5457 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5458 ( .A1(n4466), .A2(n4672), .ZN(n4451) );
  NAND2_X1 U5459 ( .A1(n4360), .A2(n7174), .ZN(n4449) );
  NAND2_X1 U5460 ( .A1(n4770), .A2(n4672), .ZN(n4448) );
  NAND3_X1 U5461 ( .A1(n4449), .A2(n4385), .A3(n4448), .ZN(n4450) );
  NAND2_X1 U5462 ( .A1(n4451), .A2(n4450), .ZN(n4687) );
  OR2_X1 U5463 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4453)
         );
  NAND2_X1 U5464 ( .A1(n4470), .A2(EBX_REG_25__SCAN_IN), .ZN(n4452) );
  OAI211_X1 U5465 ( .C1(EBX_REG_25__SCAN_IN), .C2(n4461), .A(n4453), .B(n4452), 
        .ZN(n5762) );
  INV_X1 U5466 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U5467 ( .A1(n4466), .A2(n4454), .ZN(n4458) );
  INV_X1 U5468 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U5469 ( .A1(n4360), .A2(n5855), .ZN(n4456) );
  NAND2_X1 U5470 ( .A1(n4770), .A2(n4454), .ZN(n4455) );
  NAND3_X1 U5471 ( .A1(n4456), .A2(n4385), .A3(n4455), .ZN(n4457) );
  AND2_X1 U5472 ( .A1(n4458), .A2(n4457), .ZN(n5755) );
  OR2_X1 U5473 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4460)
         );
  NAND2_X1 U5474 ( .A1(n4470), .A2(EBX_REG_27__SCAN_IN), .ZN(n4459) );
  OAI211_X1 U5475 ( .C1(EBX_REG_27__SCAN_IN), .C2(n4461), .A(n4460), .B(n4459), 
        .ZN(n5725) );
  INV_X1 U5476 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5477 ( .A1(n4360), .A2(n4576), .ZN(n4462) );
  OAI211_X1 U5478 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5657), .A(n4462), .B(n4385), 
        .ZN(n4463) );
  OAI21_X1 U5479 ( .B1(n4368), .B2(EBX_REG_28__SCAN_IN), .A(n4463), .ZN(n5712)
         );
  OR2_X1 U5480 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4465)
         );
  INV_X1 U5481 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U5482 ( .A1(n4770), .A2(n5701), .ZN(n4464) );
  NAND2_X1 U5483 ( .A1(n4465), .A2(n4464), .ZN(n4469) );
  NAND2_X1 U5484 ( .A1(n4466), .A2(n5701), .ZN(n4468) );
  OAI211_X1 U5485 ( .C1(n4470), .C2(n4469), .A(n4467), .B(n4468), .ZN(n4471)
         );
  INV_X1 U5486 ( .A(n4471), .ZN(n4472) );
  NAND2_X1 U5487 ( .A1(n4494), .A2(n4493), .ZN(n4484) );
  NAND2_X1 U5488 ( .A1(n4484), .A2(n4478), .ZN(n4509) );
  INV_X1 U5489 ( .A(n4508), .ZN(n4479) );
  XNOR2_X1 U5490 ( .A(n4509), .B(n4479), .ZN(n4480) );
  NAND2_X1 U5491 ( .A1(n4480), .A2(n4774), .ZN(n4481) );
  XNOR2_X1 U5492 ( .A(n4505), .B(n4482), .ZN(n4937) );
  XNOR2_X1 U5493 ( .A(n4484), .B(n4483), .ZN(n4485) );
  OAI21_X1 U5494 ( .B1(n4485), .B2(n6984), .A(n4487), .ZN(n4486) );
  OAI21_X1 U5495 ( .B1(n6984), .B2(n4493), .A(n4487), .ZN(n4488) );
  INV_X1 U5496 ( .A(n4488), .ZN(n4489) );
  NAND2_X1 U5497 ( .A1(n6467), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4490)
         );
  INV_X1 U5498 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4835) );
  NAND2_X1 U5499 ( .A1(n4490), .A2(n4835), .ZN(n4492) );
  AND2_X1 U5500 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5501 ( .A1(n6467), .A2(n4491), .ZN(n4501) );
  AND2_X1 U5502 ( .A1(n4492), .A2(n4501), .ZN(n4783) );
  NAND2_X1 U5503 ( .A1(n4890), .A2(n3201), .ZN(n4500) );
  XNOR2_X1 U5504 ( .A(n4494), .B(n4493), .ZN(n4497) );
  INV_X1 U5505 ( .A(n4495), .ZN(n4496) );
  OAI211_X1 U5506 ( .C1(n4497), .C2(n6984), .A(n4496), .B(n3522), .ZN(n4498)
         );
  INV_X1 U5507 ( .A(n4498), .ZN(n4499) );
  NAND2_X1 U5508 ( .A1(n4500), .A2(n4499), .ZN(n4782) );
  NAND2_X1 U5509 ( .A1(n4783), .A2(n4782), .ZN(n4502) );
  NAND2_X1 U5510 ( .A1(n4502), .A2(n4501), .ZN(n6457) );
  NAND2_X1 U5511 ( .A1(n6457), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4504)
         );
  INV_X1 U5512 ( .A(n6457), .ZN(n4503) );
  NAND2_X1 U5513 ( .A1(n4937), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5514 ( .A1(n4505), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4506)
         );
  NAND2_X1 U5515 ( .A1(n4938), .A2(n4506), .ZN(n6448) );
  NAND2_X1 U5516 ( .A1(n4507), .A2(n4534), .ZN(n4512) );
  NAND2_X1 U5517 ( .A1(n4509), .A2(n4508), .ZN(n4517) );
  XNOR2_X1 U5518 ( .A(n4517), .B(n4526), .ZN(n4510) );
  NAND2_X1 U5519 ( .A1(n4510), .A2(n4774), .ZN(n4511) );
  INV_X1 U5520 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5521 ( .A1(n6448), .A2(n6450), .ZN(n6449) );
  NAND2_X1 U5522 ( .A1(n4514), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4515)
         );
  NAND2_X1 U5523 ( .A1(n6449), .A2(n4515), .ZN(n5091) );
  NAND2_X1 U5524 ( .A1(n4516), .A2(n4534), .ZN(n4521) );
  INV_X1 U5525 ( .A(n4517), .ZN(n4528) );
  NAND2_X1 U5526 ( .A1(n4528), .A2(n4526), .ZN(n4518) );
  XNOR2_X1 U5527 ( .A(n4518), .B(n4525), .ZN(n4519) );
  NAND2_X1 U5528 ( .A1(n4519), .A2(n4774), .ZN(n4520) );
  NAND2_X1 U5529 ( .A1(n4521), .A2(n4520), .ZN(n4522) );
  INV_X1 U5530 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7294) );
  XNOR2_X1 U5531 ( .A(n4522), .B(n7294), .ZN(n5090) );
  NAND2_X1 U5532 ( .A1(n4522), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4523)
         );
  NAND2_X1 U5533 ( .A1(n5089), .A2(n4523), .ZN(n6443) );
  NAND2_X1 U5534 ( .A1(n4524), .A2(n4534), .ZN(n4531) );
  AND2_X1 U5535 ( .A1(n4526), .A2(n4525), .ZN(n4527) );
  NAND2_X1 U5536 ( .A1(n4528), .A2(n4527), .ZN(n4536) );
  XNOR2_X1 U5537 ( .A(n4536), .B(n4537), .ZN(n4529) );
  NAND2_X1 U5538 ( .A1(n4529), .A2(n4774), .ZN(n4530) );
  NAND2_X1 U5539 ( .A1(n4531), .A2(n4530), .ZN(n4532) );
  INV_X1 U5540 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U5541 ( .A(n4532), .B(n5363), .ZN(n6442) );
  NAND2_X1 U5542 ( .A1(n4532), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4533)
         );
  NAND2_X1 U5543 ( .A1(n4535), .A2(n4534), .ZN(n4542) );
  INV_X1 U5544 ( .A(n4536), .ZN(n4538) );
  NAND2_X1 U5545 ( .A1(n4538), .A2(n4537), .ZN(n4551) );
  XNOR2_X1 U5546 ( .A(n4551), .B(n4539), .ZN(n4540) );
  NAND2_X1 U5547 ( .A1(n4540), .A2(n4774), .ZN(n4541) );
  NAND2_X1 U5548 ( .A1(n4542), .A2(n4541), .ZN(n4543) );
  INV_X1 U5549 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6511) );
  XNOR2_X1 U5550 ( .A(n4543), .B(n6511), .ZN(n5261) );
  NAND2_X1 U5551 ( .A1(n5262), .A2(n5261), .ZN(n5260) );
  NAND2_X1 U5552 ( .A1(n4543), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4544)
         );
  NAND2_X1 U5553 ( .A1(n5260), .A2(n4544), .ZN(n5361) );
  INV_X1 U5554 ( .A(n4546), .ZN(n4548) );
  OR3_X1 U5555 ( .A1(n4551), .A2(n4550), .A3(n6984), .ZN(n4552) );
  NAND2_X1 U5556 ( .A1(n4561), .A2(n4552), .ZN(n4553) );
  XNOR2_X1 U5557 ( .A(n4553), .B(n5366), .ZN(n5360) );
  NAND2_X1 U5558 ( .A1(n4553), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4554)
         );
  INV_X1 U5560 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4557) );
  NAND2_X1 U5561 ( .A1(n3203), .A2(n4557), .ZN(n5535) );
  INV_X1 U5562 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4558) );
  OR2_X1 U5563 ( .A1(n3204), .A2(n4557), .ZN(n6433) );
  INV_X1 U5564 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5555) );
  NOR2_X1 U5565 ( .A1(n3203), .A2(n5555), .ZN(n5543) );
  NAND2_X1 U5566 ( .A1(n3203), .A2(n5555), .ZN(n5541) );
  XNOR2_X1 U5567 ( .A(n3204), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6167)
         );
  INV_X1 U5568 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U5569 ( .A1(n3204), .A2(n4562), .ZN(n4563) );
  NAND2_X1 U5570 ( .A1(n4564), .A2(n4563), .ZN(n5580) );
  XNOR2_X1 U5571 ( .A(n3203), .B(n7218), .ZN(n5947) );
  NAND2_X1 U5572 ( .A1(n3203), .A2(n7218), .ZN(n4565) );
  INV_X1 U5573 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U5574 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U5575 ( .A1(n3204), .A2(n5606), .ZN(n4566) );
  INV_X1 U5576 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7215) );
  INV_X1 U5577 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6053) );
  AND3_X1 U5578 ( .A1(n7215), .A2(n6053), .A3(n7164), .ZN(n4567) );
  NOR2_X1 U5579 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U5580 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6038) );
  INV_X1 U5581 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5889) );
  NAND4_X1 U5582 ( .A1(n6014), .A2(n6038), .A3(n5889), .A4(n7174), .ZN(n4569)
         );
  NAND2_X1 U5583 ( .A1(n4555), .A2(n4569), .ZN(n4570) );
  AND2_X1 U5584 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6037) );
  AND2_X1 U5585 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6013) );
  AND2_X1 U5586 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5610) );
  NAND3_X1 U5587 ( .A1(n6037), .A2(n6013), .A3(n5610), .ZN(n4571) );
  XOR2_X1 U5588 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n3204), .Z(n5878) );
  INV_X1 U5589 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U5590 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5972) );
  INV_X1 U5591 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5958) );
  INV_X1 U5592 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5630) );
  NOR2_X1 U5593 ( .A1(n5958), .A2(n5630), .ZN(n4578) );
  INV_X1 U5594 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U5595 ( .A1(n5982), .A2(n4576), .ZN(n5973) );
  OR3_X1 U5596 ( .A1(n3204), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5973), 
        .ZN(n4639) );
  NOR3_X1 U5597 ( .A1(n4639), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4577) );
  NAND2_X1 U5598 ( .A1(n4581), .A2(n3525), .ZN(n4582) );
  NAND2_X1 U5599 ( .A1(n4583), .A2(n4582), .ZN(n4721) );
  INV_X1 U5600 ( .A(n4585), .ZN(n4586) );
  NAND2_X1 U5601 ( .A1(n4586), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4628)
         );
  XNOR2_X1 U5602 ( .A(n4628), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5675)
         );
  NAND2_X1 U5603 ( .A1(n4588), .A2(n4587), .ZN(n4613) );
  INV_X1 U5604 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U5605 ( .A1(n3774), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4589), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5606 ( .A1(n4590), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4591)
         );
  OAI211_X1 U5607 ( .C1(n5039), .C2(n3629), .A(n4592), .B(n4591), .ZN(n4601)
         );
  INV_X1 U5608 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4595) );
  INV_X1 U5609 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4593) );
  OAI22_X1 U5610 ( .A1(n4596), .A2(n4595), .B1(n4594), .B2(n4593), .ZN(n4600)
         );
  OAI22_X1 U5611 ( .A1(n3440), .A2(n4598), .B1(n4597), .B2(n5242), .ZN(n4599)
         );
  OR3_X1 U5612 ( .A1(n4601), .A2(n4600), .A3(n4599), .ZN(n4611) );
  AOI22_X1 U5613 ( .A1(n4603), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4602), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4609) );
  AOI22_X1 U5614 ( .A1(n4245), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3722), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U5615 ( .A1(n3723), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5616 ( .A1(n4246), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4606) );
  NAND4_X1 U5617 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4610)
         );
  NOR2_X1 U5618 ( .A1(n4611), .A2(n4610), .ZN(n4612) );
  XOR2_X1 U5619 ( .A(n4613), .B(n4612), .Z(n4619) );
  INV_X1 U5620 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U5621 ( .A1(n3658), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4614)
         );
  OAI211_X1 U5622 ( .C1(n4616), .C2(n4615), .A(n4614), .B(n3758), .ZN(n4617)
         );
  AOI21_X1 U5623 ( .B1(n4619), .B2(n4618), .A(n4617), .ZN(n4620) );
  AOI21_X1 U5624 ( .B1(n5675), .B2(n4621), .A(n4620), .ZN(n4643) );
  NAND2_X1 U5625 ( .A1(n4644), .A2(n4643), .ZN(n4626) );
  AOI22_X1 U5626 ( .A1(n4623), .A2(EAX_REG_31__SCAN_IN), .B1(n4622), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4624) );
  XNOR2_X2 U5627 ( .A(n4626), .B(n4625), .ZN(n5812) );
  NAND3_X1 U5628 ( .A1(n6861), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6875) );
  INV_X1 U5629 ( .A(n6875), .ZN(n4627) );
  NOR2_X2 U5630 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6753) );
  NAND2_X1 U5631 ( .A1(n4627), .A2(n6753), .ZN(n6470) );
  NAND2_X1 U5632 ( .A1(n5812), .A2(n6461), .ZN(n4638) );
  INV_X1 U5633 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4645) );
  INV_X1 U5634 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U5635 ( .A1(n6658), .A2(n4634), .ZN(n6980) );
  NAND2_X1 U5636 ( .A1(n6980), .A2(n6861), .ZN(n4630) );
  NAND2_X1 U5637 ( .A1(n6861), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5638 ( .A1(n6213), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4631) );
  AND2_X1 U5639 ( .A1(n4632), .A2(n4631), .ZN(n6475) );
  INV_X1 U5640 ( .A(n6475), .ZN(n4633) );
  INV_X2 U5641 ( .A(n6556), .ZN(n6567) );
  NAND2_X1 U5642 ( .A1(n6567), .A2(REIP_REG_31__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U5643 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4635)
         );
  OAI211_X1 U5644 ( .C1(n4686), .C2(n6466), .A(n5665), .B(n4635), .ZN(n4636)
         );
  INV_X1 U5645 ( .A(n4636), .ZN(n4637) );
  OAI211_X1 U5646 ( .C1(n5669), .C2(n6468), .A(n4638), .B(n4637), .ZN(U2955)
         );
  NAND2_X1 U5647 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U5648 ( .A1(n5851), .A2(n4639), .ZN(n5843) );
  XNOR2_X1 U5649 ( .A(n4644), .B(n4643), .ZN(n5670) );
  NOR2_X1 U5650 ( .A1(n5670), .A2(n6470), .ZN(n4650) );
  NAND2_X1 U5651 ( .A1(n5675), .A2(n6438), .ZN(n4648) );
  NAND2_X1 U5652 ( .A1(n6567), .A2(REIP_REG_30__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U5653 ( .B1(n6474), .B2(n4645), .A(n5631), .ZN(n4646) );
  INV_X1 U5654 ( .A(n4646), .ZN(n4647) );
  NAND2_X1 U5655 ( .A1(n4648), .A2(n4647), .ZN(n4649) );
  NOR2_X1 U5656 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  OAI21_X1 U5657 ( .B1(n5636), .B2(n6468), .A(n4651), .ZN(U2956) );
  INV_X1 U5658 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7268) );
  INV_X1 U5659 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5467) );
  INV_X1 U5660 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4652) );
  AND2_X1 U5661 ( .A1(n4653), .A2(n4652), .ZN(n6883) );
  INV_X1 U5662 ( .A(n6883), .ZN(n6214) );
  NAND2_X1 U5663 ( .A1(n4806), .A2(n6214), .ZN(n4811) );
  NAND2_X1 U5664 ( .A1(n6981), .A2(n6213), .ZN(n4689) );
  INV_X1 U5665 ( .A(n4656), .ZN(n4661) );
  NAND3_X1 U5666 ( .A1(n4659), .A2(n4658), .A3(n4657), .ZN(n4660) );
  NAND2_X1 U5667 ( .A1(n4661), .A2(n4660), .ZN(n4663) );
  NOR2_X1 U5668 ( .A1(n6820), .A2(n6865), .ZN(n4664) );
  NAND2_X1 U5669 ( .A1(n6819), .A2(n4664), .ZN(n4698) );
  NOR3_X1 U5670 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6952), .A3(n3758), .ZN(
        n6869) );
  OR2_X1 U5671 ( .A1(n6567), .A2(n6869), .ZN(n4665) );
  NAND2_X1 U5672 ( .A1(n6952), .A2(n3658), .ZN(n6862) );
  NOR3_X1 U5673 ( .A1(n6861), .A2(n7315), .A3(n6862), .ZN(n6859) );
  OR2_X1 U5674 ( .A1(n4665), .A2(n6859), .ZN(n4666) );
  OR2_X2 U5675 ( .A1(n6979), .A2(n4666), .ZN(n6333) );
  NOR2_X1 U5676 ( .A1(n4689), .A2(n5294), .ZN(n4667) );
  AND2_X1 U5677 ( .A1(n4904), .A2(n4667), .ZN(n4668) );
  INV_X1 U5678 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7187) );
  INV_X1 U5679 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6899) );
  INV_X1 U5680 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7300) );
  INV_X1 U5681 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7306) );
  INV_X1 U5682 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6895) );
  NOR3_X1 U5683 ( .A1(n7300), .A2(n7306), .A3(n6895), .ZN(n6321) );
  NAND2_X1 U5684 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6321), .ZN(n5296) );
  NOR2_X1 U5685 ( .A1(n6899), .A2(n5296), .ZN(n5434) );
  NAND2_X1 U5686 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5434), .ZN(n5436) );
  NOR2_X1 U5687 ( .A1(n7187), .A2(n5436), .ZN(n6298) );
  NAND2_X1 U5688 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6298), .ZN(n4673) );
  NAND4_X1 U5689 ( .A1(n6289), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U5690 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6264), .ZN(n5568) );
  INV_X1 U5691 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6913) );
  INV_X1 U5692 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6912) );
  INV_X1 U5693 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7291) );
  INV_X1 U5694 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6914) );
  INV_X1 U5695 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6915) );
  NOR3_X1 U5696 ( .A1(n7291), .A2(n6914), .A3(n6915), .ZN(n4676) );
  NAND4_X1 U5697 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n6125), .ZN(n6080) );
  NOR2_X1 U5698 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6080), .ZN(n6096) );
  INV_X1 U5699 ( .A(n4689), .ZN(n4669) );
  NAND2_X1 U5700 ( .A1(n6883), .A2(n4669), .ZN(n6855) );
  NAND2_X1 U5701 ( .A1(n4774), .A2(n6855), .ZN(n5693) );
  INV_X1 U5702 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5747) );
  NAND3_X1 U5703 ( .A1(n4904), .A2(n5747), .A3(n4689), .ZN(n4670) );
  NAND2_X1 U5704 ( .A1(n5693), .A2(n4670), .ZN(n4671) );
  INV_X1 U5705 ( .A(n5294), .ZN(n5352) );
  OAI22_X1 U5706 ( .A1(n4672), .A2(n6331), .B1(n7223), .B2(n6354), .ZN(n4693)
         );
  NAND3_X1 U5707 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4675) );
  NAND3_X1 U5708 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n4674) );
  INV_X1 U5709 ( .A(n6333), .ZN(n6351) );
  NOR2_X1 U5710 ( .A1(n4674), .A2(n6277), .ZN(n6258) );
  NAND4_X1 U5711 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n6258), .ZN(n5567) );
  NOR2_X1 U5712 ( .A1(n4675), .A2(n5567), .ZN(n5737) );
  NAND2_X1 U5713 ( .A1(n5737), .A2(n4676), .ZN(n4677) );
  NAND2_X1 U5714 ( .A1(n6333), .A2(n6334), .ZN(n6278) );
  NAND2_X1 U5715 ( .A1(n4677), .A2(n6278), .ZN(n6137) );
  AND3_X1 U5716 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4678) );
  OR2_X1 U5717 ( .A1(n6334), .A2(n4678), .ZN(n4679) );
  INV_X1 U5718 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U5719 ( .A1(n6333), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4685) );
  INV_X1 U5720 ( .A(n4685), .ZN(n4680) );
  OAI22_X1 U5721 ( .A1(n6103), .A2(n6921), .B1(n5648), .B2(n6343), .ZN(n4692)
         );
  AND2_X1 U5722 ( .A1(n4682), .A2(n4683), .ZN(n4684) );
  NOR2_X1 U5723 ( .A1(n4681), .A2(n4684), .ZN(n5650) );
  INV_X1 U5724 ( .A(n5650), .ZN(n5830) );
  OR2_X1 U5725 ( .A1(n5775), .A2(n4687), .ZN(n4688) );
  NAND2_X1 U5726 ( .A1(n5763), .A2(n4688), .ZN(n5767) );
  OAI22_X1 U5727 ( .A1(n5830), .A2(n6302), .B1(n5767), .B2(n6362), .ZN(n4691)
         );
  OR4_X1 U5728 ( .A1(n6096), .A2(n4693), .A3(n4692), .A4(n4691), .ZN(U2803) );
  AND2_X1 U5729 ( .A1(n6819), .A2(n3201), .ZN(n6834) );
  OR2_X1 U5730 ( .A1(n4695), .A2(n6984), .ZN(n6856) );
  INV_X1 U5731 ( .A(n6856), .ZN(n4696) );
  OAI21_X1 U5732 ( .B1(n6834), .B2(n4696), .A(n6883), .ZN(n4697) );
  NOR2_X1 U5733 ( .A1(n6952), .A2(n3658), .ZN(n4984) );
  NAND2_X1 U5734 ( .A1(n4984), .A2(n6861), .ZN(n6419) );
  AND2_X2 U5735 ( .A1(n6422), .A2(n6419), .ZN(n6420) );
  AND2_X1 U5736 ( .A1(n6420), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U5737 ( .A(n4698), .ZN(n4700) );
  INV_X1 U5738 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7154) );
  NOR2_X1 U5739 ( .A1(n6658), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5298) );
  INV_X1 U5740 ( .A(n5298), .ZN(n4699) );
  OAI211_X1 U5741 ( .C1(n4700), .C2(n7154), .A(n4778), .B(n4699), .ZN(U2788)
         );
  INV_X1 U5742 ( .A(n6979), .ZN(n4703) );
  INV_X1 U5743 ( .A(n5353), .ZN(n4701) );
  NAND2_X1 U5744 ( .A1(n6984), .A2(n4701), .ZN(n6215) );
  OAI21_X1 U5745 ( .B1(n5298), .B2(READREQUEST_REG_SCAN_IN), .A(n4703), .ZN(
        n4702) );
  OAI21_X1 U5746 ( .B1(n4703), .B2(n6215), .A(n4702), .ZN(U3474) );
  INV_X1 U5747 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U5748 ( .A1(n6415), .A2(n4904), .ZN(n6395) );
  INV_X2 U5749 ( .A(n6419), .ZN(n6982) );
  AOI22_X1 U5750 ( .A1(n6982), .A2(UWORD_REG_3__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4704) );
  OAI21_X1 U5751 ( .B1(n4854), .B2(n6395), .A(n4704), .ZN(U2904) );
  AOI22_X1 U5752 ( .A1(n6982), .A2(UWORD_REG_5__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4705) );
  OAI21_X1 U5753 ( .B1(n4082), .B2(n6395), .A(n4705), .ZN(U2902) );
  AOI22_X1 U5754 ( .A1(n6982), .A2(UWORD_REG_6__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4706) );
  OAI21_X1 U5755 ( .B1(n4106), .B2(n6395), .A(n4706), .ZN(U2901) );
  INV_X1 U5756 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5757 ( .A1(n6982), .A2(UWORD_REG_7__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4707) );
  OAI21_X1 U5758 ( .B1(n4856), .B2(n6395), .A(n4707), .ZN(U2900) );
  AOI22_X1 U5759 ( .A1(n6982), .A2(UWORD_REG_9__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4708) );
  OAI21_X1 U5760 ( .B1(n4186), .B2(n6395), .A(n4708), .ZN(U2898) );
  AOI22_X1 U5761 ( .A1(n6982), .A2(UWORD_REG_1__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4709) );
  OAI21_X1 U5762 ( .B1(n3996), .B2(n6395), .A(n4709), .ZN(U2906) );
  AOI22_X1 U5763 ( .A1(n6982), .A2(UWORD_REG_2__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4710) );
  OAI21_X1 U5764 ( .B1(n4022), .B2(n6395), .A(n4710), .ZN(U2905) );
  AOI22_X1 U5765 ( .A1(n6982), .A2(UWORD_REG_14__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4711) );
  OAI21_X1 U5766 ( .B1(n4615), .B2(n6395), .A(n4711), .ZN(U2893) );
  AOI22_X1 U5767 ( .A1(n6982), .A2(UWORD_REG_0__SCAN_IN), .B1(
        DATAO_REG_16__SCAN_IN), .B2(n6420), .ZN(n4712) );
  OAI21_X1 U5768 ( .B1(n3976), .B2(n6395), .A(n4712), .ZN(U2907) );
  INV_X1 U5769 ( .A(n6420), .ZN(n6417) );
  INV_X1 U5770 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n7278) );
  INV_X1 U5771 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4848) );
  INV_X1 U5772 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4713) );
  OAI222_X1 U5773 ( .A1(n6417), .A2(n7278), .B1(n6395), .B2(n4848), .C1(n4713), 
        .C2(n6419), .ZN(U2896) );
  INV_X1 U5774 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n7133) );
  INV_X1 U5775 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4714) );
  OAI222_X1 U5776 ( .A1(n6417), .A2(n7133), .B1(n6395), .B2(n4062), .C1(n4714), 
        .C2(n6419), .ZN(U2903) );
  NOR2_X1 U5777 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7315), .ZN(n6943) );
  OR2_X1 U5778 ( .A1(n4721), .A2(n6204), .ZN(n6818) );
  NOR2_X1 U5779 ( .A1(n6820), .A2(READY_N), .ZN(n4805) );
  INV_X1 U5780 ( .A(n4805), .ZN(n4716) );
  OAI22_X1 U5781 ( .A1(n6822), .A2(n6818), .B1(n4715), .B2(n4716), .ZN(n4798)
         );
  NOR2_X1 U5782 ( .A1(n4770), .A2(n6883), .ZN(n4718) );
  NAND2_X1 U5783 ( .A1(n6834), .A2(n6883), .ZN(n4717) );
  OAI21_X1 U5784 ( .B1(n4718), .B2(n4695), .A(n4717), .ZN(n4719) );
  NAND2_X1 U5785 ( .A1(n4719), .A2(n6981), .ZN(n4726) );
  INV_X1 U5786 ( .A(n4720), .ZN(n4725) );
  INV_X1 U5787 ( .A(n6819), .ZN(n6205) );
  INV_X1 U5788 ( .A(n4721), .ZN(n4723) );
  NAND2_X1 U5789 ( .A1(n4723), .A2(n4722), .ZN(n4724) );
  NAND2_X1 U5790 ( .A1(n6205), .A2(n4724), .ZN(n4808) );
  OAI211_X1 U5791 ( .C1(n6822), .C2(n4726), .A(n4725), .B(n4808), .ZN(n4727)
         );
  NOR2_X1 U5792 ( .A1(n4798), .A2(n4727), .ZN(n4729) );
  NAND2_X1 U5793 ( .A1(n4729), .A2(n4728), .ZN(n6835) );
  INV_X1 U5794 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6217) );
  NAND2_X1 U5795 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4984), .ZN(n6944) );
  OAI22_X1 U5796 ( .A1(n4965), .A2(n6865), .B1(n6217), .B2(n6944), .ZN(n4745)
         );
  NOR2_X1 U5797 ( .A1(n6943), .A2(n4745), .ZN(n6959) );
  INV_X1 U5798 ( .A(n4731), .ZN(n4734) );
  AND4_X1 U5799 ( .A1(n4715), .A2(n4732), .A3(n4695), .A4(n4295), .ZN(n4733)
         );
  NAND2_X1 U5800 ( .A1(n4734), .A2(n4733), .ZN(n6832) );
  INV_X1 U5801 ( .A(n6832), .ZN(n4739) );
  AND2_X1 U5802 ( .A1(n6834), .A2(n4735), .ZN(n4751) );
  INV_X1 U5803 ( .A(n4751), .ZN(n4738) );
  INV_X1 U5804 ( .A(n4950), .ZN(n4749) );
  INV_X1 U5805 ( .A(n4736), .ZN(n4969) );
  NAND3_X1 U5806 ( .A1(n6831), .A2(n4749), .A3(n4969), .ZN(n4737) );
  OAI211_X1 U5807 ( .C1(n6074), .C2(n4739), .A(n4738), .B(n4737), .ZN(n6836)
         );
  INV_X1 U5808 ( .A(n6962), .ZN(n4762) );
  INV_X1 U5809 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6575) );
  NOR2_X1 U5810 ( .A1(n6952), .A2(n6575), .ZN(n4740) );
  AOI22_X1 U5811 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4579), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4835), .ZN(n4758) );
  NOR2_X1 U5812 ( .A1(n6953), .A2(n4950), .ZN(n4763) );
  AOI222_X1 U5813 ( .A1(n6836), .A2(n4762), .B1(n4740), .B2(n4758), .C1(n4969), 
        .C2(n4763), .ZN(n4742) );
  NAND2_X1 U5814 ( .A1(n6959), .A2(n4954), .ZN(n4741) );
  OAI21_X1 U5815 ( .B1(n6959), .B2(n4742), .A(n4741), .ZN(U3460) );
  INV_X1 U5816 ( .A(n6959), .ZN(n6957) );
  INV_X1 U5817 ( .A(n4715), .ZN(n4970) );
  INV_X1 U5818 ( .A(n6654), .ZN(n5148) );
  NOR2_X1 U5819 ( .A1(n3678), .A2(n5148), .ZN(n4744) );
  XNOR2_X1 U5820 ( .A(n4744), .B(n4743), .ZN(n6324) );
  NAND4_X1 U5821 ( .A1(n4745), .A2(n4762), .A3(n4970), .A4(n6324), .ZN(n4746)
         );
  OAI21_X1 U5822 ( .B1(n6957), .B2(n4743), .A(n4746), .ZN(U3455) );
  NAND2_X1 U5823 ( .A1(n6817), .A2(n6818), .ZN(n4962) );
  INV_X1 U5824 ( .A(n4959), .ZN(n4750) );
  MUX2_X1 U5825 ( .A(n4962), .B(n4750), .S(n4950), .Z(n4748) );
  AND2_X1 U5826 ( .A1(n6834), .A2(n4954), .ZN(n4747) );
  NOR2_X1 U5827 ( .A1(n4748), .A2(n4747), .ZN(n4754) );
  MUX2_X1 U5828 ( .A(n4962), .B(n4750), .S(n4749), .Z(n4752) );
  NOR2_X1 U5829 ( .A1(n4752), .A2(n4751), .ZN(n4753) );
  MUX2_X1 U5830 ( .A(n4754), .B(n4753), .S(n4955), .Z(n4757) );
  INV_X1 U5831 ( .A(n4755), .ZN(n5052) );
  NAND2_X1 U5832 ( .A1(n5052), .A2(n6832), .ZN(n4756) );
  NAND2_X1 U5833 ( .A1(n4757), .A2(n4756), .ZN(n4947) );
  NAND2_X1 U5834 ( .A1(n4950), .A2(n3304), .ZN(n4760) );
  OR3_X1 U5835 ( .A1(n6952), .A2(n6575), .A3(n4758), .ZN(n4759) );
  OAI21_X1 U5836 ( .B1(n6953), .B2(n4760), .A(n4759), .ZN(n4761) );
  AOI21_X1 U5837 ( .B1(n4947), .B2(n4762), .A(n4761), .ZN(n4765) );
  OAI21_X1 U5838 ( .B1(n6959), .B2(n4763), .A(n4955), .ZN(n4764) );
  OAI21_X1 U5839 ( .B1(n6959), .B2(n4765), .A(n4764), .ZN(U3459) );
  NOR2_X1 U5840 ( .A1(n4766), .A2(n4767), .ZN(n4768) );
  NOR2_X1 U5841 ( .A1(n4769), .A2(n4768), .ZN(n6347) );
  XNOR2_X1 U5842 ( .A(n6363), .B(n4770), .ZN(n4833) );
  OAI22_X1 U5843 ( .A1(n6371), .A2(n4833), .B1(n6380), .B2(n4771), .ZN(n4772)
         );
  AOI21_X1 U5844 ( .B1(n6347), .B2(n4359), .A(n4772), .ZN(n4773) );
  INV_X1 U5845 ( .A(n4773), .ZN(U2858) );
  INV_X1 U5846 ( .A(READY_N), .ZN(n6981) );
  NOR2_X1 U5847 ( .A1(n4774), .A2(n6981), .ZN(n4775) );
  NOR2_X2 U5848 ( .A1(n4778), .A2(n4775), .ZN(n4886) );
  INV_X1 U5849 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n7316) );
  AND2_X1 U5850 ( .A1(n3201), .A2(n6981), .ZN(n4776) );
  NAND2_X1 U5851 ( .A1(n4858), .A2(DATAI_12_), .ZN(n6427) );
  NOR2_X1 U5852 ( .A1(n4778), .A2(n3201), .ZN(n6429) );
  NAND2_X1 U5853 ( .A1(n6429), .A2(EAX_REG_28__SCAN_IN), .ZN(n4779) );
  OAI211_X1 U5854 ( .C1(n4886), .C2(n7316), .A(n6427), .B(n4779), .ZN(U2936)
         );
  INV_X1 U5855 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U5856 ( .A1(n4858), .A2(DATAI_13_), .ZN(n4846) );
  NAND2_X1 U5857 ( .A1(n6429), .A2(EAX_REG_29__SCAN_IN), .ZN(n4780) );
  OAI211_X1 U5858 ( .C1(n4886), .C2(n7175), .A(n4846), .B(n4780), .ZN(U2937)
         );
  INV_X1 U5859 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U5860 ( .A1(n4858), .A2(DATAI_8_), .ZN(n6423) );
  NAND2_X1 U5861 ( .A1(n6429), .A2(EAX_REG_24__SCAN_IN), .ZN(n4781) );
  OAI211_X1 U5862 ( .C1(n4886), .C2(n7151), .A(n6423), .B(n4781), .ZN(U2932)
         );
  XNOR2_X1 U5863 ( .A(n4783), .B(n4782), .ZN(n4838) );
  NAND2_X1 U5864 ( .A1(n6347), .A2(n6461), .ZN(n4786) );
  OAI22_X1 U5865 ( .A1(n6474), .A2(n6356), .B1(n6556), .B2(n6895), .ZN(n4784)
         );
  AOI21_X1 U5866 ( .B1(n6438), .B2(n6356), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5867 ( .C1(n4838), .C2(n6468), .A(n4786), .B(n4785), .ZN(U2985)
         );
  NOR2_X1 U5868 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4787)
         );
  OR2_X1 U5869 ( .A1(n4788), .A2(n4787), .ZN(n5354) );
  XOR2_X1 U5870 ( .A(n4790), .B(n4789), .Z(n6471) );
  OAI222_X1 U5871 ( .A1(n5354), .A2(n6371), .B1(n6380), .B2(n4791), .C1(n6152), 
        .C2(n6471), .ZN(U2859) );
  AOI22_X1 U5872 ( .A1(n6430), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6429), .ZN(n4792) );
  NAND2_X1 U5873 ( .A1(n4858), .A2(DATAI_10_), .ZN(n4793) );
  NAND2_X1 U5874 ( .A1(n4792), .A2(n4793), .ZN(U2949) );
  AOI22_X1 U5875 ( .A1(n6430), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6429), .ZN(n4794) );
  NAND2_X1 U5876 ( .A1(n4794), .A2(n4793), .ZN(U2934) );
  OR2_X1 U5877 ( .A1(n6204), .A2(n4353), .ZN(n4796) );
  NOR2_X1 U5878 ( .A1(n4796), .A2(n4795), .ZN(n4797) );
  OAI21_X1 U5879 ( .B1(n4798), .B2(n4797), .A(n6867), .ZN(n4799) );
  NAND2_X1 U5880 ( .A1(n3503), .A2(n3499), .ZN(n4800) );
  NAND2_X2 U5881 ( .A1(n6394), .A2(n4800), .ZN(n6156) );
  INV_X1 U5882 ( .A(n4800), .ZN(n4801) );
  INV_X1 U5883 ( .A(DATAI_0_), .ZN(n4905) );
  INV_X1 U5884 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7271) );
  OAI222_X1 U5885 ( .A1(n6156), .A2(n6471), .B1(n5577), .B2(n4905), .C1(n6394), 
        .C2(n7271), .ZN(U2891) );
  INV_X1 U5886 ( .A(n6347), .ZN(n4802) );
  INV_X1 U5887 ( .A(DATAI_1_), .ZN(n4921) );
  INV_X1 U5888 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6418) );
  OAI222_X1 U5889 ( .A1(n4802), .A2(n6156), .B1(n5577), .B2(n4921), .C1(n6394), 
        .C2(n6418), .ZN(U2890) );
  NAND2_X1 U5890 ( .A1(n6822), .A2(n4803), .ZN(n4809) );
  OAI211_X1 U5891 ( .C1(n4806), .C2(n6883), .A(n4804), .B(n4805), .ZN(n4807)
         );
  NAND3_X1 U5892 ( .A1(n4809), .A2(n4808), .A3(n4807), .ZN(n4810) );
  NAND2_X1 U5893 ( .A1(n4810), .A2(n6867), .ZN(n4818) );
  NAND2_X1 U5894 ( .A1(n4811), .A2(n6981), .ZN(n4813) );
  INV_X1 U5895 ( .A(n5684), .ZN(n4812) );
  OAI211_X1 U5896 ( .C1(n4695), .C2(n4813), .A(n4904), .B(n4812), .ZN(n4814)
         );
  NAND2_X1 U5897 ( .A1(n4814), .A2(n3511), .ZN(n4815) );
  OAI22_X1 U5898 ( .A1(n4695), .A2(n5657), .B1(n4819), .B2(n4826), .ZN(n4820)
         );
  INV_X1 U5899 ( .A(n4820), .ZN(n4821) );
  NAND4_X1 U5900 ( .A1(n4715), .A2(n4821), .A3(n6818), .A4(n6825), .ZN(n4822)
         );
  INV_X1 U5901 ( .A(n4823), .ZN(n4824) );
  INV_X1 U5902 ( .A(n6817), .ZN(n4825) );
  INV_X1 U5903 ( .A(n6558), .ZN(n5611) );
  NAND2_X1 U5904 ( .A1(n4831), .A2(n6834), .ZN(n5585) );
  NOR2_X1 U5905 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5605), .ZN(n5362)
         );
  NOR2_X1 U5906 ( .A1(n6518), .A2(n5362), .ZN(n4836) );
  NAND3_X1 U5907 ( .A1(n4827), .A2(n4826), .A3(n5684), .ZN(n4828) );
  NAND2_X1 U5908 ( .A1(n6856), .A2(n4828), .ZN(n4829) );
  INV_X1 U5909 ( .A(n5607), .ZN(n4830) );
  NOR2_X1 U5910 ( .A1(n4830), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6570)
         );
  NOR2_X1 U5911 ( .A1(n4831), .A2(n6567), .ZN(n5604) );
  NOR2_X1 U5912 ( .A1(n6570), .A2(n5604), .ZN(n5364) );
  INV_X1 U5913 ( .A(n5364), .ZN(n6516) );
  AOI22_X1 U5914 ( .A1(n6567), .A2(REIP_REG_1__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6516), .ZN(n4832) );
  OAI21_X1 U5915 ( .B1(n6551), .B2(n4833), .A(n4832), .ZN(n4834) );
  AOI21_X1 U5916 ( .B1(n4836), .B2(n4835), .A(n4834), .ZN(n4837) );
  OAI21_X1 U5917 ( .B1(n4838), .B2(n6478), .A(n4837), .ZN(U3017) );
  OAI21_X1 U5918 ( .B1(n4839), .B2(n4841), .A(n4840), .ZN(n5454) );
  AOI21_X1 U5919 ( .B1(n4842), .B2(n4879), .A(n6319), .ZN(n6544) );
  AOI22_X1 U5920 ( .A1(n4474), .A2(n6544), .B1(n5802), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4843) );
  OAI21_X1 U5921 ( .B1(n5454), .B2(n6152), .A(n4843), .ZN(U2856) );
  NAND2_X1 U5922 ( .A1(n4858), .A2(DATAI_14_), .ZN(n6431) );
  NAND2_X1 U5923 ( .A1(n6430), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4844) );
  OAI211_X1 U5924 ( .C1(n4884), .C2(n4615), .A(n6431), .B(n4844), .ZN(U2938)
         );
  NAND2_X1 U5925 ( .A1(n6430), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4845) );
  OAI211_X1 U5926 ( .C1(n4884), .C2(n3885), .A(n4846), .B(n4845), .ZN(U2952)
         );
  NAND2_X1 U5927 ( .A1(n4858), .A2(DATAI_11_), .ZN(n6425) );
  NAND2_X1 U5928 ( .A1(n6430), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4847) );
  OAI211_X1 U5929 ( .C1(n4884), .C2(n4848), .A(n6425), .B(n4847), .ZN(U2935)
         );
  AOI22_X1 U5930 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_5_), .ZN(n4849) );
  OAI21_X1 U5931 ( .B1(n4082), .B2(n4884), .A(n4849), .ZN(U2929) );
  AOI22_X1 U5932 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_4_), .ZN(n4850) );
  OAI21_X1 U5933 ( .B1(n4062), .B2(n4884), .A(n4850), .ZN(U2928) );
  AOI22_X1 U5934 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_9_), .ZN(n4851) );
  OAI21_X1 U5935 ( .B1(n4186), .B2(n4884), .A(n4851), .ZN(U2933) );
  AOI22_X1 U5936 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_0_), .ZN(n4852) );
  OAI21_X1 U5937 ( .B1(n3976), .B2(n4884), .A(n4852), .ZN(U2924) );
  AOI22_X1 U5938 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_3_), .ZN(n4853) );
  OAI21_X1 U5939 ( .B1(n4854), .B2(n4884), .A(n4853), .ZN(U2927) );
  AOI22_X1 U5940 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_7_), .ZN(n4855) );
  OAI21_X1 U5941 ( .B1(n4856), .B2(n4884), .A(n4855), .ZN(U2931) );
  AOI22_X1 U5942 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_1_), .ZN(n4857) );
  OAI21_X1 U5943 ( .B1(n3996), .B2(n4884), .A(n4857), .ZN(U2925) );
  AOI22_X1 U5944 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6430), .B1(n4858), .B2(
        DATAI_2_), .ZN(n4859) );
  OAI21_X1 U5945 ( .B1(n4022), .B2(n4884), .A(n4859), .ZN(U2926) );
  INV_X1 U5946 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4861) );
  INV_X1 U5947 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n4860) );
  INV_X1 U5948 ( .A(DATAI_2_), .ZN(n4944) );
  OAI222_X1 U5949 ( .A1(n4884), .A2(n4861), .B1(n4860), .B2(n4886), .C1(n4887), 
        .C2(n4944), .ZN(U2941) );
  INV_X1 U5950 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4862) );
  OAI222_X1 U5951 ( .A1(n4884), .A2(n6418), .B1(n4862), .B2(n4886), .C1(n4887), 
        .C2(n4921), .ZN(U2940) );
  INV_X1 U5952 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4864) );
  INV_X1 U5953 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n4863) );
  INV_X1 U5954 ( .A(DATAI_9_), .ZN(n5444) );
  OAI222_X1 U5955 ( .A1(n4884), .A2(n4864), .B1(n4863), .B2(n4886), .C1(n4887), 
        .C2(n5444), .ZN(U2948) );
  INV_X1 U5956 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4865) );
  INV_X1 U5957 ( .A(DATAI_3_), .ZN(n4917) );
  OAI222_X1 U5958 ( .A1(n4884), .A2(n7183), .B1(n4865), .B2(n4886), .C1(n4887), 
        .C2(n4917), .ZN(U2942) );
  INV_X1 U5959 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4867) );
  INV_X1 U5960 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4866) );
  INV_X1 U5961 ( .A(DATAI_4_), .ZN(n4931) );
  OAI222_X1 U5962 ( .A1(n4884), .A2(n4867), .B1(n4866), .B2(n4886), .C1(n4887), 
        .C2(n4931), .ZN(U2943) );
  INV_X1 U5963 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4868) );
  OAI222_X1 U5964 ( .A1(n4884), .A2(n7271), .B1(n4868), .B2(n4886), .C1(n4887), 
        .C2(n4905), .ZN(U2939) );
  INV_X1 U5965 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4869) );
  INV_X1 U5966 ( .A(DATAI_6_), .ZN(n4910) );
  OAI222_X1 U5967 ( .A1(n4884), .A2(n6411), .B1(n4869), .B2(n4886), .C1(n4887), 
        .C2(n4910), .ZN(U2945) );
  INV_X1 U5968 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4870) );
  INV_X1 U5969 ( .A(DATAI_7_), .ZN(n5258) );
  OAI222_X1 U5970 ( .A1(n4884), .A2(n4871), .B1(n4870), .B2(n4886), .C1(n4887), 
        .C2(n5258), .ZN(U2946) );
  INV_X1 U5971 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4873) );
  INV_X1 U5972 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4872) );
  INV_X1 U5973 ( .A(DATAI_5_), .ZN(n4993) );
  OAI222_X1 U5974 ( .A1(n4884), .A2(n4873), .B1(n4872), .B2(n4886), .C1(n4887), 
        .C2(n4993), .ZN(U2944) );
  OAI222_X1 U5975 ( .A1(n5454), .A2(n6156), .B1(n5577), .B2(n4917), .C1(n7183), 
        .C2(n6394), .ZN(U2888) );
  INV_X1 U5976 ( .A(n4874), .ZN(n4876) );
  AOI21_X1 U5977 ( .B1(n4876), .B2(n4875), .A(n4839), .ZN(n6462) );
  INV_X1 U5978 ( .A(n6462), .ZN(n4945) );
  OR2_X1 U5979 ( .A1(n4878), .A2(n4877), .ZN(n4880) );
  NAND2_X1 U5980 ( .A1(n4880), .A2(n4879), .ZN(n6552) );
  INV_X1 U5981 ( .A(n6552), .ZN(n4881) );
  AOI22_X1 U5982 ( .A1(n4881), .A2(n4474), .B1(n5802), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4882) );
  OAI21_X1 U5983 ( .B1(n4945), .B2(n6152), .A(n4882), .ZN(U2857) );
  INV_X1 U5984 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4883) );
  OAI222_X1 U5985 ( .A1(n4910), .A2(n4887), .B1(n4883), .B2(n4886), .C1(n4884), 
        .C2(n4106), .ZN(U2930) );
  INV_X1 U5986 ( .A(DATAI_15_), .ZN(n4888) );
  INV_X1 U5987 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n7217) );
  INV_X1 U5988 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4885) );
  OAI222_X1 U5989 ( .A1(n4888), .A2(n4887), .B1(n4886), .B2(n7217), .C1(n4885), 
        .C2(n4884), .ZN(U2954) );
  NAND2_X1 U5990 ( .A1(n6461), .A2(DATAI_21_), .ZN(n6788) );
  AOI21_X1 U5991 ( .B1(n4976), .B2(n6073), .A(n6470), .ZN(n4895) );
  AND2_X1 U5992 ( .A1(n6753), .A2(n6213), .ZN(n5418) );
  AND2_X1 U5993 ( .A1(n4893), .A2(n6833), .ZN(n5269) );
  NOR2_X1 U5994 ( .A1(n4755), .A2(n6074), .ZN(n5478) );
  INV_X1 U5995 ( .A(n4933), .ZN(n4894) );
  AOI21_X1 U5996 ( .B1(n5269), .B2(n5478), .A(n4894), .ZN(n4898) );
  OAI21_X1 U5997 ( .B1(n4895), .B2(n5418), .A(n4898), .ZN(n4896) );
  INV_X1 U5998 ( .A(n6862), .ZN(n6985) );
  OAI21_X1 U5999 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n7315), .A(n5054), 
        .ZN(n6586) );
  INV_X1 U6000 ( .A(n6586), .ZN(n6749) );
  OAI211_X1 U6001 ( .C1(n6753), .C2(n4899), .A(n4896), .B(n6749), .ZN(n4928)
         );
  NAND2_X1 U6002 ( .A1(n4928), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4903)
         );
  NAND2_X1 U6003 ( .A1(n6461), .A2(DATAI_29_), .ZN(n6783) );
  INV_X1 U6004 ( .A(n6783), .ZN(n6645) );
  NAND2_X1 U6005 ( .A1(n4930), .A2(n3522), .ZN(n6782) );
  INV_X1 U6006 ( .A(n4898), .ZN(n4900) );
  AOI22_X1 U6007 ( .A1(n4900), .A2(n6753), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4899), .ZN(n4932) );
  NOR2_X2 U6008 ( .A1(n4993), .A2(n5151), .ZN(n6785) );
  INV_X1 U6009 ( .A(n6785), .ZN(n5343) );
  OAI22_X1 U6010 ( .A1(n6782), .A2(n4933), .B1(n4932), .B2(n5343), .ZN(n4901)
         );
  AOI21_X1 U6011 ( .B1(n6645), .B2(n5477), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6012 ( .C1(n5246), .C2(n6788), .A(n4903), .B(n4902), .ZN(U3145)
         );
  NAND2_X1 U6013 ( .A1(n6461), .A2(DATAI_16_), .ZN(n6760) );
  NAND2_X1 U6014 ( .A1(n4928), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4908)
         );
  NAND2_X1 U6015 ( .A1(n6461), .A2(DATAI_24_), .ZN(n6742) );
  INV_X1 U6016 ( .A(n6742), .ZN(n6627) );
  NAND2_X1 U6017 ( .A1(n4930), .A2(n4904), .ZN(n6741) );
  NOR2_X2 U6018 ( .A1(n4905), .A2(n5151), .ZN(n6757) );
  INV_X1 U6019 ( .A(n6757), .ZN(n5323) );
  OAI22_X1 U6020 ( .A1(n6741), .A2(n4933), .B1(n4932), .B2(n5323), .ZN(n4906)
         );
  AOI21_X1 U6021 ( .B1(n6627), .B2(n5477), .A(n4906), .ZN(n4907) );
  OAI211_X1 U6022 ( .C1(n5246), .C2(n6760), .A(n4908), .B(n4907), .ZN(U3140)
         );
  NAND2_X1 U6023 ( .A1(n6461), .A2(DATAI_22_), .ZN(n6790) );
  NAND2_X1 U6024 ( .A1(n4928), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4913)
         );
  NAND2_X1 U6025 ( .A1(n6461), .A2(DATAI_30_), .ZN(n6804) );
  INV_X1 U6026 ( .A(n6804), .ZN(n5522) );
  NAND2_X1 U6027 ( .A1(n4930), .A2(n4909), .ZN(n6789) );
  NOR2_X2 U6028 ( .A1(n4910), .A2(n5151), .ZN(n6799) );
  INV_X1 U6029 ( .A(n6799), .ZN(n5350) );
  OAI22_X1 U6030 ( .A1(n6789), .A2(n4933), .B1(n4932), .B2(n5350), .ZN(n4911)
         );
  AOI21_X1 U6031 ( .B1(n5522), .B2(n5477), .A(n4911), .ZN(n4912) );
  OAI211_X1 U6032 ( .C1(n5246), .C2(n6790), .A(n4913), .B(n4912), .ZN(U3146)
         );
  NAND2_X1 U6033 ( .A1(n6461), .A2(DATAI_23_), .ZN(n6795) );
  NAND2_X1 U6034 ( .A1(n4928), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4916)
         );
  NAND2_X1 U6035 ( .A1(n6461), .A2(DATAI_31_), .ZN(n6814) );
  INV_X1 U6036 ( .A(n6814), .ZN(n5505) );
  NAND2_X1 U6037 ( .A1(n4930), .A2(n3499), .ZN(n6794) );
  NOR2_X2 U6038 ( .A1(n5258), .A2(n5151), .ZN(n6806) );
  INV_X1 U6039 ( .A(n6806), .ZN(n5319) );
  OAI22_X1 U6040 ( .A1(n6794), .A2(n4933), .B1(n4932), .B2(n5319), .ZN(n4914)
         );
  AOI21_X1 U6041 ( .B1(n5505), .B2(n5477), .A(n4914), .ZN(n4915) );
  OAI211_X1 U6042 ( .C1(n5246), .C2(n6795), .A(n4916), .B(n4915), .ZN(U3147)
         );
  NAND2_X1 U6043 ( .A1(n6461), .A2(DATAI_19_), .ZN(n6781) );
  NAND2_X1 U6044 ( .A1(n4928), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4920)
         );
  NAND2_X1 U6045 ( .A1(n6461), .A2(DATAI_27_), .ZN(n6776) );
  INV_X1 U6046 ( .A(n6776), .ZN(n6636) );
  NAND2_X1 U6047 ( .A1(n4930), .A2(n3514), .ZN(n6775) );
  NOR2_X2 U6048 ( .A1(n4917), .A2(n5151), .ZN(n6778) );
  INV_X1 U6049 ( .A(n6778), .ZN(n5335) );
  OAI22_X1 U6050 ( .A1(n6775), .A2(n4933), .B1(n4932), .B2(n5335), .ZN(n4918)
         );
  AOI21_X1 U6051 ( .B1(n6636), .B2(n5477), .A(n4918), .ZN(n4919) );
  OAI211_X1 U6052 ( .C1(n5246), .C2(n6781), .A(n4920), .B(n4919), .ZN(U3143)
         );
  NAND2_X1 U6053 ( .A1(n6461), .A2(DATAI_17_), .ZN(n6767) );
  NAND2_X1 U6054 ( .A1(n4928), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4924)
         );
  NAND2_X1 U6055 ( .A1(n6461), .A2(DATAI_25_), .ZN(n6762) );
  INV_X1 U6056 ( .A(n6762), .ZN(n6630) );
  NAND2_X1 U6057 ( .A1(n4930), .A2(n3201), .ZN(n6761) );
  NOR2_X2 U6058 ( .A1(n4921), .A2(n5151), .ZN(n6764) );
  INV_X1 U6059 ( .A(n6764), .ZN(n5327) );
  OAI22_X1 U6060 ( .A1(n6761), .A2(n4933), .B1(n4932), .B2(n5327), .ZN(n4922)
         );
  AOI21_X1 U6061 ( .B1(n6630), .B2(n5477), .A(n4922), .ZN(n4923) );
  OAI211_X1 U6062 ( .C1(n5246), .C2(n6767), .A(n4924), .B(n4923), .ZN(U3141)
         );
  NAND2_X1 U6063 ( .A1(n6461), .A2(DATAI_18_), .ZN(n6774) );
  NAND2_X1 U6064 ( .A1(n4928), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4927)
         );
  NAND2_X1 U6065 ( .A1(n6461), .A2(DATAI_26_), .ZN(n6769) );
  INV_X1 U6066 ( .A(n6769), .ZN(n6633) );
  NAND2_X1 U6067 ( .A1(n4930), .A2(n4804), .ZN(n6768) );
  NOR2_X2 U6068 ( .A1(n4944), .A2(n5151), .ZN(n6771) );
  INV_X1 U6069 ( .A(n6771), .ZN(n5331) );
  OAI22_X1 U6070 ( .A1(n6768), .A2(n4933), .B1(n4932), .B2(n5331), .ZN(n4925)
         );
  AOI21_X1 U6071 ( .B1(n6633), .B2(n5477), .A(n4925), .ZN(n4926) );
  OAI211_X1 U6072 ( .C1(n5246), .C2(n6774), .A(n4927), .B(n4926), .ZN(U3142)
         );
  NAND2_X1 U6073 ( .A1(n6461), .A2(DATAI_20_), .ZN(n7369) );
  NAND2_X1 U6074 ( .A1(n4928), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4936)
         );
  NAND2_X1 U6075 ( .A1(n6461), .A2(DATAI_28_), .ZN(n7378) );
  INV_X1 U6076 ( .A(n7378), .ZN(n6639) );
  NAND2_X1 U6077 ( .A1(n4930), .A2(n4929), .ZN(n7368) );
  NOR2_X2 U6078 ( .A1(n4931), .A2(n5151), .ZN(n7373) );
  INV_X1 U6079 ( .A(n7373), .ZN(n5339) );
  OAI22_X1 U6080 ( .A1(n7368), .A2(n4933), .B1(n4932), .B2(n5339), .ZN(n4934)
         );
  AOI21_X1 U6081 ( .B1(n6639), .B2(n5477), .A(n4934), .ZN(n4935) );
  OAI211_X1 U6082 ( .C1(n5246), .C2(n7369), .A(n4936), .B(n4935), .ZN(U3144)
         );
  OAI21_X1 U6083 ( .B1(n4937), .B2(n4939), .A(n4938), .ZN(n4940) );
  INV_X1 U6084 ( .A(n4940), .ZN(n6545) );
  NAND2_X1 U6085 ( .A1(n6545), .A2(n6460), .ZN(n4943) );
  AND2_X1 U6086 ( .A1(n6567), .A2(REIP_REG_3__SCAN_IN), .ZN(n6543) );
  NOR2_X1 U6087 ( .A1(n6466), .A2(n5450), .ZN(n4941) );
  AOI211_X1 U6088 ( .C1(n6456), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6543), 
        .B(n4941), .ZN(n4942) );
  OAI211_X1 U6089 ( .C1(n6470), .C2(n5454), .A(n4943), .B(n4942), .ZN(U2983)
         );
  OAI222_X1 U6090 ( .A1(n4945), .A2(n6156), .B1(n5577), .B2(n4944), .C1(n6394), 
        .C2(n4861), .ZN(U2889) );
  NAND2_X1 U6091 ( .A1(n4965), .A2(n3304), .ZN(n4946) );
  OAI21_X1 U6092 ( .B1(n4947), .B2(n4965), .A(n4946), .ZN(n6842) );
  NAND2_X1 U6093 ( .A1(n4893), .A2(n6832), .ZN(n4964) );
  NOR2_X1 U6094 ( .A1(n4950), .A2(n4955), .ZN(n4948) );
  XNOR2_X1 U6095 ( .A(n4948), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4961)
         );
  AOI21_X1 U6096 ( .B1(n4950), .B2(n4955), .A(n4949), .ZN(n4951) );
  NOR2_X1 U6097 ( .A1(n3635), .A2(n4951), .ZN(n6948) );
  NAND3_X1 U6098 ( .A1(n4953), .A2(n4955), .A3(n4954), .ZN(n4956) );
  OAI21_X1 U6099 ( .B1(n4952), .B2(n4949), .A(n4956), .ZN(n4957) );
  NAND2_X1 U6100 ( .A1(n6834), .A2(n4957), .ZN(n4958) );
  OAI21_X1 U6101 ( .B1(n6948), .B2(n4959), .A(n4958), .ZN(n4960) );
  AOI21_X1 U6102 ( .B1(n4962), .B2(n4961), .A(n4960), .ZN(n4963) );
  NAND2_X1 U6103 ( .A1(n4964), .A2(n4963), .ZN(n6947) );
  NAND2_X1 U6104 ( .A1(n6947), .A2(n6835), .ZN(n4967) );
  NAND2_X1 U6105 ( .A1(n4965), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U6106 ( .A1(n4967), .A2(n4966), .ZN(n6849) );
  NAND2_X1 U6107 ( .A1(n6849), .A2(n6952), .ZN(n4968) );
  NAND2_X1 U6108 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6217), .ZN(n4971) );
  OAI22_X1 U6109 ( .A1(n6842), .A2(n4968), .B1(n4971), .B2(n4953), .ZN(n6829)
         );
  AND2_X1 U6110 ( .A1(n6829), .A2(n4969), .ZN(n4986) );
  NAND3_X1 U6111 ( .A1(n6324), .A2(n4970), .A3(n6952), .ZN(n4974) );
  OAI21_X1 U6112 ( .B1(n6835), .B2(STATE2_REG_1__SCAN_IN), .A(n4971), .ZN(
        n4972) );
  NAND2_X1 U6113 ( .A1(n4972), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6114 ( .A1(n4974), .A2(n4973), .ZN(n6816) );
  NOR3_X1 U6115 ( .A1(n4986), .A2(n6816), .A3(FLUSH_REG_SCAN_IN), .ZN(n4975)
         );
  OAI21_X1 U6116 ( .B1(n4975), .B2(n6944), .A(n5151), .ZN(n6577) );
  INV_X1 U6117 ( .A(n5104), .ZN(n4977) );
  NAND2_X1 U6118 ( .A1(n4977), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6119 ( .A1(n5098), .A2(n5268), .ZN(n6583) );
  INV_X1 U6120 ( .A(n6583), .ZN(n4980) );
  NAND2_X1 U6121 ( .A1(n6650), .A2(n6744), .ZN(n6652) );
  AOI21_X1 U6122 ( .B1(n4980), .B2(n6652), .A(n6658), .ZN(n4982) );
  INV_X1 U6123 ( .A(n5418), .ZN(n5131) );
  INV_X1 U6124 ( .A(n4893), .ZN(n6702) );
  NOR2_X1 U6125 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6952), .ZN(n6077) );
  OAI22_X1 U6126 ( .A1(n4978), .A2(n5131), .B1(n6702), .B2(n6077), .ZN(n4981)
         );
  OAI21_X1 U6127 ( .B1(n4982), .B2(n4981), .A(n6577), .ZN(n4983) );
  OAI21_X1 U6128 ( .B1(n6577), .B2(n6850), .A(n4983), .ZN(U3462) );
  INV_X1 U6129 ( .A(n4984), .ZN(n4985) );
  NOR3_X1 U6130 ( .A1(n4986), .A2(n6816), .A3(n4985), .ZN(n6860) );
  INV_X1 U6131 ( .A(n6833), .ZN(n6653) );
  OAI22_X1 U6132 ( .A1(n4891), .A2(n6658), .B1(n6653), .B2(n6077), .ZN(n4987)
         );
  OAI21_X1 U6133 ( .B1(n6860), .B2(n4987), .A(n6577), .ZN(n4988) );
  OAI21_X1 U6134 ( .B1(n6577), .B2(n5388), .A(n4988), .ZN(U3465) );
  OR2_X1 U6135 ( .A1(n4991), .A2(n4990), .ZN(n4992) );
  NAND2_X1 U6136 ( .A1(n4989), .A2(n4992), .ZN(n5305) );
  OAI222_X1 U6137 ( .A1(n5305), .A2(n6156), .B1(n5577), .B2(n4993), .C1(n6394), 
        .C2(n4873), .ZN(U2886) );
  NAND2_X1 U6138 ( .A1(n4995), .A2(n4994), .ZN(n4998) );
  INV_X1 U6139 ( .A(n4996), .ZN(n4997) );
  NAND2_X1 U6140 ( .A1(n4998), .A2(n4997), .ZN(n6522) );
  INV_X1 U6141 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4999) );
  OAI222_X1 U6142 ( .A1(n6522), .A2(n6371), .B1(n6380), .B2(n4999), .C1(n5305), 
        .C2(n6152), .ZN(U2854) );
  XOR2_X1 U6143 ( .A(n4840), .B(n5000), .Z(n6452) );
  INV_X1 U6144 ( .A(n6452), .ZN(n5002) );
  AOI22_X1 U6145 ( .A1(n6390), .A2(DATAI_4_), .B1(n6386), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n5001) );
  OAI21_X1 U6146 ( .B1(n5002), .B2(n6156), .A(n5001), .ZN(U2887) );
  NAND2_X1 U6147 ( .A1(n5310), .A2(n6850), .ZN(n6589) );
  NOR2_X1 U6148 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6589), .ZN(n5041)
         );
  NOR2_X1 U6149 ( .A1(n6580), .A2(n6073), .ZN(n5003) );
  INV_X1 U6150 ( .A(n5416), .ZN(n5004) );
  NOR2_X1 U6151 ( .A1(n6580), .A2(n5004), .ZN(n5005) );
  INV_X1 U6152 ( .A(n6613), .ZN(n5006) );
  OAI21_X1 U6153 ( .B1(n5136), .B2(n5006), .A(n5131), .ZN(n5007) );
  AND2_X1 U6154 ( .A1(n4755), .A2(n6350), .ZN(n5307) );
  NAND2_X1 U6155 ( .A1(n6702), .A2(n5307), .ZN(n6584) );
  NAND2_X1 U6156 ( .A1(n5007), .A2(n6584), .ZN(n5008) );
  NOR2_X1 U6157 ( .A1(n5010), .A2(n3658), .ZN(n6703) );
  OAI21_X1 U6158 ( .B1(n5484), .B2(n3658), .A(n5054), .ZN(n5480) );
  NOR2_X1 U6159 ( .A1(n6703), .A2(n5480), .ZN(n5314) );
  OAI221_X1 U6160 ( .B1(n5041), .B2(n7315), .C1(n5041), .C2(n5008), .A(n5314), 
        .ZN(n5009) );
  AND2_X1 U6161 ( .A1(n5010), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6694) );
  NAND3_X1 U6162 ( .A1(n6694), .A2(n5484), .A3(n6850), .ZN(n5011) );
  OAI21_X1 U6163 ( .B1(n6584), .B2(n6658), .A(n5011), .ZN(n5040) );
  AOI22_X1 U6164 ( .A1(n6723), .A2(n5041), .B1(n7373), .B2(n5040), .ZN(n5012)
         );
  OAI21_X1 U6165 ( .B1(n7369), .B2(n6613), .A(n5012), .ZN(n5013) );
  AOI21_X1 U6166 ( .B1(n6639), .B2(n5136), .A(n5013), .ZN(n5014) );
  OAI21_X1 U6167 ( .B1(n5046), .B2(n5015), .A(n5014), .ZN(U3040) );
  AOI22_X1 U6168 ( .A1(n6715), .A2(n5041), .B1(n6771), .B2(n5040), .ZN(n5016)
         );
  OAI21_X1 U6169 ( .B1(n6774), .B2(n6613), .A(n5016), .ZN(n5017) );
  AOI21_X1 U6170 ( .B1(n6633), .B2(n5136), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6171 ( .B1(n5046), .B2(n5019), .A(n5018), .ZN(U3038) );
  AOI22_X1 U6172 ( .A1(n6711), .A2(n5041), .B1(n6764), .B2(n5040), .ZN(n5020)
         );
  OAI21_X1 U6173 ( .B1(n6767), .B2(n6613), .A(n5020), .ZN(n5021) );
  AOI21_X1 U6174 ( .B1(n6630), .B2(n5136), .A(n5021), .ZN(n5022) );
  OAI21_X1 U6175 ( .B1(n5046), .B2(n5023), .A(n5022), .ZN(U3037) );
  AOI22_X1 U6176 ( .A1(n6800), .A2(n5041), .B1(n6799), .B2(n5040), .ZN(n5024)
         );
  OAI21_X1 U6177 ( .B1(n6790), .B2(n6613), .A(n5024), .ZN(n5025) );
  AOI21_X1 U6178 ( .B1(n5522), .B2(n5136), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6179 ( .B1(n5046), .B2(n5027), .A(n5026), .ZN(U3042) );
  AOI22_X1 U6180 ( .A1(n6727), .A2(n5041), .B1(n6785), .B2(n5040), .ZN(n5028)
         );
  OAI21_X1 U6181 ( .B1(n6788), .B2(n6613), .A(n5028), .ZN(n5029) );
  AOI21_X1 U6182 ( .B1(n6645), .B2(n5136), .A(n5029), .ZN(n5030) );
  OAI21_X1 U6183 ( .B1(n5046), .B2(n5031), .A(n5030), .ZN(U3041) );
  AOI22_X1 U6184 ( .A1(n6698), .A2(n5041), .B1(n6757), .B2(n5040), .ZN(n5032)
         );
  OAI21_X1 U6185 ( .B1(n6760), .B2(n6613), .A(n5032), .ZN(n5033) );
  AOI21_X1 U6186 ( .B1(n6627), .B2(n5136), .A(n5033), .ZN(n5034) );
  OAI21_X1 U6187 ( .B1(n5046), .B2(n5035), .A(n5034), .ZN(U3036) );
  AOI22_X1 U6188 ( .A1(n6808), .A2(n5041), .B1(n6806), .B2(n5040), .ZN(n5036)
         );
  OAI21_X1 U6189 ( .B1(n6795), .B2(n6613), .A(n5036), .ZN(n5037) );
  AOI21_X1 U6190 ( .B1(n5505), .B2(n5136), .A(n5037), .ZN(n5038) );
  OAI21_X1 U6191 ( .B1(n5046), .B2(n5039), .A(n5038), .ZN(U3043) );
  AOI22_X1 U6192 ( .A1(n6719), .A2(n5041), .B1(n6778), .B2(n5040), .ZN(n5042)
         );
  OAI21_X1 U6193 ( .B1(n6781), .B2(n6613), .A(n5042), .ZN(n5043) );
  AOI21_X1 U6194 ( .B1(n6636), .B2(n5136), .A(n5043), .ZN(n5044) );
  OAI21_X1 U6195 ( .B1(n5046), .B2(n5045), .A(n5044), .ZN(U3039) );
  INV_X1 U6196 ( .A(n6649), .ZN(n5048) );
  NOR2_X1 U6197 ( .A1(n6580), .A2(n5048), .ZN(n5049) );
  INV_X1 U6198 ( .A(n6625), .ZN(n5050) );
  NOR3_X1 U6199 ( .A1(n6621), .A2(n5050), .A3(n6658), .ZN(n5051) );
  NOR2_X1 U6200 ( .A1(n5051), .A2(n5418), .ZN(n5057) );
  NAND2_X1 U6201 ( .A1(n5052), .A2(n6074), .ZN(n5147) );
  NOR2_X1 U6202 ( .A1(n5147), .A2(n6654), .ZN(n5389) );
  NAND3_X1 U6203 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6850), .A3(n6838), .ZN(n5393) );
  NOR2_X1 U6204 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5393), .ZN(n6620)
         );
  INV_X1 U6205 ( .A(n6620), .ZN(n5055) );
  INV_X1 U6206 ( .A(n5150), .ZN(n5053) );
  OR2_X1 U6207 ( .A1(n5484), .A2(n5053), .ZN(n5214) );
  INV_X1 U6208 ( .A(n5214), .ZN(n5058) );
  OAI21_X1 U6209 ( .B1(n5058), .B2(n3658), .A(n5054), .ZN(n5210) );
  AOI211_X1 U6210 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5055), .A(n6694), .B(
        n5210), .ZN(n5056) );
  OAI21_X1 U6211 ( .B1(n5057), .B2(n5389), .A(n5056), .ZN(n6622) );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5063) );
  INV_X1 U6213 ( .A(n6760), .ZN(n6708) );
  OR2_X1 U6214 ( .A1(n5147), .A2(n6658), .ZN(n5157) );
  NAND2_X1 U6215 ( .A1(n5058), .A2(n6703), .ZN(n5059) );
  OAI21_X1 U6216 ( .B1(n5157), .B2(n4893), .A(n5059), .ZN(n6619) );
  AOI22_X1 U6217 ( .A1(n6698), .A2(n6620), .B1(n6757), .B2(n6619), .ZN(n5060)
         );
  OAI21_X1 U6218 ( .B1(n6742), .B2(n6625), .A(n5060), .ZN(n5061) );
  AOI21_X1 U6219 ( .B1(n6708), .B2(n6621), .A(n5061), .ZN(n5062) );
  OAI21_X1 U6220 ( .B1(n5088), .B2(n5063), .A(n5062), .ZN(U3052) );
  INV_X1 U6221 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5067) );
  INV_X1 U6222 ( .A(n6795), .ZN(n6810) );
  AOI22_X1 U6223 ( .A1(n6808), .A2(n6620), .B1(n6806), .B2(n6619), .ZN(n5064)
         );
  OAI21_X1 U6224 ( .B1(n6814), .B2(n6625), .A(n5064), .ZN(n5065) );
  AOI21_X1 U6225 ( .B1(n6810), .B2(n6621), .A(n5065), .ZN(n5066) );
  OAI21_X1 U6226 ( .B1(n5088), .B2(n5067), .A(n5066), .ZN(U3059) );
  INV_X1 U6227 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5071) );
  INV_X1 U6228 ( .A(n6774), .ZN(n6716) );
  AOI22_X1 U6229 ( .A1(n6715), .A2(n6620), .B1(n6771), .B2(n6619), .ZN(n5068)
         );
  OAI21_X1 U6230 ( .B1(n6769), .B2(n6625), .A(n5068), .ZN(n5069) );
  AOI21_X1 U6231 ( .B1(n6716), .B2(n6621), .A(n5069), .ZN(n5070) );
  OAI21_X1 U6232 ( .B1(n5088), .B2(n5071), .A(n5070), .ZN(U3054) );
  INV_X1 U6233 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5075) );
  INV_X1 U6234 ( .A(n6788), .ZN(n6728) );
  AOI22_X1 U6235 ( .A1(n6727), .A2(n6620), .B1(n6785), .B2(n6619), .ZN(n5072)
         );
  OAI21_X1 U6236 ( .B1(n6783), .B2(n6625), .A(n5072), .ZN(n5073) );
  AOI21_X1 U6237 ( .B1(n6728), .B2(n6621), .A(n5073), .ZN(n5074) );
  OAI21_X1 U6238 ( .B1(n5088), .B2(n5075), .A(n5074), .ZN(U3057) );
  INV_X1 U6239 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5079) );
  INV_X1 U6240 ( .A(n6767), .ZN(n6712) );
  AOI22_X1 U6241 ( .A1(n6711), .A2(n6620), .B1(n6764), .B2(n6619), .ZN(n5076)
         );
  OAI21_X1 U6242 ( .B1(n6762), .B2(n6625), .A(n5076), .ZN(n5077) );
  AOI21_X1 U6243 ( .B1(n6712), .B2(n6621), .A(n5077), .ZN(n5078) );
  OAI21_X1 U6244 ( .B1(n5088), .B2(n5079), .A(n5078), .ZN(U3053) );
  INV_X1 U6245 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5083) );
  INV_X1 U6246 ( .A(n6781), .ZN(n6720) );
  AOI22_X1 U6247 ( .A1(n6719), .A2(n6620), .B1(n6778), .B2(n6619), .ZN(n5080)
         );
  OAI21_X1 U6248 ( .B1(n6776), .B2(n6625), .A(n5080), .ZN(n5081) );
  AOI21_X1 U6249 ( .B1(n6720), .B2(n6621), .A(n5081), .ZN(n5082) );
  OAI21_X1 U6250 ( .B1(n5088), .B2(n5083), .A(n5082), .ZN(U3055) );
  INV_X1 U6251 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5087) );
  INV_X1 U6252 ( .A(n7369), .ZN(n6724) );
  AOI22_X1 U6253 ( .A1(n6723), .A2(n6620), .B1(n7373), .B2(n6619), .ZN(n5084)
         );
  OAI21_X1 U6254 ( .B1(n7378), .B2(n6625), .A(n5084), .ZN(n5085) );
  AOI21_X1 U6255 ( .B1(n6724), .B2(n6621), .A(n5085), .ZN(n5086) );
  OAI21_X1 U6256 ( .B1(n5088), .B2(n5087), .A(n5086), .ZN(U3056) );
  OAI21_X1 U6257 ( .B1(n5091), .B2(n5090), .A(n5089), .ZN(n6526) );
  NAND2_X1 U6258 ( .A1(n6567), .A2(REIP_REG_5__SCAN_IN), .ZN(n6523) );
  OAI21_X1 U6259 ( .B1(n6474), .B2(n5092), .A(n6523), .ZN(n5094) );
  NOR2_X1 U6260 ( .A1(n5305), .A2(n6470), .ZN(n5093) );
  AOI211_X1 U6261 ( .C1(n6438), .C2(n5303), .A(n5094), .B(n5093), .ZN(n5095)
         );
  OAI21_X1 U6262 ( .B1(n6468), .B2(n6526), .A(n5095), .ZN(U2981) );
  XOR2_X1 U6263 ( .A(n4989), .B(n5096), .Z(n6444) );
  INV_X1 U6264 ( .A(n6444), .ZN(n5097) );
  OAI222_X1 U6265 ( .A1(n5577), .A2(n4910), .B1(n6156), .B2(n5097), .C1(n6411), 
        .C2(n6394), .ZN(U2885) );
  NAND2_X1 U6266 ( .A1(n6753), .A2(n5098), .ZN(n5102) );
  INV_X1 U6267 ( .A(n5147), .ZN(n5099) );
  NAND3_X1 U6268 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6838), .ZN(n5152) );
  NOR2_X1 U6269 ( .A1(n5388), .A2(n5152), .ZN(n5121) );
  AOI21_X1 U6270 ( .B1(n5099), .B2(n5269), .A(n5121), .ZN(n5103) );
  INV_X1 U6271 ( .A(n5103), .ZN(n5101) );
  AOI21_X1 U6272 ( .B1(n6658), .B2(n5152), .A(n6586), .ZN(n5100) );
  OAI21_X1 U6273 ( .B1(n5102), .B2(n5101), .A(n5100), .ZN(n5120) );
  OAI22_X1 U6274 ( .A1(n5103), .A2(n5102), .B1(n3658), .B2(n5152), .ZN(n5119)
         );
  AOI22_X1 U6275 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5120), .B1(n6778), 
        .B2(n5119), .ZN(n5106) );
  AOI22_X1 U6276 ( .A1(n6809), .A2(n6636), .B1(n6719), .B2(n5121), .ZN(n5105)
         );
  OAI211_X1 U6277 ( .C1(n6781), .C2(n5124), .A(n5106), .B(n5105), .ZN(U3127)
         );
  AOI22_X1 U6278 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5120), .B1(n6757), 
        .B2(n5119), .ZN(n5108) );
  AOI22_X1 U6279 ( .A1(n6809), .A2(n6627), .B1(n6698), .B2(n5121), .ZN(n5107)
         );
  OAI211_X1 U6280 ( .C1(n6760), .C2(n5124), .A(n5108), .B(n5107), .ZN(U3124)
         );
  AOI22_X1 U6281 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5120), .B1(n6764), 
        .B2(n5119), .ZN(n5110) );
  AOI22_X1 U6282 ( .A1(n6809), .A2(n6630), .B1(n6711), .B2(n5121), .ZN(n5109)
         );
  OAI211_X1 U6283 ( .C1(n6767), .C2(n5124), .A(n5110), .B(n5109), .ZN(U3125)
         );
  AOI22_X1 U6284 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5120), .B1(n6771), 
        .B2(n5119), .ZN(n5112) );
  AOI22_X1 U6285 ( .A1(n6809), .A2(n6633), .B1(n6715), .B2(n5121), .ZN(n5111)
         );
  OAI211_X1 U6286 ( .C1(n6774), .C2(n5124), .A(n5112), .B(n5111), .ZN(U3126)
         );
  AOI22_X1 U6287 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5120), .B1(n6806), 
        .B2(n5119), .ZN(n5114) );
  AOI22_X1 U6288 ( .A1(n6809), .A2(n5505), .B1(n6808), .B2(n5121), .ZN(n5113)
         );
  OAI211_X1 U6289 ( .C1(n6795), .C2(n5124), .A(n5114), .B(n5113), .ZN(U3131)
         );
  AOI22_X1 U6290 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5120), .B1(n7373), 
        .B2(n5119), .ZN(n5116) );
  AOI22_X1 U6291 ( .A1(n6809), .A2(n6639), .B1(n6723), .B2(n5121), .ZN(n5115)
         );
  OAI211_X1 U6292 ( .C1(n7369), .C2(n5124), .A(n5116), .B(n5115), .ZN(U3128)
         );
  AOI22_X1 U6293 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5120), .B1(n6799), 
        .B2(n5119), .ZN(n5118) );
  AOI22_X1 U6294 ( .A1(n6809), .A2(n5522), .B1(n6800), .B2(n5121), .ZN(n5117)
         );
  OAI211_X1 U6295 ( .C1(n6790), .C2(n5124), .A(n5118), .B(n5117), .ZN(U3130)
         );
  AOI22_X1 U6296 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5120), .B1(n6785), 
        .B2(n5119), .ZN(n5123) );
  AOI22_X1 U6297 ( .A1(n6809), .A2(n6645), .B1(n6727), .B2(n5121), .ZN(n5122)
         );
  OAI211_X1 U6298 ( .C1(n6788), .C2(n5124), .A(n5123), .B(n5122), .ZN(U3129)
         );
  XOR2_X1 U6299 ( .A(n5126), .B(n5125), .Z(n5442) );
  INV_X1 U6300 ( .A(n5442), .ZN(n5259) );
  AOI21_X1 U6301 ( .B1(n5129), .B2(n5128), .A(n5127), .ZN(n6505) );
  AOI22_X1 U6302 ( .A1(n4474), .A2(n6505), .B1(EBX_REG_7__SCAN_IN), .B2(n5802), 
        .ZN(n5130) );
  OAI21_X1 U6303 ( .B1(n5259), .B2(n6152), .A(n5130), .ZN(U2852) );
  OAI21_X1 U6304 ( .B1(n5135), .B2(n6658), .A(n5131), .ZN(n5138) );
  NAND2_X1 U6305 ( .A1(n4755), .A2(n6074), .ZN(n6701) );
  INV_X1 U6306 ( .A(n6701), .ZN(n6692) );
  NAND2_X1 U6307 ( .A1(n6702), .A2(n6692), .ZN(n5215) );
  OR2_X1 U6308 ( .A1(n5215), .A2(n6653), .ZN(n5133) );
  NAND3_X1 U6309 ( .A1(n6850), .A2(n6844), .A3(n6838), .ZN(n5209) );
  NOR2_X1 U6310 ( .A1(n5388), .A2(n5209), .ZN(n5201) );
  INV_X1 U6311 ( .A(n5201), .ZN(n5132) );
  NAND2_X1 U6312 ( .A1(n5133), .A2(n5132), .ZN(n5137) );
  INV_X1 U6313 ( .A(n5209), .ZN(n5134) );
  AOI22_X1 U6314 ( .A1(n5138), .A2(n5137), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5134), .ZN(n5206) );
  INV_X1 U6315 ( .A(n5137), .ZN(n5139) );
  AOI22_X1 U6316 ( .A1(n5139), .A2(n5138), .B1(n5209), .B2(n6658), .ZN(n5140)
         );
  NAND2_X1 U6317 ( .A1(n6749), .A2(n5140), .ZN(n5200) );
  AOI22_X1 U6318 ( .A1(n6808), .A2(n5201), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5200), .ZN(n5141) );
  OAI21_X1 U6319 ( .B1(n5203), .B2(n6795), .A(n5141), .ZN(n5142) );
  AOI21_X1 U6320 ( .B1(n5505), .B2(n5248), .A(n5142), .ZN(n5143) );
  OAI21_X1 U6321 ( .B1(n5206), .B2(n5319), .A(n5143), .ZN(U3035) );
  AOI22_X1 U6322 ( .A1(n6800), .A2(n5201), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5200), .ZN(n5144) );
  OAI21_X1 U6323 ( .B1(n5203), .B2(n6790), .A(n5144), .ZN(n5145) );
  AOI21_X1 U6324 ( .B1(n5522), .B2(n5248), .A(n5145), .ZN(n5146) );
  OAI21_X1 U6325 ( .B1(n5206), .B2(n5350), .A(n5146), .ZN(U3034) );
  NOR3_X1 U6326 ( .A1(n5181), .A2(n6809), .A3(n6658), .ZN(n5149) );
  OAI22_X1 U6327 ( .A1(n5149), .A2(n5418), .B1(n5148), .B2(n5147), .ZN(n5155)
         );
  OR2_X1 U6328 ( .A1(n5484), .A2(n5150), .ZN(n6693) );
  AOI21_X1 U6329 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6693), .A(n5151), .ZN(
        n6706) );
  INV_X1 U6330 ( .A(n6694), .ZN(n5308) );
  NOR2_X1 U6331 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5152), .ZN(n6807)
         );
  INV_X1 U6332 ( .A(n6807), .ZN(n5153) );
  NAND2_X1 U6333 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5153), .ZN(n5154) );
  NAND4_X1 U6334 ( .A1(n5155), .A2(n6706), .A3(n5308), .A4(n5154), .ZN(n6811)
         );
  INV_X1 U6335 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5161) );
  INV_X1 U6336 ( .A(n6809), .ZN(n5179) );
  INV_X1 U6337 ( .A(n6703), .ZN(n5156) );
  OAI22_X1 U6338 ( .A1(n5157), .A2(n6702), .B1(n6693), .B2(n5156), .ZN(n6805)
         );
  AOI22_X1 U6339 ( .A1(n6719), .A2(n6807), .B1(n6778), .B2(n6805), .ZN(n5158)
         );
  OAI21_X1 U6340 ( .B1(n5179), .B2(n6781), .A(n5158), .ZN(n5159) );
  AOI21_X1 U6341 ( .B1(n6636), .B2(n5181), .A(n5159), .ZN(n5160) );
  OAI21_X1 U6342 ( .B1(n5184), .B2(n5161), .A(n5160), .ZN(U3119) );
  INV_X1 U6343 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5165) );
  AOI22_X1 U6344 ( .A1(n6727), .A2(n6807), .B1(n6785), .B2(n6805), .ZN(n5162)
         );
  OAI21_X1 U6345 ( .B1(n5179), .B2(n6788), .A(n5162), .ZN(n5163) );
  AOI21_X1 U6346 ( .B1(n6645), .B2(n5181), .A(n5163), .ZN(n5164) );
  OAI21_X1 U6347 ( .B1(n5184), .B2(n5165), .A(n5164), .ZN(U3121) );
  INV_X1 U6348 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5169) );
  AOI22_X1 U6349 ( .A1(n6711), .A2(n6807), .B1(n6764), .B2(n6805), .ZN(n5166)
         );
  OAI21_X1 U6350 ( .B1(n5179), .B2(n6767), .A(n5166), .ZN(n5167) );
  AOI21_X1 U6351 ( .B1(n6630), .B2(n5181), .A(n5167), .ZN(n5168) );
  OAI21_X1 U6352 ( .B1(n5184), .B2(n5169), .A(n5168), .ZN(U3117) );
  INV_X1 U6353 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5173) );
  AOI22_X1 U6354 ( .A1(n6723), .A2(n6807), .B1(n7373), .B2(n6805), .ZN(n5170)
         );
  OAI21_X1 U6355 ( .B1(n5179), .B2(n7369), .A(n5170), .ZN(n5171) );
  AOI21_X1 U6356 ( .B1(n6639), .B2(n5181), .A(n5171), .ZN(n5172) );
  OAI21_X1 U6357 ( .B1(n5184), .B2(n5173), .A(n5172), .ZN(U3120) );
  INV_X1 U6358 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5177) );
  AOI22_X1 U6359 ( .A1(n6698), .A2(n6807), .B1(n6757), .B2(n6805), .ZN(n5174)
         );
  OAI21_X1 U6360 ( .B1(n5179), .B2(n6760), .A(n5174), .ZN(n5175) );
  AOI21_X1 U6361 ( .B1(n6627), .B2(n5181), .A(n5175), .ZN(n5176) );
  OAI21_X1 U6362 ( .B1(n5184), .B2(n5177), .A(n5176), .ZN(U3116) );
  INV_X1 U6363 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5183) );
  AOI22_X1 U6364 ( .A1(n6715), .A2(n6807), .B1(n6771), .B2(n6805), .ZN(n5178)
         );
  OAI21_X1 U6365 ( .B1(n5179), .B2(n6774), .A(n5178), .ZN(n5180) );
  AOI21_X1 U6366 ( .B1(n6633), .B2(n5181), .A(n5180), .ZN(n5182) );
  OAI21_X1 U6367 ( .B1(n5184), .B2(n5183), .A(n5182), .ZN(U3118) );
  AOI22_X1 U6368 ( .A1(n6723), .A2(n5201), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5200), .ZN(n5185) );
  OAI21_X1 U6369 ( .B1(n5203), .B2(n7369), .A(n5185), .ZN(n5186) );
  AOI21_X1 U6370 ( .B1(n6639), .B2(n5248), .A(n5186), .ZN(n5187) );
  OAI21_X1 U6371 ( .B1(n5206), .B2(n5339), .A(n5187), .ZN(U3032) );
  AOI22_X1 U6372 ( .A1(n6727), .A2(n5201), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5200), .ZN(n5188) );
  OAI21_X1 U6373 ( .B1(n5203), .B2(n6788), .A(n5188), .ZN(n5189) );
  AOI21_X1 U6374 ( .B1(n6645), .B2(n5248), .A(n5189), .ZN(n5190) );
  OAI21_X1 U6375 ( .B1(n5206), .B2(n5343), .A(n5190), .ZN(U3033) );
  AOI22_X1 U6376 ( .A1(n6698), .A2(n5201), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5200), .ZN(n5191) );
  OAI21_X1 U6377 ( .B1(n5203), .B2(n6760), .A(n5191), .ZN(n5192) );
  AOI21_X1 U6378 ( .B1(n6627), .B2(n5248), .A(n5192), .ZN(n5193) );
  OAI21_X1 U6379 ( .B1(n5206), .B2(n5323), .A(n5193), .ZN(U3028) );
  AOI22_X1 U6380 ( .A1(n6715), .A2(n5201), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5200), .ZN(n5194) );
  OAI21_X1 U6381 ( .B1(n5203), .B2(n6774), .A(n5194), .ZN(n5195) );
  AOI21_X1 U6382 ( .B1(n6633), .B2(n5248), .A(n5195), .ZN(n5196) );
  OAI21_X1 U6383 ( .B1(n5206), .B2(n5331), .A(n5196), .ZN(U3030) );
  AOI22_X1 U6384 ( .A1(n6719), .A2(n5201), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5200), .ZN(n5197) );
  OAI21_X1 U6385 ( .B1(n5203), .B2(n6781), .A(n5197), .ZN(n5198) );
  AOI21_X1 U6386 ( .B1(n6636), .B2(n5248), .A(n5198), .ZN(n5199) );
  OAI21_X1 U6387 ( .B1(n5206), .B2(n5335), .A(n5199), .ZN(U3031) );
  AOI22_X1 U6388 ( .A1(n6711), .A2(n5201), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5200), .ZN(n5202) );
  OAI21_X1 U6389 ( .B1(n5203), .B2(n6767), .A(n5202), .ZN(n5204) );
  AOI21_X1 U6390 ( .B1(n6630), .B2(n5248), .A(n5204), .ZN(n5205) );
  OAI21_X1 U6391 ( .B1(n5206), .B2(n5327), .A(n5205), .ZN(U3029) );
  OAI21_X1 U6392 ( .B1(n5248), .B2(n5207), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5208) );
  NAND3_X1 U6393 ( .A1(n5208), .A2(n6753), .A3(n5215), .ZN(n5213) );
  NOR2_X1 U6394 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5209), .ZN(n5244)
         );
  INV_X1 U6395 ( .A(n5244), .ZN(n5211) );
  AOI211_X1 U6396 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5211), .A(n6703), .B(
        n5210), .ZN(n5212) );
  OAI22_X1 U6397 ( .A1(n5215), .A2(n6658), .B1(n5308), .B2(n5214), .ZN(n5243)
         );
  AOI22_X1 U6398 ( .A1(n6711), .A2(n5244), .B1(n6764), .B2(n5243), .ZN(n5216)
         );
  OAI21_X1 U6399 ( .B1(n5246), .B2(n6762), .A(n5216), .ZN(n5217) );
  AOI21_X1 U6400 ( .B1(n6712), .B2(n5248), .A(n5217), .ZN(n5218) );
  OAI21_X1 U6401 ( .B1(n5251), .B2(n5219), .A(n5218), .ZN(U3021) );
  AOI22_X1 U6402 ( .A1(n6723), .A2(n5244), .B1(n7373), .B2(n5243), .ZN(n5220)
         );
  OAI21_X1 U6403 ( .B1(n5246), .B2(n7378), .A(n5220), .ZN(n5221) );
  AOI21_X1 U6404 ( .B1(n6724), .B2(n5248), .A(n5221), .ZN(n5222) );
  OAI21_X1 U6405 ( .B1(n5251), .B2(n5223), .A(n5222), .ZN(U3024) );
  AOI22_X1 U6406 ( .A1(n6719), .A2(n5244), .B1(n6778), .B2(n5243), .ZN(n5224)
         );
  OAI21_X1 U6407 ( .B1(n5246), .B2(n6776), .A(n5224), .ZN(n5225) );
  AOI21_X1 U6408 ( .B1(n6720), .B2(n5248), .A(n5225), .ZN(n5226) );
  OAI21_X1 U6409 ( .B1(n5251), .B2(n5227), .A(n5226), .ZN(U3023) );
  AOI22_X1 U6410 ( .A1(n6715), .A2(n5244), .B1(n6771), .B2(n5243), .ZN(n5228)
         );
  OAI21_X1 U6411 ( .B1(n5246), .B2(n6769), .A(n5228), .ZN(n5229) );
  AOI21_X1 U6412 ( .B1(n6716), .B2(n5248), .A(n5229), .ZN(n5230) );
  OAI21_X1 U6413 ( .B1(n5251), .B2(n7263), .A(n5230), .ZN(U3022) );
  AOI22_X1 U6414 ( .A1(n6698), .A2(n5244), .B1(n6757), .B2(n5243), .ZN(n5231)
         );
  OAI21_X1 U6415 ( .B1(n6742), .B2(n5246), .A(n5231), .ZN(n5232) );
  AOI21_X1 U6416 ( .B1(n6708), .B2(n5248), .A(n5232), .ZN(n5233) );
  OAI21_X1 U6417 ( .B1(n5251), .B2(n5234), .A(n5233), .ZN(U3020) );
  INV_X1 U6418 ( .A(n6790), .ZN(n6801) );
  AOI22_X1 U6419 ( .A1(n6800), .A2(n5244), .B1(n6799), .B2(n5243), .ZN(n5235)
         );
  OAI21_X1 U6420 ( .B1(n5246), .B2(n6804), .A(n5235), .ZN(n5236) );
  AOI21_X1 U6421 ( .B1(n6801), .B2(n5248), .A(n5236), .ZN(n5237) );
  OAI21_X1 U6422 ( .B1(n5251), .B2(n5238), .A(n5237), .ZN(U3026) );
  AOI22_X1 U6423 ( .A1(n6808), .A2(n5244), .B1(n6806), .B2(n5243), .ZN(n5239)
         );
  OAI21_X1 U6424 ( .B1(n5246), .B2(n6814), .A(n5239), .ZN(n5240) );
  AOI21_X1 U6425 ( .B1(n6810), .B2(n5248), .A(n5240), .ZN(n5241) );
  OAI21_X1 U6426 ( .B1(n5251), .B2(n5242), .A(n5241), .ZN(U3027) );
  AOI22_X1 U6427 ( .A1(n6727), .A2(n5244), .B1(n6785), .B2(n5243), .ZN(n5245)
         );
  OAI21_X1 U6428 ( .B1(n5246), .B2(n6783), .A(n5245), .ZN(n5247) );
  AOI21_X1 U6429 ( .B1(n6728), .B2(n5248), .A(n5247), .ZN(n5249) );
  OAI21_X1 U6430 ( .B1(n5251), .B2(n5250), .A(n5249), .ZN(U3025) );
  OAI21_X1 U6431 ( .B1(n5252), .B2(n5253), .A(n5371), .ZN(n6303) );
  OR2_X1 U6432 ( .A1(n5254), .A2(n5127), .ZN(n5255) );
  NAND2_X1 U6433 ( .A1(n5255), .A2(n5376), .ZN(n6308) );
  INV_X1 U6434 ( .A(n6308), .ZN(n5369) );
  AOI22_X1 U6435 ( .A1(n4474), .A2(n5369), .B1(n5802), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5256) );
  OAI21_X1 U6436 ( .B1(n6303), .B2(n6152), .A(n5256), .ZN(U2851) );
  AOI22_X1 U6437 ( .A1(n6390), .A2(DATAI_8_), .B1(n6386), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5257) );
  OAI21_X1 U6438 ( .B1(n6303), .B2(n6156), .A(n5257), .ZN(U2883) );
  OAI222_X1 U6439 ( .A1(n6156), .A2(n5259), .B1(n5577), .B2(n5258), .C1(n6394), 
        .C2(n4871), .ZN(U2884) );
  OAI21_X1 U6440 ( .B1(n5262), .B2(n5261), .A(n3195), .ZN(n6506) );
  NAND2_X1 U6441 ( .A1(n6567), .A2(REIP_REG_7__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U6442 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5263)
         );
  OAI211_X1 U6443 ( .C1(n6466), .C2(n5439), .A(n6503), .B(n5263), .ZN(n5264)
         );
  AOI21_X1 U6444 ( .B1(n5442), .B2(n6461), .A(n5264), .ZN(n5265) );
  OAI21_X1 U6445 ( .B1(n6506), .B2(n6468), .A(n5265), .ZN(U2979) );
  NOR2_X1 U6446 ( .A1(n6073), .A2(n6213), .ZN(n5387) );
  INV_X1 U6447 ( .A(n5387), .ZN(n5267) );
  OAI21_X1 U6448 ( .B1(n5268), .B2(n5267), .A(n6753), .ZN(n5272) );
  NAND3_X1 U6449 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6844), .A3(n6838), .ZN(n6691) );
  NOR2_X1 U6450 ( .A1(n5388), .A2(n6691), .ZN(n5291) );
  AOI21_X1 U6451 ( .B1(n5269), .B2(n6692), .A(n5291), .ZN(n5273) );
  INV_X1 U6452 ( .A(n5273), .ZN(n5271) );
  AOI21_X1 U6453 ( .B1(n6658), .B2(n6691), .A(n6586), .ZN(n5270) );
  OAI21_X1 U6454 ( .B1(n5272), .B2(n5271), .A(n5270), .ZN(n5290) );
  OAI22_X1 U6455 ( .A1(n5273), .A2(n5272), .B1(n3658), .B2(n6691), .ZN(n5289)
         );
  AOI22_X1 U6456 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5290), .B1(n7373), 
        .B2(n5289), .ZN(n5276) );
  AOI22_X1 U6457 ( .A1(n6735), .A2(n6639), .B1(n6723), .B2(n5291), .ZN(n5275)
         );
  OAI211_X1 U6458 ( .C1(n5315), .C2(n7369), .A(n5276), .B(n5275), .ZN(U3096)
         );
  AOI22_X1 U6459 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5290), .B1(n6806), 
        .B2(n5289), .ZN(n5278) );
  AOI22_X1 U6460 ( .A1(n6735), .A2(n5505), .B1(n6808), .B2(n5291), .ZN(n5277)
         );
  OAI211_X1 U6461 ( .C1(n5315), .C2(n6795), .A(n5278), .B(n5277), .ZN(U3099)
         );
  AOI22_X1 U6462 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5290), .B1(n6799), 
        .B2(n5289), .ZN(n5280) );
  AOI22_X1 U6463 ( .A1(n6735), .A2(n5522), .B1(n6800), .B2(n5291), .ZN(n5279)
         );
  OAI211_X1 U6464 ( .C1(n5315), .C2(n6790), .A(n5280), .B(n5279), .ZN(U3098)
         );
  AOI22_X1 U6465 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5290), .B1(n6785), 
        .B2(n5289), .ZN(n5282) );
  AOI22_X1 U6466 ( .A1(n6735), .A2(n6645), .B1(n6727), .B2(n5291), .ZN(n5281)
         );
  OAI211_X1 U6467 ( .C1(n5315), .C2(n6788), .A(n5282), .B(n5281), .ZN(U3097)
         );
  AOI22_X1 U6468 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5290), .B1(n6771), 
        .B2(n5289), .ZN(n5284) );
  AOI22_X1 U6469 ( .A1(n6735), .A2(n6633), .B1(n6715), .B2(n5291), .ZN(n5283)
         );
  OAI211_X1 U6470 ( .C1(n5315), .C2(n6774), .A(n5284), .B(n5283), .ZN(U3094)
         );
  AOI22_X1 U6471 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5290), .B1(n6778), 
        .B2(n5289), .ZN(n5286) );
  AOI22_X1 U6472 ( .A1(n6735), .A2(n6636), .B1(n6719), .B2(n5291), .ZN(n5285)
         );
  OAI211_X1 U6473 ( .C1(n5315), .C2(n6781), .A(n5286), .B(n5285), .ZN(U3095)
         );
  AOI22_X1 U6474 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5290), .B1(n6757), 
        .B2(n5289), .ZN(n5288) );
  AOI22_X1 U6475 ( .A1(n6735), .A2(n6627), .B1(n6698), .B2(n5291), .ZN(n5287)
         );
  OAI211_X1 U6476 ( .C1(n5315), .C2(n6760), .A(n5288), .B(n5287), .ZN(U3092)
         );
  AOI22_X1 U6477 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5290), .B1(n6764), 
        .B2(n5289), .ZN(n5293) );
  AOI22_X1 U6478 ( .A1(n6735), .A2(n6630), .B1(n6711), .B2(n5291), .ZN(n5292)
         );
  OAI211_X1 U6479 ( .C1(n5315), .C2(n6767), .A(n5293), .B(n5292), .ZN(U3093)
         );
  NOR2_X1 U6480 ( .A1(n6204), .A2(n5294), .ZN(n5295) );
  INV_X1 U6481 ( .A(n6348), .ZN(n5455) );
  OAI21_X1 U6482 ( .B1(n5434), .B2(n6334), .A(n6333), .ZN(n6310) );
  OAI21_X1 U6483 ( .B1(n6334), .B2(n5296), .A(n6899), .ZN(n5297) );
  NAND2_X1 U6484 ( .A1(n6310), .A2(n5297), .ZN(n5301) );
  NAND2_X1 U6485 ( .A1(n5298), .A2(n6333), .ZN(n6312) );
  OAI22_X1 U6486 ( .A1(n5092), .A2(n6354), .B1(n6362), .B2(n6522), .ZN(n5299)
         );
  AOI211_X1 U6487 ( .C1(n6346), .C2(EBX_REG_5__SCAN_IN), .A(n6323), .B(n5299), 
        .ZN(n5300) );
  NAND2_X1 U6488 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  AOI21_X1 U6489 ( .B1(n6357), .B2(n5303), .A(n5302), .ZN(n5304) );
  OAI21_X1 U6490 ( .B1(n5455), .B2(n5305), .A(n5304), .ZN(U2822) );
  NAND2_X1 U6491 ( .A1(n5315), .A2(n7377), .ZN(n5306) );
  AOI21_X1 U6492 ( .B1(n5306), .B2(STATEBS16_REG_SCAN_IN), .A(n6658), .ZN(
        n5312) );
  AND2_X1 U6493 ( .A1(n5307), .A2(n4893), .ZN(n6747) );
  NOR2_X1 U6494 ( .A1(n5308), .A2(n6850), .ZN(n5309) );
  AOI22_X1 U6495 ( .A1(n5312), .A2(n6747), .B1(n5484), .B2(n5309), .ZN(n5351)
         );
  INV_X1 U6496 ( .A(n6747), .ZN(n5311) );
  NAND2_X1 U6497 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5310), .ZN(n6756) );
  OR2_X1 U6498 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6756), .ZN(n5345)
         );
  AOI22_X1 U6499 ( .A1(n5312), .A2(n5311), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5345), .ZN(n5313) );
  NAND2_X1 U6500 ( .A1(n5344), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5318)
         );
  OAI22_X1 U6501 ( .A1(n7377), .A2(n6795), .B1(n5345), .B2(n6794), .ZN(n5316)
         );
  AOI21_X1 U6502 ( .B1(n5347), .B2(n5505), .A(n5316), .ZN(n5317) );
  OAI211_X1 U6503 ( .C1(n5351), .C2(n5319), .A(n5318), .B(n5317), .ZN(U3107)
         );
  NAND2_X1 U6504 ( .A1(n5344), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5322)
         );
  OAI22_X1 U6505 ( .A1(n7377), .A2(n6760), .B1(n5345), .B2(n6741), .ZN(n5320)
         );
  AOI21_X1 U6506 ( .B1(n5347), .B2(n6627), .A(n5320), .ZN(n5321) );
  OAI211_X1 U6507 ( .C1(n5351), .C2(n5323), .A(n5322), .B(n5321), .ZN(U3100)
         );
  NAND2_X1 U6508 ( .A1(n5344), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5326)
         );
  OAI22_X1 U6509 ( .A1(n7377), .A2(n6767), .B1(n5345), .B2(n6761), .ZN(n5324)
         );
  AOI21_X1 U6510 ( .B1(n5347), .B2(n6630), .A(n5324), .ZN(n5325) );
  OAI211_X1 U6511 ( .C1(n5351), .C2(n5327), .A(n5326), .B(n5325), .ZN(U3101)
         );
  NAND2_X1 U6512 ( .A1(n5344), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5330)
         );
  OAI22_X1 U6513 ( .A1(n7377), .A2(n6774), .B1(n5345), .B2(n6768), .ZN(n5328)
         );
  AOI21_X1 U6514 ( .B1(n5347), .B2(n6633), .A(n5328), .ZN(n5329) );
  OAI211_X1 U6515 ( .C1(n5351), .C2(n5331), .A(n5330), .B(n5329), .ZN(U3102)
         );
  NAND2_X1 U6516 ( .A1(n5344), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5334)
         );
  OAI22_X1 U6517 ( .A1(n7377), .A2(n6781), .B1(n5345), .B2(n6775), .ZN(n5332)
         );
  AOI21_X1 U6518 ( .B1(n5347), .B2(n6636), .A(n5332), .ZN(n5333) );
  OAI211_X1 U6519 ( .C1(n5351), .C2(n5335), .A(n5334), .B(n5333), .ZN(U3103)
         );
  NAND2_X1 U6520 ( .A1(n5344), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5338)
         );
  OAI22_X1 U6521 ( .A1(n7377), .A2(n7369), .B1(n5345), .B2(n7368), .ZN(n5336)
         );
  AOI21_X1 U6522 ( .B1(n5347), .B2(n6639), .A(n5336), .ZN(n5337) );
  OAI211_X1 U6523 ( .C1(n5351), .C2(n5339), .A(n5338), .B(n5337), .ZN(U3104)
         );
  NAND2_X1 U6524 ( .A1(n5344), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5342)
         );
  OAI22_X1 U6525 ( .A1(n7377), .A2(n6788), .B1(n5345), .B2(n6782), .ZN(n5340)
         );
  AOI21_X1 U6526 ( .B1(n5347), .B2(n6645), .A(n5340), .ZN(n5341) );
  OAI211_X1 U6527 ( .C1(n5351), .C2(n5343), .A(n5342), .B(n5341), .ZN(U3105)
         );
  NAND2_X1 U6528 ( .A1(n5344), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5349)
         );
  OAI22_X1 U6529 ( .A1(n7377), .A2(n6790), .B1(n5345), .B2(n6789), .ZN(n5346)
         );
  AOI21_X1 U6530 ( .B1(n5347), .B2(n5522), .A(n5346), .ZN(n5348) );
  OAI211_X1 U6531 ( .C1(n5351), .C2(n5350), .A(n5349), .B(n5348), .ZN(U3106)
         );
  AND2_X1 U6532 ( .A1(n5353), .A2(n5352), .ZN(n6349) );
  INV_X1 U6533 ( .A(n6349), .ZN(n6339) );
  INV_X1 U6534 ( .A(n5354), .ZN(n6568) );
  AOI22_X1 U6535 ( .A1(n6568), .A2(n6322), .B1(n6346), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5355) );
  OAI21_X1 U6536 ( .B1(n6653), .B2(n6339), .A(n5355), .ZN(n5356) );
  AOI21_X1 U6537 ( .B1(n6278), .B2(REIP_REG_0__SCAN_IN), .A(n5356), .ZN(n5358)
         );
  OAI21_X1 U6538 ( .B1(n6357), .B2(n6332), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5357) );
  OAI211_X1 U6539 ( .C1(n5455), .C2(n6471), .A(n5358), .B(n5357), .ZN(U2827)
         );
  OAI21_X1 U6540 ( .B1(n5361), .B2(n5360), .A(n5359), .ZN(n5385) );
  AND2_X1 U6541 ( .A1(n6567), .A2(REIP_REG_8__SCAN_IN), .ZN(n5379) );
  NOR2_X1 U6542 ( .A1(n6511), .A2(n5366), .ZN(n6490) );
  NAND2_X1 U6543 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6514) );
  OAI21_X1 U6544 ( .B1(n6514), .B2(n6527), .A(n6558), .ZN(n6536) );
  NAND2_X1 U6545 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U6546 ( .A1(n6564), .A2(n6553), .ZN(n6554) );
  NAND3_X1 U6547 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6554), .ZN(n5365) );
  NOR2_X1 U6548 ( .A1(n7294), .A2(n5365), .ZN(n6517) );
  NAND2_X1 U6549 ( .A1(n6536), .A2(n6517), .ZN(n6521) );
  NOR2_X1 U6550 ( .A1(n5363), .A2(n6521), .ZN(n6507) );
  OAI21_X1 U6551 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6507), .ZN(n5367) );
  NAND2_X1 U6552 ( .A1(n6558), .A2(n5364), .ZN(n5598) );
  NOR2_X1 U6553 ( .A1(n6558), .A2(n5365), .ZN(n6532) );
  NAND3_X1 U6554 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6532), .ZN(n5550) );
  INV_X1 U6555 ( .A(n5599), .ZN(n6515) );
  NAND2_X1 U6556 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U6557 ( .A1(n6537), .A2(n6514), .ZN(n6528) );
  NAND3_X1 U6558 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6528), .ZN(n5551) );
  AOI22_X1 U6559 ( .A1(n5598), .A2(n5550), .B1(n6515), .B2(n5551), .ZN(n6512)
         );
  OAI22_X1 U6560 ( .A1(n6490), .A2(n5367), .B1(n6512), .B2(n5366), .ZN(n5368)
         );
  AOI211_X1 U6561 ( .C1(n6569), .C2(n5369), .A(n5379), .B(n5368), .ZN(n5370)
         );
  OAI21_X1 U6562 ( .B1(n5385), .B2(n6478), .A(n5370), .ZN(U3010) );
  INV_X1 U6563 ( .A(n5371), .ZN(n5374) );
  NAND2_X1 U6564 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  OAI21_X1 U6565 ( .B1(n5374), .B2(n5373), .A(n5375), .ZN(n6290) );
  AOI21_X1 U6566 ( .B1(n5377), .B2(n5376), .A(n3226), .ZN(n6497) );
  AOI22_X1 U6567 ( .A1(n4474), .A2(n6497), .B1(EBX_REG_9__SCAN_IN), .B2(n5802), 
        .ZN(n5378) );
  OAI21_X1 U6568 ( .B1(n6290), .B2(n6152), .A(n5378), .ZN(U2850) );
  INV_X1 U6569 ( .A(n6303), .ZN(n5383) );
  INV_X1 U6570 ( .A(n6305), .ZN(n5381) );
  AOI21_X1 U6571 ( .B1(n6456), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5379), 
        .ZN(n5380) );
  OAI21_X1 U6572 ( .B1(n5381), .B2(n6466), .A(n5380), .ZN(n5382) );
  AOI21_X1 U6573 ( .B1(n5383), .B2(n6461), .A(n5382), .ZN(n5384) );
  OAI21_X1 U6574 ( .B1(n5385), .B2(n6468), .A(n5384), .ZN(U2978) );
  INV_X1 U6575 ( .A(n5393), .ZN(n5391) );
  AOI21_X1 U6576 ( .B1(n6650), .B2(n5387), .A(n6658), .ZN(n5392) );
  NOR2_X1 U6577 ( .A1(n5388), .A2(n5393), .ZN(n5412) );
  AOI21_X1 U6578 ( .B1(n5389), .B2(n6833), .A(n5412), .ZN(n5394) );
  NAND2_X1 U6579 ( .A1(n5392), .A2(n5394), .ZN(n5390) );
  OAI211_X1 U6580 ( .C1(n6753), .C2(n5391), .A(n6749), .B(n5390), .ZN(n5411)
         );
  INV_X1 U6581 ( .A(n5392), .ZN(n5395) );
  OAI22_X1 U6582 ( .A1(n5395), .A2(n5394), .B1(n5393), .B2(n3658), .ZN(n5410)
         );
  AOI22_X1 U6583 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n7373), .ZN(n5397) );
  AOI22_X1 U6584 ( .A1(n6621), .A2(n6639), .B1(n6723), .B2(n5412), .ZN(n5396)
         );
  OAI211_X1 U6585 ( .C1(n7369), .C2(n5415), .A(n5397), .B(n5396), .ZN(U3064)
         );
  AOI22_X1 U6586 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6806), .ZN(n5399) );
  AOI22_X1 U6587 ( .A1(n6621), .A2(n5505), .B1(n6808), .B2(n5412), .ZN(n5398)
         );
  OAI211_X1 U6588 ( .C1(n6795), .C2(n5415), .A(n5399), .B(n5398), .ZN(U3067)
         );
  AOI22_X1 U6589 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6778), .ZN(n5401) );
  AOI22_X1 U6590 ( .A1(n6621), .A2(n6636), .B1(n6719), .B2(n5412), .ZN(n5400)
         );
  OAI211_X1 U6591 ( .C1(n6781), .C2(n5415), .A(n5401), .B(n5400), .ZN(U3063)
         );
  AOI22_X1 U6592 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6785), .ZN(n5403) );
  AOI22_X1 U6593 ( .A1(n6621), .A2(n6645), .B1(n6727), .B2(n5412), .ZN(n5402)
         );
  OAI211_X1 U6594 ( .C1(n6788), .C2(n5415), .A(n5403), .B(n5402), .ZN(U3065)
         );
  AOI22_X1 U6595 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6757), .ZN(n5405) );
  AOI22_X1 U6596 ( .A1(n6621), .A2(n6627), .B1(n6698), .B2(n5412), .ZN(n5404)
         );
  OAI211_X1 U6597 ( .C1(n6760), .C2(n5415), .A(n5405), .B(n5404), .ZN(U3060)
         );
  AOI22_X1 U6598 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6799), .ZN(n5407) );
  AOI22_X1 U6599 ( .A1(n6621), .A2(n5522), .B1(n6800), .B2(n5412), .ZN(n5406)
         );
  OAI211_X1 U6600 ( .C1(n6790), .C2(n5415), .A(n5407), .B(n5406), .ZN(U3066)
         );
  AOI22_X1 U6601 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6764), .ZN(n5409) );
  AOI22_X1 U6602 ( .A1(n6621), .A2(n6630), .B1(n6711), .B2(n5412), .ZN(n5408)
         );
  OAI211_X1 U6603 ( .C1(n6767), .C2(n5415), .A(n5409), .B(n5408), .ZN(U3061)
         );
  AOI22_X1 U6604 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5411), .B1(n5410), 
        .B2(n6771), .ZN(n5414) );
  AOI22_X1 U6605 ( .A1(n6621), .A2(n6633), .B1(n6715), .B2(n5412), .ZN(n5413)
         );
  OAI211_X1 U6606 ( .C1(n6774), .C2(n5415), .A(n5414), .B(n5413), .ZN(U3062)
         );
  INV_X1 U6607 ( .A(n6685), .ZN(n5417) );
  NOR3_X1 U6608 ( .A1(n6644), .A2(n5417), .A3(n6658), .ZN(n5419) );
  INV_X1 U6609 ( .A(n5478), .ZN(n6655) );
  OAI21_X1 U6610 ( .B1(n5419), .B2(n5418), .A(n6655), .ZN(n5422) );
  NOR2_X1 U6611 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6661), .ZN(n6643)
         );
  INV_X1 U6612 ( .A(n6643), .ZN(n5420) );
  AOI211_X1 U6613 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5420), .A(n6694), .B(
        n5480), .ZN(n5421) );
  INV_X1 U6614 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5428) );
  NAND3_X1 U6615 ( .A1(n6702), .A2(n6753), .A3(n5478), .ZN(n5424) );
  NAND3_X1 U6616 ( .A1(n6703), .A2(n5484), .A3(n6850), .ZN(n5423) );
  NAND2_X1 U6617 ( .A1(n5424), .A2(n5423), .ZN(n6642) );
  AOI22_X1 U6618 ( .A1(n6808), .A2(n6643), .B1(n6806), .B2(n6642), .ZN(n5425)
         );
  OAI21_X1 U6619 ( .B1(n6795), .B2(n6685), .A(n5425), .ZN(n5426) );
  AOI21_X1 U6620 ( .B1(n5505), .B2(n6644), .A(n5426), .ZN(n5427) );
  OAI21_X1 U6621 ( .B1(n6626), .B2(n5428), .A(n5427), .ZN(U3075) );
  INV_X1 U6622 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5432) );
  AOI22_X1 U6623 ( .A1(n6800), .A2(n6643), .B1(n6799), .B2(n6642), .ZN(n5429)
         );
  OAI21_X1 U6624 ( .B1(n6790), .B2(n6685), .A(n5429), .ZN(n5430) );
  AOI21_X1 U6625 ( .B1(n5522), .B2(n6644), .A(n5430), .ZN(n5431) );
  OAI21_X1 U6626 ( .B1(n6626), .B2(n5432), .A(n5431), .ZN(U3074) );
  AOI22_X1 U6627 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6346), .B1(n6322), .B2(n6505), 
        .ZN(n5433) );
  OAI211_X1 U6628 ( .C1(n6354), .C2(n7310), .A(n5433), .B(n6312), .ZN(n5441)
         );
  INV_X1 U6629 ( .A(n6334), .ZN(n5435) );
  INV_X1 U6630 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6900) );
  AND3_X1 U6631 ( .A1(n5435), .A2(n5434), .A3(n6900), .ZN(n6309) );
  OAI21_X1 U6632 ( .B1(n6310), .B2(n6309), .A(REIP_REG_7__SCAN_IN), .ZN(n5438)
         );
  OR3_X1 U6633 ( .A1(n6334), .A2(REIP_REG_7__SCAN_IN), .A3(n5436), .ZN(n5437)
         );
  OAI211_X1 U6634 ( .C1(n6343), .C2(n5439), .A(n5438), .B(n5437), .ZN(n5440)
         );
  AOI211_X1 U6635 ( .C1(n6315), .C2(n5442), .A(n5441), .B(n5440), .ZN(n5443)
         );
  INV_X1 U6636 ( .A(n5443), .ZN(U2820) );
  OAI222_X1 U6637 ( .A1(n6290), .A2(n6156), .B1(n5577), .B2(n5444), .C1(n6394), 
        .C2(n4864), .ZN(U2882) );
  OAI21_X1 U6638 ( .B1(n6321), .B2(n6334), .A(n6333), .ZN(n6325) );
  AOI22_X1 U6639 ( .A1(n6544), .A2(n6322), .B1(n6346), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5446) );
  OR4_X1 U6640 ( .A1(n6334), .A2(n6321), .A3(n7306), .A4(n6895), .ZN(n5445) );
  NAND2_X1 U6641 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  AOI21_X1 U6642 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6325), .A(n5447), .ZN(n5448)
         );
  OAI21_X1 U6643 ( .B1(n5449), .B2(n6354), .A(n5448), .ZN(n5452) );
  NOR2_X1 U6644 ( .A1(n6343), .A2(n5450), .ZN(n5451) );
  AOI211_X1 U6645 ( .C1(n6349), .C2(n4893), .A(n5452), .B(n5451), .ZN(n5453)
         );
  OAI21_X1 U6646 ( .B1(n5455), .B2(n5454), .A(n5453), .ZN(U2824) );
  INV_X1 U6647 ( .A(n5375), .ZN(n5458) );
  OR2_X1 U6648 ( .A1(n5375), .A2(n5456), .ZN(n5529) );
  OAI21_X1 U6649 ( .B1(n5458), .B2(n5457), .A(n5529), .ZN(n6283) );
  INV_X1 U6650 ( .A(DATAI_10_), .ZN(n7205) );
  OAI222_X1 U6651 ( .A1(n6283), .A2(n6156), .B1(n5577), .B2(n7205), .C1(n6394), 
        .C2(n3862), .ZN(U2881) );
  XNOR2_X1 U6652 ( .A(n5459), .B(n3226), .ZN(n6486) );
  OAI222_X1 U6653 ( .A1(n6152), .A2(n6283), .B1(n6380), .B2(n4396), .C1(n6371), 
        .C2(n6486), .ZN(U2849) );
  XOR2_X1 U6654 ( .A(n5460), .B(n6168), .Z(n5548) );
  INV_X1 U6655 ( .A(n5548), .ZN(n5533) );
  INV_X1 U6656 ( .A(n5546), .ZN(n5469) );
  INV_X1 U6657 ( .A(n6278), .ZN(n6259) );
  OR2_X1 U6658 ( .A1(n6259), .A2(n6258), .ZN(n6271) );
  OR2_X1 U6659 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  NAND2_X1 U6660 ( .A1(n5463), .A2(n6195), .ZN(n5557) );
  OAI22_X1 U6661 ( .A1(n5464), .A2(n6354), .B1(n6362), .B2(n5557), .ZN(n5465)
         );
  AOI211_X1 U6662 ( .C1(n6346), .C2(EBX_REG_12__SCAN_IN), .A(n6323), .B(n5465), 
        .ZN(n5466) );
  OAI221_X1 U6663 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6257), .C1(n5467), .C2(
        n6271), .A(n5466), .ZN(n5468) );
  AOI21_X1 U6664 ( .B1(n6357), .B2(n5469), .A(n5468), .ZN(n5470) );
  OAI21_X1 U6665 ( .B1(n5533), .B2(n6302), .A(n5470), .ZN(U2815) );
  XNOR2_X1 U6666 ( .A(n3204), .B(n6485), .ZN(n5472) );
  XNOR2_X1 U6667 ( .A(n5471), .B(n5472), .ZN(n6499) );
  NAND2_X1 U6668 ( .A1(n6499), .A2(n6460), .ZN(n5475) );
  NAND2_X1 U6669 ( .A1(n6567), .A2(REIP_REG_9__SCAN_IN), .ZN(n6495) );
  OAI21_X1 U6670 ( .B1(n6474), .B2(n3840), .A(n6495), .ZN(n5473) );
  AOI21_X1 U6671 ( .B1(n6438), .B2(n6291), .A(n5473), .ZN(n5474) );
  OAI211_X1 U6672 ( .C1(n6470), .C2(n6290), .A(n5475), .B(n5474), .ZN(U2977)
         );
  NOR2_X1 U6673 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5476), .ZN(n5517)
         );
  OAI21_X1 U6674 ( .B1(n5521), .B2(n5477), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5479) );
  NAND2_X1 U6675 ( .A1(n5478), .A2(n4893), .ZN(n5486) );
  NOR4_X1 U6676 ( .A1(n6850), .A2(n6694), .A3(n5481), .A4(n5480), .ZN(n5482)
         );
  OAI21_X1 U6677 ( .B1(n5517), .B2(n7315), .A(n5482), .ZN(n5483) );
  NAND3_X1 U6678 ( .A1(n6703), .A2(n5484), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5485) );
  OAI21_X1 U6679 ( .B1(n5486), .B2(n6658), .A(n5485), .ZN(n5516) );
  AOI22_X1 U6680 ( .A1(n6715), .A2(n5517), .B1(n6771), .B2(n5516), .ZN(n5487)
         );
  OAI21_X1 U6681 ( .B1(n6774), .B2(n5519), .A(n5487), .ZN(n5488) );
  AOI21_X1 U6682 ( .B1(n6633), .B2(n5521), .A(n5488), .ZN(n5489) );
  OAI21_X1 U6683 ( .B1(n5525), .B2(n5490), .A(n5489), .ZN(U3134) );
  AOI22_X1 U6684 ( .A1(n6723), .A2(n5517), .B1(n7373), .B2(n5516), .ZN(n5491)
         );
  OAI21_X1 U6685 ( .B1(n7369), .B2(n5519), .A(n5491), .ZN(n5492) );
  AOI21_X1 U6686 ( .B1(n6639), .B2(n5521), .A(n5492), .ZN(n5493) );
  OAI21_X1 U6687 ( .B1(n5525), .B2(n5494), .A(n5493), .ZN(U3136) );
  AOI22_X1 U6688 ( .A1(n6727), .A2(n5517), .B1(n6785), .B2(n5516), .ZN(n5495)
         );
  OAI21_X1 U6689 ( .B1(n6788), .B2(n5519), .A(n5495), .ZN(n5496) );
  AOI21_X1 U6690 ( .B1(n6645), .B2(n5521), .A(n5496), .ZN(n5497) );
  OAI21_X1 U6691 ( .B1(n5525), .B2(n5498), .A(n5497), .ZN(U3137) );
  AOI22_X1 U6692 ( .A1(n6719), .A2(n5517), .B1(n6778), .B2(n5516), .ZN(n5499)
         );
  OAI21_X1 U6693 ( .B1(n6781), .B2(n5519), .A(n5499), .ZN(n5500) );
  AOI21_X1 U6694 ( .B1(n6636), .B2(n5521), .A(n5500), .ZN(n5501) );
  OAI21_X1 U6695 ( .B1(n5525), .B2(n5502), .A(n5501), .ZN(U3135) );
  AOI22_X1 U6696 ( .A1(n6808), .A2(n5517), .B1(n6806), .B2(n5516), .ZN(n5503)
         );
  OAI21_X1 U6697 ( .B1(n6795), .B2(n5519), .A(n5503), .ZN(n5504) );
  AOI21_X1 U6698 ( .B1(n5505), .B2(n5521), .A(n5504), .ZN(n5506) );
  OAI21_X1 U6699 ( .B1(n5525), .B2(n5507), .A(n5506), .ZN(U3139) );
  AOI22_X1 U6700 ( .A1(n6698), .A2(n5517), .B1(n6757), .B2(n5516), .ZN(n5508)
         );
  OAI21_X1 U6701 ( .B1(n6760), .B2(n5519), .A(n5508), .ZN(n5509) );
  AOI21_X1 U6702 ( .B1(n6627), .B2(n5521), .A(n5509), .ZN(n5510) );
  OAI21_X1 U6703 ( .B1(n5525), .B2(n5511), .A(n5510), .ZN(U3132) );
  AOI22_X1 U6704 ( .A1(n6711), .A2(n5517), .B1(n6764), .B2(n5516), .ZN(n5512)
         );
  OAI21_X1 U6705 ( .B1(n6767), .B2(n5519), .A(n5512), .ZN(n5513) );
  AOI21_X1 U6706 ( .B1(n6630), .B2(n5521), .A(n5513), .ZN(n5514) );
  OAI21_X1 U6707 ( .B1(n5525), .B2(n5515), .A(n5514), .ZN(U3133) );
  AOI22_X1 U6708 ( .A1(n6800), .A2(n5517), .B1(n6799), .B2(n5516), .ZN(n5518)
         );
  OAI21_X1 U6709 ( .B1(n6790), .B2(n5519), .A(n5518), .ZN(n5520) );
  AOI21_X1 U6710 ( .B1(n5522), .B2(n5521), .A(n5520), .ZN(n5523) );
  OAI21_X1 U6711 ( .B1(n5525), .B2(n5524), .A(n5523), .ZN(U3138) );
  INV_X1 U6712 ( .A(DATAI_12_), .ZN(n5527) );
  OAI222_X1 U6713 ( .A1(n5577), .A2(n5527), .B1(n6156), .B2(n5533), .C1(n5526), 
        .C2(n6394), .ZN(U2879) );
  AND2_X1 U6714 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  INV_X1 U6715 ( .A(DATAI_11_), .ZN(n5531) );
  OAI222_X1 U6716 ( .A1(n6372), .A2(n6156), .B1(n6394), .B2(n5532), .C1(n5577), 
        .C2(n5531), .ZN(U2880) );
  OAI222_X1 U6717 ( .A1(n5557), .A2(n6371), .B1(n6380), .B2(n4406), .C1(n6152), 
        .C2(n5533), .ZN(U2847) );
  NAND2_X1 U6718 ( .A1(n6433), .A2(n5535), .ZN(n5536) );
  XNOR2_X1 U6719 ( .A(n5534), .B(n5536), .ZN(n6491) );
  NAND2_X1 U6720 ( .A1(n6491), .A2(n6460), .ZN(n5539) );
  NAND2_X1 U6721 ( .A1(n6567), .A2(REIP_REG_10__SCAN_IN), .ZN(n6487) );
  OAI21_X1 U6722 ( .B1(n6474), .B2(n6280), .A(n6487), .ZN(n5537) );
  AOI21_X1 U6723 ( .B1(n6438), .B2(n6285), .A(n5537), .ZN(n5538) );
  OAI211_X1 U6724 ( .C1(n6470), .C2(n6283), .A(n5539), .B(n5538), .ZN(U2976)
         );
  INV_X1 U6725 ( .A(n5541), .ZN(n5542) );
  NOR2_X1 U6726 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  XNOR2_X1 U6727 ( .A(n5540), .B(n5544), .ZN(n5563) );
  NAND2_X1 U6728 ( .A1(n6567), .A2(REIP_REG_12__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U6729 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5545)
         );
  OAI211_X1 U6730 ( .C1(n6466), .C2(n5546), .A(n5556), .B(n5545), .ZN(n5547)
         );
  AOI21_X1 U6731 ( .B1(n5548), .B2(n6461), .A(n5547), .ZN(n5549) );
  OAI21_X1 U6732 ( .B1(n5563), .B2(n6468), .A(n5549), .ZN(U2974) );
  NAND3_X1 U6733 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6490), .ZN(n5552) );
  INV_X1 U6734 ( .A(n5597), .ZN(n5553) );
  NOR2_X1 U6735 ( .A1(n5552), .A2(n5551), .ZN(n5600) );
  INV_X1 U6736 ( .A(n5600), .ZN(n5554) );
  AOI22_X1 U6737 ( .A1(n5598), .A2(n5553), .B1(n6515), .B2(n5554), .ZN(n6476)
         );
  NOR2_X1 U6738 ( .A1(n5554), .A2(n6527), .ZN(n5624) );
  NOR2_X1 U6739 ( .A1(n5597), .A2(n5624), .ZN(n6069) );
  INV_X1 U6740 ( .A(n6069), .ZN(n6197) );
  NAND2_X1 U6741 ( .A1(n4558), .A2(n6197), .ZN(n6483) );
  AOI21_X1 U6742 ( .B1(n6476), .B2(n6483), .A(n5555), .ZN(n5561) );
  INV_X1 U6743 ( .A(n5556), .ZN(n5560) );
  NOR2_X1 U6744 ( .A1(n6551), .A2(n5557), .ZN(n5559) );
  NOR3_X1 U6745 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6069), .A3(n4558), 
        .ZN(n5558) );
  NOR4_X1 U6746 ( .A1(n5561), .A2(n5560), .A3(n5559), .A4(n5558), .ZN(n5562)
         );
  OAI21_X1 U6747 ( .B1(n5563), .B2(n6478), .A(n5562), .ZN(U3006) );
  OAI21_X1 U6748 ( .B1(n5566), .B2(n5565), .A(n5564), .ZN(n5951) );
  NAND2_X1 U6749 ( .A1(n6278), .A2(n5567), .ZN(n6249) );
  AOI21_X1 U6750 ( .B1(n7268), .B2(n5568), .A(n6249), .ZN(n5573) );
  XOR2_X1 U6751 ( .A(n6194), .B(n5569), .Z(n5590) );
  AOI22_X1 U6752 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6346), .B1(n6322), .B2(n5590), .ZN(n5570) );
  OAI211_X1 U6753 ( .C1(n6354), .C2(n5571), .A(n5570), .B(n6312), .ZN(n5572)
         );
  AOI211_X1 U6754 ( .C1(n6357), .C2(n5574), .A(n5573), .B(n5572), .ZN(n5575)
         );
  OAI21_X1 U6755 ( .B1(n5951), .B2(n6302), .A(n5575), .ZN(U2813) );
  AOI22_X1 U6756 ( .A1(n4474), .A2(n5590), .B1(EBX_REG_14__SCAN_IN), .B2(n5802), .ZN(n5576) );
  OAI21_X1 U6757 ( .B1(n5951), .B2(n6152), .A(n5576), .ZN(U2845) );
  INV_X1 U6758 ( .A(DATAI_14_), .ZN(n5578) );
  OAI222_X1 U6759 ( .A1(n5951), .A2(n6156), .B1(n6394), .B2(n5579), .C1(n5578), 
        .C2(n5577), .ZN(U2877) );
  INV_X1 U6760 ( .A(n5581), .ZN(n5583) );
  NAND2_X1 U6761 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  XNOR2_X1 U6762 ( .A(n5580), .B(n5584), .ZN(n5957) );
  NAND2_X1 U6763 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5587) );
  NOR2_X1 U6764 ( .A1(n4562), .A2(n5587), .ZN(n5596) );
  OAI21_X1 U6765 ( .B1(n5596), .B2(n5585), .A(n6476), .ZN(n5586) );
  AOI21_X1 U6766 ( .B1(n5607), .B2(n5587), .A(n5586), .ZN(n6202) );
  NOR2_X1 U6767 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5587), .ZN(n6198)
         );
  OAI21_X1 U6768 ( .B1(n5588), .B2(n5597), .A(n6198), .ZN(n5589) );
  AOI21_X1 U6769 ( .B1(n6202), .B2(n5589), .A(n7224), .ZN(n5594) );
  NAND3_X1 U6770 ( .A1(n5596), .A2(n7224), .A3(n6197), .ZN(n5592) );
  NAND2_X1 U6771 ( .A1(n6569), .A2(n5590), .ZN(n5591) );
  OAI211_X1 U6772 ( .C1(n7268), .C2(n6556), .A(n5592), .B(n5591), .ZN(n5593)
         );
  NOR2_X1 U6773 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  OAI21_X1 U6774 ( .B1(n5957), .B2(n6478), .A(n5595), .ZN(U3004) );
  NAND2_X1 U6775 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5596), .ZN(n6068) );
  NOR2_X1 U6776 ( .A1(n7218), .A2(n6068), .ZN(n6191) );
  NAND2_X1 U6777 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6191), .ZN(n6180) );
  NOR2_X1 U6778 ( .A1(n7215), .A2(n6180), .ZN(n6056) );
  NAND2_X1 U6779 ( .A1(n5597), .A2(n6056), .ZN(n5627) );
  NAND2_X1 U6780 ( .A1(n5627), .A2(n5598), .ZN(n5603) );
  INV_X1 U6781 ( .A(n6180), .ZN(n5625) );
  AOI21_X1 U6782 ( .B1(n5625), .B2(n5600), .A(n5599), .ZN(n5601) );
  INV_X1 U6783 ( .A(n5601), .ZN(n5602) );
  OR2_X1 U6784 ( .A1(n5605), .A2(n5604), .ZN(n6566) );
  INV_X1 U6785 ( .A(n5606), .ZN(n6028) );
  NAND2_X1 U6786 ( .A1(n6028), .A2(n6037), .ZN(n5626) );
  OAI21_X1 U6787 ( .B1(n5607), .B2(n6566), .A(n5626), .ZN(n5608) );
  NAND2_X1 U6788 ( .A1(n6186), .A2(n5608), .ZN(n6024) );
  NOR2_X1 U6789 ( .A1(n6518), .A2(n6013), .ZN(n5609) );
  NOR2_X1 U6790 ( .A1(n6024), .A2(n5609), .ZN(n6002) );
  INV_X1 U6791 ( .A(n5610), .ZN(n5628) );
  OAI21_X1 U6792 ( .B1(n6550), .B2(n5611), .A(n5628), .ZN(n5612) );
  NAND2_X1 U6793 ( .A1(n6002), .A2(n5612), .ZN(n5996) );
  INV_X1 U6794 ( .A(n5996), .ZN(n5615) );
  AND2_X1 U6795 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5629) );
  NOR2_X1 U6796 ( .A1(n6518), .A2(n5629), .ZN(n5613) );
  INV_X1 U6797 ( .A(n5972), .ZN(n5661) );
  OAI21_X1 U6798 ( .B1(n6518), .B2(n5661), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n5614) );
  NOR2_X1 U6799 ( .A1(n5971), .A2(n5614), .ZN(n5960) );
  AOI211_X1 U6800 ( .C1(n6518), .C2(n5615), .A(n5630), .B(n5960), .ZN(n5634)
         );
  INV_X1 U6801 ( .A(n5620), .ZN(n5619) );
  NAND2_X1 U6802 ( .A1(n5620), .A2(n4385), .ZN(n5655) );
  NAND2_X1 U6803 ( .A1(n5658), .A2(EBX_REG_30__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U6804 ( .A1(n5657), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5616) );
  AND2_X1 U6805 ( .A1(n5617), .A2(n5616), .ZN(n5653) );
  INV_X1 U6806 ( .A(n5653), .ZN(n5618) );
  OAI211_X1 U6807 ( .C1(n5619), .C2(n4467), .A(n5655), .B(n5618), .ZN(n5623)
         );
  INV_X1 U6808 ( .A(n4467), .ZN(n5621) );
  OAI211_X1 U6809 ( .C1(n5621), .C2(n4385), .A(n5653), .B(n5620), .ZN(n5622)
         );
  NAND2_X1 U6810 ( .A1(n5623), .A2(n5622), .ZN(n5688) );
  NAND2_X1 U6811 ( .A1(n5625), .A2(n5624), .ZN(n6055) );
  AOI21_X1 U6812 ( .B1(n6055), .B2(n5627), .A(n5626), .ZN(n6012) );
  NAND2_X1 U6813 ( .A1(n6012), .A2(n6013), .ZN(n6007) );
  INV_X1 U6814 ( .A(n5629), .ZN(n5990) );
  NAND4_X1 U6815 ( .A1(n5983), .A2(n5661), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5630), .ZN(n5632) );
  OAI211_X1 U6816 ( .C1(n5688), .C2(n6551), .A(n5632), .B(n5631), .ZN(n5633)
         );
  NOR2_X1 U6817 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  OAI21_X1 U6818 ( .B1(n5636), .B2(n6478), .A(n5635), .ZN(U2988) );
  XNOR2_X1 U6819 ( .A(n3204), .B(n7237), .ZN(n5919) );
  INV_X1 U6820 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5910) );
  XNOR2_X1 U6821 ( .A(n3203), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5905)
         );
  NAND2_X1 U6822 ( .A1(n5906), .A2(n5905), .ZN(n5904) );
  NAND2_X1 U6823 ( .A1(n4555), .A2(n7269), .ZN(n5894) );
  NOR2_X1 U6824 ( .A1(n5904), .A2(n5894), .ZN(n5888) );
  NAND2_X1 U6825 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5637) );
  INV_X1 U6826 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5638) );
  INV_X1 U6827 ( .A(n5895), .ZN(n5640) );
  XNOR2_X1 U6828 ( .A(n5642), .B(n7174), .ZN(n5652) );
  OAI21_X1 U6829 ( .B1(n6007), .B2(n5889), .A(n7174), .ZN(n5644) );
  NAND2_X1 U6830 ( .A1(n6567), .A2(REIP_REG_24__SCAN_IN), .ZN(n5647) );
  OAI21_X1 U6831 ( .B1(n6551), .B2(n5767), .A(n5647), .ZN(n5643) );
  AOI21_X1 U6832 ( .B1(n5644), .B2(n5996), .A(n5643), .ZN(n5645) );
  OAI21_X1 U6833 ( .B1(n5652), .B2(n6478), .A(n5645), .ZN(U2994) );
  NAND2_X1 U6834 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5646)
         );
  OAI211_X1 U6835 ( .C1(n5648), .C2(n6466), .A(n5647), .B(n5646), .ZN(n5649)
         );
  AOI21_X1 U6836 ( .B1(n5650), .B2(n6461), .A(n5649), .ZN(n5651) );
  OAI21_X1 U6837 ( .B1(n5652), .B2(n6468), .A(n5651), .ZN(U2962) );
  NAND2_X1 U6838 ( .A1(n5654), .A2(n5653), .ZN(n5656) );
  NAND2_X1 U6839 ( .A1(n5656), .A2(n5655), .ZN(n5660) );
  OAI22_X1 U6840 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5657), .ZN(n5659) );
  NAND3_X1 U6841 ( .A1(n5661), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5664) );
  INV_X1 U6842 ( .A(n5664), .ZN(n5662) );
  INV_X1 U6843 ( .A(n5971), .ZN(n5980) );
  OAI21_X1 U6844 ( .B1(n6518), .B2(n5662), .A(n5980), .ZN(n5663) );
  INV_X1 U6845 ( .A(n5983), .ZN(n5959) );
  NAND2_X1 U6846 ( .A1(n3297), .A2(n5665), .ZN(n5666) );
  AOI21_X1 U6847 ( .B1(n5663), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5666), 
        .ZN(n5667) );
  OAI21_X1 U6848 ( .B1(n5669), .B2(n6478), .A(n3294), .ZN(U2987) );
  NAND3_X1 U6849 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6850 ( .A1(n6278), .A2(n5730), .ZN(n5671) );
  NAND2_X1 U6851 ( .A1(n6103), .A2(n5671), .ZN(n6081) );
  AND2_X1 U6852 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5672) );
  NOR2_X1 U6853 ( .A1(n6334), .A2(n5672), .ZN(n5673) );
  NOR2_X1 U6854 ( .A1(n6334), .A2(REIP_REG_29__SCAN_IN), .ZN(n5674) );
  NOR2_X1 U6855 ( .A1(n5717), .A2(n5674), .ZN(n5691) );
  INV_X1 U6856 ( .A(n5691), .ZN(n5682) );
  NAND2_X1 U6857 ( .A1(n6357), .A2(n5675), .ZN(n5677) );
  AOI22_X1 U6858 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n6346), .ZN(n5676) );
  OAI211_X1 U6859 ( .C1(n6362), .C2(n5688), .A(n5677), .B(n5676), .ZN(n5681)
         );
  INV_X1 U6860 ( .A(n5730), .ZN(n5678) );
  NAND2_X1 U6861 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5678), .ZN(n5679) );
  NOR2_X1 U6862 ( .A1(n6080), .A2(n5679), .ZN(n5718) );
  NAND2_X1 U6863 ( .A1(n5718), .A2(REIP_REG_28__SCAN_IN), .ZN(n5700) );
  INV_X1 U6864 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6926) );
  NOR3_X1 U6865 ( .A1(n5700), .A2(REIP_REG_30__SCAN_IN), .A3(n6926), .ZN(n5680) );
  AOI211_X1 U6866 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5682), .A(n5681), .B(n5680), .ZN(n5683) );
  OAI21_X1 U6867 ( .B1(n5670), .B2(n6302), .A(n5683), .ZN(U2797) );
  AOI22_X1 U6868 ( .A1(n6384), .A2(DATAI_30_), .B1(n6386), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5687) );
  AND2_X1 U6869 ( .A1(n3351), .A2(n3499), .ZN(n5685) );
  NAND2_X1 U6870 ( .A1(n6387), .A2(DATAI_14_), .ZN(n5686) );
  OAI211_X1 U6871 ( .C1(n5670), .C2(n6156), .A(n5687), .B(n5686), .ZN(U2861)
         );
  INV_X1 U6872 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5689) );
  OAI222_X1 U6873 ( .A1(n6152), .A2(n5670), .B1(n5689), .B2(n6380), .C1(n5688), 
        .C2(n6371), .ZN(U2829) );
  INV_X1 U6874 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5690) );
  NAND3_X1 U6875 ( .A1(n5690), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6876 ( .A1(n5812), .A2(n6315), .ZN(n5698) );
  OAI21_X1 U6877 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6334), .A(n5691), .ZN(n5697) );
  INV_X1 U6878 ( .A(n5692), .ZN(n5694) );
  OAI22_X1 U6879 ( .A1(n6354), .A2(n5695), .B1(n5694), .B2(n5693), .ZN(n5696)
         );
  INV_X1 U6880 ( .A(n5849), .ZN(n5817) );
  INV_X1 U6881 ( .A(n5700), .ZN(n5707) );
  NAND2_X1 U6882 ( .A1(n5717), .A2(REIP_REG_29__SCAN_IN), .ZN(n5705) );
  OAI22_X1 U6883 ( .A1(n6354), .A2(n5702), .B1(n6331), .B2(n5701), .ZN(n5703)
         );
  AOI21_X1 U6884 ( .B1(n4475), .B2(n6322), .A(n5703), .ZN(n5704) );
  OAI211_X1 U6885 ( .C1(n6343), .C2(n5847), .A(n5705), .B(n5704), .ZN(n5706)
         );
  AOI21_X1 U6886 ( .B1(n5707), .B2(n6926), .A(n5706), .ZN(n5708) );
  OAI21_X1 U6887 ( .B1(n5817), .B2(n6302), .A(n5708), .ZN(U2798) );
  NAND2_X1 U6888 ( .A1(n5709), .A2(n5710), .ZN(n5711) );
  NOR2_X1 U6889 ( .A1(n6343), .A2(n5860), .ZN(n5716) );
  OR2_X1 U6890 ( .A1(n5727), .A2(n5712), .ZN(n5713) );
  NAND2_X1 U6891 ( .A1(n4467), .A2(n5713), .ZN(n5968) );
  AOI22_X1 U6892 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .B1(n6346), 
        .B2(EBX_REG_28__SCAN_IN), .ZN(n5714) );
  OAI21_X1 U6893 ( .B1(n5968), .B2(n6362), .A(n5714), .ZN(n5715) );
  AOI211_X1 U6894 ( .C1(n5717), .C2(REIP_REG_28__SCAN_IN), .A(n5716), .B(n5715), .ZN(n5720) );
  INV_X1 U6895 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U6896 ( .A1(n5718), .A2(n6928), .ZN(n5719) );
  OAI211_X1 U6897 ( .C1(n5858), .C2(n6302), .A(n5720), .B(n5719), .ZN(U2799)
         );
  INV_X1 U6898 ( .A(n5709), .ZN(n5722) );
  AOI21_X1 U6899 ( .B1(n5723), .B2(n5721), .A(n5722), .ZN(n5870) );
  INV_X1 U6900 ( .A(n5870), .ZN(n5822) );
  AOI22_X1 U6901 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6346), .B1(n5869), .B2(n6357), .ZN(n5724) );
  OAI21_X1 U6902 ( .B1(n5867), .B2(n6354), .A(n5724), .ZN(n5729) );
  AND2_X1 U6903 ( .A1(n5757), .A2(n5725), .ZN(n5726) );
  NOR2_X1 U6904 ( .A1(n5727), .A2(n5726), .ZN(n5978) );
  INV_X1 U6905 ( .A(n5978), .ZN(n5750) );
  NOR2_X1 U6906 ( .A1(n5750), .A2(n6362), .ZN(n5728) );
  AOI211_X1 U6907 ( .C1(n6081), .C2(REIP_REG_27__SCAN_IN), .A(n5729), .B(n5728), .ZN(n5732) );
  OR3_X1 U6908 ( .A1(n6080), .A2(REIP_REG_27__SCAN_IN), .A3(n5730), .ZN(n5731)
         );
  OAI211_X1 U6909 ( .C1(n5822), .C2(n6302), .A(n5732), .B(n5731), .ZN(U2800)
         );
  INV_X1 U6910 ( .A(n5734), .ZN(n5735) );
  AOI21_X1 U6911 ( .B1(n5736), .B2(n5807), .A(n5734), .ZN(n5935) );
  INV_X1 U6912 ( .A(n5935), .ZN(n5839) );
  NAND2_X1 U6913 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6243) );
  OAI21_X1 U6914 ( .B1(n6256), .B2(n6243), .A(n6913), .ZN(n5745) );
  NOR2_X1 U6915 ( .A1(n6259), .A2(n5737), .ZN(n6230) );
  INV_X1 U6916 ( .A(n5738), .ZN(n5933) );
  INV_X1 U6917 ( .A(n5796), .ZN(n5789) );
  AOI21_X1 U6918 ( .B1(n3221), .B2(n5739), .A(n5789), .ZN(n6182) );
  INV_X1 U6919 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5741) );
  OAI22_X1 U6920 ( .A1(n5741), .A2(n6331), .B1(n5740), .B2(n6354), .ZN(n5742)
         );
  AOI211_X1 U6921 ( .C1(n6182), .C2(n6322), .A(n6323), .B(n5742), .ZN(n5743)
         );
  OAI21_X1 U6922 ( .B1(n5933), .B2(n6343), .A(n5743), .ZN(n5744) );
  AOI21_X1 U6923 ( .B1(n5745), .B2(n6230), .A(n5744), .ZN(n5746) );
  OAI21_X1 U6924 ( .B1(n5839), .B2(n6302), .A(n5746), .ZN(U2810) );
  OAI22_X1 U6925 ( .A1(n5748), .A2(n6371), .B1(n6380), .B2(n5747), .ZN(U2828)
         );
  INV_X1 U6926 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5749) );
  OAI222_X1 U6927 ( .A1(n6152), .A2(n5858), .B1(n5749), .B2(n6380), .C1(n5968), 
        .C2(n6371), .ZN(U2831) );
  INV_X1 U6928 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5751) );
  OAI222_X1 U6929 ( .A1(n6152), .A2(n5822), .B1(n5751), .B2(n6380), .C1(n5750), 
        .C2(n6371), .ZN(U2832) );
  OR2_X1 U6930 ( .A1(n5752), .A2(n5753), .ZN(n5754) );
  AND2_X1 U6931 ( .A1(n5721), .A2(n5754), .ZN(n6086) );
  INV_X1 U6932 ( .A(n6086), .ZN(n5825) );
  NAND2_X1 U6933 ( .A1(n5765), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U6934 ( .A1(n5757), .A2(n5756), .ZN(n6082) );
  INV_X1 U6935 ( .A(n6082), .ZN(n5758) );
  AOI22_X1 U6936 ( .A1(n4474), .A2(n5758), .B1(EBX_REG_26__SCAN_IN), .B2(n5802), .ZN(n5759) );
  OAI21_X1 U6937 ( .B1(n5825), .B2(n6152), .A(n5759), .ZN(U2833) );
  NOR2_X1 U6938 ( .A1(n4681), .A2(n5760), .ZN(n5761) );
  OR2_X1 U6939 ( .A1(n5752), .A2(n5761), .ZN(n6093) );
  INV_X1 U6940 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U6941 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  NAND2_X1 U6942 ( .A1(n5765), .A2(n5764), .ZN(n6092) );
  OAI222_X1 U6943 ( .A1(n6093), .A2(n6152), .B1(n5766), .B2(n6380), .C1(n6371), 
        .C2(n6092), .ZN(U2834) );
  INV_X1 U6944 ( .A(n5767), .ZN(n5768) );
  AOI22_X1 U6945 ( .A1(n4474), .A2(n5768), .B1(EBX_REG_24__SCAN_IN), .B2(n5802), .ZN(n5769) );
  OAI21_X1 U6946 ( .B1(n5830), .B2(n6152), .A(n5769), .ZN(U2835) );
  NAND2_X1 U6947 ( .A1(n5770), .A2(n5771), .ZN(n5772) );
  NAND2_X1 U6948 ( .A1(n4682), .A2(n5772), .ZN(n6104) );
  NOR2_X1 U6949 ( .A1(n5780), .A2(n5773), .ZN(n5774) );
  OR2_X1 U6950 ( .A1(n5775), .A2(n5774), .ZN(n6004) );
  INV_X1 U6951 ( .A(n6004), .ZN(n6106) );
  AOI22_X1 U6952 ( .A1(n4474), .A2(n6106), .B1(EBX_REG_23__SCAN_IN), .B2(n5802), .ZN(n5776) );
  OAI21_X1 U6953 ( .B1(n6104), .B2(n6152), .A(n5776), .ZN(U2836) );
  OAI21_X1 U6954 ( .B1(n5777), .B2(n5778), .A(n5770), .ZN(n5897) );
  AND2_X1 U6955 ( .A1(n3212), .A2(n5779), .ZN(n5781) );
  OR2_X1 U6956 ( .A1(n5781), .A2(n5780), .ZN(n6120) );
  INV_X1 U6957 ( .A(n6120), .ZN(n5782) );
  AOI22_X1 U6958 ( .A1(n4474), .A2(n5782), .B1(EBX_REG_22__SCAN_IN), .B2(n5802), .ZN(n5783) );
  OAI21_X1 U6959 ( .B1(n5897), .B2(n6152), .A(n5783), .ZN(U2837) );
  AOI21_X1 U6960 ( .B1(n5785), .B2(n5784), .A(n3206), .ZN(n5786) );
  INV_X1 U6961 ( .A(n5786), .ZN(n6143) );
  NOR2_X1 U6962 ( .A1(n5787), .A2(n4385), .ZN(n5788) );
  AOI21_X1 U6963 ( .B1(n6029), .B2(n4385), .A(n5788), .ZN(n5797) );
  INV_X1 U6964 ( .A(n5797), .ZN(n5790) );
  NAND2_X1 U6965 ( .A1(n5790), .A2(n5789), .ZN(n5798) );
  XNOR2_X1 U6966 ( .A(n5798), .B(n5791), .ZN(n6142) );
  INV_X1 U6967 ( .A(n6142), .ZN(n5792) );
  AOI22_X1 U6968 ( .A1(n4474), .A2(n5792), .B1(EBX_REG_19__SCAN_IN), .B2(n5802), .ZN(n5793) );
  OAI21_X1 U6969 ( .B1(n6143), .B2(n6152), .A(n5793), .ZN(U2840) );
  NAND2_X1 U6970 ( .A1(n5735), .A2(n5794), .ZN(n5795) );
  INV_X1 U6971 ( .A(n6381), .ZN(n5801) );
  NAND2_X1 U6972 ( .A1(n5797), .A2(n5796), .ZN(n5799) );
  NAND2_X1 U6973 ( .A1(n5799), .A2(n5798), .ZN(n6237) );
  OAI222_X1 U6974 ( .A1(n5801), .A2(n6152), .B1(n5800), .B2(n6380), .C1(n6371), 
        .C2(n6237), .ZN(U2841) );
  AOI22_X1 U6975 ( .A1(n4474), .A2(n6182), .B1(EBX_REG_17__SCAN_IN), .B2(n5802), .ZN(n5803) );
  OAI21_X1 U6976 ( .B1(n5839), .B2(n6152), .A(n5803), .ZN(U2842) );
  OR2_X1 U6977 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  NAND2_X1 U6978 ( .A1(n5807), .A2(n5806), .ZN(n6238) );
  OR2_X1 U6979 ( .A1(n5808), .A2(n6064), .ZN(n5809) );
  NAND2_X1 U6980 ( .A1(n5809), .A2(n3221), .ZN(n6247) );
  OAI222_X1 U6981 ( .A1(n6238), .A2(n6152), .B1(n5810), .B2(n6380), .C1(n6247), 
        .C2(n6371), .ZN(U2843) );
  NAND3_X1 U6982 ( .A1(n5812), .A2(n5811), .A3(n6394), .ZN(n5814) );
  AOI22_X1 U6983 ( .A1(n6384), .A2(DATAI_31_), .B1(n6386), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U6984 ( .A1(n5814), .A2(n5813), .ZN(U2860) );
  AOI22_X1 U6985 ( .A1(n6384), .A2(DATAI_29_), .B1(n6386), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6986 ( .A1(n6387), .A2(DATAI_13_), .ZN(n5815) );
  OAI211_X1 U6987 ( .C1(n5817), .C2(n6156), .A(n5816), .B(n5815), .ZN(U2862)
         );
  AOI22_X1 U6988 ( .A1(n6384), .A2(DATAI_28_), .B1(n6386), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U6989 ( .A1(n6387), .A2(DATAI_12_), .ZN(n5818) );
  OAI211_X1 U6990 ( .C1(n5858), .C2(n6156), .A(n5819), .B(n5818), .ZN(U2863)
         );
  AOI22_X1 U6991 ( .A1(n6384), .A2(DATAI_27_), .B1(n6386), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U6992 ( .A1(n6387), .A2(DATAI_11_), .ZN(n5820) );
  OAI211_X1 U6993 ( .C1(n5822), .C2(n6156), .A(n5821), .B(n5820), .ZN(U2864)
         );
  AOI22_X1 U6994 ( .A1(n6387), .A2(DATAI_10_), .B1(n6386), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U6995 ( .A1(n6384), .A2(DATAI_26_), .ZN(n5823) );
  OAI211_X1 U6996 ( .C1(n5825), .C2(n6156), .A(n5824), .B(n5823), .ZN(U2865)
         );
  AOI22_X1 U6997 ( .A1(n6387), .A2(DATAI_9_), .B1(n6386), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6998 ( .A1(n6384), .A2(DATAI_25_), .ZN(n5826) );
  OAI211_X1 U6999 ( .C1(n6093), .C2(n6156), .A(n5827), .B(n5826), .ZN(U2866)
         );
  AOI22_X1 U7000 ( .A1(n6387), .A2(DATAI_8_), .B1(n6386), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7001 ( .A1(n6384), .A2(DATAI_24_), .ZN(n5828) );
  OAI211_X1 U7002 ( .C1(n5830), .C2(n6156), .A(n5829), .B(n5828), .ZN(U2867)
         );
  AOI22_X1 U7003 ( .A1(n6387), .A2(DATAI_7_), .B1(n6386), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7004 ( .A1(n6384), .A2(DATAI_23_), .ZN(n5831) );
  OAI211_X1 U7005 ( .C1(n6104), .C2(n6156), .A(n5832), .B(n5831), .ZN(U2868)
         );
  AOI22_X1 U7006 ( .A1(n6387), .A2(DATAI_6_), .B1(n6386), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7007 ( .A1(n6384), .A2(DATAI_22_), .ZN(n5833) );
  OAI211_X1 U7008 ( .C1(n5897), .C2(n6156), .A(n5834), .B(n5833), .ZN(U2869)
         );
  AOI22_X1 U7009 ( .A1(n6387), .A2(DATAI_3_), .B1(n6386), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7010 ( .A1(n6384), .A2(DATAI_19_), .ZN(n5835) );
  OAI211_X1 U7011 ( .C1(n6143), .C2(n6156), .A(n5836), .B(n5835), .ZN(U2872)
         );
  AOI22_X1 U7012 ( .A1(n6384), .A2(DATAI_17_), .B1(n6386), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7013 ( .A1(n6387), .A2(DATAI_1_), .ZN(n5837) );
  OAI211_X1 U7014 ( .C1(n5839), .C2(n6156), .A(n5838), .B(n5837), .ZN(U2874)
         );
  XOR2_X1 U7015 ( .A(n5840), .B(n5564), .Z(n6365) );
  INV_X1 U7016 ( .A(n6365), .ZN(n5842) );
  AOI22_X1 U7017 ( .A1(n6390), .A2(DATAI_15_), .B1(n6386), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5841) );
  OAI21_X1 U7018 ( .B1(n5842), .B2(n6156), .A(n5841), .ZN(U2876) );
  NOR2_X1 U7019 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  XNOR2_X1 U7020 ( .A(n5845), .B(n5958), .ZN(n5967) );
  NAND2_X1 U7021 ( .A1(n6567), .A2(REIP_REG_29__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7022 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5846)
         );
  OAI211_X1 U7023 ( .C1(n5847), .C2(n6466), .A(n5961), .B(n5846), .ZN(n5848)
         );
  AOI21_X1 U7024 ( .B1(n5849), .B2(n6461), .A(n5848), .ZN(n5850) );
  OAI21_X1 U7025 ( .B1(n5967), .B2(n6468), .A(n5850), .ZN(U2957) );
  NAND3_X1 U7026 ( .A1(n5851), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n3203), .ZN(n5856) );
  INV_X1 U7027 ( .A(n5852), .ZN(n5854) );
  NAND2_X1 U7028 ( .A1(n5997), .A2(n5855), .ZN(n5989) );
  NOR2_X1 U7029 ( .A1(n3204), .A2(n5989), .ZN(n5853) );
  NAND2_X1 U7030 ( .A1(n5854), .A2(n5853), .ZN(n5864) );
  XNOR2_X1 U7031 ( .A(n5857), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5976)
         );
  INV_X1 U7032 ( .A(n5858), .ZN(n5862) );
  NOR2_X1 U7033 ( .A1(n6556), .A2(n6928), .ZN(n5970) );
  AOI21_X1 U7034 ( .B1(n6456), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5970), 
        .ZN(n5859) );
  OAI21_X1 U7035 ( .B1(n5860), .B2(n6466), .A(n5859), .ZN(n5861) );
  AOI21_X1 U7036 ( .B1(n5862), .B2(n6461), .A(n5861), .ZN(n5863) );
  OAI21_X1 U7037 ( .B1(n5976), .B2(n6468), .A(n5863), .ZN(U2958) );
  NAND2_X1 U7038 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  XNOR2_X1 U7039 ( .A(n5866), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5985)
         );
  INV_X1 U7040 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U7041 ( .A1(n6556), .A2(n6925), .ZN(n5977) );
  NOR2_X1 U7042 ( .A1(n6474), .A2(n5867), .ZN(n5868) );
  AOI211_X1 U7043 ( .C1(n5869), .C2(n6438), .A(n5977), .B(n5868), .ZN(n5872)
         );
  NAND2_X1 U7044 ( .A1(n5870), .A2(n6461), .ZN(n5871) );
  OAI211_X1 U7045 ( .C1(n5985), .C2(n6468), .A(n5872), .B(n5871), .ZN(U2959)
         );
  XNOR2_X1 U7046 ( .A(n3204), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5873)
         );
  XNOR2_X1 U7047 ( .A(n5851), .B(n5873), .ZN(n5993) );
  AND2_X1 U7048 ( .A1(n6567), .A2(REIP_REG_26__SCAN_IN), .ZN(n5987) );
  AOI21_X1 U7049 ( .B1(n6456), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5987), 
        .ZN(n5874) );
  OAI21_X1 U7050 ( .B1(n6089), .B2(n6466), .A(n5874), .ZN(n5875) );
  AOI21_X1 U7051 ( .B1(n6086), .B2(n6461), .A(n5875), .ZN(n5876) );
  OAI21_X1 U7052 ( .B1(n5993), .B2(n6468), .A(n5876), .ZN(U2960) );
  AOI21_X1 U7053 ( .B1(n5879), .B2(n5878), .A(n3196), .ZN(n6001) );
  NAND2_X1 U7054 ( .A1(n6567), .A2(REIP_REG_25__SCAN_IN), .ZN(n5994) );
  OAI21_X1 U7055 ( .B1(n6474), .B2(n5880), .A(n5994), .ZN(n5882) );
  NOR2_X1 U7056 ( .A1(n6093), .A2(n6470), .ZN(n5881) );
  AOI211_X1 U7057 ( .C1(n6438), .C2(n6091), .A(n5882), .B(n5881), .ZN(n5883)
         );
  OAI21_X1 U7058 ( .B1(n6001), .B2(n6468), .A(n5883), .ZN(U2961) );
  INV_X1 U7059 ( .A(n6037), .ZN(n5885) );
  INV_X1 U7060 ( .A(n6013), .ZN(n5884) );
  NOR4_X1 U7061 ( .A1(n5886), .A2(n4555), .A3(n5885), .A4(n5884), .ZN(n5887)
         );
  NOR2_X1 U7062 ( .A1(n5888), .A2(n5887), .ZN(n5890) );
  XNOR2_X1 U7063 ( .A(n5890), .B(n5889), .ZN(n6010) );
  NAND2_X1 U7064 ( .A1(n6567), .A2(REIP_REG_23__SCAN_IN), .ZN(n6003) );
  OAI21_X1 U7065 ( .B1(n6474), .B2(n7299), .A(n6003), .ZN(n5892) );
  NOR2_X1 U7066 ( .A1(n6104), .A2(n6470), .ZN(n5891) );
  AOI211_X1 U7067 ( .C1(n6438), .C2(n6101), .A(n5892), .B(n5891), .ZN(n5893)
         );
  OAI21_X1 U7068 ( .B1(n6010), .B2(n6468), .A(n5893), .ZN(U2963) );
  OAI21_X1 U7069 ( .B1(n4555), .B2(n7269), .A(n5894), .ZN(n5896) );
  XOR2_X1 U7070 ( .A(n5896), .B(n5895), .Z(n6018) );
  INV_X1 U7071 ( .A(n5897), .ZN(n6115) );
  NAND2_X1 U7072 ( .A1(n6567), .A2(REIP_REG_22__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7073 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5898)
         );
  OAI211_X1 U7074 ( .C1(n5899), .C2(n6466), .A(n6011), .B(n5898), .ZN(n5900)
         );
  AOI21_X1 U7075 ( .B1(n6115), .B2(n6461), .A(n5900), .ZN(n5901) );
  OAI21_X1 U7076 ( .B1(n6018), .B2(n6468), .A(n5901), .ZN(U2964) );
  XNOR2_X1 U7077 ( .A(n5902), .B(n5903), .ZN(n6127) );
  OAI21_X1 U7078 ( .B1(n5906), .B2(n5905), .A(n5904), .ZN(n6019) );
  NAND2_X1 U7079 ( .A1(n6019), .A2(n6460), .ZN(n5909) );
  NAND2_X1 U7080 ( .A1(n6567), .A2(REIP_REG_21__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U7081 ( .B1(n6474), .B2(n6123), .A(n6022), .ZN(n5907) );
  AOI21_X1 U7082 ( .B1(n6121), .B2(n6438), .A(n5907), .ZN(n5908) );
  OAI211_X1 U7083 ( .C1(n6470), .C2(n6127), .A(n5909), .B(n5908), .ZN(U2965)
         );
  XNOR2_X1 U7084 ( .A(n3203), .B(n5910), .ZN(n5911) );
  XNOR2_X1 U7085 ( .A(n5912), .B(n5911), .ZN(n6042) );
  NOR2_X1 U7086 ( .A1(n3206), .A2(n5913), .ZN(n5914) );
  OR2_X1 U7087 ( .A1(n5902), .A2(n5914), .ZN(n6153) );
  INV_X1 U7088 ( .A(n6153), .ZN(n6160) );
  NAND2_X1 U7089 ( .A1(n6567), .A2(REIP_REG_20__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7090 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5915)
         );
  OAI211_X1 U7091 ( .C1(n6131), .C2(n6466), .A(n6035), .B(n5915), .ZN(n5916)
         );
  AOI21_X1 U7092 ( .B1(n6160), .B2(n6461), .A(n5916), .ZN(n5917) );
  OAI21_X1 U7093 ( .B1(n6042), .B2(n6468), .A(n5917), .ZN(U2966) );
  INV_X1 U7094 ( .A(n5918), .ZN(n6044) );
  NAND2_X1 U7095 ( .A1(n5920), .A2(n5919), .ZN(n6043) );
  NAND3_X1 U7096 ( .A1(n6044), .A2(n6460), .A3(n6043), .ZN(n5923) );
  NAND2_X1 U7097 ( .A1(n6567), .A2(REIP_REG_19__SCAN_IN), .ZN(n6045) );
  OAI21_X1 U7098 ( .B1(n6474), .B2(n6141), .A(n6045), .ZN(n5921) );
  AOI21_X1 U7099 ( .B1(n6139), .B2(n6438), .A(n5921), .ZN(n5922) );
  OAI211_X1 U7100 ( .C1(n6470), .C2(n6143), .A(n5923), .B(n5922), .ZN(U2967)
         );
  NAND3_X1 U7101 ( .A1(n5924), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n3203), .ZN(n6052) );
  INV_X1 U7102 ( .A(n6052), .ZN(n5931) );
  NAND2_X1 U7103 ( .A1(n4555), .A2(n7215), .ZN(n5926) );
  NOR2_X1 U7104 ( .A1(n3203), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5929)
         );
  INV_X1 U7105 ( .A(n5929), .ZN(n5938) );
  AOI22_X1 U7106 ( .A1(n5924), .A2(n5926), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5938), .ZN(n5930) );
  INV_X1 U7107 ( .A(n5928), .ZN(n5946) );
  NAND3_X1 U7108 ( .A1(n5946), .A2(n5929), .A3(n7215), .ZN(n6051) );
  OAI21_X1 U7109 ( .B1(n5931), .B2(n5930), .A(n6051), .ZN(n6183) );
  INV_X1 U7110 ( .A(n6183), .ZN(n5937) );
  AOI22_X1 U7111 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n6567), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5932) );
  OAI21_X1 U7112 ( .B1(n5933), .B2(n6466), .A(n5932), .ZN(n5934) );
  AOI21_X1 U7113 ( .B1(n5935), .B2(n6461), .A(n5934), .ZN(n5936) );
  OAI21_X1 U7114 ( .B1(n5937), .B2(n6468), .A(n5936), .ZN(U2969) );
  OAI21_X1 U7115 ( .B1(n4555), .B2(n7164), .A(n5938), .ZN(n5939) );
  XNOR2_X1 U7116 ( .A(n3220), .B(n5939), .ZN(n6187) );
  INV_X1 U7117 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5940) );
  OAI22_X1 U7118 ( .A1(n6474), .A2(n5941), .B1(n6556), .B2(n5940), .ZN(n5943)
         );
  NOR2_X1 U7119 ( .A1(n6238), .A2(n6470), .ZN(n5942) );
  AOI211_X1 U7120 ( .C1(n6438), .C2(n6239), .A(n5943), .B(n5942), .ZN(n5944)
         );
  OAI21_X1 U7121 ( .B1(n6187), .B2(n6468), .A(n5944), .ZN(U2970) );
  AOI21_X1 U7122 ( .B1(n5947), .B2(n5945), .A(n5946), .ZN(n6072) );
  NAND2_X1 U7123 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5948)
         );
  NAND2_X1 U7124 ( .A1(n6567), .A2(REIP_REG_15__SCAN_IN), .ZN(n6066) );
  OAI211_X1 U7125 ( .C1(n6466), .C2(n6252), .A(n5948), .B(n6066), .ZN(n5949)
         );
  AOI21_X1 U7126 ( .B1(n6365), .B2(n6461), .A(n5949), .ZN(n5950) );
  OAI21_X1 U7127 ( .B1(n6072), .B2(n6468), .A(n5950), .ZN(U2971) );
  INV_X1 U7128 ( .A(n5951), .ZN(n5955) );
  AOI22_X1 U7129 ( .A1(n6456), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6567), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5952) );
  OAI21_X1 U7130 ( .B1(n5953), .B2(n6466), .A(n5952), .ZN(n5954) );
  AOI21_X1 U7131 ( .B1(n5955), .B2(n6461), .A(n5954), .ZN(n5956) );
  OAI21_X1 U7132 ( .B1(n5957), .B2(n6468), .A(n5956), .ZN(U2972) );
  OAI21_X1 U7133 ( .B1(n5959), .B2(n5972), .A(n5958), .ZN(n5965) );
  INV_X1 U7134 ( .A(n5960), .ZN(n5964) );
  OAI21_X1 U7135 ( .B1(n5962), .B2(n6551), .A(n5961), .ZN(n5963) );
  AOI21_X1 U7136 ( .B1(n5965), .B2(n5964), .A(n5963), .ZN(n5966) );
  OAI21_X1 U7137 ( .B1(n5967), .B2(n6478), .A(n5966), .ZN(U2989) );
  NOR2_X1 U7138 ( .A1(n5968), .A2(n6551), .ZN(n5969) );
  AOI211_X1 U7139 ( .C1(n5971), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5970), .B(n5969), .ZN(n5975) );
  NAND3_X1 U7140 ( .A1(n5983), .A2(n5973), .A3(n5972), .ZN(n5974) );
  OAI211_X1 U7141 ( .C1(n5976), .C2(n6478), .A(n5975), .B(n5974), .ZN(U2990)
         );
  AOI21_X1 U7142 ( .B1(n5978), .B2(n6569), .A(n5977), .ZN(n5979) );
  OAI21_X1 U7143 ( .B1(n5980), .B2(n5982), .A(n5979), .ZN(n5981) );
  AOI21_X1 U7144 ( .B1(n5983), .B2(n5982), .A(n5981), .ZN(n5984) );
  OAI21_X1 U7145 ( .B1(n5985), .B2(n6478), .A(n5984), .ZN(U2991) );
  NOR2_X1 U7146 ( .A1(n6082), .A2(n6551), .ZN(n5986) );
  AOI211_X1 U7147 ( .C1(n5996), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5987), .B(n5986), .ZN(n5992) );
  INV_X1 U7148 ( .A(n5988), .ZN(n5998) );
  NAND3_X1 U7149 ( .A1(n5998), .A2(n5990), .A3(n5989), .ZN(n5991) );
  OAI211_X1 U7150 ( .C1(n5993), .C2(n6478), .A(n5992), .B(n5991), .ZN(U2992)
         );
  OAI21_X1 U7151 ( .B1(n6092), .B2(n6551), .A(n5994), .ZN(n5995) );
  AOI21_X1 U7152 ( .B1(n5996), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5995), 
        .ZN(n6000) );
  NAND2_X1 U7153 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  OAI211_X1 U7154 ( .C1(n6001), .C2(n6478), .A(n6000), .B(n5999), .ZN(U2993)
         );
  INV_X1 U7155 ( .A(n6002), .ZN(n6006) );
  OAI21_X1 U7156 ( .B1(n6551), .B2(n6004), .A(n6003), .ZN(n6005) );
  AOI21_X1 U7157 ( .B1(n6006), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6005), 
        .ZN(n6009) );
  OR2_X1 U7158 ( .A1(n6007), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6008)
         );
  OAI211_X1 U7159 ( .C1(n6010), .C2(n6478), .A(n6009), .B(n6008), .ZN(U2995)
         );
  OAI21_X1 U7160 ( .B1(n6551), .B2(n6120), .A(n6011), .ZN(n6016) );
  INV_X1 U7161 ( .A(n6012), .ZN(n6027) );
  NOR3_X1 U7162 ( .A1(n6027), .A2(n6014), .A3(n6013), .ZN(n6015) );
  AOI211_X1 U7163 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n6024), .A(n6016), .B(n6015), .ZN(n6017) );
  OAI21_X1 U7164 ( .B1(n6018), .B2(n6478), .A(n6017), .ZN(U2996) );
  NAND2_X1 U7165 ( .A1(n6019), .A2(n6571), .ZN(n6026) );
  NAND2_X1 U7166 ( .A1(n3230), .A2(n6020), .ZN(n6021) );
  NAND2_X1 U7167 ( .A1(n3212), .A2(n6021), .ZN(n6128) );
  OAI21_X1 U7168 ( .B1(n6551), .B2(n6128), .A(n6022), .ZN(n6023) );
  AOI21_X1 U7169 ( .B1(n6024), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6023), 
        .ZN(n6025) );
  OAI211_X1 U7170 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n6027), .A(n6026), .B(n6025), .ZN(U2997) );
  OAI21_X1 U7171 ( .B1(n6028), .B2(n6518), .A(n6186), .ZN(n6047) );
  NAND2_X1 U7172 ( .A1(n6031), .A2(n6029), .ZN(n6030) );
  OAI21_X1 U7173 ( .B1(n6031), .B2(n4385), .A(n6030), .ZN(n6034) );
  INV_X1 U7174 ( .A(n6032), .ZN(n6033) );
  XNOR2_X1 U7175 ( .A(n6034), .B(n6033), .ZN(n6151) );
  OAI21_X1 U7176 ( .B1(n6551), .B2(n6151), .A(n6035), .ZN(n6040) );
  NAND2_X1 U7177 ( .A1(n6056), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6036) );
  OR2_X1 U7178 ( .A1(n6069), .A2(n6036), .ZN(n6050) );
  NOR3_X1 U7179 ( .A1(n6050), .A2(n6038), .A3(n6037), .ZN(n6039) );
  AOI211_X1 U7180 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6047), .A(n6040), .B(n6039), .ZN(n6041) );
  OAI21_X1 U7181 ( .B1(n6042), .B2(n6478), .A(n6041), .ZN(U2998) );
  NAND3_X1 U7182 ( .A1(n6044), .A2(n6571), .A3(n6043), .ZN(n6049) );
  OAI21_X1 U7183 ( .B1(n6551), .B2(n6142), .A(n6045), .ZN(n6046) );
  AOI21_X1 U7184 ( .B1(n6047), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6046), 
        .ZN(n6048) );
  OAI211_X1 U7185 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6050), .A(n6049), .B(n6048), .ZN(U2999) );
  NAND2_X1 U7186 ( .A1(n6052), .A2(n6051), .ZN(n6054) );
  XNOR2_X1 U7187 ( .A(n6054), .B(n6053), .ZN(n6163) );
  OAI21_X1 U7188 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6055), .A(n6186), 
        .ZN(n6058) );
  AND2_X1 U7189 ( .A1(n6197), .A2(n6056), .ZN(n6057) );
  AOI22_X1 U7190 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6058), .B1(n6053), .B2(n6057), .ZN(n6060) );
  NAND2_X1 U7191 ( .A1(n6567), .A2(REIP_REG_18__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7192 ( .C1(n6551), .C2(n6237), .A(n6060), .B(n6059), .ZN(n6061)
         );
  AOI21_X1 U7193 ( .B1(n6163), .B2(n6571), .A(n6061), .ZN(n6062) );
  INV_X1 U7194 ( .A(n6062), .ZN(U3000) );
  INV_X1 U7195 ( .A(n6068), .ZN(n6063) );
  OAI21_X1 U7196 ( .B1(n6518), .B2(n6063), .A(n6476), .ZN(n6189) );
  AOI21_X1 U7197 ( .B1(n6065), .B2(n3231), .A(n6064), .ZN(n6364) );
  INV_X1 U7198 ( .A(n6364), .ZN(n6067) );
  OAI21_X1 U7199 ( .B1(n6551), .B2(n6067), .A(n6066), .ZN(n6070) );
  NOR3_X1 U7200 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6069), .A3(n6068), 
        .ZN(n6190) );
  AOI211_X1 U7201 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6189), .A(n6070), .B(n6190), .ZN(n6071) );
  OAI21_X1 U7202 ( .B1(n6072), .B2(n6478), .A(n6071), .ZN(U3003) );
  OAI21_X1 U7203 ( .B1(n6073), .B2(STATEBS16_REG_SCAN_IN), .A(n6753), .ZN(
        n6075) );
  OAI22_X1 U7204 ( .A1(n6075), .A2(n6744), .B1(n6074), .B2(n6077), .ZN(n6076)
         );
  MUX2_X1 U7205 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6076), .S(n6577), 
        .Z(U3464) );
  XNOR2_X1 U7206 ( .A(n6580), .B(n6744), .ZN(n6078) );
  OAI22_X1 U7207 ( .A1(n6078), .A2(n6658), .B1(n4755), .B2(n6077), .ZN(n6079)
         );
  MUX2_X1 U7208 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6079), .S(n6577), 
        .Z(U3463) );
  AOI22_X1 U7209 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6346), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6332), .ZN(n6088) );
  NOR2_X1 U7210 ( .A1(n6921), .A2(n6080), .ZN(n6090) );
  AOI21_X1 U7211 ( .B1(REIP_REG_25__SCAN_IN), .B2(n6090), .A(
        REIP_REG_26__SCAN_IN), .ZN(n6084) );
  INV_X1 U7212 ( .A(n6081), .ZN(n6083) );
  OAI22_X1 U7213 ( .A1(n6084), .A2(n6083), .B1(n6082), .B2(n6362), .ZN(n6085)
         );
  AOI21_X1 U7214 ( .B1(n6086), .B2(n6315), .A(n6085), .ZN(n6087) );
  OAI211_X1 U7215 ( .C1(n6089), .C2(n6343), .A(n6088), .B(n6087), .ZN(U2801)
         );
  INV_X1 U7216 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6923) );
  AOI22_X1 U7217 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6332), .B1(n6090), 
        .B2(n6923), .ZN(n6100) );
  AOI22_X1 U7218 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6346), .B1(n6091), .B2(n6357), .ZN(n6099) );
  OAI22_X1 U7219 ( .A1(n6093), .A2(n6302), .B1(n6362), .B2(n6092), .ZN(n6094)
         );
  INV_X1 U7220 ( .A(n6094), .ZN(n6098) );
  INV_X1 U7221 ( .A(n6103), .ZN(n6095) );
  OAI21_X1 U7222 ( .B1(n6096), .B2(n6095), .A(REIP_REG_25__SCAN_IN), .ZN(n6097) );
  NAND4_X1 U7223 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(U2802)
         );
  AOI22_X1 U7224 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6332), .B1(n6101), 
        .B2(n6357), .ZN(n6108) );
  INV_X1 U7225 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7203) );
  INV_X1 U7226 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U7227 ( .A1(n7203), .A2(n6918), .ZN(n6116) );
  AOI21_X1 U7228 ( .B1(n6125), .B2(n6116), .A(REIP_REG_23__SCAN_IN), .ZN(n6102) );
  OAI22_X1 U7229 ( .A1(n6104), .A2(n6302), .B1(n6103), .B2(n6102), .ZN(n6105)
         );
  AOI21_X1 U7230 ( .B1(n6106), .B2(n6322), .A(n6105), .ZN(n6107) );
  OAI211_X1 U7231 ( .C1(n6109), .C2(n6331), .A(n6108), .B(n6107), .ZN(U2804)
         );
  OAI22_X1 U7232 ( .A1(n6354), .A2(n4086), .B1(n6110), .B2(n6331), .ZN(n6111)
         );
  AOI21_X1 U7233 ( .B1(n6357), .B2(n6112), .A(n6111), .ZN(n6113) );
  OAI21_X1 U7234 ( .B1(n6137), .B2(n7203), .A(n6113), .ZN(n6114) );
  AOI21_X1 U7235 ( .B1(n6115), .B2(n6315), .A(n6114), .ZN(n6119) );
  INV_X1 U7236 ( .A(n6116), .ZN(n6117) );
  OAI211_X1 U7237 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n6125), .B(n6117), .ZN(n6118) );
  OAI211_X1 U7238 ( .C1(n6362), .C2(n6120), .A(n6119), .B(n6118), .ZN(U2805)
         );
  INV_X1 U7239 ( .A(n6137), .ZN(n6126) );
  AOI22_X1 U7240 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6346), .B1(n6121), .B2(n6357), .ZN(n6122) );
  OAI21_X1 U7241 ( .B1(n6123), .B2(n6354), .A(n6122), .ZN(n6124) );
  AOI221_X1 U7242 ( .B1(n6126), .B2(REIP_REG_21__SCAN_IN), .C1(n6125), .C2(
        n6918), .A(n6124), .ZN(n6130) );
  INV_X1 U7243 ( .A(n6127), .ZN(n6157) );
  INV_X1 U7244 ( .A(n6128), .ZN(n6149) );
  AOI22_X1 U7245 ( .A1(n6157), .A2(n6315), .B1(n6149), .B2(n6322), .ZN(n6129)
         );
  NAND2_X1 U7246 ( .A1(n6130), .A2(n6129), .ZN(U2806) );
  NOR2_X1 U7247 ( .A1(n6914), .A2(n6915), .ZN(n6148) );
  AOI21_X1 U7248 ( .B1(n6234), .B2(n6148), .A(REIP_REG_20__SCAN_IN), .ZN(n6138) );
  INV_X1 U7249 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6132) );
  OAI22_X1 U7250 ( .A1(n6132), .A2(n6354), .B1(n6131), .B2(n6343), .ZN(n6133)
         );
  AOI21_X1 U7251 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6346), .A(n6133), .ZN(n6136)
         );
  OAI22_X1 U7252 ( .A1(n6153), .A2(n6302), .B1(n6151), .B2(n6362), .ZN(n6134)
         );
  INV_X1 U7253 ( .A(n6134), .ZN(n6135) );
  OAI211_X1 U7254 ( .C1(n6138), .C2(n6137), .A(n6136), .B(n6135), .ZN(U2807)
         );
  OAI21_X1 U7255 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n6234), .ZN(n6147) );
  AOI22_X1 U7256 ( .A1(n6139), .A2(n6357), .B1(REIP_REG_19__SCAN_IN), .B2(
        n6230), .ZN(n6140) );
  OAI211_X1 U7257 ( .C1(n6354), .C2(n6141), .A(n6140), .B(n6312), .ZN(n6145)
         );
  OAI22_X1 U7258 ( .A1(n6143), .A2(n6302), .B1(n6142), .B2(n6362), .ZN(n6144)
         );
  AOI211_X1 U7259 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6346), .A(n6145), .B(n6144), 
        .ZN(n6146) );
  OAI21_X1 U7260 ( .B1(n6148), .B2(n6147), .A(n6146), .ZN(U2808) );
  INV_X1 U7261 ( .A(EBX_REG_21__SCAN_IN), .ZN(n7280) );
  AOI22_X1 U7262 ( .A1(n6157), .A2(n4359), .B1(n6149), .B2(n4474), .ZN(n6150)
         );
  OAI21_X1 U7263 ( .B1(n6380), .B2(n7280), .A(n6150), .ZN(U2838) );
  OAI22_X1 U7264 ( .A1(n6153), .A2(n6152), .B1(n6151), .B2(n6371), .ZN(n6154)
         );
  INV_X1 U7265 ( .A(n6154), .ZN(n6155) );
  OAI21_X1 U7266 ( .B1(n6380), .B2(n4432), .A(n6155), .ZN(U2839) );
  INV_X1 U7267 ( .A(n6156), .ZN(n6391) );
  AOI22_X1 U7268 ( .A1(n6157), .A2(n6391), .B1(n6384), .B2(DATAI_21_), .ZN(
        n6159) );
  AOI22_X1 U7269 ( .A1(n6387), .A2(DATAI_5_), .B1(n6386), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7270 ( .A1(n6159), .A2(n6158), .ZN(U2870) );
  AOI22_X1 U7271 ( .A1(n6160), .A2(n6391), .B1(n6384), .B2(DATAI_20_), .ZN(
        n6162) );
  AOI22_X1 U7272 ( .A1(n6387), .A2(DATAI_4_), .B1(n6386), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7273 ( .A1(n6162), .A2(n6161), .ZN(U2871) );
  AOI22_X1 U7274 ( .A1(n6567), .A2(REIP_REG_18__SCAN_IN), .B1(n6456), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6165) );
  AOI22_X1 U7275 ( .A1(n6163), .A2(n6460), .B1(n6461), .B2(n6381), .ZN(n6164)
         );
  OAI211_X1 U7276 ( .C1(n6466), .C2(n6232), .A(n6165), .B(n6164), .ZN(U2968)
         );
  AOI22_X1 U7277 ( .A1(n6567), .A2(REIP_REG_13__SCAN_IN), .B1(n6456), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7278 ( .A(n6166), .B(n6167), .ZN(n6199) );
  AND2_X1 U7279 ( .A1(n6169), .A2(n6168), .ZN(n6173) );
  AND2_X1 U7280 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  NOR2_X1 U7281 ( .A1(n6173), .A2(n6172), .ZN(n6175) );
  NAND2_X1 U7282 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  AND2_X1 U7283 ( .A1(n6177), .A2(n6176), .ZN(n6392) );
  AOI22_X1 U7284 ( .A1(n6199), .A2(n6460), .B1(n6461), .B2(n6392), .ZN(n6178)
         );
  OAI211_X1 U7285 ( .C1(n6466), .C2(n6267), .A(n6179), .B(n6178), .ZN(U2973)
         );
  NOR2_X1 U7286 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6180), .ZN(n6181)
         );
  AOI22_X1 U7287 ( .A1(n6567), .A2(REIP_REG_17__SCAN_IN), .B1(n6181), .B2(
        n6197), .ZN(n6185) );
  AOI22_X1 U7288 ( .A1(n6183), .A2(n6571), .B1(n6569), .B2(n6182), .ZN(n6184)
         );
  OAI211_X1 U7289 ( .C1(n6186), .C2(n7215), .A(n6185), .B(n6184), .ZN(U3001)
         );
  OAI22_X1 U7290 ( .A1(n6187), .A2(n6478), .B1(n6551), .B2(n6247), .ZN(n6188)
         );
  AOI221_X1 U7291 ( .B1(n6190), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        n6189), .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6188), .ZN(n6193) );
  NAND3_X1 U7292 ( .A1(n6191), .A2(n7164), .A3(n6197), .ZN(n6192) );
  OAI211_X1 U7293 ( .C1(n5940), .C2(n6556), .A(n6193), .B(n6192), .ZN(U3002)
         );
  AOI21_X1 U7294 ( .B1(n6196), .B2(n6195), .A(n6194), .ZN(n6367) );
  AOI22_X1 U7295 ( .A1(n6569), .A2(n6367), .B1(n6567), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n6201) );
  AOI22_X1 U7296 ( .A1(n6199), .A2(n6571), .B1(n6198), .B2(n6197), .ZN(n6200)
         );
  OAI211_X1 U7297 ( .C1(n6202), .C2(n4562), .A(n6201), .B(n6200), .ZN(U3005)
         );
  INV_X1 U7298 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6888) );
  AOI21_X1 U7299 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6888), .A(n4652), .ZN(n6211) );
  INV_X1 U7300 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6203) );
  AOI21_X1 U7301 ( .B1(n6211), .B2(n6203), .A(n3194), .ZN(U2789) );
  INV_X1 U7302 ( .A(n6868), .ZN(n6209) );
  OAI21_X1 U7303 ( .B1(n6207), .B2(n3530), .A(n6206), .ZN(n6216) );
  OAI21_X1 U7304 ( .B1(n6216), .B2(n6865), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6208) );
  OAI21_X1 U7305 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6209), .A(n6208), .ZN(
        U2790) );
  NOR2_X1 U7306 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6212) );
  OAI21_X1 U7307 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6212), .A(n6936), .ZN(n6210)
         );
  OAI21_X1 U7308 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6974), .A(n6210), .ZN(
        U2791) );
  NOR2_X1 U7309 ( .A1(n3194), .A2(n6211), .ZN(n6942) );
  OAI21_X1 U7310 ( .B1(BS16_N), .B2(n6212), .A(n6942), .ZN(n6940) );
  OAI21_X1 U7311 ( .B1(n6942), .B2(n6213), .A(n6940), .ZN(U2792) );
  AOI21_X1 U7312 ( .B1(n6215), .B2(n6214), .A(READY_N), .ZN(n6983) );
  NOR2_X1 U7313 ( .A1(n6216), .A2(n6983), .ZN(n6815) );
  NOR2_X1 U7314 ( .A1(n6815), .A2(n6865), .ZN(n6978) );
  OAI21_X1 U7315 ( .B1(n6978), .B2(n6217), .A(n6468), .ZN(U2793) );
  NOR4_X1 U7316 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6227) );
  AOI211_X1 U7317 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_3__SCAN_IN), .B(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6226) );
  NOR4_X1 U7318 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n6218) );
  INV_X1 U7319 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7246) );
  INV_X1 U7320 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n7307) );
  NAND3_X1 U7321 ( .A1(n6218), .A2(n7246), .A3(n7307), .ZN(n6224) );
  NOR4_X1 U7322 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6222) );
  NOR4_X1 U7323 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6221) );
  NOR4_X1 U7324 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6220) );
  NOR4_X1 U7325 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6219) );
  NAND4_X1 U7326 ( .A1(n6222), .A2(n6221), .A3(n6220), .A4(n6219), .ZN(n6223)
         );
  NOR4_X1 U7327 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(n6224), .A4(n6223), .ZN(n6225) );
  NAND3_X1 U7328 ( .A1(n6227), .A2(n6226), .A3(n6225), .ZN(n6966) );
  NOR2_X1 U7329 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6966), .ZN(n6963) );
  INV_X1 U7330 ( .A(n6966), .ZN(n6971) );
  INV_X1 U7331 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6964) );
  INV_X1 U7332 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6968) );
  INV_X1 U7333 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6941) );
  NAND4_X1 U7334 ( .A1(n6971), .A2(n6964), .A3(n6968), .A4(n6941), .ZN(n6228)
         );
  INV_X1 U7335 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7252) );
  AOI22_X1 U7336 ( .A1(n6963), .A2(n6228), .B1(n7252), .B2(n6966), .ZN(U2794)
         );
  INV_X1 U7337 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7338 ( .A1(n6963), .A2(n6941), .ZN(n6969) );
  OAI211_X1 U7339 ( .C1(n6971), .C2(n6229), .A(n6228), .B(n6969), .ZN(U2795)
         );
  AOI22_X1 U7340 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6346), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6230), .ZN(n6231) );
  OAI21_X1 U7341 ( .B1(n6232), .B2(n6343), .A(n6231), .ZN(n6233) );
  AOI211_X1 U7342 ( .C1(n6332), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6323), 
        .B(n6233), .ZN(n6236) );
  AOI22_X1 U7343 ( .A1(n6381), .A2(n6315), .B1(n6915), .B2(n6234), .ZN(n6235)
         );
  OAI211_X1 U7344 ( .C1(n6362), .C2(n6237), .A(n6236), .B(n6235), .ZN(U2809)
         );
  INV_X1 U7345 ( .A(n6238), .ZN(n6385) );
  AOI21_X1 U7346 ( .B1(n6332), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6323), 
        .ZN(n6241) );
  AOI22_X1 U7347 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6346), .B1(n6239), .B2(n6357), .ZN(n6240) );
  OAI211_X1 U7348 ( .C1(n5940), .C2(n6249), .A(n6241), .B(n6240), .ZN(n6242)
         );
  AOI21_X1 U7349 ( .B1(n6385), .B2(n6315), .A(n6242), .ZN(n6246) );
  OAI211_X1 U7350 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n6244), .B(n6243), .ZN(n6245) );
  OAI211_X1 U7351 ( .C1(n6247), .C2(n6362), .A(n6246), .B(n6245), .ZN(U2811)
         );
  OAI21_X1 U7352 ( .B1(n6354), .B2(n6248), .A(n6312), .ZN(n6251) );
  OAI22_X1 U7353 ( .A1(n7109), .A2(n6331), .B1(n6912), .B2(n6249), .ZN(n6250)
         );
  AOI211_X1 U7354 ( .C1(n6322), .C2(n6364), .A(n6251), .B(n6250), .ZN(n6255)
         );
  INV_X1 U7355 ( .A(n6252), .ZN(n6253) );
  AOI22_X1 U7356 ( .A1(n6365), .A2(n6315), .B1(n6357), .B2(n6253), .ZN(n6254)
         );
  OAI211_X1 U7357 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6256), .A(n6255), .B(n6254), .ZN(U2812) );
  INV_X1 U7358 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6909) );
  OAI22_X1 U7359 ( .A1(n6259), .A2(n6258), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6257), .ZN(n6263) );
  INV_X1 U7360 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6261) );
  AOI22_X1 U7361 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6346), .B1(n6322), .B2(n6367), .ZN(n6260) );
  OAI211_X1 U7362 ( .C1(n6354), .C2(n6261), .A(n6260), .B(n6312), .ZN(n6262)
         );
  AOI221_X1 U7363 ( .B1(n6264), .B2(n6909), .C1(n6263), .C2(
        REIP_REG_13__SCAN_IN), .A(n6262), .ZN(n6266) );
  NAND2_X1 U7364 ( .A1(n6392), .A2(n6315), .ZN(n6265) );
  OAI211_X1 U7365 ( .C1(n6343), .C2(n6267), .A(n6266), .B(n6265), .ZN(U2814)
         );
  AOI21_X1 U7366 ( .B1(n6269), .B2(n6268), .A(n5461), .ZN(n6370) );
  NAND2_X1 U7367 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6286) );
  NOR2_X1 U7368 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6286), .ZN(n6270) );
  AOI22_X1 U7369 ( .A1(n6322), .A2(n6370), .B1(n6289), .B2(n6270), .ZN(n6276)
         );
  INV_X1 U7370 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7240) );
  OAI22_X1 U7371 ( .A1(n6272), .A2(n6354), .B1(n7240), .B2(n6271), .ZN(n6273)
         );
  AOI211_X1 U7372 ( .C1(n6346), .C2(EBX_REG_11__SCAN_IN), .A(n6323), .B(n6273), 
        .ZN(n6275) );
  INV_X1 U7373 ( .A(n6372), .ZN(n6439) );
  AOI22_X1 U7374 ( .A1(n6439), .A2(n6315), .B1(n6357), .B2(n6437), .ZN(n6274)
         );
  NAND3_X1 U7375 ( .A1(n6276), .A2(n6275), .A3(n6274), .ZN(U2816) );
  AND2_X1 U7376 ( .A1(n6278), .A2(n6277), .ZN(n6299) );
  AOI21_X1 U7377 ( .B1(n6346), .B2(EBX_REG_10__SCAN_IN), .A(n6323), .ZN(n6279)
         );
  OAI21_X1 U7378 ( .B1(n6354), .B2(n6280), .A(n6279), .ZN(n6281) );
  AOI21_X1 U7379 ( .B1(n6299), .B2(REIP_REG_10__SCAN_IN), .A(n6281), .ZN(n6282) );
  OAI21_X1 U7380 ( .B1(n6283), .B2(n6302), .A(n6282), .ZN(n6284) );
  AOI21_X1 U7381 ( .B1(n6285), .B2(n6357), .A(n6284), .ZN(n6288) );
  OAI211_X1 U7382 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n6289), .B(n6286), .ZN(n6287) );
  OAI211_X1 U7383 ( .C1(n6486), .C2(n6362), .A(n6288), .B(n6287), .ZN(U2817)
         );
  INV_X1 U7384 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6905) );
  AOI22_X1 U7385 ( .A1(n6322), .A2(n6497), .B1(n6289), .B2(n6905), .ZN(n6296)
         );
  AOI22_X1 U7386 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6332), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6299), .ZN(n6295) );
  AOI21_X1 U7387 ( .B1(n6346), .B2(EBX_REG_9__SCAN_IN), .A(n6323), .ZN(n6294)
         );
  INV_X1 U7388 ( .A(n6290), .ZN(n6292) );
  AOI22_X1 U7389 ( .A1(n6292), .A2(n6315), .B1(n6357), .B2(n6291), .ZN(n6293)
         );
  NAND4_X1 U7390 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(U2818)
         );
  AOI21_X1 U7391 ( .B1(n6332), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6323), 
        .ZN(n6307) );
  NOR2_X1 U7392 ( .A1(n6334), .A2(REIP_REG_8__SCAN_IN), .ZN(n6297) );
  AOI22_X1 U7393 ( .A1(n6346), .A2(EBX_REG_8__SCAN_IN), .B1(n6298), .B2(n6297), 
        .ZN(n6301) );
  NAND2_X1 U7394 ( .A1(n6299), .A2(REIP_REG_8__SCAN_IN), .ZN(n6300) );
  OAI211_X1 U7395 ( .C1(n6303), .C2(n6302), .A(n6301), .B(n6300), .ZN(n6304)
         );
  AOI21_X1 U7396 ( .B1(n6305), .B2(n6357), .A(n6304), .ZN(n6306) );
  OAI211_X1 U7397 ( .C1(n6362), .C2(n6308), .A(n6307), .B(n6306), .ZN(U2819)
         );
  AOI21_X1 U7398 ( .B1(n6310), .B2(REIP_REG_6__SCAN_IN), .A(n6309), .ZN(n6317)
         );
  XOR2_X1 U7399 ( .A(n4996), .B(n6311), .Z(n6513) );
  AOI22_X1 U7400 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6332), .B1(n6322), 
        .B2(n6513), .ZN(n6313) );
  OAI211_X1 U7401 ( .C1(n6343), .C2(n6447), .A(n6313), .B(n6312), .ZN(n6314)
         );
  AOI21_X1 U7402 ( .B1(n6315), .B2(n6444), .A(n6314), .ZN(n6316) );
  OAI211_X1 U7403 ( .C1(n6377), .C2(n6331), .A(n6317), .B(n6316), .ZN(U2821)
         );
  XOR2_X1 U7404 ( .A(n6319), .B(n6318), .Z(n6538) );
  NOR2_X1 U7405 ( .A1(n6334), .A2(REIP_REG_4__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U7406 ( .A1(n6322), .A2(n6538), .B1(n6321), .B2(n6320), .ZN(n6330)
         );
  AOI21_X1 U7407 ( .B1(n6332), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6323), 
        .ZN(n6327) );
  AOI22_X1 U7408 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6325), .B1(n6324), .B2(n6349), .ZN(n6326) );
  OAI211_X1 U7409 ( .C1(n6343), .C2(n6455), .A(n6327), .B(n6326), .ZN(n6328)
         );
  AOI21_X1 U7410 ( .B1(n6452), .B2(n6348), .A(n6328), .ZN(n6329) );
  OAI211_X1 U7411 ( .C1(n6379), .C2(n6331), .A(n6330), .B(n6329), .ZN(U2823)
         );
  NOR2_X1 U7412 ( .A1(n6552), .A2(n6362), .ZN(n6341) );
  NAND2_X1 U7413 ( .A1(n6332), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6338)
         );
  OR2_X1 U7414 ( .A1(n6334), .A2(REIP_REG_1__SCAN_IN), .ZN(n6344) );
  NAND3_X1 U7415 ( .A1(n6333), .A2(REIP_REG_2__SCAN_IN), .A3(n6344), .ZN(n6336) );
  OAI21_X1 U7416 ( .B1(n6334), .B2(n6895), .A(n7306), .ZN(n6335) );
  AOI22_X1 U7417 ( .A1(n6336), .A2(n6335), .B1(n6346), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n6337) );
  OAI211_X1 U7418 ( .C1(n6339), .C2(n4755), .A(n6338), .B(n6337), .ZN(n6340)
         );
  AOI211_X1 U7419 ( .C1(n6348), .C2(n6462), .A(n6341), .B(n6340), .ZN(n6342)
         );
  OAI21_X1 U7420 ( .B1(n6465), .B2(n6343), .A(n6342), .ZN(U2825) );
  INV_X1 U7421 ( .A(n6344), .ZN(n6345) );
  AOI21_X1 U7422 ( .B1(n6346), .B2(EBX_REG_1__SCAN_IN), .A(n6345), .ZN(n6361)
         );
  NAND2_X1 U7423 ( .A1(n6348), .A2(n6347), .ZN(n6359) );
  NAND2_X1 U7424 ( .A1(n6350), .A2(n6349), .ZN(n6353) );
  NAND2_X1 U7425 ( .A1(n6351), .A2(REIP_REG_1__SCAN_IN), .ZN(n6352) );
  OAI211_X1 U7426 ( .C1(n6354), .C2(n6356), .A(n6353), .B(n6352), .ZN(n6355)
         );
  AOI21_X1 U7427 ( .B1(n6357), .B2(n6356), .A(n6355), .ZN(n6358) );
  AND2_X1 U7428 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  OAI211_X1 U7429 ( .C1(n6363), .C2(n6362), .A(n6361), .B(n6360), .ZN(U2826)
         );
  AOI22_X1 U7430 ( .A1(n6365), .A2(n4359), .B1(n4474), .B2(n6364), .ZN(n6366)
         );
  OAI21_X1 U7431 ( .B1(n6380), .B2(n7109), .A(n6366), .ZN(U2844) );
  AOI22_X1 U7432 ( .A1(n6392), .A2(n4359), .B1(n4474), .B2(n6367), .ZN(n6368)
         );
  OAI21_X1 U7433 ( .B1(n6380), .B2(n6369), .A(n6368), .ZN(U2846) );
  INV_X1 U7434 ( .A(n6370), .ZN(n6477) );
  OAI22_X1 U7435 ( .A1(n6372), .A2(n6152), .B1(n6371), .B2(n6477), .ZN(n6373)
         );
  INV_X1 U7436 ( .A(n6373), .ZN(n6374) );
  OAI21_X1 U7437 ( .B1(n6380), .B2(n6375), .A(n6374), .ZN(U2848) );
  AOI22_X1 U7438 ( .A1(n6444), .A2(n4359), .B1(n4474), .B2(n6513), .ZN(n6376)
         );
  OAI21_X1 U7439 ( .B1(n6380), .B2(n6377), .A(n6376), .ZN(U2853) );
  AOI22_X1 U7440 ( .A1(n6452), .A2(n4359), .B1(n4474), .B2(n6538), .ZN(n6378)
         );
  OAI21_X1 U7441 ( .B1(n6380), .B2(n6379), .A(n6378), .ZN(U2855) );
  AOI22_X1 U7442 ( .A1(n6381), .A2(n6391), .B1(n6384), .B2(DATAI_18_), .ZN(
        n6383) );
  AOI22_X1 U7443 ( .A1(n6387), .A2(DATAI_2_), .B1(n6386), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U7444 ( .A1(n6383), .A2(n6382), .ZN(U2873) );
  AOI22_X1 U7445 ( .A1(n6385), .A2(n6391), .B1(n6384), .B2(DATAI_16_), .ZN(
        n6389) );
  AOI22_X1 U7446 ( .A1(n6387), .A2(DATAI_0_), .B1(n6386), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U7447 ( .A1(n6389), .A2(n6388), .ZN(U2875) );
  AOI22_X1 U7448 ( .A1(n6392), .A2(n6391), .B1(DATAI_13_), .B2(n6390), .ZN(
        n6393) );
  OAI21_X1 U7449 ( .B1(n3885), .B2(n6394), .A(n6393), .ZN(U2878) );
  INV_X1 U7450 ( .A(n6395), .ZN(n6399) );
  AOI22_X1 U7451 ( .A1(n6399), .A2(EAX_REG_29__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6396) );
  OAI21_X1 U7452 ( .B1(n6419), .B2(n7175), .A(n6396), .ZN(U2894) );
  AOI22_X1 U7453 ( .A1(n6399), .A2(EAX_REG_28__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6397) );
  OAI21_X1 U7454 ( .B1(n6419), .B2(n7316), .A(n6397), .ZN(U2895) );
  INV_X1 U7455 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n7148) );
  AOI22_X1 U7456 ( .A1(n6399), .A2(EAX_REG_26__SCAN_IN), .B1(n6982), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6398) );
  OAI21_X1 U7457 ( .B1(n7148), .B2(n6417), .A(n6398), .ZN(U2897) );
  AOI22_X1 U7458 ( .A1(n6399), .A2(EAX_REG_24__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n6400) );
  OAI21_X1 U7459 ( .B1(n6419), .B2(n7151), .A(n6400), .ZN(U2899) );
  AOI22_X1 U7460 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6415), .B1(
        DATAO_REG_15__SCAN_IN), .B2(n6420), .ZN(n6401) );
  OAI21_X1 U7461 ( .B1(n6419), .B2(n7217), .A(n6401), .ZN(U2908) );
  AOI22_X1 U7462 ( .A1(n6982), .A2(LWORD_REG_14__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6402) );
  OAI21_X1 U7463 ( .B1(n5579), .B2(n6422), .A(n6402), .ZN(U2909) );
  AOI22_X1 U7464 ( .A1(n6982), .A2(LWORD_REG_13__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6403) );
  OAI21_X1 U7465 ( .B1(n3885), .B2(n6422), .A(n6403), .ZN(U2910) );
  AOI22_X1 U7466 ( .A1(n6982), .A2(LWORD_REG_12__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6404) );
  OAI21_X1 U7467 ( .B1(n5526), .B2(n6422), .A(n6404), .ZN(U2911) );
  AOI222_X1 U7468 ( .A1(n6982), .A2(LWORD_REG_11__SCAN_IN), .B1(n6415), .B2(
        EAX_REG_11__SCAN_IN), .C1(DATAO_REG_11__SCAN_IN), .C2(n6420), .ZN(
        n6405) );
  INV_X1 U7469 ( .A(n6405), .ZN(U2912) );
  AOI22_X1 U7470 ( .A1(n6982), .A2(LWORD_REG_10__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6406) );
  OAI21_X1 U7471 ( .B1(n3862), .B2(n6422), .A(n6406), .ZN(U2913) );
  AOI22_X1 U7472 ( .A1(n6982), .A2(LWORD_REG_9__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U7473 ( .B1(n4864), .B2(n6422), .A(n6407), .ZN(U2914) );
  INV_X1 U7474 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6409) );
  AOI22_X1 U7475 ( .A1(n6982), .A2(LWORD_REG_8__SCAN_IN), .B1(
        DATAO_REG_8__SCAN_IN), .B2(n6420), .ZN(n6408) );
  OAI21_X1 U7476 ( .B1(n6409), .B2(n6422), .A(n6408), .ZN(U2915) );
  AOI22_X1 U7477 ( .A1(n6982), .A2(LWORD_REG_7__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6410) );
  OAI21_X1 U7478 ( .B1(n4871), .B2(n6422), .A(n6410), .ZN(U2916) );
  INV_X1 U7479 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n7231) );
  OAI222_X1 U7480 ( .A1(n6417), .A2(n7231), .B1(n6422), .B2(n6411), .C1(n6419), 
        .C2(n4869), .ZN(U2917) );
  AOI22_X1 U7481 ( .A1(n6982), .A2(LWORD_REG_5__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6412) );
  OAI21_X1 U7482 ( .B1(n4873), .B2(n6422), .A(n6412), .ZN(U2918) );
  AOI222_X1 U7483 ( .A1(n6420), .A2(DATAO_REG_4__SCAN_IN), .B1(n6415), .B2(
        EAX_REG_4__SCAN_IN), .C1(n6982), .C2(LWORD_REG_4__SCAN_IN), .ZN(n6413)
         );
  INV_X1 U7484 ( .A(n6413), .ZN(U2919) );
  AOI22_X1 U7485 ( .A1(n6982), .A2(LWORD_REG_3__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6414) );
  OAI21_X1 U7486 ( .B1(n7183), .B2(n6422), .A(n6414), .ZN(U2920) );
  AOI222_X1 U7487 ( .A1(n6420), .A2(DATAO_REG_2__SCAN_IN), .B1(n6415), .B2(
        EAX_REG_2__SCAN_IN), .C1(n6982), .C2(LWORD_REG_2__SCAN_IN), .ZN(n6416)
         );
  INV_X1 U7488 ( .A(n6416), .ZN(U2921) );
  INV_X1 U7489 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n7230) );
  OAI222_X1 U7490 ( .A1(n6419), .A2(n4862), .B1(n6422), .B2(n6418), .C1(n7230), 
        .C2(n6417), .ZN(U2922) );
  AOI22_X1 U7491 ( .A1(n6982), .A2(LWORD_REG_0__SCAN_IN), .B1(n6420), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6421) );
  OAI21_X1 U7492 ( .B1(n7271), .B2(n6422), .A(n6421), .ZN(U2923) );
  AOI22_X1 U7493 ( .A1(n6430), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6429), .ZN(n6424) );
  NAND2_X1 U7494 ( .A1(n6424), .A2(n6423), .ZN(U2947) );
  AOI22_X1 U7495 ( .A1(n6430), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6429), .ZN(n6426) );
  NAND2_X1 U7496 ( .A1(n6426), .A2(n6425), .ZN(U2950) );
  AOI22_X1 U7497 ( .A1(n6430), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6429), .ZN(n6428) );
  NAND2_X1 U7498 ( .A1(n6428), .A2(n6427), .ZN(U2951) );
  AOI22_X1 U7499 ( .A1(n6430), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6429), .ZN(n6432) );
  NAND2_X1 U7500 ( .A1(n6432), .A2(n6431), .ZN(U2953) );
  NAND2_X1 U7501 ( .A1(n6434), .A2(n6433), .ZN(n6436) );
  XNOR2_X1 U7502 ( .A(n3203), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6435)
         );
  XNOR2_X1 U7503 ( .A(n6436), .B(n6435), .ZN(n6479) );
  AOI22_X1 U7504 ( .A1(n6567), .A2(REIP_REG_11__SCAN_IN), .B1(n6456), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6441) );
  AOI22_X1 U7505 ( .A1(n6439), .A2(n6461), .B1(n6438), .B2(n6437), .ZN(n6440)
         );
  OAI211_X1 U7506 ( .C1(n6479), .C2(n6468), .A(n6441), .B(n6440), .ZN(U2975)
         );
  AOI22_X1 U7507 ( .A1(n6567), .A2(REIP_REG_6__SCAN_IN), .B1(n6456), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6446) );
  AOI22_X1 U7508 ( .A1(n3222), .A2(n6460), .B1(n6461), .B2(n6444), .ZN(n6445)
         );
  OAI211_X1 U7509 ( .C1(n6466), .C2(n6447), .A(n6446), .B(n6445), .ZN(U2980)
         );
  AOI22_X1 U7510 ( .A1(n6567), .A2(REIP_REG_4__SCAN_IN), .B1(n6456), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6454) );
  OAI21_X1 U7511 ( .B1(n6448), .B2(n6450), .A(n6449), .ZN(n6451) );
  INV_X1 U7512 ( .A(n6451), .ZN(n6539) );
  AOI22_X1 U7513 ( .A1(n6539), .A2(n6460), .B1(n6452), .B2(n6461), .ZN(n6453)
         );
  OAI211_X1 U7514 ( .C1(n6466), .C2(n6455), .A(n6454), .B(n6453), .ZN(U2982)
         );
  AOI22_X1 U7515 ( .A1(n6567), .A2(REIP_REG_2__SCAN_IN), .B1(n6456), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6464) );
  XNOR2_X1 U7516 ( .A(n6457), .B(n6564), .ZN(n6459) );
  XNOR2_X1 U7517 ( .A(n6459), .B(n6458), .ZN(n6561) );
  AOI22_X1 U7518 ( .A1(n6462), .A2(n6461), .B1(n6460), .B2(n6561), .ZN(n6463)
         );
  OAI211_X1 U7519 ( .C1(n6466), .C2(n6465), .A(n6464), .B(n6463), .ZN(U2984)
         );
  INV_X1 U7520 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n7123) );
  XNOR2_X1 U7521 ( .A(n6467), .B(n6575), .ZN(n6572) );
  INV_X1 U7522 ( .A(n6572), .ZN(n6469) );
  OAI22_X1 U7523 ( .A1(n6471), .A2(n6470), .B1(n6469), .B2(n6468), .ZN(n6472)
         );
  AOI21_X1 U7524 ( .B1(n6567), .B2(REIP_REG_0__SCAN_IN), .A(n6472), .ZN(n6473)
         );
  OAI221_X1 U7525 ( .B1(n7123), .B2(n6475), .C1(n7123), .C2(n6474), .A(n6473), 
        .ZN(U2986) );
  INV_X1 U7526 ( .A(n6476), .ZN(n6482) );
  OAI22_X1 U7527 ( .A1(n6551), .A2(n6477), .B1(n7240), .B2(n6556), .ZN(n6481)
         );
  NOR2_X1 U7528 ( .A1(n6479), .A2(n6478), .ZN(n6480) );
  AOI211_X1 U7529 ( .C1(n6482), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n6481), .B(n6480), .ZN(n6484) );
  NAND2_X1 U7530 ( .A1(n6484), .A2(n6483), .ZN(U3007) );
  NAND2_X1 U7531 ( .A1(n6490), .A2(n6507), .ZN(n6502) );
  AOI22_X1 U7532 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n4557), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6485), .ZN(n6494) );
  INV_X1 U7533 ( .A(n6486), .ZN(n6489) );
  INV_X1 U7534 ( .A(n6487), .ZN(n6488) );
  AOI21_X1 U7535 ( .B1(n6569), .B2(n6489), .A(n6488), .ZN(n6493) );
  OAI21_X1 U7536 ( .B1(n6518), .B2(n6490), .A(n6512), .ZN(n6498) );
  AOI22_X1 U7537 ( .A1(n6491), .A2(n6571), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6498), .ZN(n6492) );
  OAI211_X1 U7538 ( .C1(n6502), .C2(n6494), .A(n6493), .B(n6492), .ZN(U3008)
         );
  INV_X1 U7539 ( .A(n6495), .ZN(n6496) );
  AOI21_X1 U7540 ( .B1(n6569), .B2(n6497), .A(n6496), .ZN(n6501) );
  AOI22_X1 U7541 ( .A1(n6499), .A2(n6571), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6498), .ZN(n6500) );
  OAI211_X1 U7542 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6502), .A(n6501), 
        .B(n6500), .ZN(U3009) );
  INV_X1 U7543 ( .A(n6503), .ZN(n6504) );
  AOI21_X1 U7544 ( .B1(n6569), .B2(n6505), .A(n6504), .ZN(n6510) );
  INV_X1 U7545 ( .A(n6506), .ZN(n6508) );
  AOI22_X1 U7546 ( .A1(n6508), .A2(n6571), .B1(n6507), .B2(n6511), .ZN(n6509)
         );
  OAI211_X1 U7547 ( .C1(n6512), .C2(n6511), .A(n6510), .B(n6509), .ZN(U3011)
         );
  AOI22_X1 U7548 ( .A1(n6569), .A2(n6513), .B1(n6567), .B2(REIP_REG_6__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U7549 ( .A1(n6558), .A2(n6516), .B1(n6515), .B2(n6514), .ZN(n6563)
         );
  OAI21_X1 U7550 ( .B1(n6518), .B2(n6517), .A(n6563), .ZN(n6531) );
  AOI22_X1 U7551 ( .A1(n3222), .A2(n6571), .B1(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .B2(n6531), .ZN(n6519) );
  OAI211_X1 U7552 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n6521), .A(n6520), 
        .B(n6519), .ZN(U3012) );
  INV_X1 U7553 ( .A(n6522), .ZN(n6525) );
  INV_X1 U7554 ( .A(n6523), .ZN(n6524) );
  AOI21_X1 U7555 ( .B1(n6569), .B2(n6525), .A(n6524), .ZN(n6535) );
  INV_X1 U7556 ( .A(n6526), .ZN(n6530) );
  NOR2_X1 U7557 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6527), .ZN(n6529)
         );
  AOI22_X1 U7558 ( .A1(n6530), .A2(n6571), .B1(n6529), .B2(n6528), .ZN(n6534)
         );
  OAI21_X1 U7559 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6532), .A(n6531), 
        .ZN(n6533) );
  NAND3_X1 U7560 ( .A1(n6535), .A2(n6534), .A3(n6533), .ZN(U3013) );
  NAND2_X1 U7561 ( .A1(n6536), .A2(n6554), .ZN(n6549) );
  OAI21_X1 U7562 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6537), .ZN(n6542) );
  AOI22_X1 U7563 ( .A1(n6569), .A2(n6538), .B1(n6567), .B2(REIP_REG_4__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U7564 ( .B1(n6554), .B2(n6558), .A(n6563), .ZN(n6546) );
  AOI22_X1 U7565 ( .A1(n6546), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6571), 
        .B2(n6539), .ZN(n6540) );
  OAI211_X1 U7566 ( .C1(n6549), .C2(n6542), .A(n6541), .B(n6540), .ZN(U3014)
         );
  AOI21_X1 U7567 ( .B1(n6569), .B2(n6544), .A(n6543), .ZN(n6548) );
  AOI22_X1 U7568 ( .A1(n6546), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6571), 
        .B2(n6545), .ZN(n6547) );
  OAI211_X1 U7569 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6549), .A(n6548), 
        .B(n6547), .ZN(U3015) );
  NAND2_X1 U7570 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6550), .ZN(n6565)
         );
  NOR2_X1 U7571 ( .A1(n6552), .A2(n6551), .ZN(n6560) );
  INV_X1 U7572 ( .A(n6554), .ZN(n6555) );
  AOI21_X1 U7573 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n4491), .A(n6555), 
        .ZN(n6557) );
  OAI22_X1 U7574 ( .A1(n6558), .A2(n6557), .B1(n7306), .B2(n6556), .ZN(n6559)
         );
  AOI211_X1 U7575 ( .C1(n6561), .C2(n6571), .A(n6560), .B(n6559), .ZN(n6562)
         );
  OAI221_X1 U7576 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6565), .C1(n6564), .C2(n6563), .A(n6562), .ZN(U3016) );
  INV_X1 U7577 ( .A(n6566), .ZN(n6576) );
  AOI22_X1 U7578 ( .A1(n6569), .A2(n6568), .B1(n6567), .B2(REIP_REG_0__SCAN_IN), .ZN(n6574) );
  AOI21_X1 U7579 ( .B1(n6572), .B2(n6571), .A(n6570), .ZN(n6573) );
  OAI211_X1 U7580 ( .C1(n6576), .C2(n6575), .A(n6574), .B(n6573), .ZN(U3018)
         );
  NOR2_X1 U7581 ( .A1(n7293), .A2(n6577), .ZN(U3019) );
  INV_X1 U7582 ( .A(n6740), .ZN(n6578) );
  NAND2_X1 U7583 ( .A1(n6578), .A2(n6850), .ZN(n6612) );
  OAI22_X1 U7584 ( .A1(n6625), .A2(n6760), .B1(n6741), .B2(n6612), .ZN(n6579)
         );
  INV_X1 U7585 ( .A(n6579), .ZN(n6593) );
  INV_X1 U7586 ( .A(n6580), .ZN(n6581) );
  NAND2_X1 U7587 ( .A1(n6581), .A2(n6744), .ZN(n6582) );
  OAI21_X1 U7588 ( .B1(n6583), .B2(n6582), .A(n6753), .ZN(n6591) );
  OR2_X1 U7589 ( .A1(n6584), .A2(n6653), .ZN(n6585) );
  AND2_X1 U7590 ( .A1(n6585), .A2(n6612), .ZN(n6590) );
  INV_X1 U7591 ( .A(n6590), .ZN(n6588) );
  AOI21_X1 U7592 ( .B1(n6589), .B2(n6658), .A(n6586), .ZN(n6587) );
  OAI21_X1 U7593 ( .B1(n6591), .B2(n6588), .A(n6587), .ZN(n6616) );
  OAI22_X1 U7594 ( .A1(n6591), .A2(n6590), .B1(n6589), .B2(n3658), .ZN(n6615)
         );
  AOI22_X1 U7595 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6616), .B1(n6757), 
        .B2(n6615), .ZN(n6592) );
  OAI211_X1 U7596 ( .C1(n6742), .C2(n6613), .A(n6593), .B(n6592), .ZN(U3044)
         );
  OAI22_X1 U7597 ( .A1(n6625), .A2(n6767), .B1(n6761), .B2(n6612), .ZN(n6594)
         );
  INV_X1 U7598 ( .A(n6594), .ZN(n6596) );
  AOI22_X1 U7599 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6616), .B1(n6764), 
        .B2(n6615), .ZN(n6595) );
  OAI211_X1 U7600 ( .C1(n6613), .C2(n6762), .A(n6596), .B(n6595), .ZN(U3045)
         );
  OAI22_X1 U7601 ( .A1(n6625), .A2(n6774), .B1(n6768), .B2(n6612), .ZN(n6597)
         );
  INV_X1 U7602 ( .A(n6597), .ZN(n6599) );
  AOI22_X1 U7603 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6616), .B1(n6771), 
        .B2(n6615), .ZN(n6598) );
  OAI211_X1 U7604 ( .C1(n6613), .C2(n6769), .A(n6599), .B(n6598), .ZN(U3046)
         );
  OAI22_X1 U7605 ( .A1(n6613), .A2(n6776), .B1(n6775), .B2(n6612), .ZN(n6600)
         );
  INV_X1 U7606 ( .A(n6600), .ZN(n6602) );
  AOI22_X1 U7607 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6616), .B1(n6778), 
        .B2(n6615), .ZN(n6601) );
  OAI211_X1 U7608 ( .C1(n6781), .C2(n6625), .A(n6602), .B(n6601), .ZN(U3047)
         );
  OAI22_X1 U7609 ( .A1(n6613), .A2(n7378), .B1(n7368), .B2(n6612), .ZN(n6603)
         );
  INV_X1 U7610 ( .A(n6603), .ZN(n6605) );
  AOI22_X1 U7611 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6616), .B1(n7373), 
        .B2(n6615), .ZN(n6604) );
  OAI211_X1 U7612 ( .C1(n7369), .C2(n6625), .A(n6605), .B(n6604), .ZN(U3048)
         );
  OAI22_X1 U7613 ( .A1(n6625), .A2(n6788), .B1(n6782), .B2(n6612), .ZN(n6606)
         );
  INV_X1 U7614 ( .A(n6606), .ZN(n6608) );
  AOI22_X1 U7615 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6616), .B1(n6785), 
        .B2(n6615), .ZN(n6607) );
  OAI211_X1 U7616 ( .C1(n6613), .C2(n6783), .A(n6608), .B(n6607), .ZN(U3049)
         );
  OAI22_X1 U7617 ( .A1(n6625), .A2(n6790), .B1(n6789), .B2(n6612), .ZN(n6609)
         );
  INV_X1 U7618 ( .A(n6609), .ZN(n6611) );
  AOI22_X1 U7619 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6616), .B1(n6799), 
        .B2(n6615), .ZN(n6610) );
  OAI211_X1 U7620 ( .C1(n6613), .C2(n6804), .A(n6611), .B(n6610), .ZN(U3050)
         );
  OAI22_X1 U7621 ( .A1(n6613), .A2(n6814), .B1(n6794), .B2(n6612), .ZN(n6614)
         );
  INV_X1 U7622 ( .A(n6614), .ZN(n6618) );
  AOI22_X1 U7623 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6616), .B1(n6806), 
        .B2(n6615), .ZN(n6617) );
  OAI211_X1 U7624 ( .C1(n6795), .C2(n6625), .A(n6618), .B(n6617), .ZN(U3051)
         );
  AOI22_X1 U7625 ( .A1(n6800), .A2(n6620), .B1(n6799), .B2(n6619), .ZN(n6624)
         );
  AOI22_X1 U7626 ( .A1(n6622), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6801), 
        .B2(n6621), .ZN(n6623) );
  OAI211_X1 U7627 ( .C1(n6804), .C2(n6625), .A(n6624), .B(n6623), .ZN(U3058)
         );
  AOI22_X1 U7628 ( .A1(n6698), .A2(n6643), .B1(n6757), .B2(n6642), .ZN(n6629)
         );
  AOI22_X1 U7629 ( .A1(n6646), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6627), 
        .B2(n6644), .ZN(n6628) );
  OAI211_X1 U7630 ( .C1(n6760), .C2(n6685), .A(n6629), .B(n6628), .ZN(U3068)
         );
  AOI22_X1 U7631 ( .A1(n6711), .A2(n6643), .B1(n6764), .B2(n6642), .ZN(n6632)
         );
  AOI22_X1 U7632 ( .A1(n6646), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6630), 
        .B2(n6644), .ZN(n6631) );
  OAI211_X1 U7633 ( .C1(n6767), .C2(n6685), .A(n6632), .B(n6631), .ZN(U3069)
         );
  AOI22_X1 U7634 ( .A1(n6715), .A2(n6643), .B1(n6771), .B2(n6642), .ZN(n6635)
         );
  AOI22_X1 U7635 ( .A1(n6646), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6633), 
        .B2(n6644), .ZN(n6634) );
  OAI211_X1 U7636 ( .C1(n6774), .C2(n6685), .A(n6635), .B(n6634), .ZN(U3070)
         );
  AOI22_X1 U7637 ( .A1(n6719), .A2(n6643), .B1(n6778), .B2(n6642), .ZN(n6638)
         );
  AOI22_X1 U7638 ( .A1(n6646), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6636), 
        .B2(n6644), .ZN(n6637) );
  OAI211_X1 U7639 ( .C1(n6781), .C2(n6685), .A(n6638), .B(n6637), .ZN(U3071)
         );
  AOI22_X1 U7640 ( .A1(n6723), .A2(n6643), .B1(n7373), .B2(n6642), .ZN(n6641)
         );
  AOI22_X1 U7641 ( .A1(n6646), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6639), 
        .B2(n6644), .ZN(n6640) );
  OAI211_X1 U7642 ( .C1(n7369), .C2(n6685), .A(n6641), .B(n6640), .ZN(U3072)
         );
  AOI22_X1 U7643 ( .A1(n6727), .A2(n6643), .B1(n6785), .B2(n6642), .ZN(n6648)
         );
  AOI22_X1 U7644 ( .A1(n6646), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6645), 
        .B2(n6644), .ZN(n6647) );
  OAI211_X1 U7645 ( .C1(n6788), .C2(n6685), .A(n6648), .B(n6647), .ZN(U3073)
         );
  OAI22_X1 U7646 ( .A1(n6685), .A2(n6742), .B1(n6741), .B2(n6684), .ZN(n6651)
         );
  INV_X1 U7647 ( .A(n6651), .ZN(n6665) );
  NOR3_X1 U7648 ( .A1(n6655), .A2(n6654), .A3(n6653), .ZN(n6657) );
  INV_X1 U7649 ( .A(n6684), .ZN(n6656) );
  NOR2_X1 U7650 ( .A1(n6657), .A2(n6656), .ZN(n6663) );
  AOI22_X1 U7651 ( .A1(n6660), .A2(n6663), .B1(n6661), .B2(n6658), .ZN(n6659)
         );
  NAND2_X1 U7652 ( .A1(n6749), .A2(n6659), .ZN(n6688) );
  INV_X1 U7653 ( .A(n6660), .ZN(n6662) );
  OAI22_X1 U7654 ( .A1(n6663), .A2(n6662), .B1(n3658), .B2(n6661), .ZN(n6687)
         );
  AOI22_X1 U7655 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6688), .B1(n6757), 
        .B2(n6687), .ZN(n6664) );
  OAI211_X1 U7656 ( .C1(n6760), .C2(n6739), .A(n6665), .B(n6664), .ZN(U3076)
         );
  OAI22_X1 U7657 ( .A1(n6685), .A2(n6762), .B1(n6761), .B2(n6684), .ZN(n6666)
         );
  INV_X1 U7658 ( .A(n6666), .ZN(n6668) );
  AOI22_X1 U7659 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6688), .B1(n6764), 
        .B2(n6687), .ZN(n6667) );
  OAI211_X1 U7660 ( .C1(n6767), .C2(n6739), .A(n6668), .B(n6667), .ZN(U3077)
         );
  OAI22_X1 U7661 ( .A1(n6739), .A2(n6774), .B1(n6768), .B2(n6684), .ZN(n6669)
         );
  INV_X1 U7662 ( .A(n6669), .ZN(n6671) );
  AOI22_X1 U7663 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6688), .B1(n6771), 
        .B2(n6687), .ZN(n6670) );
  OAI211_X1 U7664 ( .C1(n6769), .C2(n6685), .A(n6671), .B(n6670), .ZN(U3078)
         );
  OAI22_X1 U7665 ( .A1(n6685), .A2(n6776), .B1(n6775), .B2(n6684), .ZN(n6672)
         );
  INV_X1 U7666 ( .A(n6672), .ZN(n6674) );
  AOI22_X1 U7667 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6688), .B1(n6778), 
        .B2(n6687), .ZN(n6673) );
  OAI211_X1 U7668 ( .C1(n6781), .C2(n6739), .A(n6674), .B(n6673), .ZN(U3079)
         );
  OAI22_X1 U7669 ( .A1(n6685), .A2(n7378), .B1(n7368), .B2(n6684), .ZN(n6675)
         );
  INV_X1 U7670 ( .A(n6675), .ZN(n6677) );
  AOI22_X1 U7671 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6688), .B1(n7373), 
        .B2(n6687), .ZN(n6676) );
  OAI211_X1 U7672 ( .C1(n7369), .C2(n6739), .A(n6677), .B(n6676), .ZN(U3080)
         );
  OAI22_X1 U7673 ( .A1(n6685), .A2(n6783), .B1(n6782), .B2(n6684), .ZN(n6678)
         );
  INV_X1 U7674 ( .A(n6678), .ZN(n6680) );
  AOI22_X1 U7675 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6688), .B1(n6785), 
        .B2(n6687), .ZN(n6679) );
  OAI211_X1 U7676 ( .C1(n6788), .C2(n6739), .A(n6680), .B(n6679), .ZN(U3081)
         );
  OAI22_X1 U7677 ( .A1(n6685), .A2(n6804), .B1(n6789), .B2(n6684), .ZN(n6681)
         );
  INV_X1 U7678 ( .A(n6681), .ZN(n6683) );
  AOI22_X1 U7679 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6688), .B1(n6799), 
        .B2(n6687), .ZN(n6682) );
  OAI211_X1 U7680 ( .C1(n6790), .C2(n6739), .A(n6683), .B(n6682), .ZN(U3082)
         );
  OAI22_X1 U7681 ( .A1(n6685), .A2(n6814), .B1(n6794), .B2(n6684), .ZN(n6686)
         );
  INV_X1 U7682 ( .A(n6686), .ZN(n6690) );
  AOI22_X1 U7683 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6688), .B1(n6806), 
        .B2(n6687), .ZN(n6689) );
  OAI211_X1 U7684 ( .C1(n6795), .C2(n6739), .A(n6690), .B(n6689), .ZN(U3083)
         );
  NOR2_X1 U7685 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6691), .ZN(n6734)
         );
  NAND3_X1 U7686 ( .A1(n6692), .A2(n6753), .A3(n4893), .ZN(n6697) );
  INV_X1 U7687 ( .A(n6693), .ZN(n6695) );
  NAND2_X1 U7688 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  NAND2_X1 U7689 ( .A1(n6697), .A2(n6696), .ZN(n6733) );
  AOI22_X1 U7690 ( .A1(n6698), .A2(n6734), .B1(n6757), .B2(n6733), .ZN(n6710)
         );
  INV_X1 U7691 ( .A(n6739), .ZN(n6699) );
  OAI21_X1 U7692 ( .B1(n6735), .B2(n6699), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6700) );
  OAI211_X1 U7693 ( .C1(n6702), .C2(n6701), .A(n6700), .B(n6753), .ZN(n6707)
         );
  INV_X1 U7694 ( .A(n6734), .ZN(n6704) );
  AOI21_X1 U7695 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6704), .A(n6703), .ZN(
        n6705) );
  NAND3_X1 U7696 ( .A1(n6707), .A2(n6706), .A3(n6705), .ZN(n6736) );
  AOI22_X1 U7697 ( .A1(n6736), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6708), 
        .B2(n6735), .ZN(n6709) );
  OAI211_X1 U7698 ( .C1(n6742), .C2(n6739), .A(n6710), .B(n6709), .ZN(U3084)
         );
  AOI22_X1 U7699 ( .A1(n6711), .A2(n6734), .B1(n6764), .B2(n6733), .ZN(n6714)
         );
  AOI22_X1 U7700 ( .A1(n6736), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6712), 
        .B2(n6735), .ZN(n6713) );
  OAI211_X1 U7701 ( .C1(n6762), .C2(n6739), .A(n6714), .B(n6713), .ZN(U3085)
         );
  AOI22_X1 U7702 ( .A1(n6715), .A2(n6734), .B1(n6771), .B2(n6733), .ZN(n6718)
         );
  AOI22_X1 U7703 ( .A1(n6736), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6716), 
        .B2(n6735), .ZN(n6717) );
  OAI211_X1 U7704 ( .C1(n6769), .C2(n6739), .A(n6718), .B(n6717), .ZN(U3086)
         );
  AOI22_X1 U7705 ( .A1(n6719), .A2(n6734), .B1(n6778), .B2(n6733), .ZN(n6722)
         );
  AOI22_X1 U7706 ( .A1(n6736), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6720), 
        .B2(n6735), .ZN(n6721) );
  OAI211_X1 U7707 ( .C1(n6776), .C2(n6739), .A(n6722), .B(n6721), .ZN(U3087)
         );
  AOI22_X1 U7708 ( .A1(n6723), .A2(n6734), .B1(n7373), .B2(n6733), .ZN(n6726)
         );
  AOI22_X1 U7709 ( .A1(n6736), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6724), 
        .B2(n6735), .ZN(n6725) );
  OAI211_X1 U7710 ( .C1(n7378), .C2(n6739), .A(n6726), .B(n6725), .ZN(U3088)
         );
  AOI22_X1 U7711 ( .A1(n6727), .A2(n6734), .B1(n6785), .B2(n6733), .ZN(n6730)
         );
  AOI22_X1 U7712 ( .A1(n6736), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6728), 
        .B2(n6735), .ZN(n6729) );
  OAI211_X1 U7713 ( .C1(n6783), .C2(n6739), .A(n6730), .B(n6729), .ZN(U3089)
         );
  AOI22_X1 U7714 ( .A1(n6800), .A2(n6734), .B1(n6799), .B2(n6733), .ZN(n6732)
         );
  AOI22_X1 U7715 ( .A1(n6736), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6801), 
        .B2(n6735), .ZN(n6731) );
  OAI211_X1 U7716 ( .C1(n6804), .C2(n6739), .A(n6732), .B(n6731), .ZN(U3090)
         );
  AOI22_X1 U7717 ( .A1(n6808), .A2(n6734), .B1(n6806), .B2(n6733), .ZN(n6738)
         );
  AOI22_X1 U7718 ( .A1(n6736), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6810), 
        .B2(n6735), .ZN(n6737) );
  OAI211_X1 U7719 ( .C1(n6814), .C2(n6739), .A(n6738), .B(n6737), .ZN(U3091)
         );
  NOR2_X1 U7720 ( .A1(n6850), .A2(n6740), .ZN(n6746) );
  INV_X1 U7721 ( .A(n6746), .ZN(n7367) );
  OAI22_X1 U7722 ( .A1(n7377), .A2(n6742), .B1(n6741), .B2(n7367), .ZN(n6743)
         );
  INV_X1 U7723 ( .A(n6743), .ZN(n6759) );
  INV_X1 U7724 ( .A(n6756), .ZN(n6750) );
  NAND2_X1 U7725 ( .A1(n6745), .A2(n6744), .ZN(n6754) );
  AOI21_X1 U7726 ( .B1(n6747), .B2(n6833), .A(n6746), .ZN(n6751) );
  NAND3_X1 U7727 ( .A1(n6754), .A2(n6753), .A3(n6751), .ZN(n6748) );
  OAI211_X1 U7728 ( .C1(n6753), .C2(n6750), .A(n6749), .B(n6748), .ZN(n7374)
         );
  INV_X1 U7729 ( .A(n6751), .ZN(n6752) );
  NAND3_X1 U7730 ( .A1(n6754), .A2(n6753), .A3(n6752), .ZN(n6755) );
  OAI21_X1 U7731 ( .B1(n6756), .B2(n3658), .A(n6755), .ZN(n7372) );
  AOI22_X1 U7732 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n7374), .B1(n6757), 
        .B2(n7372), .ZN(n6758) );
  OAI211_X1 U7733 ( .C1(n6760), .C2(n7370), .A(n6759), .B(n6758), .ZN(U3108)
         );
  OAI22_X1 U7734 ( .A1(n7377), .A2(n6762), .B1(n6761), .B2(n7367), .ZN(n6763)
         );
  INV_X1 U7735 ( .A(n6763), .ZN(n6766) );
  AOI22_X1 U7736 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n7374), .B1(n6764), 
        .B2(n7372), .ZN(n6765) );
  OAI211_X1 U7737 ( .C1(n6767), .C2(n7370), .A(n6766), .B(n6765), .ZN(U3109)
         );
  OAI22_X1 U7738 ( .A1(n7377), .A2(n6769), .B1(n6768), .B2(n7367), .ZN(n6770)
         );
  INV_X1 U7739 ( .A(n6770), .ZN(n6773) );
  AOI22_X1 U7740 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n7374), .B1(n6771), 
        .B2(n7372), .ZN(n6772) );
  OAI211_X1 U7741 ( .C1(n6774), .C2(n7370), .A(n6773), .B(n6772), .ZN(U3110)
         );
  OAI22_X1 U7742 ( .A1(n7377), .A2(n6776), .B1(n6775), .B2(n7367), .ZN(n6777)
         );
  INV_X1 U7743 ( .A(n6777), .ZN(n6780) );
  AOI22_X1 U7744 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n7374), .B1(n6778), 
        .B2(n7372), .ZN(n6779) );
  OAI211_X1 U7745 ( .C1(n6781), .C2(n7370), .A(n6780), .B(n6779), .ZN(U3111)
         );
  OAI22_X1 U7746 ( .A1(n7377), .A2(n6783), .B1(n6782), .B2(n7367), .ZN(n6784)
         );
  INV_X1 U7747 ( .A(n6784), .ZN(n6787) );
  AOI22_X1 U7748 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n7374), .B1(n6785), 
        .B2(n7372), .ZN(n6786) );
  OAI211_X1 U7749 ( .C1(n6788), .C2(n7370), .A(n6787), .B(n6786), .ZN(U3113)
         );
  OAI22_X1 U7750 ( .A1(n7370), .A2(n6790), .B1(n6789), .B2(n7367), .ZN(n6791)
         );
  INV_X1 U7751 ( .A(n6791), .ZN(n6793) );
  AOI22_X1 U7752 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n7374), .B1(n6799), 
        .B2(n7372), .ZN(n6792) );
  OAI211_X1 U7753 ( .C1(n6804), .C2(n7377), .A(n6793), .B(n6792), .ZN(U3114)
         );
  OAI22_X1 U7754 ( .A1(n7370), .A2(n6795), .B1(n6794), .B2(n7367), .ZN(n6796)
         );
  INV_X1 U7755 ( .A(n6796), .ZN(n6798) );
  AOI22_X1 U7756 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n7374), .B1(n6806), 
        .B2(n7372), .ZN(n6797) );
  OAI211_X1 U7757 ( .C1(n6814), .C2(n7377), .A(n6798), .B(n6797), .ZN(U3115)
         );
  AOI22_X1 U7758 ( .A1(n6800), .A2(n6807), .B1(n6799), .B2(n6805), .ZN(n6803)
         );
  AOI22_X1 U7759 ( .A1(n6811), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6801), 
        .B2(n6809), .ZN(n6802) );
  OAI211_X1 U7760 ( .C1(n6804), .C2(n7370), .A(n6803), .B(n6802), .ZN(U3122)
         );
  AOI22_X1 U7761 ( .A1(n6808), .A2(n6807), .B1(n6806), .B2(n6805), .ZN(n6813)
         );
  AOI22_X1 U7762 ( .A1(n6811), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6810), 
        .B2(n6809), .ZN(n6812) );
  OAI211_X1 U7763 ( .C1(n6814), .C2(n7370), .A(n6813), .B(n6812), .ZN(U3123)
         );
  OAI21_X1 U7764 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6815), 
        .ZN(n6827) );
  INV_X1 U7765 ( .A(n6816), .ZN(n6826) );
  OR2_X1 U7766 ( .A1(n6817), .A2(n6822), .ZN(n6824) );
  AOI22_X1 U7767 ( .A1(n6822), .A2(n6821), .B1(n6820), .B2(n6819), .ZN(n6823)
         );
  AND2_X1 U7768 ( .A1(n6824), .A2(n6823), .ZN(n6977) );
  NAND4_X1 U7769 ( .A1(n6827), .A2(n6826), .A3(n6977), .A4(n6825), .ZN(n6828)
         );
  NOR2_X1 U7770 ( .A1(n6829), .A2(n6828), .ZN(n6852) );
  AOI22_X1 U7771 ( .A1(n6833), .A2(n6832), .B1(n6831), .B2(n6830), .ZN(n6956)
         );
  NAND2_X1 U7772 ( .A1(n6834), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6961) );
  NAND3_X1 U7773 ( .A1(n6956), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6961), .ZN(n6837) );
  OAI211_X1 U7774 ( .C1(n6838), .C2(n6837), .A(n6836), .B(n6835), .ZN(n6840)
         );
  NAND2_X1 U7775 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  NAND2_X1 U7776 ( .A1(n6840), .A2(n6839), .ZN(n6845) );
  NAND2_X1 U7777 ( .A1(n6844), .A2(n6845), .ZN(n6841) );
  NAND2_X1 U7778 ( .A1(n6842), .A2(n6841), .ZN(n6843) );
  OAI21_X1 U7779 ( .B1(n6845), .B2(n6844), .A(n6843), .ZN(n6847) );
  NAND2_X1 U7780 ( .A1(n6849), .A2(n6850), .ZN(n6846) );
  NAND2_X1 U7781 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  OAI211_X1 U7782 ( .C1(n6850), .C2(n6849), .A(n6848), .B(n7293), .ZN(n6851)
         );
  AND2_X1 U7783 ( .A1(n6852), .A2(n6851), .ZN(n6866) );
  NAND2_X1 U7784 ( .A1(n6866), .A2(n6867), .ZN(n6854) );
  NAND2_X1 U7785 ( .A1(READY_N), .A2(n6982), .ZN(n6853) );
  NAND2_X1 U7786 ( .A1(n6854), .A2(n6853), .ZN(n6858) );
  OR2_X1 U7787 ( .A1(n6856), .A2(n6855), .ZN(n6857) );
  OAI21_X1 U7788 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6981), .A(n6946), .ZN(
        n6870) );
  AOI221_X1 U7789 ( .B1(n6860), .B2(STATE2_REG_0__SCAN_IN), .C1(n6870), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6859), .ZN(n6864) );
  OAI211_X1 U7790 ( .C1(n6862), .C2(n6953), .A(n6861), .B(n6946), .ZN(n6863)
         );
  OAI211_X1 U7791 ( .C1(n6866), .C2(n6865), .A(n6864), .B(n6863), .ZN(U3148)
         );
  AOI21_X1 U7792 ( .B1(n6868), .B2(n6981), .A(n6867), .ZN(n6873) );
  INV_X1 U7793 ( .A(n6869), .ZN(n6872) );
  OAI211_X1 U7794 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6870), .ZN(n6871) );
  OAI211_X1 U7795 ( .C1(n6874), .C2(n6873), .A(n6872), .B(n6871), .ZN(U3149)
         );
  OAI221_X1 U7796 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6981), .A(n6944), .ZN(n6876) );
  OAI21_X1 U7797 ( .B1(n6985), .B2(n6876), .A(n6875), .ZN(U3150) );
  AND2_X1 U7798 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6939), .ZN(U3151) );
  AND2_X1 U7799 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6939), .ZN(U3152) );
  AND2_X1 U7800 ( .A1(n6939), .A2(DATAWIDTH_REG_29__SCAN_IN), .ZN(U3153) );
  AND2_X1 U7801 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6939), .ZN(U3154) );
  INV_X1 U7802 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n7201) );
  NOR2_X1 U7803 ( .A1(n6942), .A2(n7201), .ZN(U3155) );
  AND2_X1 U7804 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6939), .ZN(U3156) );
  AND2_X1 U7805 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6939), .ZN(U3157) );
  AND2_X1 U7806 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6939), .ZN(U3158) );
  NOR2_X1 U7807 ( .A1(n6942), .A2(n7307), .ZN(U3159) );
  AND2_X1 U7808 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6939), .ZN(U3160) );
  AND2_X1 U7809 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6939), .ZN(U3161) );
  AND2_X1 U7810 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6939), .ZN(U3162) );
  AND2_X1 U7811 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6939), .ZN(U3163) );
  INV_X1 U7812 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7239) );
  NOR2_X1 U7813 ( .A1(n6942), .A2(n7239), .ZN(U3164) );
  AND2_X1 U7814 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6939), .ZN(U3165) );
  NOR2_X1 U7815 ( .A1(n6942), .A2(n7246), .ZN(U3166) );
  INV_X1 U7816 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7135) );
  NOR2_X1 U7817 ( .A1(n6942), .A2(n7135), .ZN(U3167) );
  AND2_X1 U7818 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6939), .ZN(U3168) );
  AND2_X1 U7819 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6939), .ZN(U3169) );
  AND2_X1 U7820 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6939), .ZN(U3170) );
  AND2_X1 U7821 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6939), .ZN(U3171) );
  AND2_X1 U7822 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6939), .ZN(U3172) );
  AND2_X1 U7823 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6939), .ZN(U3173) );
  AND2_X1 U7824 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6939), .ZN(U3174) );
  AND2_X1 U7825 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6939), .ZN(U3175) );
  AND2_X1 U7826 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6939), .ZN(U3176) );
  INV_X1 U7827 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7137) );
  NOR2_X1 U7828 ( .A1(n6942), .A2(n7137), .ZN(U3177) );
  AND2_X1 U7829 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6939), .ZN(U3178) );
  AND2_X1 U7830 ( .A1(n6939), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7831 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6939), .ZN(U3180) );
  NAND2_X1 U7832 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6885) );
  NAND2_X1 U7833 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6880) );
  NAND2_X1 U7834 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6882) );
  OAI21_X1 U7835 ( .B1(n6877), .B2(n6981), .A(n6882), .ZN(n6879) );
  INV_X1 U7836 ( .A(NA_N), .ZN(n6878) );
  AOI221_X1 U7837 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6878), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6893) );
  AOI21_X1 U7838 ( .B1(n6880), .B2(n6879), .A(n6893), .ZN(n6881) );
  OAI221_X1 U7839 ( .B1(n3194), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n3194), 
        .C2(n6885), .A(n6881), .ZN(U3181) );
  INV_X1 U7840 ( .A(n6882), .ZN(n6886) );
  NAND2_X1 U7841 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6889) );
  AOI21_X1 U7842 ( .B1(STATE_REG_1__SCAN_IN), .B2(READY_N), .A(n6883), .ZN(
        n6884) );
  OAI221_X1 U7843 ( .B1(n6886), .B2(n6889), .C1(n6886), .C2(n6885), .A(n6884), 
        .ZN(U3182) );
  AOI221_X1 U7844 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6981), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6887) );
  OAI21_X1 U7845 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6887), .A(HOLD), .ZN(n6892)
         );
  OAI21_X1 U7846 ( .B1(NA_N), .B2(n6889), .A(n6888), .ZN(n6890) );
  NAND3_X1 U7847 ( .A1(READY_N), .A2(n6890), .A3(STATE_REG_1__SCAN_IN), .ZN(
        n6891) );
  OAI221_X1 U7848 ( .B1(n6893), .B2(STATE_REG_0__SCAN_IN), .C1(n6893), .C2(
        n6892), .A(n6891), .ZN(U3183) );
  NAND2_X1 U7849 ( .A1(STATE_REG_2__SCAN_IN), .A2(n3194), .ZN(n6934) );
  NOR2_X1 U7850 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6936), .ZN(n6932) );
  AOI22_X1 U7851 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6936), .ZN(n6894) );
  OAI21_X1 U7852 ( .B1(n6895), .B2(n6934), .A(n6894), .ZN(U3184) );
  AOI22_X1 U7853 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6936), .ZN(n6896) );
  OAI21_X1 U7854 ( .B1(n7306), .B2(n6934), .A(n6896), .ZN(U3185) );
  AOI22_X1 U7855 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6936), .ZN(n6897) );
  OAI21_X1 U7856 ( .B1(n7300), .B2(n6934), .A(n6897), .ZN(U3186) );
  INV_X1 U7857 ( .A(n6934), .ZN(n6929) );
  AOI22_X1 U7858 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6974), .ZN(n6898) );
  OAI21_X1 U7859 ( .B1(n6899), .B2(n6931), .A(n6898), .ZN(U3187) );
  INV_X1 U7860 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7283) );
  OAI222_X1 U7861 ( .A1(n6934), .A2(n6899), .B1(n7283), .B2(n3194), .C1(n6900), 
        .C2(n6931), .ZN(U3188) );
  INV_X1 U7862 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7161) );
  OAI222_X1 U7863 ( .A1(n6934), .A2(n6900), .B1(n7161), .B2(n3194), .C1(n7187), 
        .C2(n6931), .ZN(U3189) );
  INV_X1 U7864 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6902) );
  AOI22_X1 U7865 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6974), .ZN(n6901) );
  OAI21_X1 U7866 ( .B1(n6902), .B2(n6931), .A(n6901), .ZN(U3190) );
  AOI22_X1 U7867 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6974), .ZN(n6903) );
  OAI21_X1 U7868 ( .B1(n6905), .B2(n6931), .A(n6903), .ZN(U3191) );
  AOI22_X1 U7869 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6974), .ZN(n6904) );
  OAI21_X1 U7870 ( .B1(n6905), .B2(n6934), .A(n6904), .ZN(U3192) );
  AOI22_X1 U7871 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6974), .ZN(n6906) );
  OAI21_X1 U7872 ( .B1(n7240), .B2(n6931), .A(n6906), .ZN(U3193) );
  AOI22_X1 U7873 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6974), .ZN(n6907) );
  OAI21_X1 U7874 ( .B1(n7240), .B2(n6934), .A(n6907), .ZN(U3194) );
  AOI22_X1 U7875 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6974), .ZN(n6908) );
  OAI21_X1 U7876 ( .B1(n6909), .B2(n6931), .A(n6908), .ZN(U3195) );
  AOI22_X1 U7877 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6936), .ZN(n6910) );
  OAI21_X1 U7878 ( .B1(n7268), .B2(n6931), .A(n6910), .ZN(U3196) );
  AOI22_X1 U7879 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6936), .ZN(n6911) );
  OAI21_X1 U7880 ( .B1(n7268), .B2(n6934), .A(n6911), .ZN(U3197) );
  INV_X1 U7881 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7282) );
  OAI222_X1 U7882 ( .A1(n6934), .A2(n6912), .B1(n7282), .B2(n3194), .C1(n5940), 
        .C2(n6931), .ZN(U3198) );
  INV_X1 U7883 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7149) );
  OAI222_X1 U7884 ( .A1(n6934), .A2(n5940), .B1(n7149), .B2(n3194), .C1(n6913), 
        .C2(n6931), .ZN(U3199) );
  INV_X1 U7885 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7245) );
  OAI222_X1 U7886 ( .A1(n6931), .A2(n6915), .B1(n7245), .B2(n3194), .C1(n6913), 
        .C2(n6934), .ZN(U3200) );
  INV_X1 U7887 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7115) );
  OAI222_X1 U7888 ( .A1(n6934), .A2(n6915), .B1(n7115), .B2(n3194), .C1(n6914), 
        .C2(n6931), .ZN(U3201) );
  AOI22_X1 U7889 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6936), .ZN(n6916) );
  OAI21_X1 U7890 ( .B1(n7291), .B2(n6931), .A(n6916), .ZN(U3202) );
  AOI22_X1 U7891 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6936), .ZN(n6917) );
  OAI21_X1 U7892 ( .B1(n7291), .B2(n6934), .A(n6917), .ZN(U3203) );
  INV_X1 U7893 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7172) );
  OAI222_X1 U7894 ( .A1(n6934), .A2(n6918), .B1(n7172), .B2(n3194), .C1(n7203), 
        .C2(n6931), .ZN(U3204) );
  AOI22_X1 U7895 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6936), .ZN(n6919) );
  OAI21_X1 U7896 ( .B1(n7203), .B2(n6934), .A(n6919), .ZN(U3205) );
  AOI22_X1 U7897 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6936), .ZN(n6920) );
  OAI21_X1 U7898 ( .B1(n6921), .B2(n6931), .A(n6920), .ZN(U3206) );
  INV_X1 U7899 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7285) );
  OAI222_X1 U7900 ( .A1(n6931), .A2(n6923), .B1(n7285), .B2(n3194), .C1(n6921), 
        .C2(n6934), .ZN(U3207) );
  AOI22_X1 U7901 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6974), .ZN(n6922) );
  OAI21_X1 U7902 ( .B1(n6923), .B2(n6934), .A(n6922), .ZN(U3208) );
  AOI22_X1 U7903 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6936), .ZN(n6924) );
  OAI21_X1 U7904 ( .B1(n6925), .B2(n6931), .A(n6924), .ZN(U3209) );
  INV_X1 U7905 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7177) );
  OAI222_X1 U7906 ( .A1(n6934), .A2(n6925), .B1(n7177), .B2(n3194), .C1(n6928), 
        .C2(n6931), .ZN(U3210) );
  INV_X1 U7907 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6927) );
  OAI222_X1 U7908 ( .A1(n6934), .A2(n6928), .B1(n6927), .B2(n3194), .C1(n6926), 
        .C2(n6931), .ZN(U3211) );
  INV_X1 U7909 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6935) );
  AOI22_X1 U7910 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6929), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6936), .ZN(n6930) );
  OAI21_X1 U7911 ( .B1(n6935), .B2(n6931), .A(n6930), .ZN(U3212) );
  AOI22_X1 U7912 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6932), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6936), .ZN(n6933) );
  OAI21_X1 U7913 ( .B1(n6935), .B2(n6934), .A(n6933), .ZN(U3213) );
  MUX2_X1 U7914 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n3194), .Z(U3445) );
  MUX2_X1 U7915 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n3194), .Z(U3446) );
  MUX2_X1 U7916 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n3194), .Z(U3447) );
  OAI22_X1 U7917 ( .A1(n6936), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n3194), .ZN(n6937) );
  INV_X1 U7918 ( .A(n6937), .ZN(U3448) );
  INV_X1 U7919 ( .A(n6940), .ZN(n6938) );
  AOI21_X1 U7920 ( .B1(n6968), .B2(n6939), .A(n6938), .ZN(U3451) );
  OAI21_X1 U7921 ( .B1(n6942), .B2(n6941), .A(n6940), .ZN(U3452) );
  INV_X1 U7922 ( .A(n6943), .ZN(n6945) );
  OAI211_X1 U7923 ( .C1(n7315), .C2(n6946), .A(n6945), .B(n6944), .ZN(U3453)
         );
  INV_X1 U7924 ( .A(n6947), .ZN(n6949) );
  OAI22_X1 U7925 ( .A1(n6949), .A2(n6962), .B1(n6948), .B2(n6953), .ZN(n6950)
         );
  OAI22_X1 U7926 ( .A1(n6957), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n6950), .B2(n6959), .ZN(n6951) );
  INV_X1 U7927 ( .A(n6951), .ZN(U3456) );
  OAI22_X1 U7928 ( .A1(n6953), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6952), .ZN(n6954) );
  INV_X1 U7929 ( .A(n6954), .ZN(n6955) );
  OAI21_X1 U7930 ( .B1(n6956), .B2(n6962), .A(n6955), .ZN(n6958) );
  AOI22_X1 U7931 ( .A1(n6959), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n6958), .B2(n6957), .ZN(n6960) );
  OAI21_X1 U7932 ( .B1(n6962), .B2(n6961), .A(n6960), .ZN(U3461) );
  NAND2_X1 U7933 ( .A1(n6963), .A2(n6964), .ZN(n6970) );
  NOR2_X1 U7934 ( .A1(n6966), .A2(n6964), .ZN(n6965) );
  AOI22_X1 U7935 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6966), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6965), .ZN(n6967) );
  OAI221_X1 U7936 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6969), .C1(n6968), 
        .C2(n6970), .A(n6967), .ZN(U3468) );
  OAI21_X1 U7937 ( .B1(n6971), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6970), .ZN(
        n6972) );
  INV_X1 U7938 ( .A(n6972), .ZN(U3469) );
  NAND2_X1 U7939 ( .A1(n6974), .A2(W_R_N_REG_SCAN_IN), .ZN(n6973) );
  OAI21_X1 U7940 ( .B1(n6974), .B2(READREQUEST_REG_SCAN_IN), .A(n6973), .ZN(
        U3470) );
  INV_X1 U7941 ( .A(MORE_REG_SCAN_IN), .ZN(n6976) );
  INV_X1 U7942 ( .A(n6978), .ZN(n6975) );
  AOI22_X1 U7943 ( .A1(n6978), .A2(n6977), .B1(n6976), .B2(n6975), .ZN(U3471)
         );
  AOI211_X1 U7944 ( .C1(n6982), .C2(n6981), .A(n6980), .B(n6979), .ZN(n6989)
         );
  OAI211_X1 U7945 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6984), .A(n6983), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6986) );
  AOI21_X1 U7946 ( .B1(n6986), .B2(STATE2_REG_0__SCAN_IN), .A(n6985), .ZN(
        n6988) );
  NAND2_X1 U7947 ( .A1(n6989), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6987) );
  OAI21_X1 U7948 ( .B1(n6989), .B2(n6988), .A(n6987), .ZN(U3472) );
  MUX2_X1 U7949 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n3194), .Z(U3473) );
  OAI22_X1 U7950 ( .A1(EBX_REG_25__SCAN_IN), .A2(keyinput27), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput44), .ZN(n6991) );
  AOI221_X1 U7951 ( .B1(EBX_REG_25__SCAN_IN), .B2(keyinput27), .C1(keyinput44), 
        .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n6991), .ZN(n6998) );
  OAI22_X1 U7952 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput99), .B1(
        keyinput84), .B2(DATAO_REG_16__SCAN_IN), .ZN(n6992) );
  AOI221_X1 U7953 ( .B1(INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput99), .C1(
        DATAO_REG_16__SCAN_IN), .C2(keyinput84), .A(n6992), .ZN(n6997) );
  OAI22_X1 U7954 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(keyinput71), .B1(
        keyinput62), .B2(ADDRESS_REG_27__SCAN_IN), .ZN(n6993) );
  AOI221_X1 U7955 ( .B1(INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput71), .C1(
        ADDRESS_REG_27__SCAN_IN), .C2(keyinput62), .A(n6993), .ZN(n6996) );
  OAI22_X1 U7956 ( .A1(DATAI_2_), .A2(keyinput56), .B1(keyinput121), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n6994) );
  AOI221_X1 U7957 ( .B1(DATAI_2_), .B2(keyinput56), .C1(DATAO_REG_20__SCAN_IN), 
        .C2(keyinput121), .A(n6994), .ZN(n6995) );
  NAND4_X1 U7958 ( .A1(n6998), .A2(n6997), .A3(n6996), .A4(n6995), .ZN(n7026)
         );
  OAI22_X1 U7959 ( .A1(EBX_REG_12__SCAN_IN), .A2(keyinput47), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput46), .ZN(n6999) );
  AOI221_X1 U7960 ( .B1(EBX_REG_12__SCAN_IN), .B2(keyinput47), .C1(keyinput46), 
        .C2(ADDRESS_REG_15__SCAN_IN), .A(n6999), .ZN(n7006) );
  OAI22_X1 U7961 ( .A1(UWORD_REG_11__SCAN_IN), .A2(keyinput49), .B1(keyinput38), .B2(UWORD_REG_13__SCAN_IN), .ZN(n7000) );
  AOI221_X1 U7962 ( .B1(UWORD_REG_11__SCAN_IN), .B2(keyinput49), .C1(
        UWORD_REG_13__SCAN_IN), .C2(keyinput38), .A(n7000), .ZN(n7005) );
  OAI22_X1 U7963 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(keyinput67), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput61), .ZN(n7001) );
  AOI221_X1 U7964 ( .B1(INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput67), .C1(
        keyinput61), .C2(BE_N_REG_0__SCAN_IN), .A(n7001), .ZN(n7004) );
  OAI22_X1 U7965 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput9), .B1(
        keyinput29), .B2(ADDRESS_REG_5__SCAN_IN), .ZN(n7002) );
  AOI221_X1 U7966 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput9), .C1(
        ADDRESS_REG_5__SCAN_IN), .C2(keyinput29), .A(n7002), .ZN(n7003) );
  NAND4_X1 U7967 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .ZN(n7025)
         );
  OAI22_X1 U7968 ( .A1(LWORD_REG_0__SCAN_IN), .A2(keyinput104), .B1(
        UWORD_REG_6__SCAN_IN), .B2(keyinput82), .ZN(n7007) );
  AOI221_X1 U7969 ( .B1(LWORD_REG_0__SCAN_IN), .B2(keyinput104), .C1(
        keyinput82), .C2(UWORD_REG_6__SCAN_IN), .A(n7007), .ZN(n7014) );
  OAI22_X1 U7970 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(keyinput24), .B1(
        keyinput13), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7008) );
  AOI221_X1 U7971 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput24), 
        .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(keyinput13), .A(n7008), .ZN(
        n7013) );
  OAI22_X1 U7972 ( .A1(n7151), .A2(keyinput6), .B1(keyinput14), .B2(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n7009) );
  AOI221_X1 U7973 ( .B1(n7151), .B2(keyinput6), .C1(DATAWIDTH_REG_29__SCAN_IN), 
        .C2(keyinput14), .A(n7009), .ZN(n7012) );
  OAI22_X1 U7974 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(keyinput12), .B1(
        REIP_REG_7__SCAN_IN), .B2(keyinput74), .ZN(n7010) );
  AOI221_X1 U7975 ( .B1(INSTQUEUE_REG_10__3__SCAN_IN), .B2(keyinput12), .C1(
        keyinput74), .C2(REIP_REG_7__SCAN_IN), .A(n7010), .ZN(n7011) );
  NAND4_X1 U7976 ( .A1(n7014), .A2(n7013), .A3(n7012), .A4(n7011), .ZN(n7024)
         );
  OAI22_X1 U7977 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(keyinput113), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(keyinput70), .ZN(n7015) );
  AOI221_X1 U7978 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput113), .C1(
        keyinput70), .C2(ADDRESS_REG_26__SCAN_IN), .A(n7015), .ZN(n7022) );
  OAI22_X1 U7979 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(keyinput51), .B1(
        keyinput101), .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n7016) );
  AOI221_X1 U7980 ( .B1(INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput51), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput101), .A(n7016), .ZN(n7021)
         );
  OAI22_X1 U7981 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput10), .B1(
        keyinput31), .B2(DATAO_REG_26__SCAN_IN), .ZN(n7017) );
  AOI221_X1 U7982 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput10), 
        .C1(DATAO_REG_26__SCAN_IN), .C2(keyinput31), .A(n7017), .ZN(n7020) );
  OAI22_X1 U7983 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(keyinput5), .B1(
        keyinput98), .B2(EBX_REG_15__SCAN_IN), .ZN(n7018) );
  AOI221_X1 U7984 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput5), .C1(
        EBX_REG_15__SCAN_IN), .C2(keyinput98), .A(n7018), .ZN(n7019) );
  NAND4_X1 U7985 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n7023)
         );
  NOR4_X1 U7986 ( .A1(n7026), .A2(n7025), .A3(n7024), .A4(n7023), .ZN(n7366)
         );
  AOI22_X1 U7987 ( .A1(DATAI_2_), .A2(keyinput184), .B1(
        INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput145), .ZN(n7027) );
  OAI221_X1 U7988 ( .B1(DATAI_2_), .B2(keyinput184), .C1(
        INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput145), .A(n7027), .ZN(n7034)
         );
  AOI22_X1 U7989 ( .A1(DATAO_REG_15__SCAN_IN), .A2(keyinput186), .B1(
        EAX_REG_20__SCAN_IN), .B2(keyinput246), .ZN(n7028) );
  OAI221_X1 U7990 ( .B1(DATAO_REG_15__SCAN_IN), .B2(keyinput186), .C1(
        EAX_REG_20__SCAN_IN), .C2(keyinput246), .A(n7028), .ZN(n7033) );
  AOI22_X1 U7991 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput153), .B1(
        INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput199), .ZN(n7029) );
  OAI221_X1 U7992 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput153), .C1(
        INSTQUEUE_REG_7__7__SCAN_IN), .C2(keyinput199), .A(n7029), .ZN(n7032)
         );
  AOI22_X1 U7993 ( .A1(UWORD_REG_11__SCAN_IN), .A2(keyinput177), .B1(
        REIP_REG_2__SCAN_IN), .B2(keyinput196), .ZN(n7030) );
  OAI221_X1 U7994 ( .B1(UWORD_REG_11__SCAN_IN), .B2(keyinput177), .C1(
        REIP_REG_2__SCAN_IN), .C2(keyinput196), .A(n7030), .ZN(n7031) );
  NOR4_X1 U7995 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n7062)
         );
  AOI22_X1 U7996 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(keyinput251), .B1(
        n4955), .B2(keyinput158), .ZN(n7035) );
  OAI221_X1 U7997 ( .B1(INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput251), .C1(
        n4955), .C2(keyinput158), .A(n7035), .ZN(n7042) );
  AOI22_X1 U7998 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput180), .B1(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput200), .ZN(n7036) );
  OAI221_X1 U7999 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput180), .C1(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(keyinput200), .A(n7036), .ZN(
        n7041) );
  AOI22_X1 U8000 ( .A1(ADDRESS_REG_4__SCAN_IN), .A2(keyinput250), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput234), .ZN(n7037) );
  OAI221_X1 U8001 ( .B1(ADDRESS_REG_4__SCAN_IN), .B2(keyinput250), .C1(
        DATAWIDTH_REG_18__SCAN_IN), .C2(keyinput234), .A(n7037), .ZN(n7040) );
  AOI22_X1 U8002 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput214), 
        .B1(INSTQUEUE_REG_6__3__SCAN_IN), .B2(keyinput168), .ZN(n7038) );
  OAI221_X1 U8003 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput214), 
        .C1(INSTQUEUE_REG_6__3__SCAN_IN), .C2(keyinput168), .A(n7038), .ZN(
        n7039) );
  NOR4_X1 U8004 ( .A1(n7042), .A2(n7041), .A3(n7040), .A4(n7039), .ZN(n7061)
         );
  AOI22_X1 U8005 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput205), .B1(
        INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput179), .ZN(n7043) );
  OAI221_X1 U8006 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput205), .C1(
        INSTQUEUE_REG_4__1__SCAN_IN), .C2(keyinput179), .A(n7043), .ZN(n7050)
         );
  AOI22_X1 U8007 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput150), 
        .B1(INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput192), .ZN(n7044) );
  OAI221_X1 U8008 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput150), 
        .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(keyinput192), .A(n7044), .ZN(
        n7049) );
  AOI22_X1 U8009 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput238), .B1(
        INSTQUEUE_REG_10__3__SCAN_IN), .B2(keyinput140), .ZN(n7045) );
  OAI221_X1 U8010 ( .B1(PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput238), 
        .C1(INSTQUEUE_REG_10__3__SCAN_IN), .C2(keyinput140), .A(n7045), .ZN(
        n7048) );
  AOI22_X1 U8011 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(keyinput195), .B1(
        INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput149), .ZN(n7046) );
  OAI221_X1 U8012 ( .B1(INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput195), .C1(
        INSTQUEUE_REG_11__5__SCAN_IN), .C2(keyinput149), .A(n7046), .ZN(n7047)
         );
  NOR4_X1 U8013 ( .A1(n7050), .A2(n7049), .A3(n7048), .A4(n7047), .ZN(n7060)
         );
  AOI22_X1 U8014 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput220), .B1(
        INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput165), .ZN(n7051) );
  OAI221_X1 U8015 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput220), .C1(
        INSTQUEUE_REG_5__1__SCAN_IN), .C2(keyinput165), .A(n7051), .ZN(n7058)
         );
  AOI22_X1 U8016 ( .A1(DATAI_19_), .A2(keyinput144), .B1(
        INSTQUEUE_REG_13__1__SCAN_IN), .B2(keyinput203), .ZN(n7052) );
  OAI221_X1 U8017 ( .B1(DATAI_19_), .B2(keyinput144), .C1(
        INSTQUEUE_REG_13__1__SCAN_IN), .C2(keyinput203), .A(n7052), .ZN(n7057)
         );
  AOI22_X1 U8018 ( .A1(LWORD_REG_0__SCAN_IN), .A2(keyinput232), .B1(
        DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput131), .ZN(n7053) );
  OAI221_X1 U8019 ( .B1(LWORD_REG_0__SCAN_IN), .B2(keyinput232), .C1(
        DATAWIDTH_REG_3__SCAN_IN), .C2(keyinput131), .A(n7053), .ZN(n7056) );
  AOI22_X1 U8020 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(keyinput219), .B1(
        DATAO_REG_27__SCAN_IN), .B2(keyinput240), .ZN(n7054) );
  OAI221_X1 U8021 ( .B1(ADDRESS_REG_14__SCAN_IN), .B2(keyinput219), .C1(
        DATAO_REG_27__SCAN_IN), .C2(keyinput240), .A(n7054), .ZN(n7055) );
  NOR4_X1 U8022 ( .A1(n7058), .A2(n7057), .A3(n7056), .A4(n7055), .ZN(n7059)
         );
  NAND4_X1 U8023 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n7199)
         );
  AOI22_X1 U8024 ( .A1(EAX_REG_0__SCAN_IN), .A2(keyinput239), .B1(
        INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput201), .ZN(n7063) );
  OAI221_X1 U8025 ( .B1(EAX_REG_0__SCAN_IN), .B2(keyinput239), .C1(
        INSTQUEUE_REG_1__6__SCAN_IN), .C2(keyinput201), .A(n7063), .ZN(n7070)
         );
  AOI22_X1 U8026 ( .A1(LWORD_REG_1__SCAN_IN), .A2(keyinput162), .B1(
        INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput227), .ZN(n7064) );
  OAI221_X1 U8027 ( .B1(LWORD_REG_1__SCAN_IN), .B2(keyinput162), .C1(
        INSTQUEUE_REG_13__0__SCAN_IN), .C2(keyinput227), .A(n7064), .ZN(n7069)
         );
  AOI22_X1 U8028 ( .A1(DATAI_31_), .A2(keyinput181), .B1(
        INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput148), .ZN(n7065) );
  OAI221_X1 U8029 ( .B1(DATAI_31_), .B2(keyinput181), .C1(
        INSTQUEUE_REG_4__7__SCAN_IN), .C2(keyinput148), .A(n7065), .ZN(n7068)
         );
  AOI22_X1 U8030 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput235), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput247), .ZN(n7066) );
  OAI221_X1 U8031 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput235), .C1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .C2(keyinput247), .A(n7066), .ZN(
        n7067) );
  NOR4_X1 U8032 ( .A1(n7070), .A2(n7069), .A3(n7068), .A4(n7067), .ZN(n7098)
         );
  AOI22_X1 U8033 ( .A1(DATAI_30_), .A2(keyinput171), .B1(
        INSTADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput187), .ZN(n7071) );
  OAI221_X1 U8034 ( .B1(DATAI_30_), .B2(keyinput171), .C1(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput187), .A(n7071), .ZN(
        n7078) );
  AOI22_X1 U8035 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput217), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput188), .ZN(n7072) );
  OAI221_X1 U8036 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput217), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput188), .A(n7072), .ZN(n7077) );
  AOI22_X1 U8037 ( .A1(REIP_REG_11__SCAN_IN), .A2(keyinput228), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput154), .ZN(n7073) );
  OAI221_X1 U8038 ( .B1(REIP_REG_11__SCAN_IN), .B2(keyinput228), .C1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput154), .A(n7073), .ZN(
        n7076) );
  AOI22_X1 U8039 ( .A1(EAX_REG_4__SCAN_IN), .A2(keyinput230), .B1(
        INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput139), .ZN(n7074) );
  OAI221_X1 U8040 ( .B1(EAX_REG_4__SCAN_IN), .B2(keyinput230), .C1(
        INSTQUEUE_REG_8__0__SCAN_IN), .C2(keyinput139), .A(n7074), .ZN(n7075)
         );
  NOR4_X1 U8041 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7097)
         );
  AOI22_X1 U8042 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput224), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput172), .ZN(n7079) );
  OAI221_X1 U8043 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput224), .C1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .C2(keyinput172), .A(n7079), .ZN(
        n7086) );
  AOI22_X1 U8044 ( .A1(DATAI_10_), .A2(keyinput209), .B1(EBX_REG_25__SCAN_IN), 
        .B2(keyinput155), .ZN(n7080) );
  OAI221_X1 U8045 ( .B1(DATAI_10_), .B2(keyinput209), .C1(EBX_REG_25__SCAN_IN), 
        .C2(keyinput155), .A(n7080), .ZN(n7085) );
  AOI22_X1 U8046 ( .A1(LWORD_REG_11__SCAN_IN), .A2(keyinput178), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput161), .ZN(n7081) );
  OAI221_X1 U8047 ( .B1(LWORD_REG_11__SCAN_IN), .B2(keyinput178), .C1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .C2(keyinput161), .A(n7081), .ZN(
        n7084) );
  AOI22_X1 U8048 ( .A1(REIP_REG_3__SCAN_IN), .A2(keyinput182), .B1(
        INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput204), .ZN(n7082) );
  OAI221_X1 U8049 ( .B1(REIP_REG_3__SCAN_IN), .B2(keyinput182), .C1(
        INSTQUEUE_REG_4__3__SCAN_IN), .C2(keyinput204), .A(n7082), .ZN(n7083)
         );
  NOR4_X1 U8050 ( .A1(n7086), .A2(n7085), .A3(n7084), .A4(n7083), .ZN(n7096)
         );
  AOI22_X1 U8051 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput191), .B1(
        INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput248), .ZN(n7087) );
  OAI221_X1 U8052 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput191), .C1(
        INSTQUEUE_REG_6__5__SCAN_IN), .C2(keyinput248), .A(n7087), .ZN(n7094)
         );
  AOI22_X1 U8053 ( .A1(BS16_N), .A2(keyinput215), .B1(STATE2_REG_3__SCAN_IN), 
        .B2(keyinput193), .ZN(n7088) );
  OAI221_X1 U8054 ( .B1(BS16_N), .B2(keyinput215), .C1(STATE2_REG_3__SCAN_IN), 
        .C2(keyinput193), .A(n7088), .ZN(n7093) );
  AOI22_X1 U8055 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(keyinput142), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput212), .ZN(n7089) );
  OAI221_X1 U8056 ( .B1(DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput142), .C1(
        DATAO_REG_16__SCAN_IN), .C2(keyinput212), .A(n7089), .ZN(n7092) );
  AOI22_X1 U8057 ( .A1(LWORD_REG_15__SCAN_IN), .A2(keyinput129), .B1(
        INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput229), .ZN(n7090) );
  OAI221_X1 U8058 ( .B1(LWORD_REG_15__SCAN_IN), .B2(keyinput129), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput229), .A(n7090), .ZN(n7091)
         );
  NOR4_X1 U8059 ( .A1(n7094), .A2(n7093), .A3(n7092), .A4(n7091), .ZN(n7095)
         );
  NAND4_X1 U8060 ( .A1(n7098), .A2(n7097), .A3(n7096), .A4(n7095), .ZN(n7198)
         );
  AOI22_X1 U8061 ( .A1(UWORD_REG_6__SCAN_IN), .A2(keyinput210), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput237), .ZN(n7099) );
  OAI221_X1 U8062 ( .B1(UWORD_REG_6__SCAN_IN), .B2(keyinput210), .C1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput237), .A(n7099), .ZN(
        n7106) );
  AOI22_X1 U8063 ( .A1(BE_N_REG_0__SCAN_IN), .A2(keyinput189), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput152), .ZN(n7100) );
  OAI221_X1 U8064 ( .B1(BE_N_REG_0__SCAN_IN), .B2(keyinput189), .C1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(keyinput152), .A(n7100), .ZN(
        n7105) );
  AOI22_X1 U8065 ( .A1(ADDRESS_REG_27__SCAN_IN), .A2(keyinput190), .B1(
        EBX_REG_21__SCAN_IN), .B2(keyinput231), .ZN(n7101) );
  OAI221_X1 U8066 ( .B1(ADDRESS_REG_27__SCAN_IN), .B2(keyinput190), .C1(
        EBX_REG_21__SCAN_IN), .C2(keyinput231), .A(n7101), .ZN(n7104) );
  AOI22_X1 U8067 ( .A1(DATAO_REG_8__SCAN_IN), .A2(keyinput236), .B1(n7310), 
        .B2(keyinput222), .ZN(n7102) );
  OAI221_X1 U8068 ( .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput236), .C1(n7310), 
        .C2(keyinput222), .A(n7102), .ZN(n7103) );
  NOR4_X1 U8069 ( .A1(n7106), .A2(n7105), .A3(n7104), .A4(n7103), .ZN(n7146)
         );
  INV_X1 U8070 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n7108) );
  AOI22_X1 U8071 ( .A1(n7254), .A2(keyinput130), .B1(keyinput173), .B2(n7108), 
        .ZN(n7107) );
  OAI221_X1 U8072 ( .B1(n7254), .B2(keyinput130), .C1(n7108), .C2(keyinput173), 
        .A(n7107), .ZN(n7112) );
  XOR2_X1 U8073 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput255), .Z(n7111)
         );
  XNOR2_X1 U8074 ( .A(n7109), .B(keyinput226), .ZN(n7110) );
  OR3_X1 U8075 ( .A1(n7112), .A2(n7111), .A3(n7110), .ZN(n7118) );
  AOI22_X1 U8076 ( .A1(n5494), .A2(keyinput243), .B1(keyinput147), .B2(n7285), 
        .ZN(n7113) );
  OAI221_X1 U8077 ( .B1(n5494), .B2(keyinput243), .C1(n7285), .C2(keyinput147), 
        .A(n7113), .ZN(n7117) );
  AOI22_X1 U8078 ( .A1(n7115), .A2(keyinput194), .B1(n6356), .B2(keyinput253), 
        .ZN(n7114) );
  OAI221_X1 U8079 ( .B1(n7115), .B2(keyinput194), .C1(n6356), .C2(keyinput253), 
        .A(n7114), .ZN(n7116) );
  NOR3_X1 U8080 ( .A1(n7118), .A2(n7117), .A3(n7116), .ZN(n7145) );
  AOI22_X1 U8081 ( .A1(n7252), .A2(keyinput183), .B1(n4406), .B2(keyinput175), 
        .ZN(n7119) );
  OAI221_X1 U8082 ( .B1(n7252), .B2(keyinput183), .C1(n4406), .C2(keyinput175), 
        .A(n7119), .ZN(n7121) );
  XNOR2_X1 U8083 ( .A(n7307), .B(keyinput207), .ZN(n7120) );
  NOR2_X1 U8084 ( .A1(n7121), .A2(n7120), .ZN(n7130) );
  AOI22_X1 U8085 ( .A1(n7123), .A2(keyinput241), .B1(keyinput156), .B2(n3976), 
        .ZN(n7122) );
  OAI221_X1 U8086 ( .B1(n7123), .B2(keyinput241), .C1(n3976), .C2(keyinput156), 
        .A(n7122), .ZN(n7124) );
  INV_X1 U8087 ( .A(n7124), .ZN(n7129) );
  INV_X1 U8088 ( .A(DATAI_26_), .ZN(n7207) );
  AOI22_X1 U8089 ( .A1(n7245), .A2(keyinput128), .B1(n7207), .B2(keyinput167), 
        .ZN(n7125) );
  OAI221_X1 U8090 ( .B1(n7245), .B2(keyinput128), .C1(n7207), .C2(keyinput167), 
        .A(n7125), .ZN(n7126) );
  INV_X1 U8091 ( .A(n7126), .ZN(n7128) );
  XNOR2_X1 U8092 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .B(keyinput197), .ZN(n7127) );
  AND4_X1 U8093 ( .A1(n7130), .A2(n7129), .A3(n7128), .A4(n7127), .ZN(n7144)
         );
  AOI22_X1 U8094 ( .A1(n7294), .A2(keyinput164), .B1(keyinput170), .B2(n7299), 
        .ZN(n7131) );
  OAI221_X1 U8095 ( .B1(n7294), .B2(keyinput164), .C1(n7299), .C2(keyinput170), 
        .A(n7131), .ZN(n7142) );
  INV_X1 U8096 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n7251) );
  AOI22_X1 U8097 ( .A1(n7133), .A2(keyinput249), .B1(n7251), .B2(keyinput160), 
        .ZN(n7132) );
  OAI221_X1 U8098 ( .B1(n7133), .B2(keyinput249), .C1(n7251), .C2(keyinput160), 
        .A(n7132), .ZN(n7141) );
  AOI22_X1 U8099 ( .A1(n7135), .A2(keyinput233), .B1(n5234), .B2(keyinput151), 
        .ZN(n7134) );
  OAI221_X1 U8100 ( .B1(n7135), .B2(keyinput233), .C1(n5234), .C2(keyinput151), 
        .A(n7134), .ZN(n7140) );
  INV_X1 U8101 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n7138) );
  AOI22_X1 U8102 ( .A1(n7138), .A2(keyinput242), .B1(keyinput244), .B2(n7137), 
        .ZN(n7136) );
  OAI221_X1 U8103 ( .B1(n7138), .B2(keyinput242), .C1(n7137), .C2(keyinput244), 
        .A(n7136), .ZN(n7139) );
  NOR4_X1 U8104 ( .A1(n7142), .A2(n7141), .A3(n7140), .A4(n7139), .ZN(n7143)
         );
  NAND4_X1 U8105 ( .A1(n7146), .A2(n7145), .A3(n7144), .A4(n7143), .ZN(n7197)
         );
  AOI22_X1 U8106 ( .A1(n7149), .A2(keyinput174), .B1(keyinput159), .B2(n7148), 
        .ZN(n7147) );
  OAI221_X1 U8107 ( .B1(n7149), .B2(keyinput174), .C1(n7148), .C2(keyinput159), 
        .A(n7147), .ZN(n7159) );
  AOI22_X1 U8108 ( .A1(n3984), .A2(keyinput169), .B1(keyinput134), .B2(n7151), 
        .ZN(n7150) );
  OAI221_X1 U8109 ( .B1(n3984), .B2(keyinput169), .C1(n7151), .C2(keyinput134), 
        .A(n7150), .ZN(n7158) );
  AOI22_X1 U8110 ( .A1(n7224), .A2(keyinput213), .B1(keyinput143), .B2(n3862), 
        .ZN(n7152) );
  OAI221_X1 U8111 ( .B1(n7224), .B2(keyinput213), .C1(n3862), .C2(keyinput143), 
        .A(n7152), .ZN(n7157) );
  INV_X1 U8112 ( .A(DATAI_16_), .ZN(n7155) );
  AOI22_X1 U8113 ( .A1(n7155), .A2(keyinput185), .B1(keyinput137), .B2(n7154), 
        .ZN(n7153) );
  OAI221_X1 U8114 ( .B1(n7155), .B2(keyinput185), .C1(n7154), .C2(keyinput137), 
        .A(n7153), .ZN(n7156) );
  NOR4_X1 U8115 ( .A1(n7159), .A2(n7158), .A3(n7157), .A4(n7156), .ZN(n7195)
         );
  AOI22_X1 U8116 ( .A1(n7268), .A2(keyinput245), .B1(keyinput157), .B2(n7161), 
        .ZN(n7160) );
  OAI221_X1 U8117 ( .B1(n7268), .B2(keyinput245), .C1(n7161), .C2(keyinput157), 
        .A(n7160), .ZN(n7169) );
  INV_X1 U8118 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n7232) );
  INV_X1 U8119 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n7264) );
  AOI22_X1 U8120 ( .A1(n7232), .A2(keyinput252), .B1(n7264), .B2(keyinput132), 
        .ZN(n7162) );
  OAI221_X1 U8121 ( .B1(n7232), .B2(keyinput252), .C1(n7264), .C2(keyinput132), 
        .A(n7162), .ZN(n7168) );
  AOI22_X1 U8122 ( .A1(n7201), .A2(keyinput135), .B1(n7164), .B2(keyinput141), 
        .ZN(n7163) );
  OAI221_X1 U8123 ( .B1(n7201), .B2(keyinput135), .C1(n7164), .C2(keyinput141), 
        .A(n7163), .ZN(n7167) );
  AOI22_X1 U8124 ( .A1(n4864), .A2(keyinput146), .B1(n3688), .B2(keyinput223), 
        .ZN(n7165) );
  OAI221_X1 U8125 ( .B1(n4864), .B2(keyinput146), .C1(n3688), .C2(keyinput223), 
        .A(n7165), .ZN(n7166) );
  NOR4_X1 U8126 ( .A1(n7169), .A2(n7168), .A3(n7167), .A4(n7166), .ZN(n7194)
         );
  AOI22_X1 U8127 ( .A1(n4432), .A2(keyinput254), .B1(n7263), .B2(keyinput225), 
        .ZN(n7170) );
  OAI221_X1 U8128 ( .B1(n4432), .B2(keyinput254), .C1(n7263), .C2(keyinput225), 
        .A(n7170), .ZN(n7181) );
  AOI22_X1 U8129 ( .A1(n7172), .A2(keyinput218), .B1(n3885), .B2(keyinput208), 
        .ZN(n7171) );
  OAI221_X1 U8130 ( .B1(n7172), .B2(keyinput218), .C1(n3885), .C2(keyinput208), 
        .A(n7171), .ZN(n7180) );
  AOI22_X1 U8131 ( .A1(n7175), .A2(keyinput166), .B1(n7174), .B2(keyinput136), 
        .ZN(n7173) );
  OAI221_X1 U8132 ( .B1(n7175), .B2(keyinput166), .C1(n7174), .C2(keyinput136), 
        .A(n7173), .ZN(n7179) );
  AOI22_X1 U8133 ( .A1(n6053), .A2(keyinput138), .B1(keyinput198), .B2(n7177), 
        .ZN(n7176) );
  OAI221_X1 U8134 ( .B1(n6053), .B2(keyinput138), .C1(n7177), .C2(keyinput198), 
        .A(n7176), .ZN(n7178) );
  NOR4_X1 U8135 ( .A1(n7181), .A2(n7180), .A3(n7179), .A4(n7178), .ZN(n7193)
         );
  AOI22_X1 U8136 ( .A1(n7183), .A2(keyinput206), .B1(keyinput221), .B2(n5940), 
        .ZN(n7182) );
  OAI221_X1 U8137 ( .B1(n7183), .B2(keyinput206), .C1(n5940), .C2(keyinput221), 
        .A(n7182), .ZN(n7191) );
  AOI22_X1 U8138 ( .A1(n3627), .A2(keyinput133), .B1(keyinput163), .B2(n7316), 
        .ZN(n7184) );
  OAI221_X1 U8139 ( .B1(n3627), .B2(keyinput133), .C1(n7316), .C2(keyinput163), 
        .A(n7184), .ZN(n7190) );
  INV_X1 U8140 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n7296) );
  AOI22_X1 U8141 ( .A1(n7296), .A2(keyinput211), .B1(n5177), .B2(keyinput216), 
        .ZN(n7185) );
  OAI221_X1 U8142 ( .B1(n7296), .B2(keyinput211), .C1(n5177), .C2(keyinput216), 
        .A(n7185), .ZN(n7189) );
  AOI22_X1 U8143 ( .A1(n7187), .A2(keyinput202), .B1(n5023), .B2(keyinput176), 
        .ZN(n7186) );
  OAI221_X1 U8144 ( .B1(n7187), .B2(keyinput202), .C1(n5023), .C2(keyinput176), 
        .A(n7186), .ZN(n7188) );
  NOR4_X1 U8145 ( .A1(n7191), .A2(n7190), .A3(n7189), .A4(n7188), .ZN(n7192)
         );
  NAND4_X1 U8146 ( .A1(n7195), .A2(n7194), .A3(n7193), .A4(n7192), .ZN(n7196)
         );
  NOR4_X1 U8147 ( .A1(n7199), .A2(n7198), .A3(n7197), .A4(n7196), .ZN(n7327)
         );
  AOI22_X1 U8148 ( .A1(n4062), .A2(keyinput118), .B1(keyinput7), .B2(n7201), 
        .ZN(n7200) );
  OAI221_X1 U8149 ( .B1(n4062), .B2(keyinput118), .C1(n7201), .C2(keyinput7), 
        .A(n7200), .ZN(n7213) );
  AOI22_X1 U8150 ( .A1(n5023), .A2(keyinput48), .B1(keyinput96), .B2(n7203), 
        .ZN(n7202) );
  OAI221_X1 U8151 ( .B1(n5023), .B2(keyinput48), .C1(n7203), .C2(keyinput96), 
        .A(n7202), .ZN(n7212) );
  INV_X1 U8152 ( .A(BS16_N), .ZN(n7206) );
  AOI22_X1 U8153 ( .A1(n7206), .A2(keyinput87), .B1(n7205), .B2(keyinput81), 
        .ZN(n7204) );
  OAI221_X1 U8154 ( .B1(n7206), .B2(keyinput87), .C1(n7205), .C2(keyinput81), 
        .A(n7204), .ZN(n7211) );
  XOR2_X1 U8155 ( .A(n7207), .B(keyinput39), .Z(n7209) );
  XNOR2_X1 U8156 ( .A(n4955), .B(keyinput30), .ZN(n7208) );
  NAND2_X1 U8157 ( .A1(n7209), .A2(n7208), .ZN(n7210) );
  NOR4_X1 U8158 ( .A1(n7213), .A2(n7212), .A3(n7211), .A4(n7210), .ZN(n7261)
         );
  AOI22_X1 U8159 ( .A1(n3984), .A2(keyinput41), .B1(keyinput22), .B2(n7215), 
        .ZN(n7214) );
  OAI221_X1 U8160 ( .B1(n3984), .B2(keyinput41), .C1(n7215), .C2(keyinput22), 
        .A(n7214), .ZN(n7228) );
  AOI22_X1 U8161 ( .A1(n7218), .A2(keyinput59), .B1(keyinput1), .B2(n7217), 
        .ZN(n7216) );
  OAI221_X1 U8162 ( .B1(n7218), .B2(keyinput59), .C1(n7217), .C2(keyinput1), 
        .A(n7216), .ZN(n7227) );
  INV_X1 U8163 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n7221) );
  INV_X1 U8164 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7220) );
  AOI22_X1 U8165 ( .A1(n7221), .A2(keyinput11), .B1(keyinput89), .B2(n7220), 
        .ZN(n7219) );
  OAI221_X1 U8166 ( .B1(n7221), .B2(keyinput11), .C1(n7220), .C2(keyinput89), 
        .A(n7219), .ZN(n7226) );
  AOI22_X1 U8167 ( .A1(n7224), .A2(keyinput85), .B1(keyinput33), .B2(n7223), 
        .ZN(n7222) );
  OAI221_X1 U8168 ( .B1(n7224), .B2(keyinput85), .C1(n7223), .C2(keyinput33), 
        .A(n7222), .ZN(n7225) );
  NOR4_X1 U8169 ( .A1(n7228), .A2(n7227), .A3(n7226), .A4(n7225), .ZN(n7260)
         );
  AOI22_X1 U8170 ( .A1(n7231), .A2(keyinput25), .B1(keyinput107), .B2(n7230), 
        .ZN(n7229) );
  OAI221_X1 U8171 ( .B1(n7231), .B2(keyinput25), .C1(n7230), .C2(keyinput107), 
        .A(n7229), .ZN(n7235) );
  XOR2_X1 U8172 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .B(keyinput69), .Z(n7234)
         );
  XNOR2_X1 U8173 ( .A(n7232), .B(keyinput124), .ZN(n7233) );
  OR3_X1 U8174 ( .A1(n7235), .A2(n7234), .A3(n7233), .ZN(n7243) );
  AOI22_X1 U8175 ( .A1(n7237), .A2(keyinput26), .B1(keyinput28), .B2(n3976), 
        .ZN(n7236) );
  OAI221_X1 U8176 ( .B1(n7237), .B2(keyinput26), .C1(n3976), .C2(keyinput28), 
        .A(n7236), .ZN(n7242) );
  AOI22_X1 U8177 ( .A1(n7240), .A2(keyinput100), .B1(keyinput106), .B2(n7239), 
        .ZN(n7238) );
  OAI221_X1 U8178 ( .B1(n7240), .B2(keyinput100), .C1(n7239), .C2(keyinput106), 
        .A(n7238), .ZN(n7241) );
  NOR3_X1 U8179 ( .A1(n7243), .A2(n7242), .A3(n7241), .ZN(n7259) );
  AOI22_X1 U8180 ( .A1(n7245), .A2(keyinput0), .B1(n3688), .B2(keyinput95), 
        .ZN(n7244) );
  OAI221_X1 U8181 ( .B1(n7245), .B2(keyinput0), .C1(n3688), .C2(keyinput95), 
        .A(n7244), .ZN(n7249) );
  XOR2_X1 U8182 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .B(keyinput123), .Z(n7248)
         );
  XNOR2_X1 U8183 ( .A(n7246), .B(keyinput60), .ZN(n7247) );
  OR3_X1 U8184 ( .A1(n7249), .A2(n7248), .A3(n7247), .ZN(n7257) );
  AOI22_X1 U8185 ( .A1(n7252), .A2(keyinput55), .B1(n7251), .B2(keyinput32), 
        .ZN(n7250) );
  OAI221_X1 U8186 ( .B1(n7252), .B2(keyinput55), .C1(n7251), .C2(keyinput32), 
        .A(n7250), .ZN(n7256) );
  AOI22_X1 U8187 ( .A1(n7254), .A2(keyinput2), .B1(n5177), .B2(keyinput88), 
        .ZN(n7253) );
  OAI221_X1 U8188 ( .B1(n7254), .B2(keyinput2), .C1(n5177), .C2(keyinput88), 
        .A(n7253), .ZN(n7255) );
  NOR3_X1 U8189 ( .A1(n7257), .A2(n7256), .A3(n7255), .ZN(n7258) );
  NAND4_X1 U8190 ( .A1(n7261), .A2(n7260), .A3(n7259), .A4(n7258), .ZN(n7326)
         );
  AOI22_X1 U8191 ( .A1(n7264), .A2(keyinput4), .B1(n7263), .B2(keyinput97), 
        .ZN(n7262) );
  OAI221_X1 U8192 ( .B1(n7264), .B2(keyinput4), .C1(n7263), .C2(keyinput97), 
        .A(n7262), .ZN(n7275) );
  AOI22_X1 U8193 ( .A1(n4094), .A2(keyinput73), .B1(n7266), .B2(keyinput64), 
        .ZN(n7265) );
  OAI221_X1 U8194 ( .B1(n4094), .B2(keyinput73), .C1(n7266), .C2(keyinput64), 
        .A(n7265), .ZN(n7274) );
  AOI22_X1 U8195 ( .A1(n7269), .A2(keyinput109), .B1(keyinput117), .B2(n7268), 
        .ZN(n7267) );
  OAI221_X1 U8196 ( .B1(n7269), .B2(keyinput109), .C1(n7268), .C2(keyinput117), 
        .A(n7267), .ZN(n7273) );
  AOI22_X1 U8197 ( .A1(n7271), .A2(keyinput111), .B1(n5083), .B2(keyinput76), 
        .ZN(n7270) );
  OAI221_X1 U8198 ( .B1(n7271), .B2(keyinput111), .C1(n5083), .C2(keyinput76), 
        .A(n7270), .ZN(n7272) );
  NOR4_X1 U8199 ( .A1(n7275), .A2(n7274), .A3(n7273), .A4(n7272), .ZN(n7324)
         );
  INV_X1 U8200 ( .A(DATAI_30_), .ZN(n7277) );
  AOI22_X1 U8201 ( .A1(n7278), .A2(keyinput112), .B1(n7277), .B2(keyinput43), 
        .ZN(n7276) );
  OAI221_X1 U8202 ( .B1(n7278), .B2(keyinput112), .C1(n7277), .C2(keyinput43), 
        .A(n7276), .ZN(n7289) );
  AOI22_X1 U8203 ( .A1(n7280), .A2(keyinput103), .B1(keyinput18), .B2(n4864), 
        .ZN(n7279) );
  OAI221_X1 U8204 ( .B1(n7280), .B2(keyinput103), .C1(n4864), .C2(keyinput18), 
        .A(n7279), .ZN(n7288) );
  AOI22_X1 U8205 ( .A1(n7283), .A2(keyinput122), .B1(keyinput91), .B2(n7282), 
        .ZN(n7281) );
  OAI221_X1 U8206 ( .B1(n7283), .B2(keyinput122), .C1(n7282), .C2(keyinput91), 
        .A(n7281), .ZN(n7287) );
  AOI22_X1 U8207 ( .A1(n5940), .A2(keyinput93), .B1(keyinput19), .B2(n7285), 
        .ZN(n7284) );
  OAI221_X1 U8208 ( .B1(n5940), .B2(keyinput93), .C1(n7285), .C2(keyinput19), 
        .A(n7284), .ZN(n7286) );
  NOR4_X1 U8209 ( .A1(n7289), .A2(n7288), .A3(n7287), .A4(n7286), .ZN(n7323)
         );
  AOI22_X1 U8210 ( .A1(n7291), .A2(keyinput52), .B1(keyinput34), .B2(n4862), 
        .ZN(n7290) );
  OAI221_X1 U8211 ( .B1(n7291), .B2(keyinput52), .C1(n4862), .C2(keyinput34), 
        .A(n7290), .ZN(n7304) );
  AOI22_X1 U8212 ( .A1(n7294), .A2(keyinput36), .B1(n7293), .B2(keyinput72), 
        .ZN(n7292) );
  OAI221_X1 U8213 ( .B1(n7294), .B2(keyinput36), .C1(n7293), .C2(keyinput72), 
        .A(n7292), .ZN(n7303) );
  INV_X1 U8214 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n7297) );
  AOI22_X1 U8215 ( .A1(n7297), .A2(keyinput77), .B1(keyinput83), .B2(n7296), 
        .ZN(n7295) );
  OAI221_X1 U8216 ( .B1(n7297), .B2(keyinput77), .C1(n7296), .C2(keyinput83), 
        .A(n7295), .ZN(n7302) );
  AOI22_X1 U8217 ( .A1(n7300), .A2(keyinput54), .B1(n7299), .B2(keyinput42), 
        .ZN(n7298) );
  OAI221_X1 U8218 ( .B1(n7300), .B2(keyinput54), .C1(n7299), .C2(keyinput42), 
        .A(n7298), .ZN(n7301) );
  NOR4_X1 U8219 ( .A1(n7304), .A2(n7303), .A3(n7302), .A4(n7301), .ZN(n7322)
         );
  AOI22_X1 U8220 ( .A1(n7307), .A2(keyinput79), .B1(n7306), .B2(keyinput68), 
        .ZN(n7305) );
  OAI221_X1 U8221 ( .B1(n7307), .B2(keyinput79), .C1(n7306), .C2(keyinput68), 
        .A(n7305), .ZN(n7320) );
  INV_X1 U8222 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n7309) );
  AOI22_X1 U8223 ( .A1(n7310), .A2(keyinput94), .B1(n7309), .B2(keyinput75), 
        .ZN(n7308) );
  OAI221_X1 U8224 ( .B1(n7310), .B2(keyinput94), .C1(n7309), .C2(keyinput75), 
        .A(n7308), .ZN(n7319) );
  INV_X1 U8225 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n7313) );
  INV_X1 U8226 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n7312) );
  AOI22_X1 U8227 ( .A1(n7313), .A2(keyinput92), .B1(n7312), .B2(keyinput120), 
        .ZN(n7311) );
  OAI221_X1 U8228 ( .B1(n7313), .B2(keyinput92), .C1(n7312), .C2(keyinput120), 
        .A(n7311), .ZN(n7318) );
  AOI22_X1 U8229 ( .A1(n7316), .A2(keyinput35), .B1(n7315), .B2(keyinput65), 
        .ZN(n7314) );
  OAI221_X1 U8230 ( .B1(n7316), .B2(keyinput35), .C1(n7315), .C2(keyinput65), 
        .A(n7314), .ZN(n7317) );
  NOR4_X1 U8231 ( .A1(n7320), .A2(n7319), .A3(n7318), .A4(n7317), .ZN(n7321)
         );
  NAND4_X1 U8232 ( .A1(n7324), .A2(n7323), .A3(n7322), .A4(n7321), .ZN(n7325)
         );
  NOR3_X1 U8233 ( .A1(n7327), .A2(n7326), .A3(n7325), .ZN(n7365) );
  OAI22_X1 U8234 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(keyinput20), .B1(
        keyinput58), .B2(DATAO_REG_15__SCAN_IN), .ZN(n7328) );
  AOI221_X1 U8235 ( .B1(INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput20), .C1(
        DATAO_REG_15__SCAN_IN), .C2(keyinput58), .A(n7328), .ZN(n7335) );
  OAI22_X1 U8236 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput15), .B1(
        LWORD_REG_11__SCAN_IN), .B2(keyinput50), .ZN(n7329) );
  AOI221_X1 U8237 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput15), .C1(keyinput50), 
        .C2(LWORD_REG_11__SCAN_IN), .A(n7329), .ZN(n7334) );
  OAI22_X1 U8238 ( .A1(DATAI_31_), .A2(keyinput53), .B1(DATAI_16_), .B2(
        keyinput57), .ZN(n7330) );
  AOI221_X1 U8239 ( .B1(DATAI_31_), .B2(keyinput53), .C1(keyinput57), .C2(
        DATAI_16_), .A(n7330), .ZN(n7333) );
  OAI22_X1 U8240 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(keyinput40), .B1(
        EAX_REG_3__SCAN_IN), .B2(keyinput78), .ZN(n7331) );
  AOI221_X1 U8241 ( .B1(INSTQUEUE_REG_6__3__SCAN_IN), .B2(keyinput40), .C1(
        keyinput78), .C2(EAX_REG_3__SCAN_IN), .A(n7331), .ZN(n7332) );
  NAND4_X1 U8242 ( .A1(n7335), .A2(n7334), .A3(n7333), .A4(n7332), .ZN(n7363)
         );
  OAI22_X1 U8243 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(keyinput125), .B1(
        DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput105), .ZN(n7336) );
  AOI221_X1 U8244 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(keyinput125), .C1(
        keyinput105), .C2(DATAWIDTH_REG_15__SCAN_IN), .A(n7336), .ZN(n7343) );
  OAI22_X1 U8245 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput37), .B1(
        keyinput119), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n7337) );
  AOI221_X1 U8246 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput37), .C1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .C2(keyinput119), .A(n7337), .ZN(
        n7342) );
  OAI22_X1 U8247 ( .A1(EBX_REG_20__SCAN_IN), .A2(keyinput126), .B1(
        EAX_REG_4__SCAN_IN), .B2(keyinput102), .ZN(n7338) );
  AOI221_X1 U8248 ( .B1(EBX_REG_20__SCAN_IN), .B2(keyinput126), .C1(
        keyinput102), .C2(EAX_REG_4__SCAN_IN), .A(n7338), .ZN(n7341) );
  OAI22_X1 U8249 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput115), .B1(
        DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput3), .ZN(n7339) );
  AOI221_X1 U8250 ( .B1(INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput115), .C1(
        keyinput3), .C2(DATAWIDTH_REG_3__SCAN_IN), .A(n7339), .ZN(n7340) );
  NAND4_X1 U8251 ( .A1(n7343), .A2(n7342), .A3(n7341), .A4(n7340), .ZN(n7362)
         );
  OAI22_X1 U8252 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput8), .B1(
        keyinput90), .B2(ADDRESS_REG_20__SCAN_IN), .ZN(n7344) );
  AOI221_X1 U8253 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput8), .C1(
        ADDRESS_REG_20__SCAN_IN), .C2(keyinput90), .A(n7344), .ZN(n7351) );
  OAI22_X1 U8254 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(keyinput21), .B1(
        DATAO_REG_11__SCAN_IN), .B2(keyinput45), .ZN(n7345) );
  AOI221_X1 U8255 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput21), .C1(
        keyinput45), .C2(DATAO_REG_11__SCAN_IN), .A(n7345), .ZN(n7350) );
  OAI22_X1 U8256 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(keyinput127), .B1(
        INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput86), .ZN(n7346) );
  AOI221_X1 U8257 ( .B1(INSTQUEUE_REG_0__1__SCAN_IN), .B2(keyinput127), .C1(
        keyinput86), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n7346), .ZN(
        n7349) );
  OAI22_X1 U8258 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(keyinput114), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput110), .ZN(n7347) );
  AOI221_X1 U8259 ( .B1(INSTQUEUE_REG_15__3__SCAN_IN), .B2(keyinput114), .C1(
        keyinput110), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n7347), .ZN(
        n7348) );
  NAND4_X1 U8260 ( .A1(n7351), .A2(n7350), .A3(n7349), .A4(n7348), .ZN(n7361)
         );
  OAI22_X1 U8261 ( .A1(EAX_REG_13__SCAN_IN), .A2(keyinput80), .B1(DATAI_19_), 
        .B2(keyinput16), .ZN(n7352) );
  AOI221_X1 U8262 ( .B1(EAX_REG_13__SCAN_IN), .B2(keyinput80), .C1(keyinput16), 
        .C2(DATAI_19_), .A(n7352), .ZN(n7359) );
  OAI22_X1 U8263 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput63), .B1(keyinput108), .B2(DATAO_REG_8__SCAN_IN), .ZN(n7353) );
  AOI221_X1 U8264 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput63), .C1(
        DATAO_REG_8__SCAN_IN), .C2(keyinput108), .A(n7353), .ZN(n7358) );
  OAI22_X1 U8265 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(keyinput17), .B1(
        keyinput116), .B2(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7354) );
  AOI221_X1 U8266 ( .B1(INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput17), .C1(
        DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput116), .A(n7354), .ZN(n7357) );
  OAI22_X1 U8267 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(keyinput23), .B1(
        keyinput66), .B2(ADDRESS_REG_17__SCAN_IN), .ZN(n7355) );
  AOI221_X1 U8268 ( .B1(INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput23), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput66), .A(n7355), .ZN(n7356) );
  NAND4_X1 U8269 ( .A1(n7359), .A2(n7358), .A3(n7357), .A4(n7356), .ZN(n7360)
         );
  NOR4_X1 U8270 ( .A1(n7363), .A2(n7362), .A3(n7361), .A4(n7360), .ZN(n7364)
         );
  NAND3_X1 U8271 ( .A1(n7366), .A2(n7365), .A3(n7364), .ZN(n7380) );
  OAI22_X1 U8272 ( .A1(n7370), .A2(n7369), .B1(n7368), .B2(n7367), .ZN(n7371)
         );
  INV_X1 U8273 ( .A(n7371), .ZN(n7376) );
  AOI22_X1 U8274 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n7374), .B1(n7373), 
        .B2(n7372), .ZN(n7375) );
  OAI211_X1 U8275 ( .C1(n7378), .C2(n7377), .A(n7376), .B(n7375), .ZN(n7379)
         );
  XNOR2_X1 U8276 ( .A(n7380), .B(n7379), .ZN(U3112) );
  NOR2_X1 U4303 ( .A1(n4953), .A2(n4735), .ZN(n4952) );
  AND2_X2 U3794 ( .A1(n3309), .A2(n3314), .ZN(n3430) );
  CLKBUF_X2 U3676 ( .A(n3510), .Z(n4904) );
  BUF_X1 U3646 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4955) );
  CLKBUF_X2 U3693 ( .A(n4561), .Z(n3204) );
  CLKBUF_X1 U3669 ( .A(n4156), .Z(n4590) );
  NAND2_X1 U3677 ( .A1(n3563), .A2(n3562), .ZN(n3609) );
  CLKBUF_X1 U3685 ( .A(n3468), .Z(n3200) );
  CLKBUF_X1 U3687 ( .A(n3617), .Z(n3199) );
  NAND2_X2 U3691 ( .A1(n4470), .A2(n4770), .ZN(n4368) );
  CLKBUF_X2 U3694 ( .A(n4561), .Z(n3203) );
  OR2_X2 U3697 ( .A1(n3622), .A2(n3621), .ZN(n3678) );
  CLKBUF_X1 U3711 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n4954) );
  INV_X1 U4115 ( .A(n4561), .ZN(n4555) );
endmodule

