

module b14_C_AntiSAT_k_256_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2226, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079;

  INV_X1 U2468 ( .A(n2537), .ZN(n2750) );
  CLKBUF_X1 U2469 ( .A(n4480), .Z(n2230) );
  INV_X2 U2470 ( .A(n3733), .ZN(n2908) );
  INV_X1 U2472 ( .A(n2537), .ZN(n2226) );
  NOR2_X1 U2473 ( .A1(n4469), .A2(n2501), .ZN(n2549) );
  NOR2_X1 U2475 ( .A1(n4469), .A2(n2998), .ZN(n2550) );
  XNOR2_X1 U2477 ( .A(n4087), .B(n4116), .ZN(n4602) );
  OAI21_X1 U2478 ( .B1(n4655), .B2(n4698), .A(n4545), .ZN(n4081) );
  NAND2_X1 U2479 ( .A1(n4524), .A2(n4078), .ZN(n4079) );
  AND2_X2 U2480 ( .A1(n2980), .A2(n4261), .ZN(n4491) );
  INV_X2 U2481 ( .A(n4507), .ZN(n2229) );
  OR2_X1 U2482 ( .A1(n3039), .A2(n3040), .ZN(n2347) );
  XNOR2_X1 U2483 ( .A(n3098), .B(n2348), .ZN(n3039) );
  NAND2_X2 U2484 ( .A1(n2322), .A2(n2899), .ZN(n3733) );
  NAND4_X1 U2485 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n4058)
         );
  NAND2_X2 U2486 ( .A1(n2899), .A2(n3146), .ZN(n3732) );
  CLKBUF_X1 U2487 ( .A(n2826), .Z(n3873) );
  CLKBUF_X1 U2488 ( .A(n2537), .Z(n3876) );
  XNOR2_X1 U2489 ( .A(n2418), .B(IR_REG_30__SCAN_IN), .ZN(n4469) );
  INV_X1 U2490 ( .A(n2343), .ZN(n2566) );
  NAND2_X1 U2491 ( .A1(n2342), .A2(n2341), .ZN(n2343) );
  NOR2_X1 U2492 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2480)
         );
  NOR2_X1 U2493 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2477)
         );
  INV_X1 U2494 ( .A(IR_REG_23__SCAN_IN), .ZN(n4936) );
  XNOR2_X1 U2495 ( .A(n2354), .B(n2353), .ZN(n4480) );
  INV_X1 U2496 ( .A(n2428), .ZN(n2423) );
  NOR2_X1 U2497 ( .A1(n2472), .A2(n2490), .ZN(n2471) );
  NAND2_X1 U2498 ( .A1(n2491), .A2(n2487), .ZN(n2472) );
  AND2_X1 U2499 ( .A1(n2475), .A2(n2575), .ZN(n2476) );
  NOR2_X1 U2500 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2475)
         );
  AND2_X1 U2501 ( .A1(n2566), .A2(n2478), .ZN(n2452) );
  NOR2_X1 U2502 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2478)
         );
  AND4_X1 U2503 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n2485)
         );
  NOR2_X1 U2504 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2484)
         );
  NOR2_X1 U2505 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2483)
         );
  NOR2_X1 U2506 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2482)
         );
  INV_X1 U2507 ( .A(n2699), .ZN(n2374) );
  INV_X1 U2508 ( .A(n3003), .ZN(n2862) );
  NAND2_X1 U2509 ( .A1(n2317), .A2(n2315), .ZN(n3329) );
  AOI21_X1 U2510 ( .B1(n2318), .B2(n2933), .A(n2316), .ZN(n2315) );
  NOR2_X1 U2511 ( .A1(n3280), .A2(n2246), .ZN(n2318) );
  INV_X1 U2512 ( .A(n3791), .ZN(n2449) );
  AND2_X1 U2513 ( .A1(n3769), .A2(n2414), .ZN(n2413) );
  NAND2_X1 U2514 ( .A1(n3840), .A2(n2415), .ZN(n2414) );
  INV_X1 U2515 ( .A(n3356), .ZN(n2426) );
  NAND2_X1 U2516 ( .A1(n2429), .A2(n2434), .ZN(n2428) );
  NAND2_X1 U2517 ( .A1(n2430), .A2(n3354), .ZN(n2429) );
  INV_X1 U2518 ( .A(n3379), .ZN(n2430) );
  OR2_X1 U2519 ( .A1(n2757), .A2(n3813), .ZN(n2527) );
  INV_X1 U2520 ( .A(n3078), .ZN(n2288) );
  NAND2_X1 U2522 ( .A1(n2326), .A2(IR_REG_31__SCAN_IN), .ZN(n2884) );
  AND2_X1 U2523 ( .A1(n2471), .A2(n2328), .ZN(n2327) );
  INV_X1 U2524 ( .A(IR_REG_26__SCAN_IN), .ZN(n2328) );
  XNOR2_X1 U2525 ( .A(n4103), .B(n2355), .ZN(n4516) );
  XNOR2_X1 U2526 ( .A(n4106), .B(n2344), .ZN(n4537) );
  NAND2_X1 U2527 ( .A1(n4608), .A2(n2350), .ZN(n4120) );
  NAND2_X1 U2528 ( .A1(n4646), .A2(n2351), .ZN(n2350) );
  INV_X1 U2529 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2351) );
  NOR2_X1 U2530 ( .A1(n4120), .A2(n4121), .ZN(n4128) );
  OR2_X1 U2531 ( .A1(n2527), .A2(n4955), .ZN(n2519) );
  AND2_X1 U2533 ( .A1(n2471), .A2(n2496), .ZN(n2469) );
  NOR2_X1 U2534 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2496)
         );
  NAND2_X1 U2535 ( .A1(n2733), .A2(n2732), .ZN(n2773) );
  INV_X1 U2536 ( .A(n4566), .ZN(n2279) );
  INV_X1 U2537 ( .A(IR_REG_16__SCAN_IN), .ZN(n4933) );
  INV_X1 U2538 ( .A(IR_REG_13__SCAN_IN), .ZN(n2674) );
  NOR2_X1 U2539 ( .A1(n2432), .A2(n3379), .ZN(n2431) );
  NOR2_X1 U2540 ( .A1(n2460), .A2(n2456), .ZN(n2455) );
  AND2_X1 U2541 ( .A1(n3651), .A2(n2461), .ZN(n2460) );
  INV_X1 U2542 ( .A(n3644), .ZN(n2456) );
  AND2_X1 U2543 ( .A1(n2458), .A2(n2294), .ZN(n2293) );
  AND2_X1 U2544 ( .A1(n4496), .A2(n2459), .ZN(n2458) );
  NAND2_X1 U2545 ( .A1(n2455), .A2(n2295), .ZN(n2294) );
  OR2_X1 U2546 ( .A1(n3651), .A2(n2461), .ZN(n2459) );
  INV_X1 U2547 ( .A(n2906), .ZN(n3741) );
  AOI21_X1 U2548 ( .B1(n3038), .B2(REG1_REG_5__SCAN_IN), .A(n3088), .ZN(n3098)
         );
  NAND2_X1 U2549 ( .A1(n4548), .A2(n4108), .ZN(n4109) );
  AND2_X1 U2550 ( .A1(n4160), .A2(n3740), .ZN(n3898) );
  AND2_X1 U2551 ( .A1(n4280), .A2(n4258), .ZN(n2409) );
  OR2_X1 U2552 ( .A1(n4231), .A2(n4230), .ZN(n4292) );
  OAI21_X1 U2553 ( .B1(n3942), .B2(n2374), .A(n2712), .ZN(n2373) );
  NOR2_X1 U2554 ( .A1(n2374), .A2(n2371), .ZN(n2370) );
  INV_X1 U2555 ( .A(n2687), .ZN(n2371) );
  AND2_X1 U2556 ( .A1(n4471), .A2(n3955), .ZN(n3012) );
  NAND2_X1 U2557 ( .A1(n4026), .A2(n3955), .ZN(n3146) );
  NAND2_X1 U2558 ( .A1(n4247), .A2(n4200), .ZN(n2332) );
  AND2_X1 U2559 ( .A1(n2235), .A2(n3333), .ZN(n2333) );
  AND2_X1 U2560 ( .A1(n3190), .A2(n3206), .ZN(n3189) );
  NAND2_X1 U2561 ( .A1(n2546), .A2(DATAI_2_), .ZN(n2557) );
  NAND2_X1 U2562 ( .A1(n2324), .A2(n4479), .ZN(n2323) );
  INV_X1 U2563 ( .A(n2546), .ZN(n2324) );
  NAND2_X1 U2564 ( .A1(n2489), .A2(n4936), .ZN(n2490) );
  NAND2_X1 U2565 ( .A1(n2451), .A2(n2452), .ZN(n2454) );
  AND2_X1 U2566 ( .A1(n2450), .A2(n2476), .ZN(n2451) );
  AND3_X1 U2567 ( .A1(n2479), .A2(n2477), .A3(n2480), .ZN(n2450) );
  OR3_X1 U2568 ( .A1(n2628), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2638) );
  AOI21_X1 U2569 ( .B1(n2448), .B2(n2303), .A(n2260), .ZN(n2302) );
  INV_X1 U2570 ( .A(n3790), .ZN(n2303) );
  AOI22_X1 U2571 ( .A1(n3625), .A2(n3624), .B1(n3623), .B2(n3622), .ZN(n3643)
         );
  NAND2_X1 U2572 ( .A1(n2307), .A2(n2313), .ZN(n2305) );
  INV_X1 U2573 ( .A(n2431), .ZN(n2425) );
  NAND2_X1 U2574 ( .A1(n2423), .A2(n2427), .ZN(n2422) );
  AOI21_X1 U2575 ( .B1(n2446), .B2(n2445), .A(n2444), .ZN(n2443) );
  NOR2_X1 U2576 ( .A1(n3737), .A2(n3738), .ZN(n2444) );
  NOR2_X1 U2577 ( .A1(n2448), .A2(n2260), .ZN(n2445) );
  NOR2_X1 U2578 ( .A1(n2601), .A2(n2600), .ZN(n2611) );
  INV_X1 U2579 ( .A(n2230), .ZN(n2368) );
  AND2_X1 U2580 ( .A1(n3471), .A2(n3470), .ZN(n3552) );
  NAND2_X1 U2581 ( .A1(n2466), .A2(n2465), .ZN(n3809) );
  AOI21_X1 U2582 ( .B1(n3329), .B2(n3330), .A(n2944), .ZN(n3356) );
  NAND2_X1 U2583 ( .A1(n2314), .A2(n2311), .ZN(n2310) );
  INV_X1 U2584 ( .A(n3820), .ZN(n2311) );
  NOR2_X1 U2585 ( .A1(n2463), .A2(n2308), .ZN(n2307) );
  INV_X1 U2586 ( .A(n2310), .ZN(n2308) );
  NAND2_X1 U2587 ( .A1(n3702), .A2(n2464), .ZN(n2463) );
  INV_X1 U2588 ( .A(n3699), .ZN(n2464) );
  NAND2_X1 U2589 ( .A1(n3682), .A2(n2312), .ZN(n2309) );
  OR2_X1 U2590 ( .A1(n2640), .A2(n4879), .ZN(n2652) );
  NAND2_X1 U2591 ( .A1(n3839), .A2(n3841), .ZN(n3838) );
  NAND2_X1 U2592 ( .A1(n3666), .A2(n3798), .ZN(n3839) );
  NAND2_X1 U2593 ( .A1(n2663), .A2(REG3_REG_13__SCAN_IN), .ZN(n2680) );
  AND2_X1 U2594 ( .A1(n2908), .A2(n2974), .ZN(n4033) );
  NOR2_X1 U2595 ( .A1(n2992), .A2(n2859), .ZN(n2844) );
  NAND2_X1 U2596 ( .A1(n3115), .A2(n3034), .ZN(n3035) );
  NOR2_X1 U2597 ( .A1(n2285), .A2(n2243), .ZN(n3022) );
  NAND2_X1 U2598 ( .A1(n4100), .A2(n2261), .ZN(n4103) );
  NAND2_X1 U2599 ( .A1(n4516), .A2(REG2_REG_8__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U2600 ( .A1(n4527), .A2(n4105), .ZN(n4106) );
  NAND2_X1 U2601 ( .A1(n4537), .A2(REG2_REG_10__SCAN_IN), .ZN(n4536) );
  OR2_X1 U2602 ( .A1(n4580), .A2(n4113), .ZN(n2273) );
  OAI21_X1 U2603 ( .B1(n4580), .B2(n2271), .A(n2270), .ZN(n4117) );
  NAND2_X1 U2604 ( .A1(n4588), .A2(n2274), .ZN(n2270) );
  OR2_X1 U2605 ( .A1(n4113), .A2(n2356), .ZN(n2271) );
  NAND2_X1 U2606 ( .A1(n4592), .A2(n4086), .ZN(n4087) );
  NOR2_X1 U2607 ( .A1(n4616), .A2(n4089), .ZN(n4124) );
  NAND2_X1 U2608 ( .A1(n2763), .A2(n2762), .ZN(n2875) );
  NAND2_X1 U2609 ( .A1(n4180), .A2(n4162), .ZN(n2762) );
  OR2_X1 U2610 ( .A1(n3898), .A2(n3895), .ZN(n3948) );
  NAND2_X1 U2611 ( .A1(n2378), .A2(n2377), .ZN(n4172) );
  OR2_X1 U2612 ( .A1(n4178), .A2(n4200), .ZN(n2377) );
  NAND2_X1 U2613 ( .A1(n4191), .A2(n2262), .ZN(n2378) );
  OAI21_X1 U2614 ( .B1(n4185), .B2(n2832), .A(n2517), .ZN(n4197) );
  NAND2_X1 U2615 ( .A1(n2407), .A2(n2403), .ZN(n2402) );
  INV_X1 U2616 ( .A(n2409), .ZN(n2403) );
  NOR2_X1 U2617 ( .A1(n2409), .A2(n2405), .ZN(n2404) );
  INV_X1 U2618 ( .A(n2754), .ZN(n2405) );
  AND2_X1 U2619 ( .A1(n2408), .A2(n2241), .ZN(n4255) );
  NAND2_X1 U2620 ( .A1(n4276), .A2(n2754), .ZN(n2408) );
  NOR2_X1 U2621 ( .A1(n2744), .A2(n4983), .ZN(n2746) );
  AND2_X1 U2622 ( .A1(n2746), .A2(REG3_REG_22__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U2623 ( .A1(n3597), .A2(n2726), .ZN(n4317) );
  NAND2_X1 U2624 ( .A1(n2688), .A2(n2687), .ZN(n3543) );
  NAND2_X1 U2625 ( .A1(n3543), .A2(n3942), .ZN(n3542) );
  AOI21_X1 U2626 ( .B1(n2396), .B2(n2394), .A(n2248), .ZN(n2393) );
  AND2_X1 U2627 ( .A1(n2242), .A2(n2662), .ZN(n2394) );
  NAND2_X1 U2628 ( .A1(n3516), .A2(n3515), .ZN(n2396) );
  AOI21_X1 U2629 ( .B1(n2381), .B2(n2237), .A(n2247), .ZN(n2380) );
  NOR2_X1 U2630 ( .A1(n2622), .A2(n2387), .ZN(n2386) );
  INV_X1 U2631 ( .A(n2359), .ZN(n2358) );
  OAI21_X1 U2632 ( .B1(n2240), .B2(n2360), .A(n2599), .ZN(n2359) );
  NAND2_X1 U2633 ( .A1(n3283), .A2(n3313), .ZN(n2364) );
  AND2_X1 U2634 ( .A1(n4482), .A2(n3012), .ZN(n4328) );
  OR2_X1 U2635 ( .A1(n2233), .A2(n4162), .ZN(n4164) );
  OR2_X1 U2636 ( .A1(n4482), .A2(n2964), .ZN(n4406) );
  NAND2_X1 U2637 ( .A1(n2842), .A2(n3006), .ZN(n3003) );
  INV_X1 U2638 ( .A(IR_REG_21__SCAN_IN), .ZN(n2486) );
  NOR2_X1 U2639 ( .A1(n2490), .A2(IR_REG_22__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U2640 ( .A1(n2286), .A2(IR_REG_31__SCAN_IN), .ZN(n2733) );
  INV_X1 U2641 ( .A(IR_REG_19__SCAN_IN), .ZN(n2732) );
  AND2_X1 U2642 ( .A1(n2519), .A2(n2518), .ZN(n4203) );
  NAND2_X1 U2643 ( .A1(n3058), .A2(n3057), .ZN(n3056) );
  OR2_X1 U2644 ( .A1(n2916), .A2(n2917), .ZN(n2290) );
  OAI21_X1 U2645 ( .B1(n4150), .B2(n2832), .A(n2831), .ZN(n4044) );
  INV_X1 U2646 ( .A(n4407), .ZN(n4048) );
  NAND2_X1 U2647 ( .A1(n4549), .A2(n4550), .ZN(n4548) );
  NAND2_X1 U2648 ( .A1(n4593), .A2(n4594), .ZN(n4592) );
  XNOR2_X1 U2649 ( .A(n4117), .B(n4116), .ZN(n4599) );
  NAND2_X1 U2650 ( .A1(n4599), .A2(n4597), .ZN(n4598) );
  NOR2_X1 U2651 ( .A1(n4602), .A2(REG1_REG_16__SCAN_IN), .ZN(n4603) );
  NOR2_X1 U2652 ( .A1(n4615), .A2(n4614), .ZN(n4616) );
  XNOR2_X1 U2653 ( .A(n4124), .B(n2340), .ZN(n2339) );
  INV_X1 U2654 ( .A(n4123), .ZN(n2340) );
  INV_X1 U2655 ( .A(n4128), .ZN(n2284) );
  AOI21_X1 U2656 ( .B1(n4120), .B2(n4121), .A(n4606), .ZN(n2283) );
  XNOR2_X1 U2657 ( .A(n2349), .B(n4130), .ZN(n4135) );
  NOR2_X1 U2658 ( .A1(n4128), .A2(n2269), .ZN(n2349) );
  INV_X1 U2659 ( .A(IR_REG_29__SCAN_IN), .ZN(n2417) );
  INV_X1 U2660 ( .A(n4495), .ZN(n2461) );
  INV_X1 U2661 ( .A(n3642), .ZN(n2295) );
  NOR2_X1 U2662 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2481)
         );
  AOI22_X1 U2663 ( .A1(n2468), .A2(n3307), .B1(n2940), .B2(n2232), .ZN(n2467)
         );
  OR2_X1 U2664 ( .A1(n2232), .A2(n2940), .ZN(n2468) );
  INV_X1 U2665 ( .A(n3841), .ZN(n2415) );
  NOR2_X1 U2666 ( .A1(n2416), .A2(n2412), .ZN(n2411) );
  INV_X1 U2667 ( .A(n3798), .ZN(n2412) );
  INV_X1 U2668 ( .A(n3830), .ZN(n3702) );
  INV_X1 U2669 ( .A(n3732), .ZN(n3739) );
  NAND2_X1 U2670 ( .A1(n3645), .A2(n3644), .ZN(n2462) );
  NAND2_X1 U2671 ( .A1(n3643), .A2(n3642), .ZN(n3645) );
  INV_X1 U2672 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U2673 ( .A1(n2281), .A2(n2280), .ZN(n4112) );
  NAND2_X1 U2674 ( .A1(n4653), .A2(n4567), .ZN(n2280) );
  NAND2_X1 U2675 ( .A1(n4557), .A2(n2245), .ZN(n2281) );
  AND2_X1 U2676 ( .A1(n3748), .A2(n4162), .ZN(n3897) );
  OR2_X1 U2677 ( .A1(n3603), .A2(n3602), .ZN(n4231) );
  INV_X1 U2678 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U2679 ( .A1(n2590), .A2(n2364), .ZN(n2360) );
  NOR2_X1 U2680 ( .A1(n2240), .A2(n2363), .ZN(n2362) );
  INV_X1 U2681 ( .A(n2364), .ZN(n2363) );
  NAND2_X1 U2682 ( .A1(n3180), .A2(n3222), .ZN(n3958) );
  AND4_X1 U2683 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n2905)
         );
  OR2_X1 U2684 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  AND2_X1 U2685 ( .A1(n2336), .A2(n4335), .ZN(n2335) );
  NOR2_X1 U2686 ( .A1(n2809), .A2(n3668), .ZN(n2336) );
  NOR2_X1 U2687 ( .A1(n3432), .A2(n2901), .ZN(n2329) );
  NAND2_X1 U2688 ( .A1(n3175), .A2(n3174), .ZN(n3217) );
  NOR2_X1 U2689 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2479)
         );
  INV_X1 U2690 ( .A(n2485), .ZN(n2453) );
  INV_X1 U2691 ( .A(IR_REG_20__SCAN_IN), .ZN(n2774) );
  AND2_X1 U2692 ( .A1(n2709), .A2(n2674), .ZN(n2321) );
  AND3_X1 U2693 ( .A1(n4933), .A2(n2708), .A3(n2707), .ZN(n2709) );
  INV_X1 U2694 ( .A(IR_REG_14__SCAN_IN), .ZN(n2708) );
  INV_X1 U2695 ( .A(IR_REG_15__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U2696 ( .A1(n2675), .A2(n2674), .ZN(n2706) );
  INV_X1 U2697 ( .A(n2454), .ZN(n2675) );
  NOR2_X1 U2698 ( .A1(n2638), .A2(IR_REG_9__SCAN_IN), .ZN(n2647) );
  OR2_X1 U2699 ( .A1(n3755), .A2(n2260), .ZN(n2447) );
  INV_X1 U2700 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4983) );
  AOI21_X1 U2701 ( .B1(n2421), .B2(n2423), .A(n3465), .ZN(n2420) );
  NOR2_X1 U2702 ( .A1(n2431), .A2(n2968), .ZN(n2421) );
  INV_X1 U2703 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2651) );
  OR2_X1 U2704 ( .A1(n3207), .A2(n2933), .ZN(n2320) );
  NAND2_X1 U2705 ( .A1(n2292), .A2(n2291), .ZN(n3800) );
  AOI21_X1 U2706 ( .B1(n2293), .B2(n2296), .A(n3658), .ZN(n2291) );
  INV_X1 U2707 ( .A(n2455), .ZN(n2296) );
  INV_X1 U2708 ( .A(n3146), .ZN(n2322) );
  INV_X1 U2709 ( .A(n3467), .ZN(n3742) );
  INV_X1 U2710 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3813) );
  AOI21_X1 U2711 ( .B1(n3067), .B2(n3068), .A(n2913), .ZN(n3063) );
  NAND2_X1 U2712 ( .A1(n3682), .A2(n3681), .ZN(n3821) );
  INV_X1 U2713 ( .A(n3552), .ZN(n3555) );
  AND2_X1 U2714 ( .A1(n2320), .A2(n2319), .ZN(n3279) );
  INV_X1 U2715 ( .A(n3280), .ZN(n2319) );
  NAND2_X1 U2716 ( .A1(n2462), .A2(n3651), .ZN(n4494) );
  INV_X1 U2717 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2679) );
  AND4_X1 U2718 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(n3368)
         );
  INV_X1 U2719 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U2720 ( .A1(n3048), .A2(n3036), .ZN(n3037) );
  NAND2_X1 U2721 ( .A1(n3124), .A2(REG1_REG_4__SCAN_IN), .ZN(n3127) );
  NOR2_X1 U2722 ( .A1(n2278), .A2(n2277), .ZN(n2276) );
  NAND2_X1 U2723 ( .A1(n2347), .A2(n2346), .ZN(n4072) );
  NAND2_X1 U2724 ( .A1(n3100), .A2(n4476), .ZN(n2346) );
  NAND2_X1 U2725 ( .A1(n4520), .A2(n4077), .ZN(n4525) );
  NAND2_X1 U2726 ( .A1(n4525), .A2(n4526), .ZN(n4524) );
  XNOR2_X1 U2727 ( .A(n4109), .B(n2352), .ZN(n4558) );
  NAND2_X1 U2728 ( .A1(n4558), .A2(REG2_REG_12__SCAN_IN), .ZN(n4557) );
  XNOR2_X1 U2729 ( .A(n4112), .B(n4651), .ZN(n4581) );
  NAND2_X1 U2730 ( .A1(n4574), .A2(n4083), .ZN(n4084) );
  INV_X1 U2731 ( .A(n2375), .ZN(n4157) );
  OAI21_X1 U2732 ( .B1(n4172), .B2(n2258), .A(n2376), .ZN(n2375) );
  NAND2_X1 U2733 ( .A1(n5076), .A2(n4186), .ZN(n2376) );
  NOR2_X1 U2734 ( .A1(n4017), .A2(n3897), .ZN(n4159) );
  OAI21_X1 U2735 ( .B1(n4276), .B2(n2400), .A(n2397), .ZN(n4208) );
  AOI21_X1 U2736 ( .B1(n2399), .B2(n2398), .A(n2263), .ZN(n2397) );
  INV_X1 U2737 ( .A(n2404), .ZN(n2398) );
  NAND2_X1 U2738 ( .A1(n2546), .A2(DATAI_22_), .ZN(n4270) );
  OR2_X1 U2739 ( .A1(n4007), .A2(n4234), .ZN(n4275) );
  AND3_X1 U2740 ( .A1(n2753), .A2(n2752), .A3(n2751), .ZN(n4297) );
  INV_X1 U2741 ( .A(n2373), .ZN(n2372) );
  NAND2_X1 U2742 ( .A1(n2884), .A2(IR_REG_28__SCAN_IN), .ZN(n2365) );
  OR2_X1 U2743 ( .A1(n2884), .A2(IR_REG_27__SCAN_IN), .ZN(n2366) );
  AND4_X1 U2744 ( .A1(n2720), .A2(n2719), .A3(n2718), .A4(n2717), .ZN(n4332)
         );
  OR3_X1 U2745 ( .A1(n2680), .A2(n2679), .A3(n2678), .ZN(n2689) );
  INV_X1 U2746 ( .A(n2390), .ZN(n2389) );
  OAI21_X1 U2747 ( .B1(n2393), .B2(n2391), .A(n2677), .ZN(n2390) );
  INV_X1 U2748 ( .A(n3416), .ZN(n3628) );
  AOI21_X1 U2749 ( .B1(n2383), .B2(n2382), .A(n2252), .ZN(n2381) );
  INV_X1 U2750 ( .A(n2386), .ZN(n2382) );
  AND2_X1 U2751 ( .A1(n2611), .A2(REG3_REG_8__SCAN_IN), .ZN(n2630) );
  AND2_X1 U2752 ( .A1(n4030), .A2(n2823), .ZN(n4182) );
  AND2_X1 U2753 ( .A1(n4058), .A2(n3071), .ZN(n3170) );
  CLKBUF_X1 U2754 ( .A(n2905), .Z(n3224) );
  INV_X1 U2755 ( .A(n4328), .ZN(n4296) );
  INV_X1 U2756 ( .A(n3071), .ZN(n3175) );
  AND2_X1 U2757 ( .A1(n4034), .A2(n3949), .ZN(n3135) );
  AOI21_X1 U2758 ( .B1(n2862), .B2(n3008), .A(n2861), .ZN(n2962) );
  NOR2_X1 U2759 ( .A1(n4347), .A2(n4348), .ZN(n4346) );
  NOR2_X1 U2760 ( .A1(n4164), .A2(n3740), .ZN(n2892) );
  NAND2_X1 U2761 ( .A1(n4368), .A2(n4186), .ZN(n2331) );
  NAND2_X1 U2762 ( .A1(n2546), .A2(DATAI_25_), .ZN(n4200) );
  NOR3_X1 U2763 ( .A1(n4260), .A2(n2822), .A3(n4240), .ZN(n4218) );
  NOR2_X1 U2764 ( .A1(n4260), .A2(n4240), .ZN(n4245) );
  OR2_X1 U2765 ( .A1(n4283), .A2(n4258), .ZN(n4260) );
  NAND2_X1 U2766 ( .A1(n4308), .A2(n4384), .ZN(n4283) );
  INV_X1 U2767 ( .A(n4329), .ZN(n4385) );
  AND2_X1 U2768 ( .A1(n3579), .A2(n2334), .ZN(n4308) );
  AND2_X1 U2769 ( .A1(n2335), .A2(n4391), .ZN(n2334) );
  NAND2_X1 U2770 ( .A1(n3579), .A2(n2336), .ZN(n4333) );
  NAND2_X1 U2771 ( .A1(n3579), .A2(n4404), .ZN(n3599) );
  AND2_X1 U2772 ( .A1(n3544), .A2(n4490), .ZN(n3579) );
  NOR2_X1 U2773 ( .A1(n4415), .A2(n3648), .ZN(n3544) );
  AND4_X1 U2774 ( .A1(n2673), .A2(n2672), .A3(n2671), .A4(n2670), .ZN(n3864)
         );
  INV_X1 U2775 ( .A(n3415), .ZN(n3529) );
  NAND2_X1 U2776 ( .A1(n3426), .A2(n3529), .ZN(n3455) );
  NAND2_X1 U2777 ( .A1(n2329), .A2(n3474), .ZN(n3406) );
  NOR2_X1 U2778 ( .A1(n3406), .A2(n3516), .ZN(n3426) );
  INV_X1 U2779 ( .A(n2329), .ZN(n3433) );
  AND2_X1 U2780 ( .A1(n2239), .A2(n3189), .ZN(n3363) );
  NAND2_X1 U2781 ( .A1(n3189), .A2(n2235), .ZN(n3297) );
  NAND2_X1 U2782 ( .A1(n3189), .A2(n3283), .ZN(n3299) );
  NOR2_X1 U2783 ( .A1(n4670), .A2(n3261), .ZN(n3190) );
  NAND2_X1 U2784 ( .A1(n3245), .A2(n4664), .ZN(n4681) );
  NAND2_X1 U2785 ( .A1(n2325), .A2(n3080), .ZN(n4670) );
  INV_X1 U2786 ( .A(n3217), .ZN(n2325) );
  AND2_X1 U2787 ( .A1(n4026), .A2(n3135), .ZN(n4669) );
  AND3_X1 U2788 ( .A1(n2858), .A2(n2857), .A3(n2960), .ZN(n2869) );
  AND2_X1 U2789 ( .A1(n2899), .A2(n4645), .ZN(n3139) );
  XNOR2_X1 U2790 ( .A(n2775), .B(n2774), .ZN(n4026) );
  NAND2_X1 U2791 ( .A1(n2773), .A2(IR_REG_31__SCAN_IN), .ZN(n2775) );
  NOR2_X1 U2792 ( .A1(n2721), .A2(IR_REG_17__SCAN_IN), .ZN(n2722) );
  XNOR2_X1 U2793 ( .A(n2659), .B(IR_REG_11__SCAN_IN), .ZN(n4097) );
  XNOR2_X1 U2794 ( .A(n2629), .B(IR_REG_9__SCAN_IN), .ZN(n4098) );
  INV_X1 U2795 ( .A(IR_REG_3__SCAN_IN), .ZN(n2575) );
  INV_X1 U2796 ( .A(IR_REG_2__SCAN_IN), .ZN(n2565) );
  OAI21_X1 U2797 ( .B1(n3755), .B2(n2302), .A(n2299), .ZN(n2298) );
  NAND2_X1 U2798 ( .A1(n2302), .A2(n2300), .ZN(n2299) );
  NAND2_X1 U2799 ( .A1(n2304), .A2(n2446), .ZN(n2300) );
  NAND2_X1 U2800 ( .A1(n2448), .A2(n3755), .ZN(n2301) );
  INV_X1 U2801 ( .A(n2307), .ZN(n2306) );
  AND4_X1 U2802 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n3562)
         );
  NOR2_X1 U2803 ( .A1(n2424), .A2(n2422), .ZN(n3466) );
  NOR2_X1 U2804 ( .A1(n2426), .A2(n2425), .ZN(n2424) );
  AND2_X1 U2805 ( .A1(n2289), .A2(n2256), .ZN(n3152) );
  NAND2_X1 U2806 ( .A1(n3838), .A2(n3840), .ZN(n3770) );
  NOR2_X1 U2807 ( .A1(n3746), .A2(n2437), .ZN(n2436) );
  INV_X1 U2808 ( .A(n2443), .ZN(n2437) );
  OAI21_X1 U2809 ( .B1(n3746), .B2(n2440), .A(n2439), .ZN(n2438) );
  AND2_X1 U2810 ( .A1(n2443), .A2(n2447), .ZN(n2440) );
  NAND2_X1 U2811 ( .A1(n3746), .A2(n2443), .ZN(n2439) );
  NAND2_X1 U2812 ( .A1(n3746), .A2(n2442), .ZN(n2441) );
  INV_X1 U2813 ( .A(n2447), .ZN(n2442) );
  INV_X1 U2814 ( .A(n3174), .ZN(n3177) );
  AND2_X1 U2815 ( .A1(n2532), .A2(n2531), .ZN(n4244) );
  INV_X1 U2816 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4955) );
  INV_X1 U2817 ( .A(n3653), .ZN(n4490) );
  AND4_X1 U2818 ( .A1(n2695), .A2(n2694), .A3(n2693), .A4(n2692), .ZN(n4407)
         );
  INV_X1 U2819 ( .A(n3193), .ZN(n3206) );
  AOI21_X1 U2820 ( .B1(n3356), .B2(n3353), .A(n3354), .ZN(n3380) );
  NAND2_X1 U2821 ( .A1(n2309), .A2(n2310), .ZN(n3700) );
  AND4_X1 U2822 ( .A1(n2705), .A2(n2704), .A3(n2703), .A4(n2702), .ZN(n3845)
         );
  NAND2_X1 U2823 ( .A1(n2982), .A2(n2978), .ZN(n3863) );
  INV_X1 U2824 ( .A(n3858), .ZN(n4498) );
  AND2_X1 U2825 ( .A1(n2976), .A2(n3054), .ZN(n4503) );
  NAND2_X1 U2826 ( .A1(n2525), .A2(n2524), .ZN(n4215) );
  INV_X1 U2827 ( .A(n4244), .ZN(n4045) );
  OAI211_X1 U2828 ( .C1(n4262), .C2(n2832), .A(n2535), .B(n2534), .ZN(n4280)
         );
  INV_X1 U2829 ( .A(n3845), .ZN(n4484) );
  OR2_X1 U2830 ( .A1(n2899), .A2(n3005), .ZN(n4057) );
  NAND3_X1 U2831 ( .A1(n4062), .A2(REG2_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n4061) );
  AOI21_X1 U2832 ( .B1(n4061), .B2(n3112), .A(n3113), .ZN(n2285) );
  XNOR2_X1 U2833 ( .A(n3035), .B(n3046), .ZN(n3049) );
  AOI22_X1 U2834 ( .A1(n3123), .A2(REG2_REG_4__SCAN_IN), .B1(n4477), .B2(n3025), .ZN(n3087) );
  NOR2_X1 U2835 ( .A1(n3087), .A2(n3086), .ZN(n3085) );
  NOR2_X1 U2836 ( .A1(n3090), .A2(n3089), .ZN(n3088) );
  AND2_X1 U2837 ( .A1(n3127), .A2(n2345), .ZN(n3090) );
  NAND2_X1 U2838 ( .A1(n3037), .A2(n4477), .ZN(n2345) );
  XNOR2_X1 U2839 ( .A(n2275), .B(n2348), .ZN(n3095) );
  INV_X1 U2840 ( .A(n2347), .ZN(n3099) );
  AOI22_X1 U2841 ( .A1(n3095), .A2(REG2_REG_6__SCAN_IN), .B1(n2275), .B2(n4476), .ZN(n3097) );
  NOR2_X1 U2842 ( .A1(n3097), .A2(n3096), .ZN(n4099) );
  INV_X1 U2843 ( .A(n4072), .ZN(n4075) );
  NAND2_X1 U2844 ( .A1(n4515), .A2(n4104), .ZN(n4528) );
  XNOR2_X1 U2845 ( .A(n4079), .B(n2344), .ZN(n4542) );
  NAND2_X1 U2846 ( .A1(n4536), .A2(n4107), .ZN(n4549) );
  NAND2_X1 U2847 ( .A1(n4562), .A2(n4082), .ZN(n4575) );
  NAND2_X1 U2848 ( .A1(n4575), .A2(n4576), .ZN(n4574) );
  NAND2_X1 U2849 ( .A1(n4557), .A2(n4110), .ZN(n4570) );
  XNOR2_X1 U2850 ( .A(n4084), .B(n4651), .ZN(n4585) );
  INV_X1 U2851 ( .A(n4588), .ZN(n2272) );
  INV_X1 U2852 ( .A(n2273), .ZN(n4589) );
  NAND2_X1 U2853 ( .A1(n4598), .A2(n4118), .ZN(n4607) );
  NOR2_X1 U2854 ( .A1(n4088), .A2(n4603), .ZN(n4615) );
  AOI21_X1 U2855 ( .B1(n2875), .B2(n3948), .A(n2874), .ZN(n2876) );
  OR2_X1 U2856 ( .A1(n2513), .A2(n2512), .ZN(n4185) );
  NAND2_X1 U2857 ( .A1(n2401), .A2(n2402), .ZN(n4228) );
  NAND2_X1 U2858 ( .A1(n4276), .A2(n2404), .ZN(n2401) );
  AND2_X1 U2859 ( .A1(n2408), .A2(n2406), .ZN(n4257) );
  INV_X1 U2860 ( .A(n3691), .ZN(n4384) );
  NAND4_X1 U2861 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(n4312)
         );
  AND2_X1 U2862 ( .A1(n4507), .A2(n4241), .ZN(n4313) );
  NAND2_X1 U2863 ( .A1(n3542), .A2(n2699), .ZN(n3577) );
  OR2_X1 U2864 ( .A1(n3455), .A2(n3613), .ZN(n4415) );
  NAND2_X1 U2865 ( .A1(n3449), .A2(n3932), .ZN(n3448) );
  NAND2_X1 U2866 ( .A1(n2395), .A2(n2393), .ZN(n3449) );
  NAND2_X1 U2867 ( .A1(n3405), .A2(n2231), .ZN(n2395) );
  NAND2_X1 U2868 ( .A1(n2392), .A2(n2396), .ZN(n3425) );
  OR2_X1 U2869 ( .A1(n3405), .A2(n2662), .ZN(n2392) );
  NAND2_X1 U2870 ( .A1(n2610), .A2(n2386), .ZN(n2385) );
  NAND2_X1 U2871 ( .A1(n2357), .A2(n2364), .ZN(n3289) );
  OR2_X1 U2872 ( .A1(n3232), .A2(n2590), .ZN(n2357) );
  INV_X1 U2873 ( .A(n4339), .ZN(n4637) );
  AND4_X1 U2874 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(n3254)
         );
  INV_X1 U2875 ( .A(n4261), .ZN(n4634) );
  AND2_X2 U2876 ( .A1(n2869), .A2(n2962), .ZN(n4700) );
  INV_X1 U2877 ( .A(n4700), .ZN(n4697) );
  AND2_X2 U2878 ( .A1(n2869), .A2(n3143), .ZN(n4690) );
  NAND2_X1 U2879 ( .A1(n3003), .A2(n3139), .ZN(n4643) );
  NAND2_X1 U2880 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2418) );
  XNOR2_X1 U2881 ( .A(n2841), .B(IR_REG_26__SCAN_IN), .ZN(n3006) );
  OR2_X1 U2882 ( .A1(n2255), .A2(n3000), .ZN(n2841) );
  OR2_X1 U2883 ( .A1(n2837), .A2(n2255), .ZN(n2992) );
  MUX2_X1 U2884 ( .A(n3000), .B(n2836), .S(IR_REG_25__SCAN_IN), .Z(n2837) );
  XNOR2_X1 U2885 ( .A(n2839), .B(IR_REG_24__SCAN_IN), .ZN(n3004) );
  AND2_X1 U2886 ( .A1(n3011), .A2(STATE_REG_SCAN_IN), .ZN(n4645) );
  AND2_X1 U2887 ( .A1(n2781), .A2(n2780), .ZN(n4471) );
  INV_X1 U2888 ( .A(n3949), .ZN(n3955) );
  AND2_X1 U2889 ( .A1(n2773), .A2(n2734), .ZN(n4473) );
  NAND2_X1 U2890 ( .A1(n2343), .A2(IR_REG_31__SCAN_IN), .ZN(n2555) );
  INV_X1 U2891 ( .A(IR_REG_1__SCAN_IN), .ZN(n2353) );
  AND2_X1 U2892 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2354)
         );
  NAND2_X1 U2893 ( .A1(n3056), .A2(n2290), .ZN(n3077) );
  NAND2_X1 U2894 ( .A1(n2338), .A2(n2282), .ZN(U3258) );
  AOI21_X1 U2895 ( .B1(n2284), .B2(n2283), .A(n4122), .ZN(n2282) );
  NAND2_X1 U2896 ( .A1(n2339), .A2(n4613), .ZN(n2338) );
  NAND3_X4 U2897 ( .A1(n2366), .A2(n2365), .A3(n2492), .ZN(n2546) );
  AND2_X1 U2898 ( .A1(n2396), .A2(n2242), .ZN(n2231) );
  AND2_X1 U2899 ( .A1(n2938), .A2(n2937), .ZN(n2232) );
  OR3_X1 U2900 ( .A1(n4260), .A2(n2332), .A3(n2331), .ZN(n2233) );
  AND2_X1 U2901 ( .A1(n2309), .A2(n2307), .ZN(n2234) );
  INV_X1 U2902 ( .A(n3250), .ZN(n3283) );
  AND2_X1 U2903 ( .A1(n3283), .A2(n3310), .ZN(n2235) );
  NAND2_X1 U2904 ( .A1(n4050), .A2(n2901), .ZN(n2236) );
  AND2_X1 U2905 ( .A1(n2384), .A2(n2236), .ZN(n2237) );
  AND2_X1 U2906 ( .A1(n2497), .A2(n2417), .ZN(n2238) );
  INV_X1 U2907 ( .A(n4051), .ZN(n3438) );
  AND2_X1 U2908 ( .A1(n2333), .A2(n3367), .ZN(n2239) );
  INV_X1 U2909 ( .A(n4476), .ZN(n2348) );
  AND2_X1 U2910 ( .A1(n4318), .A2(n4319), .ZN(n3923) );
  INV_X1 U2911 ( .A(n4186), .ZN(n2864) );
  NAND2_X1 U2912 ( .A1(n2546), .A2(DATAI_26_), .ZN(n4186) );
  NOR2_X1 U2913 ( .A1(n4052), .A2(n3300), .ZN(n2240) );
  INV_X1 U2914 ( .A(n2384), .ZN(n2383) );
  NAND2_X1 U2915 ( .A1(n2621), .A2(n2244), .ZN(n2384) );
  OR2_X1 U2916 ( .A1(n3085), .A2(n2276), .ZN(n2275) );
  OR2_X1 U2917 ( .A1(n4046), .A2(n3691), .ZN(n2241) );
  NAND2_X1 U2918 ( .A1(n3416), .A2(n3415), .ZN(n2242) );
  AND2_X1 U2919 ( .A1(n4479), .A2(REG2_REG_2__SCAN_IN), .ZN(n2243) );
  OR2_X1 U2920 ( .A1(n4051), .A2(n3342), .ZN(n2244) );
  INV_X1 U2921 ( .A(n2968), .ZN(n2427) );
  AND2_X1 U2922 ( .A1(n4110), .A2(n2279), .ZN(n2245) );
  NOR2_X1 U2923 ( .A1(n2940), .A2(n3307), .ZN(n2246) );
  INV_X1 U2924 ( .A(n3342), .ZN(n3383) );
  AND2_X1 U2925 ( .A1(n3476), .A2(n3437), .ZN(n2247) );
  AND2_X1 U2926 ( .A1(n3628), .A2(n3529), .ZN(n2248) );
  AND2_X1 U2927 ( .A1(n2273), .A2(n2272), .ZN(n2249) );
  OR2_X1 U2928 ( .A1(n2454), .A2(n2453), .ZN(n2250) );
  AND4_X1 U2929 ( .A1(n2479), .A2(n2480), .A3(n2477), .A4(n2486), .ZN(n2251)
         );
  INV_X1 U2930 ( .A(n2400), .ZN(n2399) );
  NAND2_X1 U2931 ( .A1(n2402), .A2(n2259), .ZN(n2400) );
  AND2_X1 U2932 ( .A1(n3342), .A2(n4051), .ZN(n2252) );
  INV_X1 U2933 ( .A(n2407), .ZN(n2406) );
  NAND2_X1 U2934 ( .A1(n4265), .A2(n2241), .ZN(n2407) );
  INV_X1 U2935 ( .A(IR_REG_31__SCAN_IN), .ZN(n3000) );
  AND2_X1 U2936 ( .A1(n2381), .A2(n2236), .ZN(n2253) );
  OR2_X1 U2937 ( .A1(n3700), .A2(n3699), .ZN(n2254) );
  AND2_X1 U2938 ( .A1(n2488), .A2(n2471), .ZN(n2255) );
  NAND2_X1 U2939 ( .A1(n2924), .A2(n2923), .ZN(n2256) );
  AND2_X1 U2940 ( .A1(n2231), .A2(n3932), .ZN(n2257) );
  INV_X1 U2941 ( .A(IR_REG_28__SCAN_IN), .ZN(n2497) );
  INV_X1 U2942 ( .A(n3755), .ZN(n2446) );
  INV_X1 U2943 ( .A(n3932), .ZN(n2391) );
  NAND2_X1 U2944 ( .A1(n2844), .A2(n3006), .ZN(n2899) );
  AND2_X1 U2945 ( .A1(n2510), .A2(n2509), .ZN(n3748) );
  INV_X1 U2946 ( .A(n3748), .ZN(n4180) );
  INV_X1 U2947 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2277) );
  OAI211_X1 U2948 ( .C1(n3876), .C2(n4250), .A(n2759), .B(n2758), .ZN(n4267)
         );
  INV_X1 U2949 ( .A(IR_REG_6__SCAN_IN), .ZN(n2607) );
  AND2_X1 U2950 ( .A1(n4197), .A2(n2864), .ZN(n2258) );
  OR2_X1 U2951 ( .A1(n4267), .A2(n4240), .ZN(n2259) );
  AND2_X1 U2952 ( .A1(n3731), .A2(n3730), .ZN(n2260) );
  AND2_X1 U2953 ( .A1(n2772), .A2(n2771), .ZN(n4160) );
  NAND2_X1 U2954 ( .A1(n2557), .A2(n2323), .ZN(n3222) );
  INV_X1 U2955 ( .A(n2433), .ZN(n3553) );
  INV_X1 U2956 ( .A(n2330), .ZN(n4202) );
  NOR3_X1 U2957 ( .A1(n4260), .A2(n2332), .A3(n2822), .ZN(n2330) );
  OR2_X1 U2958 ( .A1(n4102), .A2(n4101), .ZN(n2261) );
  OR2_X1 U2959 ( .A1(n4215), .A2(n2761), .ZN(n2262) );
  INV_X1 U2960 ( .A(n2457), .ZN(n4493) );
  NOR2_X1 U2961 ( .A1(n2462), .A2(n3651), .ZN(n2457) );
  NAND2_X1 U2962 ( .A1(n3579), .A2(n2335), .ZN(n2337) );
  INV_X1 U2963 ( .A(n2949), .ZN(n3367) );
  INV_X1 U2964 ( .A(n2313), .ZN(n2312) );
  NAND2_X1 U2965 ( .A1(n2314), .A2(n3681), .ZN(n2313) );
  INV_X1 U2966 ( .A(n2448), .ZN(n2304) );
  NOR2_X1 U2967 ( .A1(n3851), .A2(n2449), .ZN(n2448) );
  AND2_X1 U2968 ( .A1(n4267), .A2(n4240), .ZN(n2263) );
  AND2_X1 U2969 ( .A1(n2302), .A2(n2446), .ZN(n2264) );
  OR2_X1 U2970 ( .A1(n2424), .A2(n2428), .ZN(n2265) );
  AND2_X1 U2971 ( .A1(n2305), .A2(n3711), .ZN(n2266) );
  INV_X1 U2972 ( .A(n2785), .ZN(n3220) );
  NAND2_X1 U2973 ( .A1(n3961), .A2(n3958), .ZN(n2785) );
  OAI21_X1 U2974 ( .B1(n2610), .B2(n2384), .A(n2381), .ZN(n3435) );
  NAND2_X1 U2975 ( .A1(n2385), .A2(n2621), .ZN(n3323) );
  INV_X1 U2976 ( .A(n3840), .ZN(n2416) );
  NAND2_X1 U2977 ( .A1(n2361), .A2(n2358), .ZN(n3274) );
  NOR2_X1 U2978 ( .A1(n3279), .A2(n2232), .ZN(n2267) );
  INV_X1 U2979 ( .A(n3353), .ZN(n2432) );
  INV_X1 U2980 ( .A(n3686), .ZN(n4391) );
  AND2_X1 U2981 ( .A1(n3189), .A2(n2333), .ZN(n2268) );
  AND2_X1 U2982 ( .A1(n2546), .A2(DATAI_24_), .ZN(n2822) );
  INV_X1 U2983 ( .A(n4247), .ZN(n4240) );
  NAND2_X1 U2984 ( .A1(n2546), .A2(DATAI_23_), .ZN(n4247) );
  INV_X1 U2985 ( .A(n2822), .ZN(n4368) );
  INV_X1 U2986 ( .A(n2356), .ZN(n2274) );
  AND2_X1 U2987 ( .A1(n4115), .A2(REG2_REG_15__SCAN_IN), .ZN(n2356) );
  INV_X1 U2988 ( .A(n4556), .ZN(n2352) );
  INV_X1 U2989 ( .A(n4514), .ZN(n2355) );
  INV_X1 U2990 ( .A(n4119), .ZN(n4646) );
  XNOR2_X1 U2991 ( .A(n2639), .B(IR_REG_10__SCAN_IN), .ZN(n4535) );
  INV_X1 U2992 ( .A(n4535), .ZN(n2344) );
  INV_X1 U2993 ( .A(DATAI_1_), .ZN(n2367) );
  AND2_X1 U2994 ( .A1(n4474), .A2(REG2_REG_18__SCAN_IN), .ZN(n2269) );
  AND2_X1 U2995 ( .A1(n2589), .A2(n2588), .ZN(n3038) );
  INV_X1 U2996 ( .A(n3038), .ZN(n2278) );
  NOR3_X1 U2997 ( .A1(n4606), .A2(n2285), .A3(n3114), .ZN(n3122) );
  INV_X1 U2998 ( .A(n2722), .ZN(n2731) );
  NAND2_X1 U2999 ( .A1(n2722), .A2(n2287), .ZN(n2286) );
  INV_X1 U3000 ( .A(IR_REG_18__SCAN_IN), .ZN(n2287) );
  NAND3_X1 U3001 ( .A1(n3056), .A2(n2290), .A3(n2288), .ZN(n2289) );
  INV_X1 U3002 ( .A(n2289), .ZN(n3076) );
  NAND2_X1 U3003 ( .A1(n3643), .A2(n2293), .ZN(n2292) );
  NAND2_X1 U3004 ( .A1(n3792), .A2(n2264), .ZN(n2297) );
  OAI211_X1 U3005 ( .C1(n3792), .C2(n2301), .A(n2298), .B(n2297), .ZN(n3761)
         );
  NAND2_X1 U3006 ( .A1(n3792), .A2(n3790), .ZN(n3725) );
  OAI21_X1 U3007 ( .B1(n3682), .B2(n2306), .A(n2266), .ZN(n2466) );
  INV_X1 U3008 ( .A(n3696), .ZN(n2314) );
  INV_X1 U3009 ( .A(n2467), .ZN(n2316) );
  NAND2_X1 U3010 ( .A1(n3207), .A2(n2318), .ZN(n2317) );
  INV_X1 U3011 ( .A(n2320), .ZN(n3281) );
  NAND2_X1 U3012 ( .A1(n2675), .A2(n2321), .ZN(n2721) );
  AND4_X2 U3013 ( .A1(n2452), .A2(n2251), .A3(n2485), .A4(n2476), .ZN(n2488)
         );
  NAND2_X1 U3014 ( .A1(n2327), .A2(n2488), .ZN(n2326) );
  INV_X1 U3015 ( .A(n2488), .ZN(n2777) );
  INV_X1 U3016 ( .A(n2337), .ZN(n4334) );
  INV_X1 U3017 ( .A(IR_REG_1__SCAN_IN), .ZN(n2341) );
  INV_X1 U3018 ( .A(IR_REG_0__SCAN_IN), .ZN(n2342) );
  MUX2_X1 U3019 ( .A(REG2_REG_1__SCAN_IN), .B(n2536), .S(n2230), .Z(n4062) );
  NOR2_X1 U3020 ( .A1(n3457), .A2(n4581), .ZN(n4580) );
  AOI21_X1 U3021 ( .B1(n4135), .B2(n4568), .A(n4134), .ZN(n4136) );
  XOR2_X1 U3022 ( .A(n4081), .B(n4556), .Z(n4563) );
  OAI21_X1 U3023 ( .B1(n4072), .B2(REG1_REG_7__SCAN_IN), .A(n4475), .ZN(n4073)
         );
  XOR2_X1 U3024 ( .A(n4514), .B(n4076), .Z(n4521) );
  XNOR2_X2 U3025 ( .A(n2555), .B(IR_REG_2__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U3026 ( .A1(n3232), .A2(n2362), .ZN(n2361) );
  MUX2_X1 U3027 ( .A(n2368), .B(n2367), .S(n2546), .Z(n3174) );
  NAND2_X1 U3028 ( .A1(n2369), .A2(n2372), .ZN(n2714) );
  NAND2_X1 U3029 ( .A1(n2688), .A2(n2370), .ZN(n2369) );
  NAND2_X1 U3030 ( .A1(n2610), .A2(n2253), .ZN(n2379) );
  NAND2_X1 U3031 ( .A1(n2379), .A2(n2380), .ZN(n3390) );
  NAND2_X1 U3032 ( .A1(n2610), .A2(n2609), .ZN(n3365) );
  INV_X1 U3033 ( .A(n2609), .ZN(n2387) );
  NAND2_X1 U3034 ( .A1(n3405), .A2(n2257), .ZN(n2388) );
  NAND2_X1 U3035 ( .A1(n2388), .A2(n2389), .ZN(n3499) );
  NAND2_X1 U3036 ( .A1(n2410), .A2(n2413), .ZN(n3682) );
  NAND2_X1 U3037 ( .A1(n3666), .A2(n2411), .ZN(n2410) );
  NAND2_X1 U3038 ( .A1(n2498), .A2(n2497), .ZN(n2499) );
  NAND2_X1 U3039 ( .A1(n2498), .A2(n2238), .ZN(n2419) );
  OAI21_X1 U3040 ( .B1(n3356), .B2(n2422), .A(n2420), .ZN(n2433) );
  OR2_X1 U3041 ( .A1(n2959), .A2(n2958), .ZN(n2434) );
  NAND2_X1 U3042 ( .A1(n3725), .A2(n2436), .ZN(n2435) );
  OAI211_X1 U3043 ( .C1(n3725), .C2(n2441), .A(n2438), .B(n2435), .ZN(n3754)
         );
  NAND2_X1 U3044 ( .A1(n3725), .A2(n3791), .ZN(n3853) );
  NAND2_X1 U3045 ( .A1(n2476), .A2(n2566), .ZN(n2587) );
  NOR2_X1 U3046 ( .A1(n3715), .A2(n3717), .ZN(n2465) );
  AND2_X1 U3047 ( .A1(n2488), .A2(n2470), .ZN(n2835) );
  NAND2_X1 U3048 ( .A1(n2488), .A2(n2469), .ZN(n2824) );
  NAND2_X1 U3049 ( .A1(n2488), .A2(n2487), .ZN(n2780) );
  AND2_X1 U3050 ( .A1(n2546), .A2(n3013), .ZN(n3026) );
  AND2_X1 U3051 ( .A1(n2546), .A2(DATAI_21_), .ZN(n3691) );
  AND2_X1 U3052 ( .A1(n2546), .A2(DATAI_20_), .ZN(n3686) );
  XNOR2_X1 U3053 ( .A(n2915), .B(n2917), .ZN(n3058) );
  INV_X1 U3054 ( .A(n2905), .ZN(n2547) );
  NOR2_X1 U3055 ( .A1(n2587), .A2(IR_REG_5__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U3056 ( .A1(n2499), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  NAND2_X2 U3057 ( .A1(n3145), .A2(n4261), .ZN(n4507) );
  INV_X1 U3058 ( .A(n4479), .ZN(n2556) );
  INV_X1 U3059 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2678) );
  OR2_X1 U3060 ( .A1(n4486), .A2(n3648), .ZN(n2473) );
  NOR2_X1 U3061 ( .A1(n2865), .A2(n2892), .ZN(n2474) );
  AND2_X1 U3062 ( .A1(n2546), .A2(DATAI_28_), .ZN(n3740) );
  INV_X1 U3063 ( .A(IR_REG_24__SCAN_IN), .ZN(n2489) );
  INV_X1 U3064 ( .A(IR_REG_25__SCAN_IN), .ZN(n2491) );
  AND2_X1 U3065 ( .A1(n4291), .A2(n2813), .ZN(n4233) );
  OR2_X1 U3066 ( .A1(n4473), .A2(n4034), .ZN(n2973) );
  AND2_X1 U3067 ( .A1(n3908), .A2(n4301), .ZN(n2742) );
  INV_X1 U3068 ( .A(n3923), .ZN(n2724) );
  NOR2_X1 U3069 ( .A1(n4160), .A2(n3747), .ZN(n2874) );
  OAI21_X1 U3070 ( .B1(n3161), .B2(n2569), .A(n2568), .ZN(n3191) );
  NAND2_X1 U3071 ( .A1(n2905), .A2(n3177), .ZN(n3957) );
  INV_X1 U3072 ( .A(IR_REG_22__SCAN_IN), .ZN(n2487) );
  AND2_X1 U3073 ( .A1(n2943), .A2(n2942), .ZN(n2944) );
  AND2_X1 U3074 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  INV_X1 U3075 ( .A(n2947), .ZN(n3467) );
  NAND2_X1 U3076 ( .A1(n3680), .A2(n3679), .ZN(n3681) );
  INV_X1 U3077 ( .A(n2549), .ZN(n2504) );
  NOR2_X1 U3078 ( .A1(n2519), .A2(n2511), .ZN(n2512) );
  NAND2_X1 U3079 ( .A1(n2686), .A2(n2473), .ZN(n2688) );
  AND2_X1 U3080 ( .A1(REG3_REG_10__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2493) );
  INV_X1 U3081 ( .A(n3004), .ZN(n2859) );
  NOR2_X1 U3082 ( .A1(n2652), .A2(n2651), .ZN(n2663) );
  AND3_X1 U3083 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2591) );
  OR2_X1 U3084 ( .A1(n2736), .A2(n2494), .ZN(n2744) );
  INV_X1 U3085 ( .A(n3515), .ZN(n3531) );
  NAND2_X1 U3086 ( .A1(n2715), .A2(REG3_REG_18__SCAN_IN), .ZN(n2736) );
  INV_X1 U3087 ( .A(n4471), .ZN(n4034) );
  OR2_X1 U3088 ( .A1(n4220), .A2(n2832), .ZN(n2532) );
  INV_X1 U3089 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4879) );
  INV_X1 U3090 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4483) );
  INV_X1 U3091 ( .A(n4405), .ZN(n4327) );
  INV_X1 U3092 ( .A(n4162), .ZN(n4355) );
  AOI21_X1 U3093 ( .B1(n4244), .B2(n4368), .A(n2760), .ZN(n4191) );
  NAND2_X1 U3094 ( .A1(n2630), .A2(n2493), .ZN(n2640) );
  AND2_X1 U3095 ( .A1(n2860), .A2(n2859), .ZN(n2861) );
  AND2_X1 U3096 ( .A1(n2546), .A2(DATAI_27_), .ZN(n4162) );
  INV_X1 U3097 ( .A(n4270), .ZN(n4258) );
  INV_X1 U3098 ( .A(n4052), .ZN(n3332) );
  NAND2_X1 U3099 ( .A1(n4472), .A2(n3135), .ZN(n4405) );
  AND2_X1 U3100 ( .A1(n2495), .A2(n2764), .ZN(n4165) );
  NAND2_X1 U3101 ( .A1(n2755), .A2(REG3_REG_23__SCAN_IN), .ZN(n2757) );
  AND2_X1 U3102 ( .A1(n4150), .A2(n2765), .ZN(n3752) );
  NOR2_X1 U3103 ( .A1(n2689), .A2(n4483), .ZN(n2700) );
  AND2_X1 U3104 ( .A1(n2700), .A2(REG3_REG_17__SCAN_IN), .ZN(n2715) );
  INV_X1 U3105 ( .A(n2975), .ZN(n2982) );
  OR2_X1 U3106 ( .A1(n2764), .A2(n4780), .ZN(n4150) );
  INV_X1 U3107 ( .A(n2747), .ZN(n2832) );
  INV_X1 U3108 ( .A(n3368), .ZN(n3292) );
  NOR2_X1 U3109 ( .A1(n4513), .A2(n4037), .ZN(n4568) );
  NAND3_X1 U3110 ( .A1(n3139), .A2(n4688), .A3(n3949), .ZN(n4261) );
  INV_X1 U3111 ( .A(n4182), .ZN(n4324) );
  INV_X1 U3112 ( .A(n4473), .ZN(n4133) );
  INV_X1 U3113 ( .A(n4342), .ZN(n4304) );
  INV_X1 U3114 ( .A(n4412), .ZN(n2866) );
  OR2_X1 U3115 ( .A1(n3138), .A2(n4471), .ZN(n4664) );
  INV_X1 U3116 ( .A(n4466), .ZN(n4423) );
  INV_X1 U3117 ( .A(n4664), .ZN(n4688) );
  INV_X1 U3118 ( .A(n4645), .ZN(n3005) );
  XNOR2_X1 U3119 ( .A(n2661), .B(IR_REG_12__SCAN_IN), .ZN(n4556) );
  AND2_X1 U3120 ( .A1(n3027), .A2(n3014), .ZN(n4612) );
  NAND2_X1 U3121 ( .A1(n2982), .A2(n2967), .ZN(n3858) );
  INV_X1 U3122 ( .A(n4160), .ZN(n4149) );
  INV_X1 U3123 ( .A(n3180), .ZN(n4056) );
  INV_X1 U3124 ( .A(n4568), .ZN(n4606) );
  NAND2_X1 U3125 ( .A1(n3028), .A2(n4482), .ZN(n4619) );
  NAND2_X1 U3126 ( .A1(n4507), .A2(n3173), .ZN(n4339) );
  NAND2_X1 U3127 ( .A1(n4507), .A2(n3246), .ZN(n4342) );
  OR2_X1 U3128 ( .A1(n4151), .A2(n4412), .ZN(n2893) );
  NAND2_X1 U3129 ( .A1(n4700), .A2(n4669), .ZN(n4412) );
  OR2_X1 U3130 ( .A1(n4151), .A2(n4466), .ZN(n2897) );
  NAND2_X1 U3131 ( .A1(n4690), .A2(n4669), .ZN(n4466) );
  INV_X1 U3132 ( .A(n4690), .ZN(n4689) );
  INV_X1 U3133 ( .A(n4643), .ZN(n4644) );
  XNOR2_X1 U3134 ( .A(n2825), .B(n2497), .ZN(n4482) );
  INV_X1 U3135 ( .A(n4097), .ZN(n4655) );
  INV_X2 U3136 ( .A(n4057), .ZN(U4043) );
  NAND2_X1 U3137 ( .A1(n2497), .A2(IR_REG_27__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3138 ( .A1(n2591), .A2(REG3_REG_6__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U3139 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2494) );
  INV_X1 U3140 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2511) );
  OR2_X1 U3141 ( .A1(n2512), .A2(REG3_REG_27__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3142 ( .A1(n2512), .A2(REG3_REG_27__SCAN_IN), .ZN(n2764) );
  INV_X1 U3143 ( .A(n2824), .ZN(n2498) );
  XNOR2_X2 U3144 ( .A(n2500), .B(IR_REG_29__SCAN_IN), .ZN(n2998) );
  AND2_X4 U3145 ( .A1(n4469), .A2(n2998), .ZN(n2747) );
  NAND2_X1 U3146 ( .A1(n4165), .A2(n2747), .ZN(n2510) );
  INV_X1 U3147 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2507) );
  INV_X1 U31480 ( .A(n2998), .ZN(n2501) );
  NAND2_X1 U31490 ( .A1(n4469), .A2(n2501), .ZN(n2537) );
  NAND2_X1 U3150 ( .A1(n2766), .A2(REG0_REG_27__SCAN_IN), .ZN(n2506) );
  INV_X2 U3152 ( .A(n2504), .ZN(n2826) );
  NAND2_X1 U3153 ( .A1(n3873), .A2(REG1_REG_27__SCAN_IN), .ZN(n2505) );
  OAI211_X1 U3154 ( .C1(n2507), .C2(n3876), .A(n2506), .B(n2505), .ZN(n2508)
         );
  INV_X1 U3155 ( .A(n2508), .ZN(n2509) );
  AND2_X1 U3156 ( .A1(n2519), .A2(n2511), .ZN(n2513) );
  INV_X1 U3157 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U3158 ( .A1(n2766), .A2(REG0_REG_26__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U3159 ( .A1(n2826), .A2(REG1_REG_26__SCAN_IN), .ZN(n2514) );
  OAI211_X1 U3160 ( .C1(n4184), .C2(n3876), .A(n2515), .B(n2514), .ZN(n2516)
         );
  INV_X1 U3161 ( .A(n2516), .ZN(n2517) );
  INV_X1 U3162 ( .A(n4197), .ZN(n5076) );
  NAND2_X1 U3163 ( .A1(n2527), .A2(n4955), .ZN(n2518) );
  NAND2_X1 U3164 ( .A1(n4203), .A2(n2747), .ZN(n2525) );
  INV_X1 U3165 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3166 ( .A1(n2766), .A2(REG0_REG_25__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U3167 ( .A1(n3873), .A2(REG1_REG_25__SCAN_IN), .ZN(n2520) );
  OAI211_X1 U3168 ( .C1(n2522), .C2(n3876), .A(n2521), .B(n2520), .ZN(n2523)
         );
  INV_X1 U3169 ( .A(n2523), .ZN(n2524) );
  INV_X1 U3170 ( .A(n4215), .ZN(n4178) );
  INV_X1 U3171 ( .A(n4200), .ZN(n2761) );
  NAND2_X1 U3172 ( .A1(n2757), .A2(n3813), .ZN(n2526) );
  NAND2_X1 U3173 ( .A1(n2527), .A2(n2526), .ZN(n4220) );
  INV_X1 U3174 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4221) );
  NAND2_X1 U3175 ( .A1(n2766), .A2(REG0_REG_24__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U3176 ( .A1(n3873), .A2(REG1_REG_24__SCAN_IN), .ZN(n2528) );
  OAI211_X1 U3177 ( .C1(n4221), .C2(n3876), .A(n2529), .B(n2528), .ZN(n2530)
         );
  INV_X1 U3178 ( .A(n2530), .ZN(n2531) );
  NOR2_X1 U3179 ( .A1(n2746), .A2(REG3_REG_22__SCAN_IN), .ZN(n2533) );
  OR2_X1 U3180 ( .A1(n2755), .A2(n2533), .ZN(n4262) );
  AOI22_X1 U3181 ( .A1(n2766), .A2(REG0_REG_22__SCAN_IN), .B1(n2826), .B2(
        REG1_REG_22__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U3182 ( .A1(n2827), .A2(REG2_REG_22__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U3183 ( .A1(n2550), .A2(REG0_REG_1__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U3184 ( .A1(n2747), .A2(REG3_REG_1__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U3185 ( .A1(n2549), .A2(REG1_REG_1__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U3186 ( .A1(n2547), .A2(n3174), .ZN(n3953) );
  NAND2_X1 U3187 ( .A1(n3953), .A2(n3957), .ZN(n2783) );
  NAND2_X1 U3188 ( .A1(n2226), .A2(REG2_REG_0__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U3189 ( .A1(n2747), .A2(REG3_REG_0__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U3190 ( .A1(n2549), .A2(REG1_REG_0__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U3191 ( .A1(n2550), .A2(REG0_REG_0__SCAN_IN), .ZN(n2542) );
  MUX2_X1 U3192 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2546), .Z(n3071) );
  NAND2_X1 U3193 ( .A1(n2783), .A2(n3170), .ZN(n3172) );
  NAND2_X1 U3194 ( .A1(n2547), .A2(n3177), .ZN(n2548) );
  NAND2_X1 U3195 ( .A1(n3172), .A2(n2548), .ZN(n3215) );
  INV_X1 U3196 ( .A(n3215), .ZN(n2558) );
  NAND2_X1 U3197 ( .A1(n2750), .A2(REG2_REG_2__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U3198 ( .A1(n2747), .A2(REG3_REG_2__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U3199 ( .A1(n2549), .A2(REG1_REG_2__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U3200 ( .A1(n2550), .A2(REG0_REG_2__SCAN_IN), .ZN(n2551) );
  AND4_X2 U3201 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(n3180)
         );
  INV_X1 U3202 ( .A(n3222), .ZN(n3080) );
  NAND2_X1 U3203 ( .A1(n4056), .A2(n3080), .ZN(n3961) );
  NAND2_X1 U3204 ( .A1(n2558), .A2(n2785), .ZN(n3214) );
  NAND2_X1 U3205 ( .A1(n3180), .A2(n3080), .ZN(n2559) );
  NAND2_X1 U3206 ( .A1(n3214), .A2(n2559), .ZN(n3161) );
  NAND2_X1 U3207 ( .A1(n2750), .A2(REG2_REG_3__SCAN_IN), .ZN(n2564) );
  INV_X1 U3208 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U3209 ( .A1(n2747), .A2(n2560), .ZN(n2563) );
  NAND2_X1 U32100 ( .A1(n2826), .A2(REG1_REG_3__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32110 ( .A1(n2766), .A2(REG0_REG_3__SCAN_IN), .ZN(n2561) );
  NAND4_X1 U32120 ( .A1(n2564), .A2(n2563), .A3(n2562), .A4(n2561), .ZN(n4055)
         );
  NAND2_X1 U32130 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  NAND2_X1 U32140 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  XNOR2_X1 U32150 ( .A(n2576), .B(IR_REG_3__SCAN_IN), .ZN(n4478) );
  MUX2_X1 U32160 ( .A(n4478), .B(DATAI_3_), .S(n2546), .Z(n3261) );
  NOR2_X1 U32170 ( .A1(n2228), .A2(n3261), .ZN(n2569) );
  NAND2_X1 U32180 ( .A1(n2228), .A2(n3261), .ZN(n2568) );
  NAND2_X1 U32190 ( .A1(n2750), .A2(REG2_REG_4__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U32200 ( .A1(n2766), .A2(REG0_REG_4__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32210 ( .A1(n2826), .A2(REG1_REG_4__SCAN_IN), .ZN(n2572) );
  INV_X1 U32220 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2570) );
  XNOR2_X1 U32230 ( .A(n2570), .B(REG3_REG_3__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U32240 ( .A1(n2747), .A2(n3212), .ZN(n2571) );
  NAND2_X1 U32250 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  NAND2_X1 U32260 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U32270 ( .A(n2578), .B(IR_REG_4__SCAN_IN), .ZN(n4477) );
  MUX2_X1 U32280 ( .A(n4477), .B(DATAI_4_), .S(n2546), .Z(n3193) );
  NAND2_X1 U32290 ( .A1(n3254), .A2(n3193), .ZN(n3964) );
  INV_X1 U32300 ( .A(n3254), .ZN(n4054) );
  NAND2_X1 U32310 ( .A1(n4054), .A2(n3206), .ZN(n3967) );
  NAND2_X1 U32320 ( .A1(n3964), .A2(n3967), .ZN(n3938) );
  NAND2_X1 U32330 ( .A1(n3191), .A2(n3938), .ZN(n2580) );
  NAND2_X1 U32340 ( .A1(n4054), .A2(n3193), .ZN(n2579) );
  NAND2_X1 U32350 ( .A1(n2580), .A2(n2579), .ZN(n3232) );
  NAND2_X1 U32360 ( .A1(n2750), .A2(REG2_REG_5__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32370 ( .A1(n2766), .A2(REG0_REG_5__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32380 ( .A1(n2826), .A2(REG1_REG_5__SCAN_IN), .ZN(n2583) );
  AOI21_X1 U32390 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2581) );
  NOR2_X1 U32400 ( .A1(n2581), .A2(n2591), .ZN(n3248) );
  NAND2_X1 U32410 ( .A1(n2747), .A2(n3248), .ZN(n2582) );
  NAND4_X1 U32420 ( .A1(n2585), .A2(n2584), .A3(n2583), .A4(n2582), .ZN(n4053)
         );
  NAND2_X1 U32430 ( .A1(n2587), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  MUX2_X1 U32440 ( .A(IR_REG_31__SCAN_IN), .B(n2586), .S(IR_REG_5__SCAN_IN), 
        .Z(n2589) );
  INV_X1 U32450 ( .A(n2608), .ZN(n2588) );
  MUX2_X1 U32460 ( .A(n3038), .B(DATAI_5_), .S(n2546), .Z(n3250) );
  AND2_X1 U32470 ( .A1(n4053), .A2(n3250), .ZN(n2590) );
  NAND2_X1 U32480 ( .A1(n2750), .A2(REG2_REG_6__SCAN_IN), .ZN(n2597) );
  INV_X1 U32490 ( .A(n2591), .ZN(n2592) );
  INV_X1 U32500 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U32510 ( .A1(n2592), .A2(n3029), .ZN(n2593) );
  AND2_X1 U32520 ( .A1(n2593), .A2(n2601), .ZN(n4635) );
  NAND2_X1 U32530 ( .A1(n2747), .A2(n4635), .ZN(n2596) );
  NAND2_X1 U32540 ( .A1(n2826), .A2(REG1_REG_6__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U32550 ( .A1(n2766), .A2(REG0_REG_6__SCAN_IN), .ZN(n2594) );
  NAND4_X1 U32560 ( .A1(n2597), .A2(n2596), .A3(n2595), .A4(n2594), .ZN(n4052)
         );
  OR2_X1 U32570 ( .A1(n2608), .A2(n3000), .ZN(n2598) );
  XNOR2_X1 U32580 ( .A(n2598), .B(IR_REG_6__SCAN_IN), .ZN(n4476) );
  MUX2_X1 U32590 ( .A(n4476), .B(DATAI_6_), .S(n2546), .Z(n3300) );
  NAND2_X1 U32600 ( .A1(n4052), .A2(n3300), .ZN(n2599) );
  NAND2_X1 U32610 ( .A1(n2750), .A2(REG2_REG_7__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U32620 ( .A1(n2766), .A2(REG0_REG_7__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U32630 ( .A1(n2826), .A2(REG1_REG_7__SCAN_IN), .ZN(n2604) );
  AND2_X1 U32640 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  NOR2_X1 U32650 ( .A1(n2611), .A2(n2602), .ZN(n3275) );
  NAND2_X1 U32660 ( .A1(n2747), .A2(n3275), .ZN(n2603) );
  NAND2_X1 U32670 ( .A1(n2608), .A2(n2607), .ZN(n2628) );
  NAND2_X1 U32680 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2618) );
  XNOR2_X1 U32690 ( .A(n2618), .B(IR_REG_7__SCAN_IN), .ZN(n4475) );
  MUX2_X1 U32700 ( .A(n4475), .B(DATAI_7_), .S(n2546), .Z(n3271) );
  NAND2_X1 U32710 ( .A1(n3368), .A2(n3271), .ZN(n2791) );
  INV_X1 U32720 ( .A(n3271), .ZN(n3333) );
  NAND2_X1 U32730 ( .A1(n3292), .A2(n3333), .ZN(n3973) );
  NAND2_X1 U32740 ( .A1(n2791), .A2(n3973), .ZN(n3924) );
  NAND2_X1 U32750 ( .A1(n3274), .A2(n3924), .ZN(n2610) );
  NAND2_X1 U32760 ( .A1(n3292), .A2(n3271), .ZN(n2609) );
  NAND2_X1 U32770 ( .A1(n2750), .A2(REG2_REG_8__SCAN_IN), .ZN(n2616) );
  NOR2_X1 U32780 ( .A1(n2611), .A2(REG3_REG_8__SCAN_IN), .ZN(n2612) );
  OR2_X1 U32790 ( .A1(n2630), .A2(n2612), .ZN(n3362) );
  INV_X1 U32800 ( .A(n3362), .ZN(n4627) );
  NAND2_X1 U32810 ( .A1(n2747), .A2(n4627), .ZN(n2615) );
  NAND2_X1 U32820 ( .A1(n2826), .A2(REG1_REG_8__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U32830 ( .A1(n2766), .A2(REG0_REG_8__SCAN_IN), .ZN(n2613) );
  NAND4_X1 U32840 ( .A1(n2616), .A2(n2615), .A3(n2614), .A4(n2613), .ZN(n3343)
         );
  INV_X1 U32850 ( .A(IR_REG_7__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U32860 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  NAND2_X1 U32870 ( .A1(n2619), .A2(IR_REG_31__SCAN_IN), .ZN(n2620) );
  XNOR2_X1 U32880 ( .A(n2620), .B(IR_REG_8__SCAN_IN), .ZN(n4514) );
  MUX2_X1 U32890 ( .A(n4514), .B(DATAI_8_), .S(n2546), .Z(n2949) );
  AND2_X1 U32900 ( .A1(n3343), .A2(n2949), .ZN(n2622) );
  INV_X1 U32910 ( .A(n3343), .ZN(n3382) );
  NAND2_X1 U32920 ( .A1(n3382), .A2(n3367), .ZN(n2621) );
  NAND2_X1 U32930 ( .A1(n2750), .A2(REG2_REG_9__SCAN_IN), .ZN(n2627) );
  XNOR2_X1 U32940 ( .A(n2630), .B(REG3_REG_9__SCAN_IN), .ZN(n3389) );
  INV_X1 U32950 ( .A(n3389), .ZN(n2623) );
  NAND2_X1 U32960 ( .A1(n2747), .A2(n2623), .ZN(n2626) );
  NAND2_X1 U32970 ( .A1(n2826), .A2(REG1_REG_9__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U32980 ( .A1(n2766), .A2(REG0_REG_9__SCAN_IN), .ZN(n2624) );
  NAND4_X1 U32990 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n4051)
         );
  NAND2_X1 U33000 ( .A1(n2638), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  MUX2_X1 U33010 ( .A(n4098), .B(DATAI_9_), .S(n2546), .Z(n3342) );
  NAND2_X1 U33020 ( .A1(n2750), .A2(REG2_REG_10__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U33030 ( .A1(n2766), .A2(REG0_REG_10__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U33040 ( .A1(n2826), .A2(REG1_REG_10__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U33050 ( .A1(n2630), .A2(REG3_REG_9__SCAN_IN), .ZN(n2632) );
  INV_X1 U33060 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U33070 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  AND2_X1 U33080 ( .A1(n2633), .A2(n2640), .ZN(n4620) );
  NAND2_X1 U33090 ( .A1(n2747), .A2(n4620), .ZN(n2634) );
  NAND4_X1 U33100 ( .A1(n2637), .A2(n2636), .A3(n2635), .A4(n2634), .ZN(n4050)
         );
  OR2_X1 U33110 ( .A1(n2647), .A2(n3000), .ZN(n2639) );
  MUX2_X1 U33120 ( .A(n4535), .B(DATAI_10_), .S(n2546), .Z(n2901) );
  INV_X1 U33130 ( .A(n4050), .ZN(n3476) );
  INV_X1 U33140 ( .A(n2901), .ZN(n3437) );
  NAND2_X1 U33150 ( .A1(n2827), .A2(REG2_REG_11__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U33160 ( .A1(n2766), .A2(REG0_REG_11__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U33170 ( .A1(n2826), .A2(REG1_REG_11__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U33180 ( .A1(n2640), .A2(n4879), .ZN(n2641) );
  AND2_X1 U33190 ( .A1(n2652), .A2(n2641), .ZN(n3461) );
  NAND2_X1 U33200 ( .A1(n2747), .A2(n3461), .ZN(n2642) );
  INV_X1 U33210 ( .A(IR_REG_10__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U33220 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U33230 ( .A1(n2648), .A2(IR_REG_31__SCAN_IN), .ZN(n2659) );
  MUX2_X1 U33240 ( .A(n4097), .B(DATAI_11_), .S(n2546), .Z(n3469) );
  NAND2_X1 U33250 ( .A1(n3562), .A2(n3469), .ZN(n3400) );
  INV_X1 U33260 ( .A(n3562), .ZN(n3440) );
  INV_X1 U33270 ( .A(n3469), .ZN(n3474) );
  NAND2_X1 U33280 ( .A1(n3440), .A2(n3474), .ZN(n3402) );
  NAND2_X1 U33290 ( .A1(n3400), .A2(n3402), .ZN(n3925) );
  NAND2_X1 U33300 ( .A1(n3390), .A2(n3925), .ZN(n2650) );
  NAND2_X1 U33310 ( .A1(n3562), .A2(n3474), .ZN(n2649) );
  NAND2_X1 U33320 ( .A1(n2650), .A2(n2649), .ZN(n3405) );
  NAND2_X1 U33330 ( .A1(n2827), .A2(REG2_REG_12__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U33340 ( .A1(n2766), .A2(REG0_REG_12__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U33350 ( .A1(n2826), .A2(REG1_REG_12__SCAN_IN), .ZN(n2655) );
  AND2_X1 U33360 ( .A1(n2652), .A2(n2651), .ZN(n2653) );
  NOR2_X1 U33370 ( .A1(n2663), .A2(n2653), .ZN(n3550) );
  NAND2_X1 U33380 ( .A1(n2747), .A2(n3550), .ZN(n2654) );
  NAND4_X1 U33390 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n3515)
         );
  INV_X1 U33400 ( .A(IR_REG_11__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U33410 ( .A1(n2659), .A2(n2658), .ZN(n2660) );
  NAND2_X1 U33420 ( .A1(n2660), .A2(IR_REG_31__SCAN_IN), .ZN(n2661) );
  MUX2_X1 U33430 ( .A(n4556), .B(DATAI_12_), .S(n2546), .Z(n3516) );
  NOR2_X1 U33440 ( .A1(n3515), .A2(n3516), .ZN(n2662) );
  INV_X1 U33450 ( .A(n3516), .ZN(n3561) );
  NAND2_X1 U33460 ( .A1(n2827), .A2(REG2_REG_13__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U33470 ( .A1(n2766), .A2(REG0_REG_13__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U33480 ( .A1(n2826), .A2(REG1_REG_13__SCAN_IN), .ZN(n2666) );
  OR2_X1 U33490 ( .A1(n2663), .A2(REG3_REG_13__SCAN_IN), .ZN(n2664) );
  AND2_X1 U33500 ( .A1(n2680), .A2(n2664), .ZN(n3511) );
  NAND2_X1 U33510 ( .A1(n2747), .A2(n3511), .ZN(n2665) );
  NAND4_X1 U33520 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n3416)
         );
  OR2_X1 U3353 ( .A1(n2675), .A2(n3000), .ZN(n2669) );
  XNOR2_X1 U33540 ( .A(n2669), .B(IR_REG_13__SCAN_IN), .ZN(n4111) );
  MUX2_X1 U3355 ( .A(n4111), .B(DATAI_13_), .S(n2546), .Z(n3415) );
  NAND2_X1 U3356 ( .A1(n2827), .A2(REG2_REG_14__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3357 ( .A1(n2766), .A2(REG0_REG_14__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3358 ( .A1(n2826), .A2(REG1_REG_14__SCAN_IN), .ZN(n2671) );
  XNOR2_X1 U3359 ( .A(n2680), .B(REG3_REG_14__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U3360 ( .A1(n2747), .A2(n3456), .ZN(n2670) );
  NAND2_X1 U3361 ( .A1(n2706), .A2(IR_REG_31__SCAN_IN), .ZN(n2676) );
  XNOR2_X1 U3362 ( .A(n2676), .B(IR_REG_14__SCAN_IN), .ZN(n4096) );
  MUX2_X1 U3363 ( .A(n4096), .B(DATAI_14_), .S(n2546), .Z(n3613) );
  NAND2_X1 U3364 ( .A1(n3864), .A2(n3613), .ZN(n3878) );
  INV_X1 U3365 ( .A(n3864), .ZN(n4049) );
  INV_X1 U3366 ( .A(n3613), .ZN(n3629) );
  NAND2_X1 U3367 ( .A1(n4049), .A2(n3629), .ZN(n3879) );
  NAND2_X1 U3368 ( .A1(n3878), .A2(n3879), .ZN(n3932) );
  NAND2_X1 U3369 ( .A1(n3864), .A2(n3629), .ZN(n2677) );
  INV_X1 U3370 ( .A(n3499), .ZN(n2686) );
  NAND2_X1 U3371 ( .A1(n2827), .A2(REG2_REG_15__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U3372 ( .A1(n2766), .A2(REG0_REG_15__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3373 ( .A1(n2826), .A2(REG1_REG_15__SCAN_IN), .ZN(n2683) );
  OAI21_X1 U3374 ( .B1(n2680), .B2(n2679), .A(n2678), .ZN(n2681) );
  AND2_X1 U3375 ( .A1(n2681), .A2(n2689), .ZN(n3860) );
  NAND2_X1 U3376 ( .A1(n2747), .A2(n3860), .ZN(n2682) );
  NAND4_X1 U3377 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n4486)
         );
  OAI21_X1 U3378 ( .B1(n2706), .B2(IR_REG_14__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2696) );
  XNOR2_X1 U3379 ( .A(n2696), .B(IR_REG_15__SCAN_IN), .ZN(n4115) );
  MUX2_X1 U3380 ( .A(n4115), .B(DATAI_15_), .S(n2546), .Z(n3648) );
  NAND2_X1 U3381 ( .A1(n4486), .A2(n3648), .ZN(n2687) );
  NAND2_X1 U3382 ( .A1(n2827), .A2(REG2_REG_16__SCAN_IN), .ZN(n2695) );
  AND2_X1 U3383 ( .A1(n2689), .A2(n4483), .ZN(n2690) );
  OR2_X1 U3384 ( .A1(n2690), .A2(n2700), .ZN(n4502) );
  INV_X1 U3385 ( .A(n4502), .ZN(n2691) );
  NAND2_X1 U3386 ( .A1(n2747), .A2(n2691), .ZN(n2694) );
  NAND2_X1 U3387 ( .A1(n3873), .A2(REG1_REG_16__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3388 ( .A1(n2766), .A2(REG0_REG_16__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3389 ( .A1(n2696), .A2(n2707), .ZN(n2697) );
  NAND2_X1 U3390 ( .A1(n2697), .A2(IR_REG_31__SCAN_IN), .ZN(n2698) );
  XNOR2_X1 U3391 ( .A(n2698), .B(IR_REG_16__SCAN_IN), .ZN(n4116) );
  MUX2_X1 U3392 ( .A(n4116), .B(DATAI_16_), .S(n2546), .Z(n3653) );
  NAND2_X1 U3393 ( .A1(n4407), .A2(n3653), .ZN(n4002) );
  NAND2_X1 U3394 ( .A1(n4048), .A2(n4490), .ZN(n3883) );
  NAND2_X1 U3395 ( .A1(n4002), .A2(n3883), .ZN(n3942) );
  NAND2_X1 U3396 ( .A1(n4048), .A2(n3653), .ZN(n2699) );
  NAND2_X1 U3397 ( .A1(n2827), .A2(REG2_REG_17__SCAN_IN), .ZN(n2705) );
  NOR2_X1 U3398 ( .A1(n2700), .A2(REG3_REG_17__SCAN_IN), .ZN(n2701) );
  OR2_X1 U3399 ( .A1(n2715), .A2(n2701), .ZN(n3808) );
  INV_X1 U3400 ( .A(n3808), .ZN(n3580) );
  NAND2_X1 U3401 ( .A1(n2747), .A2(n3580), .ZN(n2704) );
  NAND2_X1 U3402 ( .A1(n3873), .A2(REG1_REG_17__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U3403 ( .A1(n2766), .A2(REG0_REG_17__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U3404 ( .A1(n2721), .A2(IR_REG_31__SCAN_IN), .ZN(n2710) );
  XNOR2_X1 U3405 ( .A(n2710), .B(IR_REG_17__SCAN_IN), .ZN(n4119) );
  INV_X1 U3406 ( .A(DATAI_17_), .ZN(n2711) );
  MUX2_X1 U3407 ( .A(n4646), .B(n2711), .S(n2546), .Z(n4404) );
  NAND2_X1 U3408 ( .A1(n3845), .A2(n4404), .ZN(n2712) );
  INV_X1 U3409 ( .A(n4404), .ZN(n2809) );
  NAND2_X1 U3410 ( .A1(n4484), .A2(n2809), .ZN(n2713) );
  NAND2_X1 U3411 ( .A1(n2714), .A2(n2713), .ZN(n3596) );
  INV_X1 U3412 ( .A(n3596), .ZN(n2725) );
  NAND2_X1 U3413 ( .A1(n2827), .A2(REG2_REG_18__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3414 ( .A1(n2766), .A2(REG0_REG_18__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3415 ( .A1(n3873), .A2(REG1_REG_18__SCAN_IN), .ZN(n2718) );
  OR2_X1 U3416 ( .A1(n2715), .A2(REG3_REG_18__SCAN_IN), .ZN(n2716) );
  AND2_X1 U3417 ( .A1(n2736), .A2(n2716), .ZN(n3608) );
  NAND2_X1 U3418 ( .A1(n2747), .A2(n3608), .ZN(n2717) );
  NAND2_X1 U3419 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2723) );
  XNOR2_X1 U3420 ( .A(n2723), .B(IR_REG_18__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U3421 ( .A(n4474), .B(DATAI_18_), .S(n2546), .Z(n3668) );
  NAND2_X1 U3422 ( .A1(n4332), .A2(n3668), .ZN(n4318) );
  INV_X1 U3423 ( .A(n4332), .ZN(n4047) );
  INV_X1 U3424 ( .A(n3668), .ZN(n3844) );
  NAND2_X1 U3425 ( .A1(n4047), .A2(n3844), .ZN(n4319) );
  NAND2_X1 U3426 ( .A1(n2725), .A2(n2724), .ZN(n3597) );
  NAND2_X1 U3427 ( .A1(n4332), .A2(n3844), .ZN(n2726) );
  NAND2_X1 U3428 ( .A1(n2827), .A2(REG2_REG_19__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3429 ( .A1(n2766), .A2(REG0_REG_19__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U3430 ( .A1(n3873), .A2(REG1_REG_19__SCAN_IN), .ZN(n2728) );
  XNOR2_X1 U3431 ( .A(n2736), .B(REG3_REG_19__SCAN_IN), .ZN(n4337) );
  NAND2_X1 U3432 ( .A1(n2747), .A2(n4337), .ZN(n2727) );
  OR2_X1 U3433 ( .A1(n2733), .A2(n2732), .ZN(n2734) );
  MUX2_X1 U3434 ( .A(n4473), .B(DATAI_19_), .S(n2546), .Z(n4326) );
  NOR2_X1 U3435 ( .A1(n4312), .A2(n4326), .ZN(n4300) );
  NAND2_X1 U3436 ( .A1(n2827), .A2(REG2_REG_20__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U3437 ( .A1(n2766), .A2(REG0_REG_20__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U3438 ( .A1(n3873), .A2(REG1_REG_20__SCAN_IN), .ZN(n2739) );
  INV_X1 U3439 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2735) );
  INV_X1 U3440 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3824) );
  OAI21_X1 U3441 ( .B1(n2736), .B2(n2735), .A(n3824), .ZN(n2737) );
  AND2_X1 U3442 ( .A1(n2737), .A2(n2744), .ZN(n4305) );
  NAND2_X1 U3443 ( .A1(n2747), .A2(n4305), .ZN(n2738) );
  NAND4_X1 U3444 ( .A1(n2741), .A2(n2740), .A3(n2739), .A4(n2738), .ZN(n4329)
         );
  NAND2_X1 U3445 ( .A1(n4329), .A2(n3686), .ZN(n3908) );
  NAND2_X1 U3446 ( .A1(n4312), .A2(n4326), .ZN(n4301) );
  OAI21_X1 U3447 ( .B1(n4317), .B2(n4300), .A(n2742), .ZN(n2743) );
  NAND2_X1 U3448 ( .A1(n4385), .A2(n4391), .ZN(n3909) );
  NAND2_X1 U3449 ( .A1(n2743), .A2(n3909), .ZN(n4276) );
  AND2_X1 U3450 ( .A1(n2744), .A2(n4983), .ZN(n2745) );
  NOR2_X1 U3451 ( .A1(n2746), .A2(n2745), .ZN(n4284) );
  NAND2_X1 U3452 ( .A1(n4284), .A2(n2747), .ZN(n2753) );
  NAND2_X1 U3453 ( .A1(n2766), .A2(REG0_REG_21__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U3454 ( .A1(n3873), .A2(REG1_REG_21__SCAN_IN), .ZN(n2748) );
  AND2_X1 U3455 ( .A1(n2749), .A2(n2748), .ZN(n2752) );
  NAND2_X1 U3456 ( .A1(n2827), .A2(REG2_REG_21__SCAN_IN), .ZN(n2751) );
  INV_X1 U3457 ( .A(n4297), .ZN(n4046) );
  NAND2_X1 U34580 ( .A1(n4046), .A2(n3691), .ZN(n2754) );
  OR2_X1 U34590 ( .A1(n4280), .A2(n4270), .ZN(n4235) );
  NAND2_X1 U3460 ( .A1(n4280), .A2(n4270), .ZN(n2817) );
  NAND2_X1 U3461 ( .A1(n4235), .A2(n2817), .ZN(n4265) );
  INV_X1 U3462 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4250) );
  OR2_X1 U3463 ( .A1(n2755), .A2(REG3_REG_23__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U3464 ( .A1(n2757), .A2(n2756), .ZN(n4249) );
  OR2_X1 U3465 ( .A1(n4249), .A2(n2832), .ZN(n2759) );
  AOI22_X1 U3466 ( .A1(n2766), .A2(REG0_REG_23__SCAN_IN), .B1(n2826), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n2758) );
  INV_X1 U34670 ( .A(n4267), .ZN(n4369) );
  AOI21_X1 U3468 ( .B1(n2822), .B2(n4045), .A(n4208), .ZN(n2760) );
  OAI21_X1 U34690 ( .B1(n4162), .B2(n4180), .A(n4157), .ZN(n2763) );
  NAND2_X1 U3470 ( .A1(n2764), .A2(n4780), .ZN(n2765) );
  NAND2_X1 U34710 ( .A1(n3752), .A2(n2747), .ZN(n2772) );
  INV_X1 U3472 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U34730 ( .A1(n2766), .A2(REG0_REG_28__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U3474 ( .A1(n3873), .A2(REG1_REG_28__SCAN_IN), .ZN(n2767) );
  OAI211_X1 U34750 ( .C1(n2769), .C2(n3876), .A(n2768), .B(n2767), .ZN(n2770)
         );
  INV_X1 U3476 ( .A(n2770), .ZN(n2771) );
  NOR2_X1 U34770 ( .A1(n4160), .A2(n3740), .ZN(n3895) );
  XNOR2_X1 U3478 ( .A(n2875), .B(n3948), .ZN(n3641) );
  NAND2_X1 U34790 ( .A1(n2250), .A2(IR_REG_31__SCAN_IN), .ZN(n2776) );
  MUX2_X1 U3480 ( .A(IR_REG_31__SCAN_IN), .B(n2776), .S(IR_REG_21__SCAN_IN), 
        .Z(n2778) );
  NAND2_X1 U34810 ( .A1(n2778), .A2(n2777), .ZN(n3949) );
  NAND2_X1 U3482 ( .A1(n2777), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  MUX2_X1 U34830 ( .A(IR_REG_31__SCAN_IN), .B(n2779), .S(IR_REG_22__SCAN_IN), 
        .Z(n2781) );
  XNOR2_X1 U3484 ( .A(n3146), .B(n4471), .ZN(n2782) );
  NAND2_X1 U34850 ( .A1(n2782), .A2(n4133), .ZN(n3245) );
  NAND2_X1 U3486 ( .A1(n4026), .A2(n4473), .ZN(n3138) );
  INV_X1 U34870 ( .A(n4681), .ZN(n4402) );
  INV_X1 U3488 ( .A(n4058), .ZN(n3059) );
  NAND2_X1 U34890 ( .A1(n3059), .A2(n3071), .ZN(n3952) );
  OR2_X1 U3490 ( .A1(n2783), .A2(n3952), .ZN(n2784) );
  NAND2_X1 U34910 ( .A1(n2784), .A2(n3957), .ZN(n3221) );
  NAND2_X1 U3492 ( .A1(n3221), .A2(n3220), .ZN(n2786) );
  NAND2_X1 U34930 ( .A1(n2786), .A2(n3958), .ZN(n3163) );
  INV_X1 U3494 ( .A(n4055), .ZN(n3195) );
  NAND2_X1 U34950 ( .A1(n3195), .A2(n3261), .ZN(n3963) );
  INV_X1 U3496 ( .A(n3261), .ZN(n3162) );
  NAND2_X1 U34970 ( .A1(n2228), .A2(n3162), .ZN(n3960) );
  AND2_X1 U3498 ( .A1(n3963), .A2(n3960), .ZN(n3160) );
  NAND2_X1 U34990 ( .A1(n3163), .A2(n3160), .ZN(n2787) );
  NAND2_X1 U3500 ( .A1(n2787), .A2(n3963), .ZN(n3192) );
  INV_X1 U35010 ( .A(n3964), .ZN(n2788) );
  OR2_X1 U3502 ( .A1(n3192), .A2(n2788), .ZN(n2789) );
  NAND2_X1 U35030 ( .A1(n2789), .A2(n3967), .ZN(n3235) );
  AND2_X1 U3504 ( .A1(n4053), .A2(n3283), .ZN(n3233) );
  INV_X1 U35050 ( .A(n4053), .ZN(n3313) );
  NAND2_X1 U35060 ( .A1(n3313), .A2(n3250), .ZN(n3981) );
  OAI21_X1 U35070 ( .B1(n3235), .B2(n3233), .A(n3981), .ZN(n3290) );
  INV_X1 U35080 ( .A(n3300), .ZN(n3310) );
  NAND2_X1 U35090 ( .A1(n4052), .A2(n3310), .ZN(n3979) );
  NAND2_X1 U35100 ( .A1(n3290), .A2(n3979), .ZN(n2790) );
  NAND2_X1 U35110 ( .A1(n3332), .A2(n3300), .ZN(n3969) );
  NAND2_X1 U35120 ( .A1(n2790), .A2(n3969), .ZN(n3269) );
  INV_X1 U35130 ( .A(n2791), .ZN(n2792) );
  OR2_X1 U35140 ( .A1(n3269), .A2(n2792), .ZN(n2793) );
  NAND2_X1 U35150 ( .A1(n2793), .A2(n3973), .ZN(n3366) );
  NAND2_X1 U35160 ( .A1(n3382), .A2(n2949), .ZN(n3975) );
  NAND2_X1 U35170 ( .A1(n3366), .A2(n3975), .ZN(n2794) );
  NAND2_X1 U35180 ( .A1(n3343), .A2(n3367), .ZN(n3972) );
  NAND2_X1 U35190 ( .A1(n2794), .A2(n3972), .ZN(n3320) );
  AND2_X1 U35200 ( .A1(n4051), .A2(n3383), .ZN(n3989) );
  OR2_X1 U35210 ( .A1(n3320), .A2(n3989), .ZN(n2795) );
  NAND2_X1 U35220 ( .A1(n3438), .A2(n3342), .ZN(n3974) );
  NAND2_X1 U35230 ( .A1(n2795), .A2(n3974), .ZN(n3436) );
  NAND2_X1 U35240 ( .A1(n4050), .A2(n3437), .ZN(n3992) );
  NAND2_X1 U35250 ( .A1(n3436), .A2(n3992), .ZN(n2796) );
  NAND2_X1 U35260 ( .A1(n3476), .A2(n2901), .ZN(n3990) );
  NAND2_X1 U35270 ( .A1(n2796), .A2(n3990), .ZN(n3403) );
  NAND2_X1 U35280 ( .A1(n3515), .A2(n3561), .ZN(n3417) );
  NAND2_X1 U35290 ( .A1(n3416), .A2(n3529), .ZN(n2797) );
  NAND2_X1 U35300 ( .A1(n3417), .A2(n2797), .ZN(n2799) );
  INV_X1 U35310 ( .A(n3402), .ZN(n2798) );
  NOR2_X1 U35320 ( .A1(n2799), .A2(n2798), .ZN(n3993) );
  NAND2_X1 U35330 ( .A1(n3403), .A2(n3993), .ZN(n2803) );
  NAND2_X1 U35340 ( .A1(n3531), .A2(n3516), .ZN(n3419) );
  NAND2_X1 U35350 ( .A1(n3400), .A2(n3419), .ZN(n2802) );
  INV_X1 U35360 ( .A(n2799), .ZN(n2801) );
  NOR2_X1 U35370 ( .A1(n3416), .A2(n3529), .ZN(n2800) );
  AOI21_X1 U35380 ( .B1(n2802), .B2(n2801), .A(n2800), .ZN(n3995) );
  NAND2_X1 U35390 ( .A1(n2803), .A2(n3995), .ZN(n3882) );
  NAND2_X1 U35400 ( .A1(n3882), .A2(n2391), .ZN(n3500) );
  INV_X1 U35410 ( .A(n4486), .ZN(n3646) );
  NAND2_X1 U35420 ( .A1(n3646), .A2(n3648), .ZN(n3881) );
  INV_X1 U35430 ( .A(n3648), .ZN(n3865) );
  NAND2_X1 U35440 ( .A1(n4486), .A2(n3865), .ZN(n3880) );
  NAND2_X1 U35450 ( .A1(n3881), .A2(n3880), .ZN(n3931) );
  INV_X1 U35460 ( .A(n3878), .ZN(n2804) );
  NOR2_X1 U35470 ( .A1(n3931), .A2(n2804), .ZN(n2805) );
  NAND2_X1 U35480 ( .A1(n3500), .A2(n2805), .ZN(n2806) );
  NAND2_X1 U35490 ( .A1(n2806), .A2(n3880), .ZN(n3537) );
  INV_X1 U35500 ( .A(n3942), .ZN(n2807) );
  NAND2_X1 U35510 ( .A1(n3537), .A2(n2807), .ZN(n2808) );
  NAND2_X1 U35520 ( .A1(n2808), .A2(n3883), .ZN(n3603) );
  NAND2_X1 U35530 ( .A1(n3845), .A2(n2809), .ZN(n3604) );
  NAND2_X1 U35540 ( .A1(n4318), .A2(n3604), .ZN(n2812) );
  INV_X1 U35550 ( .A(n4326), .ZN(n4335) );
  NAND2_X1 U35560 ( .A1(n4312), .A2(n4335), .ZN(n2810) );
  AND2_X1 U35570 ( .A1(n4319), .A2(n2810), .ZN(n4229) );
  NOR2_X1 U35580 ( .A1(n4312), .A2(n4335), .ZN(n2811) );
  AOI21_X1 U35590 ( .B1(n2812), .B2(n4229), .A(n2811), .ZN(n4291) );
  NAND2_X1 U35600 ( .A1(n4385), .A2(n3686), .ZN(n2813) );
  NAND2_X1 U35610 ( .A1(n3603), .A2(n4233), .ZN(n2814) );
  NAND2_X1 U35620 ( .A1(n4484), .A2(n4404), .ZN(n3601) );
  NAND2_X1 U35630 ( .A1(n4229), .A2(n3601), .ZN(n4003) );
  AND2_X1 U35640 ( .A1(n4329), .A2(n4391), .ZN(n4232) );
  AOI21_X1 U35650 ( .B1(n4233), .B2(n4003), .A(n4232), .ZN(n3885) );
  NAND2_X1 U35660 ( .A1(n2814), .A2(n3885), .ZN(n2816) );
  NAND2_X1 U35670 ( .A1(n4297), .A2(n3691), .ZN(n3937) );
  NAND2_X1 U35680 ( .A1(n4235), .A2(n3937), .ZN(n4009) );
  INV_X1 U35690 ( .A(n4009), .ZN(n2815) );
  NAND2_X1 U35700 ( .A1(n2816), .A2(n2815), .ZN(n2821) );
  NAND2_X1 U35710 ( .A1(n4267), .A2(n4247), .ZN(n2818) );
  NAND2_X1 U35720 ( .A1(n2818), .A2(n2817), .ZN(n4012) );
  INV_X1 U35730 ( .A(n4012), .ZN(n2820) );
  NOR2_X1 U35740 ( .A1(n4297), .A2(n3691), .ZN(n4007) );
  NAND2_X1 U35750 ( .A1(n4007), .A2(n4235), .ZN(n2819) );
  AND2_X1 U35760 ( .A1(n2820), .A2(n2819), .ZN(n3889) );
  NAND2_X1 U35770 ( .A1(n2821), .A2(n3889), .ZN(n4210) );
  NAND2_X1 U35780 ( .A1(n4244), .A2(n2822), .ZN(n3906) );
  NAND2_X1 U35790 ( .A1(n4369), .A2(n4240), .ZN(n4209) );
  AND2_X1 U35800 ( .A1(n3906), .A2(n4209), .ZN(n4011) );
  AND2_X1 U35810 ( .A1(n4045), .A2(n4368), .ZN(n3877) );
  AOI21_X1 U3582 ( .B1(n4210), .B2(n4011), .A(n3877), .ZN(n4194) );
  NAND2_X1 U3583 ( .A1(n4215), .A2(n4200), .ZN(n3929) );
  NAND2_X1 U3584 ( .A1(n4194), .A2(n3929), .ZN(n4175) );
  NOR2_X1 U3585 ( .A1(n4197), .A2(n4186), .ZN(n3935) );
  NOR2_X1 U3586 ( .A1(n4215), .A2(n4200), .ZN(n4173) );
  NOR2_X1 U3587 ( .A1(n3935), .A2(n4173), .ZN(n4019) );
  NAND2_X1 U3588 ( .A1(n4197), .A2(n4186), .ZN(n3896) );
  INV_X1 U3589 ( .A(n3896), .ZN(n3936) );
  AOI21_X1 U3590 ( .B1(n4175), .B2(n4019), .A(n3936), .ZN(n4158) );
  NOR2_X1 U3591 ( .A1(n3748), .A2(n4162), .ZN(n4017) );
  AOI21_X1 U3592 ( .B1(n4158), .B2(n4159), .A(n3897), .ZN(n2878) );
  XNOR2_X1 U3593 ( .A(n2878), .B(n3948), .ZN(n2833) );
  INV_X1 U3594 ( .A(n4026), .ZN(n4472) );
  NAND2_X1 U3595 ( .A1(n4472), .A2(n3955), .ZN(n4030) );
  OR2_X1 U3596 ( .A1(n4133), .A2(n4034), .ZN(n2823) );
  NAND2_X1 U3597 ( .A1(n2824), .A2(IR_REG_31__SCAN_IN), .ZN(n2825) );
  INV_X1 U3598 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3599 ( .A1(n2766), .A2(REG0_REG_29__SCAN_IN), .ZN(n2829) );
  NAND2_X1 U3600 ( .A1(n2827), .A2(REG2_REG_29__SCAN_IN), .ZN(n2828) );
  OAI211_X1 U3601 ( .C1(n2891), .C2(n2504), .A(n2829), .B(n2828), .ZN(n2830)
         );
  INV_X1 U3602 ( .A(n2830), .ZN(n2831) );
  AOI22_X1 U3603 ( .A1(n2833), .A2(n4324), .B1(n4328), .B2(n4044), .ZN(n3637)
         );
  INV_X1 U3604 ( .A(n3012), .ZN(n2964) );
  INV_X1 U3605 ( .A(n4406), .ZN(n4241) );
  AOI22_X1 U3606 ( .A1(n4180), .A2(n4241), .B1(n3740), .B2(n4327), .ZN(n2834)
         );
  OAI211_X1 U3607 ( .C1(n3641), .C2(n4402), .A(n3637), .B(n2834), .ZN(n2870)
         );
  NOR2_X1 U3608 ( .A1(n2835), .A2(n3000), .ZN(n2836) );
  NAND2_X1 U3609 ( .A1(n2992), .A2(B_REG_SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3610 ( .A1(n2780), .A2(IR_REG_31__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3611 ( .A1(n2845), .A2(n4936), .ZN(n2838) );
  NAND2_X1 U3612 ( .A1(n2838), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  MUX2_X1 U3613 ( .A(n2840), .B(B_REG_SCAN_IN), .S(n3004), .Z(n2842) );
  INV_X1 U3614 ( .A(D_REG_1__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3615 ( .A1(n2862), .A2(n2843), .ZN(n2961) );
  INV_X1 U3616 ( .A(n3006), .ZN(n2860) );
  NAND2_X1 U3617 ( .A1(n2860), .A2(n2992), .ZN(n3009) );
  NAND2_X1 U3618 ( .A1(n2961), .A2(n3009), .ZN(n2858) );
  XNOR2_X1 U3619 ( .A(n2845), .B(n4936), .ZN(n3011) );
  NAND2_X1 U3620 ( .A1(n4026), .A2(n4133), .ZN(n2963) );
  NAND2_X1 U3621 ( .A1(n2963), .A2(n3012), .ZN(n3142) );
  OAI211_X1 U3622 ( .C1(n3955), .C2(n4664), .A(n3139), .B(n3142), .ZN(n2846)
         );
  INV_X1 U3623 ( .A(n2846), .ZN(n2857) );
  NOR4_X1 U3624 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2850) );
  NOR4_X1 U3625 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2849) );
  NOR4_X1 U3626 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2848) );
  NOR4_X1 U3627 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2847) );
  NAND4_X1 U3628 ( .A1(n2850), .A2(n2849), .A3(n2848), .A4(n2847), .ZN(n2856)
         );
  NOR2_X1 U3629 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_10__SCAN_IN), .ZN(n2854) );
  NOR4_X1 U3630 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2853) );
  NOR4_X1 U3631 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2852) );
  NOR4_X1 U3632 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2851) );
  NAND4_X1 U3633 ( .A1(n2854), .A2(n2853), .A3(n2852), .A4(n2851), .ZN(n2855)
         );
  OAI21_X1 U3634 ( .B1(n2856), .B2(n2855), .A(n2862), .ZN(n2960) );
  INV_X1 U3635 ( .A(D_REG_0__SCAN_IN), .ZN(n3008) );
  MUX2_X1 U3636 ( .A(REG1_REG_28__SCAN_IN), .B(n2870), .S(n4700), .Z(n2863) );
  INV_X1 U3637 ( .A(n2863), .ZN(n2868) );
  NAND2_X1 U3638 ( .A1(n3363), .A2(n3383), .ZN(n3432) );
  AND2_X1 U3639 ( .A1(n4164), .A2(n3740), .ZN(n2865) );
  NAND2_X1 U3640 ( .A1(n2474), .A2(n2866), .ZN(n2867) );
  NAND2_X1 U3641 ( .A1(n2868), .A2(n2867), .ZN(U3546) );
  INV_X1 U3642 ( .A(n2962), .ZN(n3143) );
  MUX2_X1 U3643 ( .A(REG0_REG_28__SCAN_IN), .B(n2870), .S(n4690), .Z(n2871) );
  INV_X1 U3644 ( .A(n2871), .ZN(n2873) );
  NAND2_X1 U3645 ( .A1(n2474), .A2(n4423), .ZN(n2872) );
  NAND2_X1 U3646 ( .A1(n2873), .A2(n2872), .ZN(U3514) );
  NAND2_X1 U3647 ( .A1(n2546), .A2(DATAI_29_), .ZN(n4147) );
  XNOR2_X1 U3648 ( .A(n4044), .B(n4147), .ZN(n3950) );
  XNOR2_X1 U3649 ( .A(n2876), .B(n3950), .ZN(n4145) );
  INV_X1 U3650 ( .A(n3898), .ZN(n2877) );
  OAI21_X1 U3651 ( .B1(n2878), .B2(n3895), .A(n2877), .ZN(n2879) );
  XNOR2_X1 U3652 ( .A(n2879), .B(n3950), .ZN(n2886) );
  INV_X1 U3653 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3654 ( .A1(n3873), .A2(REG1_REG_30__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3655 ( .A1(n2766), .A2(REG0_REG_30__SCAN_IN), .ZN(n2880) );
  OAI211_X1 U3656 ( .C1(n3876), .C2(n2882), .A(n2881), .B(n2880), .ZN(n4043)
         );
  INV_X1 U3657 ( .A(n4043), .ZN(n2885) );
  INV_X1 U3658 ( .A(B_REG_SCAN_IN), .ZN(n4967) );
  INV_X1 U3659 ( .A(IR_REG_27__SCAN_IN), .ZN(n2883) );
  XNOR2_X1 U3660 ( .A(n2884), .B(n2883), .ZN(n4509) );
  OAI21_X1 U3661 ( .B1(n4967), .B2(n4509), .A(n4328), .ZN(n4140) );
  OAI22_X1 U3662 ( .A1(n2886), .A2(n4182), .B1(n2885), .B2(n4140), .ZN(n4153)
         );
  INV_X1 U3663 ( .A(n4153), .ZN(n2889) );
  OAI22_X1 U3664 ( .A1(n4160), .A2(n4406), .B1(n4147), .B2(n4405), .ZN(n2887)
         );
  INV_X1 U3665 ( .A(n2887), .ZN(n2888) );
  NAND2_X1 U3666 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  AOI21_X1 U3667 ( .B1(n4145), .B2(n4681), .A(n2890), .ZN(n2895) );
  MUX2_X1 U3668 ( .A(n2891), .B(n2895), .S(n4700), .Z(n2894) );
  NAND2_X1 U3669 ( .A1(n2892), .A2(n4147), .ZN(n4347) );
  OAI21_X1 U3670 ( .B1(n2892), .B2(n4147), .A(n4347), .ZN(n4151) );
  NAND2_X1 U3671 ( .A1(n2894), .A2(n2893), .ZN(U3547) );
  INV_X1 U3672 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2896) );
  MUX2_X1 U3673 ( .A(n2896), .B(n2895), .S(n4690), .Z(n2898) );
  NAND2_X1 U3674 ( .A1(n2898), .A2(n2897), .ZN(U3515) );
  INV_X2 U3675 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  OR2_X2 U3676 ( .A1(n3732), .A2(n4669), .ZN(n2906) );
  AND2_X1 U3677 ( .A1(n2901), .A2(n2908), .ZN(n2900) );
  AOI21_X1 U3678 ( .B1(n4050), .B2(n3741), .A(n2900), .ZN(n3463) );
  NAND2_X1 U3679 ( .A1(n4050), .A2(n2908), .ZN(n2903) );
  NAND2_X1 U3680 ( .A1(n2901), .A2(n3739), .ZN(n2902) );
  NAND2_X1 U3681 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  NAND2_X1 U3682 ( .A1(n3146), .A2(n2973), .ZN(n2947) );
  XNOR2_X1 U3683 ( .A(n2904), .B(n2947), .ZN(n3462) );
  XOR2_X1 U3684 ( .A(n3463), .B(n3462), .Z(n2968) );
  OAI22_X1 U3685 ( .A1(n3224), .A2(n2906), .B1(n3733), .B2(n3174), .ZN(n2914)
         );
  INV_X1 U3686 ( .A(n2914), .ZN(n2917) );
  OAI22_X1 U3687 ( .A1(n3224), .A2(n3733), .B1(n3732), .B2(n3174), .ZN(n2907)
         );
  XNOR2_X1 U3688 ( .A(n2907), .B(n2947), .ZN(n2915) );
  INV_X1 U3689 ( .A(n2915), .ZN(n2916) );
  NAND2_X1 U3690 ( .A1(n4058), .A2(n2908), .ZN(n2910) );
  NAND2_X1 U3691 ( .A1(n3071), .A2(n3739), .ZN(n2909) );
  NAND2_X1 U3692 ( .A1(n2910), .A2(n2909), .ZN(n3068) );
  NAND2_X1 U3693 ( .A1(n4058), .A2(n3741), .ZN(n2912) );
  NAND2_X1 U3694 ( .A1(n3071), .A2(n2908), .ZN(n2911) );
  NAND2_X1 U3695 ( .A1(n2912), .A2(n2911), .ZN(n3067) );
  NAND2_X1 U3696 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3032) );
  NOR2_X1 U3697 ( .A1(n2899), .A2(n3032), .ZN(n2913) );
  OAI21_X1 U3698 ( .B1(n2947), .B2(n3068), .A(n3063), .ZN(n3057) );
  OAI22_X1 U3699 ( .A1(n3180), .A2(n3733), .B1(n3080), .B2(n3732), .ZN(n2918)
         );
  XNOR2_X1 U3700 ( .A(n2918), .B(n2947), .ZN(n2921) );
  OR2_X1 U3701 ( .A1(n3180), .A2(n2906), .ZN(n2920) );
  NAND2_X1 U3702 ( .A1(n3222), .A2(n2908), .ZN(n2919) );
  NAND2_X1 U3703 ( .A1(n2920), .A2(n2919), .ZN(n2922) );
  XNOR2_X1 U3704 ( .A(n2921), .B(n2922), .ZN(n3078) );
  INV_X1 U3705 ( .A(n2921), .ZN(n2924) );
  INV_X1 U3706 ( .A(n2922), .ZN(n2923) );
  NAND2_X1 U3707 ( .A1(n2228), .A2(n2908), .ZN(n2926) );
  NAND2_X1 U3708 ( .A1(n3261), .A2(n3739), .ZN(n2925) );
  NAND2_X1 U3709 ( .A1(n2926), .A2(n2925), .ZN(n2927) );
  XNOR2_X1 U3710 ( .A(n2927), .B(n3742), .ZN(n2929) );
  OAI22_X1 U3711 ( .A1(n3195), .A2(n2906), .B1(n3733), .B2(n3162), .ZN(n2928)
         );
  XNOR2_X1 U3712 ( .A(n2929), .B(n2928), .ZN(n3151) );
  OAI22_X1 U3713 ( .A1(n3152), .A2(n3151), .B1(n2929), .B2(n2928), .ZN(n3208)
         );
  OAI22_X1 U3714 ( .A1(n3254), .A2(n3733), .B1(n3732), .B2(n3206), .ZN(n2930)
         );
  XNOR2_X1 U3715 ( .A(n2930), .B(n2947), .ZN(n2932) );
  OAI22_X1 U3716 ( .A1(n3254), .A2(n2906), .B1(n3733), .B2(n3206), .ZN(n2931)
         );
  XNOR2_X1 U3717 ( .A(n2932), .B(n2931), .ZN(n3209) );
  NOR2_X1 U3718 ( .A1(n3208), .A2(n3209), .ZN(n3207) );
  AND2_X1 U3719 ( .A1(n3250), .A2(n2908), .ZN(n2934) );
  AOI21_X1 U3720 ( .B1(n4053), .B2(n3741), .A(n2934), .ZN(n2936) );
  OAI22_X1 U3721 ( .A1(n3313), .A2(n3733), .B1(n3732), .B2(n3283), .ZN(n2935)
         );
  XNOR2_X1 U3722 ( .A(n2935), .B(n3742), .ZN(n2938) );
  XOR2_X1 U3723 ( .A(n2936), .B(n2938), .Z(n3280) );
  INV_X1 U3724 ( .A(n2936), .ZN(n2937) );
  OAI22_X1 U3725 ( .A1(n3332), .A2(n2906), .B1(n3310), .B2(n3733), .ZN(n2940)
         );
  INV_X1 U3726 ( .A(n2940), .ZN(n3306) );
  OAI22_X1 U3727 ( .A1(n3332), .A2(n3733), .B1(n3310), .B2(n3732), .ZN(n2939)
         );
  XNOR2_X1 U3728 ( .A(n2939), .B(n2947), .ZN(n3307) );
  OAI22_X1 U3729 ( .A1(n3368), .A2(n2906), .B1(n3733), .B2(n3333), .ZN(n2942)
         );
  OAI22_X1 U3730 ( .A1(n3368), .A2(n3733), .B1(n3732), .B2(n3333), .ZN(n2941)
         );
  XNOR2_X1 U3731 ( .A(n2941), .B(n2947), .ZN(n2943) );
  XOR2_X1 U3732 ( .A(n2942), .B(n2943), .Z(n3330) );
  NAND2_X1 U3733 ( .A1(n3343), .A2(n2908), .ZN(n2946) );
  NAND2_X1 U3734 ( .A1(n2949), .A2(n3739), .ZN(n2945) );
  NAND2_X1 U3735 ( .A1(n2946), .A2(n2945), .ZN(n2948) );
  XNOR2_X1 U3736 ( .A(n2948), .B(n3467), .ZN(n2954) );
  INV_X1 U3737 ( .A(n2954), .ZN(n2952) );
  AND2_X1 U3738 ( .A1(n2949), .A2(n2908), .ZN(n2950) );
  AOI21_X1 U3739 ( .B1(n3343), .B2(n3741), .A(n2950), .ZN(n2953) );
  INV_X1 U3740 ( .A(n2953), .ZN(n2951) );
  NAND2_X1 U3741 ( .A1(n2952), .A2(n2951), .ZN(n3353) );
  AND2_X1 U3742 ( .A1(n2954), .A2(n2953), .ZN(n3354) );
  NAND2_X1 U3743 ( .A1(n4051), .A2(n2908), .ZN(n2956) );
  NAND2_X1 U3744 ( .A1(n3342), .A2(n3739), .ZN(n2955) );
  NAND2_X1 U3745 ( .A1(n2956), .A2(n2955), .ZN(n2957) );
  XNOR2_X1 U3746 ( .A(n2957), .B(n2947), .ZN(n2959) );
  OAI22_X1 U3747 ( .A1(n3438), .A2(n2906), .B1(n3733), .B2(n3383), .ZN(n2958)
         );
  XNOR2_X1 U3748 ( .A(n2959), .B(n2958), .ZN(n3379) );
  AND2_X1 U3749 ( .A1(n2960), .A2(n3009), .ZN(n3144) );
  NAND3_X1 U3750 ( .A1(n3144), .A2(n2962), .A3(n2961), .ZN(n2975) );
  NAND2_X1 U3751 ( .A1(n2963), .A2(n3135), .ZN(n2965) );
  NAND2_X1 U3752 ( .A1(n2965), .A2(n2964), .ZN(n2969) );
  INV_X1 U3753 ( .A(n2969), .ZN(n2966) );
  AND2_X1 U3754 ( .A1(n3139), .A2(n2966), .ZN(n2967) );
  AOI211_X1 U3755 ( .C1(n2968), .C2(n2265), .A(n3858), .B(n3466), .ZN(n2986)
         );
  NAND2_X1 U3756 ( .A1(n2969), .A2(n4405), .ZN(n2970) );
  NAND2_X1 U3757 ( .A1(n2975), .A2(n2970), .ZN(n2971) );
  NAND2_X1 U3758 ( .A1(n2971), .A2(n3142), .ZN(n3053) );
  NAND2_X1 U3759 ( .A1(n2899), .A2(n3011), .ZN(n2972) );
  OAI21_X1 U3760 ( .B1(n3053), .B2(n2972), .A(STATE_REG_SCAN_IN), .ZN(n2976)
         );
  NOR2_X1 U3761 ( .A1(n3005), .A2(n2973), .ZN(n2974) );
  NAND2_X1 U3762 ( .A1(n2975), .A2(n4033), .ZN(n3054) );
  INV_X1 U3763 ( .A(n4620), .ZN(n2977) );
  NOR2_X1 U3764 ( .A1(n4503), .A2(n2977), .ZN(n2985) );
  INV_X1 U3765 ( .A(n4482), .ZN(n3108) );
  AND2_X1 U3766 ( .A1(n4033), .A2(n3108), .ZN(n2978) );
  NAND2_X1 U3767 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4538) );
  OAI21_X1 U3768 ( .B1(n3863), .B2(n3438), .A(n4538), .ZN(n2984) );
  AND2_X1 U3769 ( .A1(n3139), .A2(n4327), .ZN(n2979) );
  NAND2_X1 U3770 ( .A1(n2982), .A2(n2979), .ZN(n2980) );
  AND2_X1 U3771 ( .A1(n4033), .A2(n4482), .ZN(n2981) );
  NAND2_X2 U3772 ( .A1(n2982), .A2(n2981), .ZN(n3867) );
  OAI22_X1 U3773 ( .A1(n4491), .A2(n3437), .B1(n3562), .B2(n3867), .ZN(n2983)
         );
  OR4_X1 U3774 ( .A1(n2986), .A2(n2985), .A3(n2984), .A4(n2983), .ZN(U3214) );
  INV_X1 U3775 ( .A(DATAI_21_), .ZN(n4916) );
  NAND2_X1 U3776 ( .A1(n3955), .A2(STATE_REG_SCAN_IN), .ZN(n2987) );
  OAI21_X1 U3777 ( .B1(STATE_REG_SCAN_IN), .B2(n4916), .A(n2987), .ZN(U3331)
         );
  INV_X1 U3778 ( .A(DATAI_5_), .ZN(n2988) );
  MUX2_X1 U3779 ( .A(n2278), .B(n2988), .S(U3149), .Z(n2989) );
  INV_X1 U3780 ( .A(n2989), .ZN(U3347) );
  INV_X1 U3781 ( .A(DATAI_24_), .ZN(n2991) );
  NAND2_X1 U3782 ( .A1(n3004), .A2(STATE_REG_SCAN_IN), .ZN(n2990) );
  OAI21_X1 U3783 ( .B1(STATE_REG_SCAN_IN), .B2(n2991), .A(n2990), .ZN(U3328)
         );
  INV_X1 U3784 ( .A(DATAI_25_), .ZN(n2995) );
  INV_X1 U3785 ( .A(n2992), .ZN(n2993) );
  NAND2_X1 U3786 ( .A1(n2993), .A2(STATE_REG_SCAN_IN), .ZN(n2994) );
  OAI21_X1 U3787 ( .B1(STATE_REG_SCAN_IN), .B2(n2995), .A(n2994), .ZN(U3327)
         );
  INV_X1 U3788 ( .A(DATAI_26_), .ZN(n2997) );
  NAND2_X1 U3789 ( .A1(n3006), .A2(STATE_REG_SCAN_IN), .ZN(n2996) );
  OAI21_X1 U3790 ( .B1(STATE_REG_SCAN_IN), .B2(n2997), .A(n2996), .ZN(U3326)
         );
  INV_X1 U3791 ( .A(DATAI_29_), .ZN(n4762) );
  NAND2_X1 U3792 ( .A1(n2998), .A2(STATE_REG_SCAN_IN), .ZN(n2999) );
  OAI21_X1 U3793 ( .B1(STATE_REG_SCAN_IN), .B2(n4762), .A(n2999), .ZN(U3323)
         );
  INV_X1 U3794 ( .A(DATAI_31_), .ZN(n3002) );
  OR4_X1 U3795 ( .A1(n2419), .A2(IR_REG_30__SCAN_IN), .A3(n3000), .A4(U3149), 
        .ZN(n3001) );
  OAI21_X1 U3796 ( .B1(STATE_REG_SCAN_IN), .B2(n3002), .A(n3001), .ZN(U3321)
         );
  NOR3_X1 U3797 ( .A1(n3006), .A2(n3005), .A3(n3004), .ZN(n3007) );
  AOI21_X1 U3798 ( .B1(n4643), .B2(n3008), .A(n3007), .ZN(U3458) );
  INV_X1 U3799 ( .A(n3009), .ZN(n3010) );
  AOI22_X1 U3800 ( .A1(n4643), .A2(n2843), .B1(n3010), .B2(n4645), .ZN(U3459)
         );
  OR2_X1 U3801 ( .A1(n3011), .A2(U3149), .ZN(n4040) );
  INV_X1 U3802 ( .A(n4040), .ZN(n4035) );
  OR2_X1 U3803 ( .A1(n3139), .A2(n4035), .ZN(n3027) );
  NAND2_X1 U3804 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  INV_X1 U3805 ( .A(n3026), .ZN(n3014) );
  NOR2_X1 U3806 ( .A1(n4612), .A2(U4043), .ZN(U3148) );
  INV_X1 U3807 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U3808 ( .A1(n3515), .A2(U4043), .ZN(n3015) );
  OAI21_X1 U3809 ( .B1(U4043), .B2(n4968), .A(n3015), .ZN(U3562) );
  INV_X1 U3810 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3017) );
  NAND2_X1 U3811 ( .A1(n3343), .A2(U4043), .ZN(n3016) );
  OAI21_X1 U3812 ( .B1(U4043), .B2(n3017), .A(n3016), .ZN(U3558) );
  INV_X1 U3813 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U3814 ( .A1(n3416), .A2(U4043), .ZN(n3018) );
  OAI21_X1 U3815 ( .B1(U4043), .B2(n4934), .A(n3018), .ZN(U3563) );
  INV_X1 U3816 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4860) );
  NAND2_X1 U3817 ( .A1(n4329), .A2(U4043), .ZN(n3019) );
  OAI21_X1 U3818 ( .B1(U4043), .B2(n4860), .A(n3019), .ZN(U3570) );
  INV_X1 U3819 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U3820 ( .A1(n3440), .A2(U4043), .ZN(n3020) );
  OAI21_X1 U3821 ( .B1(U4043), .B2(n4893), .A(n3020), .ZN(U3561) );
  INV_X1 U3822 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U3823 ( .A1(n3292), .A2(U4043), .ZN(n3021) );
  OAI21_X1 U3824 ( .B1(U4043), .B2(n4851), .A(n3021), .ZN(U3557) );
  NAND2_X1 U3825 ( .A1(n2230), .A2(REG2_REG_1__SCAN_IN), .ZN(n3112) );
  MUX2_X1 U3826 ( .A(n4944), .B(REG2_REG_2__SCAN_IN), .S(n4479), .Z(n3113) );
  XNOR2_X1 U3827 ( .A(n3022), .B(n4478), .ZN(n3045) );
  INV_X1 U3828 ( .A(n3022), .ZN(n3023) );
  AOI22_X1 U3829 ( .A1(n3045), .A2(REG2_REG_3__SCAN_IN), .B1(n4478), .B2(n3023), .ZN(n3024) );
  XNOR2_X1 U3830 ( .A(n3024), .B(n4477), .ZN(n3123) );
  INV_X1 U3831 ( .A(n3024), .ZN(n3025) );
  MUX2_X1 U3832 ( .A(n2277), .B(REG2_REG_5__SCAN_IN), .S(n3038), .Z(n3086) );
  XNOR2_X1 U3833 ( .A(n3095), .B(REG2_REG_6__SCAN_IN), .ZN(n3044) );
  NAND2_X1 U3834 ( .A1(n3027), .A2(n3026), .ZN(n4513) );
  OR2_X1 U3835 ( .A1(n4482), .A2(n4509), .ZN(n4037) );
  INV_X1 U3836 ( .A(n4513), .ZN(n3028) );
  INV_X1 U3837 ( .A(n4619), .ZN(n4059) );
  NOR2_X1 U3838 ( .A1(STATE_REG_SCAN_IN), .A2(n3029), .ZN(n3311) );
  AOI21_X1 U3839 ( .B1(n4612), .B2(ADDR_REG_6__SCAN_IN), .A(n3311), .ZN(n3030)
         );
  INV_X1 U3840 ( .A(n3030), .ZN(n3042) );
  INV_X1 U3841 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3040) );
  INV_X1 U3842 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4905) );
  MUX2_X1 U3843 ( .A(REG1_REG_2__SCAN_IN), .B(n4905), .S(n4479), .Z(n3117) );
  INV_X1 U3844 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3031) );
  XNOR2_X1 U3845 ( .A(n4480), .B(n3031), .ZN(n4066) );
  INV_X1 U3846 ( .A(n3032), .ZN(n4065) );
  NAND2_X1 U3847 ( .A1(n4066), .A2(n4065), .ZN(n4064) );
  NAND2_X1 U3848 ( .A1(n2230), .A2(REG1_REG_1__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U3849 ( .A1(n4064), .A2(n3033), .ZN(n3116) );
  NAND2_X1 U3850 ( .A1(n3117), .A2(n3116), .ZN(n3115) );
  NAND2_X1 U3851 ( .A1(n4479), .A2(REG1_REG_2__SCAN_IN), .ZN(n3034) );
  INV_X1 U3852 ( .A(n4478), .ZN(n3046) );
  NAND2_X1 U3853 ( .A1(n3049), .A2(REG1_REG_3__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U3854 ( .A1(n3035), .A2(n4478), .ZN(n3036) );
  INV_X1 U3855 ( .A(n4477), .ZN(n3130) );
  XNOR2_X1 U3856 ( .A(n3037), .B(n3130), .ZN(n3124) );
  XNOR2_X1 U3857 ( .A(n3038), .B(REG1_REG_5__SCAN_IN), .ZN(n3089) );
  INV_X1 U3858 ( .A(n4509), .ZN(n4470) );
  NOR2_X2 U3859 ( .A1(n4513), .A2(n4470), .ZN(n4613) );
  INV_X1 U3860 ( .A(n4613), .ZN(n4138) );
  AOI211_X1 U3861 ( .C1(n3040), .C2(n3039), .A(n4138), .B(n3099), .ZN(n3041)
         );
  AOI211_X1 U3862 ( .C1(n4059), .C2(n4476), .A(n3042), .B(n3041), .ZN(n3043)
         );
  OAI21_X1 U3863 ( .B1(n3044), .B2(n4606), .A(n3043), .ZN(U3246) );
  XNOR2_X1 U3864 ( .A(n3045), .B(REG2_REG_3__SCAN_IN), .ZN(n3052) );
  NOR2_X1 U3865 ( .A1(STATE_REG_SCAN_IN), .A2(n2560), .ZN(n3154) );
  NOR2_X1 U3866 ( .A1(n4619), .A2(n3046), .ZN(n3047) );
  AOI211_X1 U3867 ( .C1(n4612), .C2(ADDR_REG_3__SCAN_IN), .A(n3154), .B(n3047), 
        .ZN(n3051) );
  OAI211_X1 U3868 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3049), .A(n4613), .B(n3048), 
        .ZN(n3050) );
  OAI211_X1 U3869 ( .C1(n3052), .C2(n4606), .A(n3051), .B(n3050), .ZN(U3243)
         );
  INV_X1 U3870 ( .A(n3053), .ZN(n3055) );
  NAND3_X1 U3871 ( .A1(n3055), .A2(n3139), .A3(n3054), .ZN(n3082) );
  INV_X1 U3872 ( .A(n3082), .ZN(n3075) );
  INV_X1 U3873 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3176) );
  OAI211_X1 U3874 ( .C1(n3058), .C2(n3057), .A(n3056), .B(n4498), .ZN(n3062)
         );
  INV_X1 U3875 ( .A(n4491), .ZN(n3756) );
  OAI22_X1 U3876 ( .A1(n3059), .A2(n3863), .B1(n3867), .B2(n3180), .ZN(n3060)
         );
  AOI21_X1 U3877 ( .B1(n3177), .B2(n3756), .A(n3060), .ZN(n3061) );
  OAI211_X1 U3878 ( .C1(n3075), .C2(n3176), .A(n3062), .B(n3061), .ZN(U3219)
         );
  INV_X1 U3879 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3074) );
  INV_X1 U3880 ( .A(n3063), .ZN(n3070) );
  INV_X1 U3881 ( .A(IR_REG_0__SCAN_IN), .ZN(n3065) );
  INV_X1 U3882 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3064) );
  AOI21_X1 U3883 ( .B1(n3065), .B2(n3064), .A(n2899), .ZN(n3066) );
  NOR3_X1 U3884 ( .A1(n3068), .A2(n3067), .A3(n3066), .ZN(n3069) );
  NOR2_X1 U3885 ( .A1(n3070), .A2(n3069), .ZN(n3109) );
  NAND2_X1 U3886 ( .A1(n3109), .A2(n4498), .ZN(n3073) );
  INV_X1 U3887 ( .A(n3867), .ZN(n4485) );
  AOI22_X1 U3888 ( .A1(n3756), .A2(n3071), .B1(n4485), .B2(n2547), .ZN(n3072)
         );
  OAI211_X1 U3889 ( .C1(n3075), .C2(n3074), .A(n3073), .B(n3072), .ZN(U3229)
         );
  AOI21_X1 U3890 ( .B1(n3078), .B2(n3077), .A(n3076), .ZN(n3084) );
  INV_X1 U3891 ( .A(n3863), .ZN(n4487) );
  AOI22_X1 U3892 ( .A1(n4487), .A2(n2547), .B1(n4485), .B2(n2228), .ZN(n3079)
         );
  OAI21_X1 U3893 ( .B1(n4491), .B2(n3080), .A(n3079), .ZN(n3081) );
  AOI21_X1 U3894 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3082), .A(n3081), .ZN(n3083)
         );
  OAI21_X1 U3895 ( .B1(n3084), .B2(n3858), .A(n3083), .ZN(U3234) );
  AOI211_X1 U3896 ( .C1(n3087), .C2(n3086), .A(n4606), .B(n3085), .ZN(n3094)
         );
  AOI211_X1 U3897 ( .C1(n3090), .C2(n3089), .A(n3088), .B(n4138), .ZN(n3093)
         );
  AND2_X1 U3898 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3285) );
  AOI21_X1 U3899 ( .B1(n4612), .B2(ADDR_REG_5__SCAN_IN), .A(n3285), .ZN(n3091)
         );
  OAI21_X1 U3900 ( .B1(n4619), .B2(n2278), .A(n3091), .ZN(n3092) );
  OR3_X1 U3901 ( .A1(n3094), .A2(n3093), .A3(n3092), .ZN(U3245) );
  MUX2_X1 U3902 ( .A(n4101), .B(REG2_REG_7__SCAN_IN), .S(n4475), .Z(n3096) );
  AOI211_X1 U3903 ( .C1(n3097), .C2(n3096), .A(n4606), .B(n4099), .ZN(n3106)
         );
  INV_X1 U3904 ( .A(n3098), .ZN(n3100) );
  XNOR2_X1 U3905 ( .A(n4475), .B(REG1_REG_7__SCAN_IN), .ZN(n3102) );
  OAI21_X1 U3906 ( .B1(n4075), .B2(n3102), .A(n4613), .ZN(n3101) );
  AOI21_X1 U3907 ( .B1(n4075), .B2(n3102), .A(n3101), .ZN(n3105) );
  INV_X1 U3908 ( .A(n4475), .ZN(n4102) );
  AND2_X1 U3909 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3334) );
  AOI21_X1 U3910 ( .B1(n4612), .B2(ADDR_REG_7__SCAN_IN), .A(n3334), .ZN(n3103)
         );
  OAI21_X1 U3911 ( .B1(n4619), .B2(n4102), .A(n3103), .ZN(n3104) );
  OR3_X1 U3912 ( .A1(n3106), .A2(n3105), .A3(n3104), .ZN(U3247) );
  OR2_X1 U3913 ( .A1(n4509), .A2(REG2_REG_0__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3914 ( .A1(n3108), .A2(n3107), .ZN(n4508) );
  NAND2_X1 U3915 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4060) );
  OAI21_X1 U3916 ( .B1(n4060), .B2(n4037), .A(U4043), .ZN(n3111) );
  NOR3_X1 U3917 ( .A1(n3109), .A2(n4470), .A3(n4482), .ZN(n3110) );
  AOI211_X1 U3918 ( .C1(n3065), .C2(n4508), .A(n3111), .B(n3110), .ZN(n3131)
         );
  AND3_X1 U3919 ( .A1(n3113), .A2(n4061), .A3(n3112), .ZN(n3114) );
  OAI211_X1 U3920 ( .C1(n3117), .C2(n3116), .A(n4613), .B(n3115), .ZN(n3118)
         );
  INV_X1 U3921 ( .A(n3118), .ZN(n3121) );
  AOI22_X1 U3922 ( .A1(n4612), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3119) );
  OAI21_X1 U3923 ( .B1(n4619), .B2(n2556), .A(n3119), .ZN(n3120) );
  OR4_X1 U3924 ( .A1(n3131), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(U3242) );
  XOR2_X1 U3925 ( .A(REG2_REG_4__SCAN_IN), .B(n3123), .Z(n3133) );
  INV_X1 U3926 ( .A(n3124), .ZN(n3125) );
  INV_X1 U3927 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U3928 ( .A1(n3125), .A2(n4694), .ZN(n3126) );
  NAND3_X1 U3929 ( .A1(n4613), .A2(n3127), .A3(n3126), .ZN(n3129) );
  AND2_X1 U3930 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3203) );
  AOI21_X1 U3931 ( .B1(n4612), .B2(ADDR_REG_4__SCAN_IN), .A(n3203), .ZN(n3128)
         );
  OAI211_X1 U3932 ( .C1(n4619), .C2(n3130), .A(n3129), .B(n3128), .ZN(n3132)
         );
  AOI211_X1 U3933 ( .C1(n4568), .C2(n3133), .A(n3132), .B(n3131), .ZN(n3134)
         );
  INV_X1 U3934 ( .A(n3134), .ZN(U3244) );
  INV_X1 U3935 ( .A(n3135), .ZN(n3136) );
  NOR2_X1 U3936 ( .A1(n3175), .A2(n3136), .ZN(n4661) );
  NAND2_X1 U3937 ( .A1(n4058), .A2(n3175), .ZN(n3954) );
  AND2_X1 U3938 ( .A1(n3952), .A2(n3954), .ZN(n3916) );
  INV_X1 U3939 ( .A(n3245), .ZN(n3454) );
  NOR2_X1 U3940 ( .A1(n3454), .A2(n4324), .ZN(n3137) );
  OAI22_X1 U3941 ( .A1(n3916), .A2(n3137), .B1(n3224), .B2(n4296), .ZN(n4660)
         );
  AOI21_X1 U3942 ( .B1(n4661), .B2(n3138), .A(n4660), .ZN(n3150) );
  NAND2_X1 U3943 ( .A1(n3139), .A2(D_REG_1__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U3944 ( .A1(n4643), .A2(n3140), .ZN(n3141) );
  NAND4_X1 U3945 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3145)
         );
  AOI22_X1 U3946 ( .A1(n2229), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4634), .ZN(n3149) );
  INV_X1 U3947 ( .A(n3916), .ZN(n4662) );
  OR2_X1 U3948 ( .A1(n3146), .A2(n4133), .ZN(n3244) );
  INV_X1 U3949 ( .A(n3244), .ZN(n3147) );
  AND2_X1 U3950 ( .A1(n4507), .A2(n3147), .ZN(n4638) );
  NAND2_X1 U3951 ( .A1(n4662), .A2(n4638), .ZN(n3148) );
  OAI211_X1 U3952 ( .C1(n3150), .C2(n2229), .A(n3149), .B(n3148), .ZN(U3290)
         );
  XNOR2_X1 U3953 ( .A(n3152), .B(n3151), .ZN(n3153) );
  NAND2_X1 U3954 ( .A1(n3153), .A2(n4498), .ZN(n3159) );
  OAI22_X1 U3955 ( .A1(n4491), .A2(n3162), .B1(n3180), .B2(n3863), .ZN(n3157)
         );
  INV_X1 U3956 ( .A(n3154), .ZN(n3155) );
  OAI21_X1 U3957 ( .B1(n3867), .B2(n3254), .A(n3155), .ZN(n3156) );
  NOR2_X1 U3958 ( .A1(n3157), .A2(n3156), .ZN(n3158) );
  OAI211_X1 U3959 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4503), .A(n3159), .B(n3158), 
        .ZN(U3215) );
  INV_X1 U3960 ( .A(n3160), .ZN(n3939) );
  XNOR2_X1 U3961 ( .A(n3161), .B(n3939), .ZN(n3266) );
  OAI22_X1 U3962 ( .A1(n3180), .A2(n4406), .B1(n3162), .B2(n4405), .ZN(n3165)
         );
  XNOR2_X1 U3963 ( .A(n3163), .B(n3939), .ZN(n3164) );
  OAI22_X1 U3964 ( .A1(n3164), .A2(n4182), .B1(n3254), .B2(n4296), .ZN(n3259)
         );
  AOI211_X1 U3965 ( .C1(n4681), .C2(n3266), .A(n3165), .B(n3259), .ZN(n3169)
         );
  AND2_X1 U3966 ( .A1(n4670), .A2(n3261), .ZN(n3166) );
  NOR2_X1 U3967 ( .A1(n3190), .A2(n3166), .ZN(n3260) );
  AOI22_X1 U3968 ( .A1(n3260), .A2(n4423), .B1(REG0_REG_3__SCAN_IN), .B2(n4689), .ZN(n3167) );
  OAI21_X1 U3969 ( .B1(n3169), .B2(n4689), .A(n3167), .ZN(U3473) );
  AOI22_X1 U3970 ( .A1(n3260), .A2(n2866), .B1(REG1_REG_3__SCAN_IN), .B2(n4697), .ZN(n3168) );
  OAI21_X1 U3971 ( .B1(n3169), .B2(n4697), .A(n3168), .ZN(U3521) );
  OR2_X1 U3972 ( .A1(n2783), .A2(n3170), .ZN(n3171) );
  NAND2_X1 U3973 ( .A1(n3172), .A2(n3171), .ZN(n4665) );
  INV_X1 U3974 ( .A(n4665), .ZN(n3187) );
  AND2_X1 U3975 ( .A1(n4669), .A2(n4133), .ZN(n3173) );
  OAI21_X1 U3976 ( .B1(n3175), .B2(n3174), .A(n3217), .ZN(n4663) );
  OAI22_X1 U3977 ( .A1(n4339), .A2(n4663), .B1(n3176), .B2(n4261), .ZN(n3186)
         );
  NAND2_X1 U3978 ( .A1(n3177), .A2(n4327), .ZN(n3179) );
  NAND2_X1 U3979 ( .A1(n4058), .A2(n4241), .ZN(n3178) );
  OAI211_X1 U3980 ( .C1(n3180), .C2(n4296), .A(n3179), .B(n3178), .ZN(n3181)
         );
  INV_X1 U3981 ( .A(n3181), .ZN(n3184) );
  XNOR2_X1 U3982 ( .A(n2783), .B(n3952), .ZN(n3182) );
  NAND2_X1 U3983 ( .A1(n3182), .A2(n4324), .ZN(n3183) );
  OAI211_X1 U3984 ( .C1(n4665), .C2(n3245), .A(n3184), .B(n3183), .ZN(n4667)
         );
  MUX2_X1 U3985 ( .A(REG2_REG_1__SCAN_IN), .B(n4667), .S(n4507), .Z(n3185) );
  AOI211_X1 U3986 ( .C1(n3187), .C2(n4638), .A(n3186), .B(n3185), .ZN(n3188)
         );
  INV_X1 U3987 ( .A(n3188), .ZN(U3289) );
  INV_X1 U3988 ( .A(n3189), .ZN(n3239) );
  OAI211_X1 U3989 ( .C1(n3190), .C2(n3206), .A(n3239), .B(n4669), .ZN(n4674)
         );
  NOR2_X1 U3990 ( .A1(n4674), .A2(n4473), .ZN(n3199) );
  XNOR2_X1 U3991 ( .A(n3191), .B(n3938), .ZN(n3200) );
  XOR2_X1 U3992 ( .A(n3938), .B(n3192), .Z(n3197) );
  AOI22_X1 U3993 ( .A1(n4053), .A2(n4328), .B1(n4327), .B2(n3193), .ZN(n3194)
         );
  OAI21_X1 U3994 ( .B1(n3195), .B2(n4406), .A(n3194), .ZN(n3196) );
  AOI21_X1 U3995 ( .B1(n3197), .B2(n4324), .A(n3196), .ZN(n3198) );
  OAI21_X1 U3996 ( .B1(n3245), .B2(n3200), .A(n3198), .ZN(n4675) );
  AOI211_X1 U3997 ( .C1(n4634), .C2(n3212), .A(n3199), .B(n4675), .ZN(n3202)
         );
  INV_X1 U3998 ( .A(n3200), .ZN(n4677) );
  AOI22_X1 U3999 ( .A1(n4677), .A2(n4638), .B1(REG2_REG_4__SCAN_IN), .B2(n2229), .ZN(n3201) );
  OAI21_X1 U4000 ( .B1(n3202), .B2(n2229), .A(n3201), .ZN(U3286) );
  INV_X1 U4001 ( .A(n4503), .ZN(n3834) );
  AOI21_X1 U4002 ( .B1(n4485), .B2(n4053), .A(n3203), .ZN(n3205) );
  NAND2_X1 U4003 ( .A1(n4487), .A2(n2228), .ZN(n3204) );
  OAI211_X1 U4004 ( .C1(n4491), .C2(n3206), .A(n3205), .B(n3204), .ZN(n3211)
         );
  AOI211_X1 U4005 ( .C1(n3209), .C2(n3208), .A(n3858), .B(n3207), .ZN(n3210)
         );
  AOI211_X1 U4006 ( .C1(n3212), .C2(n3834), .A(n3211), .B(n3210), .ZN(n3213)
         );
  INV_X1 U4007 ( .A(n3213), .ZN(U3227) );
  NAND2_X1 U4008 ( .A1(n3215), .A2(n3220), .ZN(n3216) );
  NAND2_X1 U4009 ( .A1(n3214), .A2(n3216), .ZN(n4673) );
  INV_X1 U4010 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4011 ( .A1(n3217), .A2(n3222), .ZN(n4668) );
  NAND3_X1 U4012 ( .A1(n4637), .A2(n4670), .A3(n4668), .ZN(n3218) );
  OAI21_X1 U4013 ( .B1(n4261), .B2(n3219), .A(n3218), .ZN(n3230) );
  XNOR2_X1 U4014 ( .A(n3221), .B(n2785), .ZN(n3228) );
  NAND2_X1 U4015 ( .A1(n4673), .A2(n3454), .ZN(n3227) );
  AOI22_X1 U4016 ( .A1(n2228), .A2(n4328), .B1(n4327), .B2(n3222), .ZN(n3223)
         );
  OAI21_X1 U4017 ( .B1(n3224), .B2(n4406), .A(n3223), .ZN(n3225) );
  INV_X1 U4018 ( .A(n3225), .ZN(n3226) );
  OAI211_X1 U4019 ( .C1(n3228), .C2(n4182), .A(n3227), .B(n3226), .ZN(n4671)
         );
  MUX2_X1 U4020 ( .A(n4671), .B(REG2_REG_2__SCAN_IN), .S(n2229), .Z(n3229) );
  AOI211_X1 U4021 ( .C1(n4638), .C2(n4673), .A(n3230), .B(n3229), .ZN(n3231)
         );
  INV_X1 U4022 ( .A(n3231), .ZN(U3288) );
  INV_X1 U4023 ( .A(n3233), .ZN(n3966) );
  NAND2_X1 U4024 ( .A1(n3966), .A2(n3981), .ZN(n3921) );
  INV_X1 U4025 ( .A(n3921), .ZN(n3234) );
  XNOR2_X1 U4026 ( .A(n3232), .B(n3234), .ZN(n3256) );
  OAI22_X1 U4027 ( .A1(n3254), .A2(n4406), .B1(n3283), .B2(n4405), .ZN(n3237)
         );
  XOR2_X1 U4028 ( .A(n3921), .B(n3235), .Z(n3236) );
  OAI22_X1 U4029 ( .A1(n3236), .A2(n4182), .B1(n3332), .B2(n4296), .ZN(n3243)
         );
  AOI211_X1 U4030 ( .C1(n3256), .C2(n4681), .A(n3237), .B(n3243), .ZN(n3242)
         );
  INV_X1 U4031 ( .A(n3299), .ZN(n3238) );
  AOI21_X1 U4032 ( .B1(n3250), .B2(n3239), .A(n3238), .ZN(n3247) );
  AOI22_X1 U4033 ( .A1(n3247), .A2(n2866), .B1(REG1_REG_5__SCAN_IN), .B2(n4697), .ZN(n3240) );
  OAI21_X1 U4034 ( .B1(n3242), .B2(n4697), .A(n3240), .ZN(U3523) );
  AOI22_X1 U4035 ( .A1(n3247), .A2(n4423), .B1(REG0_REG_5__SCAN_IN), .B2(n4689), .ZN(n3241) );
  OAI21_X1 U4036 ( .B1(n3242), .B2(n4689), .A(n3241), .ZN(U3477) );
  INV_X1 U4037 ( .A(n3243), .ZN(n3258) );
  NAND2_X1 U4038 ( .A1(n3245), .A2(n3244), .ZN(n3246) );
  INV_X1 U4039 ( .A(n4313), .ZN(n3253) );
  NAND2_X1 U4040 ( .A1(n3247), .A2(n4637), .ZN(n3252) );
  NAND2_X1 U4041 ( .A1(n4507), .A2(n4327), .ZN(n4307) );
  INV_X1 U4042 ( .A(n4307), .ZN(n3324) );
  INV_X1 U40430 ( .A(n3248), .ZN(n3288) );
  OAI22_X1 U4044 ( .A1(n4507), .A2(n2277), .B1(n3288), .B2(n4261), .ZN(n3249)
         );
  AOI21_X1 U4045 ( .B1(n3250), .B2(n3324), .A(n3249), .ZN(n3251) );
  OAI211_X1 U4046 ( .C1(n3254), .C2(n3253), .A(n3252), .B(n3251), .ZN(n3255)
         );
  AOI21_X1 U4047 ( .B1(n3256), .B2(n4304), .A(n3255), .ZN(n3257) );
  OAI21_X1 U4048 ( .B1(n3258), .B2(n2229), .A(n3257), .ZN(U3285) );
  INV_X1 U4049 ( .A(n3259), .ZN(n3268) );
  INV_X1 U4050 ( .A(n3260), .ZN(n3264) );
  AOI22_X1 U4051 ( .A1(n2229), .A2(REG2_REG_3__SCAN_IN), .B1(n4634), .B2(n2560), .ZN(n3263) );
  AOI22_X1 U4052 ( .A1(n3324), .A2(n3261), .B1(n4313), .B2(n4056), .ZN(n3262)
         );
  OAI211_X1 U4053 ( .C1(n3264), .C2(n4339), .A(n3263), .B(n3262), .ZN(n3265)
         );
  AOI21_X1 U4054 ( .B1(n3266), .B2(n4304), .A(n3265), .ZN(n3267) );
  OAI21_X1 U4055 ( .B1(n3268), .B2(n2229), .A(n3267), .ZN(U3287) );
  INV_X1 U4056 ( .A(n4669), .ZN(n4683) );
  AOI211_X1 U4057 ( .C1(n3271), .C2(n3297), .A(n4683), .B(n2268), .ZN(n4680)
         );
  INV_X1 U4058 ( .A(n3924), .ZN(n3970) );
  XNOR2_X1 U4059 ( .A(n3269), .B(n3970), .ZN(n3270) );
  NAND2_X1 U4060 ( .A1(n3270), .A2(n4324), .ZN(n3273) );
  AOI22_X1 U4061 ( .A1(n3343), .A2(n4328), .B1(n4327), .B2(n3271), .ZN(n3272)
         );
  OAI211_X1 U4062 ( .C1(n3332), .C2(n4406), .A(n3273), .B(n3272), .ZN(n4679)
         );
  AOI21_X1 U4063 ( .B1(n4680), .B2(n4133), .A(n4679), .ZN(n3278) );
  XOR2_X1 U4064 ( .A(n3274), .B(n3924), .Z(n4682) );
  INV_X1 U4065 ( .A(n3275), .ZN(n3340) );
  OAI22_X1 U4066 ( .A1(n4507), .A2(n4101), .B1(n3340), .B2(n4261), .ZN(n3276)
         );
  AOI21_X1 U4067 ( .B1(n4682), .B2(n4304), .A(n3276), .ZN(n3277) );
  OAI21_X1 U4068 ( .B1(n3278), .B2(n2229), .A(n3277), .ZN(U3283) );
  AOI211_X1 U4069 ( .C1(n3281), .C2(n3280), .A(n3858), .B(n3279), .ZN(n3282)
         );
  INV_X1 U4070 ( .A(n3282), .ZN(n3287) );
  OAI22_X1 U4071 ( .A1(n4491), .A2(n3283), .B1(n3332), .B2(n3867), .ZN(n3284)
         );
  AOI211_X1 U4072 ( .C1(n4487), .C2(n4054), .A(n3285), .B(n3284), .ZN(n3286)
         );
  OAI211_X1 U4073 ( .C1(n4503), .C2(n3288), .A(n3287), .B(n3286), .ZN(U3224)
         );
  NAND2_X1 U4074 ( .A1(n3969), .A2(n3979), .ZN(n3940) );
  XNOR2_X1 U4075 ( .A(n3289), .B(n3940), .ZN(n4639) );
  XNOR2_X1 U4076 ( .A(n3290), .B(n3940), .ZN(n3294) );
  OAI22_X1 U4077 ( .A1(n3313), .A2(n4406), .B1(n3310), .B2(n4405), .ZN(n3291)
         );
  AOI21_X1 U4078 ( .B1(n4328), .B2(n3292), .A(n3291), .ZN(n3293) );
  OAI21_X1 U4079 ( .B1(n3294), .B2(n4182), .A(n3293), .ZN(n3295) );
  AOI21_X1 U4080 ( .B1(n3454), .B2(n4639), .A(n3295), .ZN(n4642) );
  INV_X1 U4081 ( .A(n4642), .ZN(n3296) );
  AOI21_X1 U4082 ( .B1(n4688), .B2(n4639), .A(n3296), .ZN(n3305) );
  INV_X1 U4083 ( .A(n3297), .ZN(n3298) );
  AOI21_X1 U4084 ( .B1(n3300), .B2(n3299), .A(n3298), .ZN(n4636) );
  INV_X1 U4085 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3301) );
  NOR2_X1 U4086 ( .A1(n4690), .A2(n3301), .ZN(n3302) );
  AOI21_X1 U4087 ( .B1(n4636), .B2(n4423), .A(n3302), .ZN(n3303) );
  OAI21_X1 U4088 ( .B1(n3305), .B2(n4689), .A(n3303), .ZN(U3479) );
  AOI22_X1 U4089 ( .A1(n4636), .A2(n2866), .B1(n4697), .B2(REG1_REG_6__SCAN_IN), .ZN(n3304) );
  OAI21_X1 U4090 ( .B1(n3305), .B2(n4697), .A(n3304), .ZN(U3524) );
  INV_X1 U4091 ( .A(n4635), .ZN(n3318) );
  XNOR2_X1 U4092 ( .A(n3307), .B(n3306), .ZN(n3308) );
  XNOR2_X1 U4093 ( .A(n2267), .B(n3308), .ZN(n3309) );
  NAND2_X1 U4094 ( .A1(n3309), .A2(n4498), .ZN(n3317) );
  OAI22_X1 U4095 ( .A1(n4491), .A2(n3310), .B1(n3368), .B2(n3867), .ZN(n3315)
         );
  INV_X1 U4096 ( .A(n3311), .ZN(n3312) );
  OAI21_X1 U4097 ( .B1(n3863), .B2(n3313), .A(n3312), .ZN(n3314) );
  NOR2_X1 U4098 ( .A1(n3315), .A2(n3314), .ZN(n3316) );
  OAI211_X1 U4099 ( .C1(n4503), .C2(n3318), .A(n3317), .B(n3316), .ZN(U3236)
         );
  INV_X1 U4100 ( .A(n3989), .ZN(n3319) );
  NAND2_X1 U4101 ( .A1(n3319), .A2(n3974), .ZN(n3922) );
  XNOR2_X1 U4102 ( .A(n3320), .B(n3922), .ZN(n3322) );
  AND2_X1 U4103 ( .A1(n4050), .A2(n4328), .ZN(n3321) );
  AOI21_X1 U4104 ( .B1(n3322), .B2(n4324), .A(n3321), .ZN(n3346) );
  XNOR2_X1 U4105 ( .A(n3323), .B(n3922), .ZN(n3341) );
  INV_X1 U4106 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4902) );
  OAI22_X1 U4107 ( .A1(n3389), .A2(n4261), .B1(n4902), .B2(n4507), .ZN(n3327)
         );
  OAI21_X1 U4108 ( .B1(n3363), .B2(n3383), .A(n3432), .ZN(n3352) );
  AOI22_X1 U4109 ( .A1(n3324), .A2(n3342), .B1(n4313), .B2(n3343), .ZN(n3325)
         );
  OAI21_X1 U4110 ( .B1(n3352), .B2(n4339), .A(n3325), .ZN(n3326) );
  AOI211_X1 U4111 ( .C1(n3341), .C2(n4304), .A(n3327), .B(n3326), .ZN(n3328)
         );
  OAI21_X1 U4112 ( .B1(n2229), .B2(n3346), .A(n3328), .ZN(U3281) );
  XOR2_X1 U4113 ( .A(n3330), .B(n3329), .Z(n3331) );
  NAND2_X1 U4114 ( .A1(n3331), .A2(n4498), .ZN(n3339) );
  OAI22_X1 U4115 ( .A1(n4491), .A2(n3333), .B1(n3332), .B2(n3863), .ZN(n3337)
         );
  INV_X1 U4116 ( .A(n3334), .ZN(n3335) );
  OAI21_X1 U4117 ( .B1(n3867), .B2(n3382), .A(n3335), .ZN(n3336) );
  NOR2_X1 U4118 ( .A1(n3337), .A2(n3336), .ZN(n3338) );
  OAI211_X1 U4119 ( .C1(n4503), .C2(n3340), .A(n3339), .B(n3338), .ZN(U3210)
         );
  NAND2_X1 U4120 ( .A1(n3341), .A2(n4681), .ZN(n3345) );
  AOI22_X1 U4121 ( .A1(n3343), .A2(n4241), .B1(n3342), .B2(n4327), .ZN(n3344)
         );
  NAND3_X1 U4122 ( .A1(n3346), .A2(n3345), .A3(n3344), .ZN(n3349) );
  MUX2_X1 U4123 ( .A(n3349), .B(REG0_REG_9__SCAN_IN), .S(n4689), .Z(n3347) );
  INV_X1 U4124 ( .A(n3347), .ZN(n3348) );
  OAI21_X1 U4125 ( .B1(n3352), .B2(n4466), .A(n3348), .ZN(U3485) );
  MUX2_X1 U4126 ( .A(REG1_REG_9__SCAN_IN), .B(n3349), .S(n4700), .Z(n3350) );
  INV_X1 U4127 ( .A(n3350), .ZN(n3351) );
  OAI21_X1 U4128 ( .B1(n4412), .B2(n3352), .A(n3351), .ZN(U3527) );
  NOR2_X1 U4129 ( .A1(n2432), .A2(n3354), .ZN(n3355) );
  XNOR2_X1 U4130 ( .A(n3356), .B(n3355), .ZN(n3357) );
  NAND2_X1 U4131 ( .A1(n3357), .A2(n4498), .ZN(n3361) );
  OAI22_X1 U4132 ( .A1(n4491), .A2(n3367), .B1(n3368), .B2(n3863), .ZN(n3359)
         );
  NAND2_X1 U4133 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4518) );
  OAI21_X1 U4134 ( .B1(n3867), .B2(n3438), .A(n4518), .ZN(n3358) );
  NOR2_X1 U4135 ( .A1(n3359), .A2(n3358), .ZN(n3360) );
  OAI211_X1 U4136 ( .C1(n4503), .C2(n3362), .A(n3361), .B(n3360), .ZN(U3218)
         );
  INV_X1 U4137 ( .A(n3363), .ZN(n3364) );
  OAI21_X1 U4138 ( .B1(n2268), .B2(n3367), .A(n3364), .ZN(n4628) );
  INV_X1 U4139 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U4140 ( .A1(n3975), .A2(n3972), .ZN(n3919) );
  XOR2_X1 U4141 ( .A(n3919), .B(n3365), .Z(n4630) );
  XOR2_X1 U4142 ( .A(n3919), .B(n3366), .Z(n3371) );
  OAI22_X1 U4143 ( .A1(n3368), .A2(n4406), .B1(n3367), .B2(n4405), .ZN(n3369)
         );
  AOI21_X1 U4144 ( .B1(n4328), .B2(n4051), .A(n3369), .ZN(n3370) );
  OAI21_X1 U4145 ( .B1(n3371), .B2(n4182), .A(n3370), .ZN(n3372) );
  AOI21_X1 U4146 ( .B1(n3454), .B2(n4630), .A(n3372), .ZN(n4633) );
  INV_X1 U4147 ( .A(n4633), .ZN(n3373) );
  AOI21_X1 U4148 ( .B1(n4688), .B2(n4630), .A(n3373), .ZN(n3376) );
  MUX2_X1 U4149 ( .A(n3374), .B(n3376), .S(n4690), .Z(n3375) );
  OAI21_X1 U4150 ( .B1(n4628), .B2(n4466), .A(n3375), .ZN(U3483) );
  INV_X1 U4151 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3377) );
  MUX2_X1 U4152 ( .A(n3377), .B(n3376), .S(n4700), .Z(n3378) );
  OAI21_X1 U4153 ( .B1(n4628), .B2(n4412), .A(n3378), .ZN(U3526) );
  XNOR2_X1 U4154 ( .A(n3380), .B(n3379), .ZN(n3381) );
  NAND2_X1 U4155 ( .A1(n3381), .A2(n4498), .ZN(n3388) );
  OAI22_X1 U4156 ( .A1(n4491), .A2(n3383), .B1(n3382), .B2(n3863), .ZN(n3386)
         );
  INV_X1 U4157 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4987) );
  NOR2_X1 U4158 ( .A1(STATE_REG_SCAN_IN), .A2(n4987), .ZN(n4533) );
  INV_X1 U4159 ( .A(n4533), .ZN(n3384) );
  OAI21_X1 U4160 ( .B1(n3867), .B2(n3476), .A(n3384), .ZN(n3385) );
  NOR2_X1 U4161 ( .A1(n3386), .A2(n3385), .ZN(n3387) );
  OAI211_X1 U4162 ( .C1(n4503), .C2(n3389), .A(n3388), .B(n3387), .ZN(U3228)
         );
  XNOR2_X1 U4163 ( .A(n3403), .B(n3925), .ZN(n3394) );
  XNOR2_X1 U4164 ( .A(n3390), .B(n3925), .ZN(n4687) );
  NAND2_X1 U4165 ( .A1(n4687), .A2(n3454), .ZN(n3393) );
  OAI22_X1 U4166 ( .A1(n3531), .A2(n4296), .B1(n4405), .B2(n3474), .ZN(n3391)
         );
  AOI21_X1 U4167 ( .B1(n4241), .B2(n4050), .A(n3391), .ZN(n3392) );
  OAI211_X1 U4168 ( .C1(n4182), .C2(n3394), .A(n3393), .B(n3392), .ZN(n4685)
         );
  INV_X1 U4169 ( .A(n4685), .ZN(n3399) );
  NAND2_X1 U4170 ( .A1(n3433), .A2(n3469), .ZN(n3395) );
  NAND2_X1 U4171 ( .A1(n3406), .A2(n3395), .ZN(n4684) );
  AOI22_X1 U4172 ( .A1(n2229), .A2(REG2_REG_11__SCAN_IN), .B1(n3461), .B2(
        n4634), .ZN(n3396) );
  OAI21_X1 U4173 ( .B1(n4684), .B2(n4339), .A(n3396), .ZN(n3397) );
  AOI21_X1 U4174 ( .B1(n4687), .B2(n4638), .A(n3397), .ZN(n3398) );
  OAI21_X1 U4175 ( .B1(n3399), .B2(n2229), .A(n3398), .ZN(U3279) );
  NAND2_X1 U4176 ( .A1(n3419), .A2(n3417), .ZN(n3920) );
  INV_X1 U4177 ( .A(n3400), .ZN(n3401) );
  AOI21_X1 U4178 ( .B1(n3403), .B2(n3402), .A(n3401), .ZN(n3420) );
  XOR2_X1 U4179 ( .A(n3920), .B(n3420), .Z(n3404) );
  OAI22_X1 U4180 ( .A1(n3404), .A2(n4182), .B1(n3628), .B2(n4296), .ZN(n3482)
         );
  INV_X1 U4181 ( .A(n3482), .ZN(n3414) );
  XNOR2_X1 U4182 ( .A(n3405), .B(n3920), .ZN(n3484) );
  INV_X1 U4183 ( .A(n3406), .ZN(n3408) );
  INV_X1 U4184 ( .A(n3426), .ZN(n3407) );
  OAI21_X1 U4185 ( .B1(n3408), .B2(n3561), .A(n3407), .ZN(n3490) );
  NOR2_X1 U4186 ( .A1(n3490), .A2(n4339), .ZN(n3412) );
  AOI22_X1 U4187 ( .A1(n2229), .A2(REG2_REG_12__SCAN_IN), .B1(n3550), .B2(
        n4634), .ZN(n3410) );
  NAND2_X1 U4188 ( .A1(n4313), .A2(n3440), .ZN(n3409) );
  OAI211_X1 U4189 ( .C1(n4307), .C2(n3561), .A(n3410), .B(n3409), .ZN(n3411)
         );
  AOI211_X1 U4190 ( .C1(n3484), .C2(n4304), .A(n3412), .B(n3411), .ZN(n3413)
         );
  OAI21_X1 U4191 ( .B1(n3414), .B2(n2229), .A(n3413), .ZN(U3278) );
  XNOR2_X1 U4192 ( .A(n3416), .B(n3415), .ZN(n3934) );
  INV_X1 U4193 ( .A(n3417), .ZN(n3418) );
  AOI21_X1 U4194 ( .B1(n3420), .B2(n3419), .A(n3418), .ZN(n3421) );
  XOR2_X1 U4195 ( .A(n3934), .B(n3421), .Z(n3424) );
  OAI22_X1 U4196 ( .A1(n3864), .A2(n4296), .B1(n4405), .B2(n3529), .ZN(n3422)
         );
  AOI21_X1 U4197 ( .B1(n4241), .B2(n3515), .A(n3422), .ZN(n3423) );
  OAI21_X1 U4198 ( .B1(n3424), .B2(n4182), .A(n3423), .ZN(n3491) );
  INV_X1 U4199 ( .A(n3491), .ZN(n3431) );
  XNOR2_X1 U4200 ( .A(n3425), .B(n3934), .ZN(n3492) );
  OR2_X1 U4201 ( .A1(n3426), .A2(n3529), .ZN(n3427) );
  NAND2_X1 U4202 ( .A1(n3455), .A2(n3427), .ZN(n3498) );
  AOI22_X1 U4203 ( .A1(n2229), .A2(REG2_REG_13__SCAN_IN), .B1(n3511), .B2(
        n4634), .ZN(n3428) );
  OAI21_X1 U4204 ( .B1(n3498), .B2(n4339), .A(n3428), .ZN(n3429) );
  AOI21_X1 U4205 ( .B1(n3492), .B2(n4304), .A(n3429), .ZN(n3430) );
  OAI21_X1 U4206 ( .B1(n3431), .B2(n2229), .A(n3430), .ZN(U3277) );
  INV_X1 U4207 ( .A(n3432), .ZN(n3434) );
  OAI21_X1 U4208 ( .B1(n3434), .B2(n3437), .A(n3433), .ZN(n4621) );
  INV_X1 U4209 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4816) );
  NAND2_X1 U4210 ( .A1(n3990), .A2(n3992), .ZN(n3941) );
  XOR2_X1 U4211 ( .A(n3941), .B(n3435), .Z(n4623) );
  XNOR2_X1 U4212 ( .A(n3436), .B(n3941), .ZN(n3442) );
  OAI22_X1 U4213 ( .A1(n3438), .A2(n4406), .B1(n3437), .B2(n4405), .ZN(n3439)
         );
  AOI21_X1 U4214 ( .B1(n4328), .B2(n3440), .A(n3439), .ZN(n3441) );
  OAI21_X1 U4215 ( .B1(n3442), .B2(n4182), .A(n3441), .ZN(n3443) );
  AOI21_X1 U4216 ( .B1(n4623), .B2(n3454), .A(n3443), .ZN(n4626) );
  INV_X1 U4217 ( .A(n4626), .ZN(n3444) );
  AOI21_X1 U4218 ( .B1(n4688), .B2(n4623), .A(n3444), .ZN(n3446) );
  MUX2_X1 U4219 ( .A(n4816), .B(n3446), .S(n4700), .Z(n3445) );
  OAI21_X1 U4220 ( .B1(n4621), .B2(n4412), .A(n3445), .ZN(U3528) );
  INV_X1 U4221 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4970) );
  MUX2_X1 U4222 ( .A(n4970), .B(n3446), .S(n4690), .Z(n3447) );
  OAI21_X1 U4223 ( .B1(n4621), .B2(n4466), .A(n3447), .ZN(U3487) );
  OAI21_X1 U4224 ( .B1(n3449), .B2(n3932), .A(n3448), .ZN(n4413) );
  OAI21_X1 U4225 ( .B1(n2391), .B2(n3882), .A(n3500), .ZN(n3450) );
  NAND2_X1 U4226 ( .A1(n3450), .A2(n4324), .ZN(n3452) );
  AOI22_X1 U4227 ( .A1(n4486), .A2(n4328), .B1(n4327), .B2(n3613), .ZN(n3451)
         );
  OAI211_X1 U4228 ( .C1(n3628), .C2(n4406), .A(n3452), .B(n3451), .ZN(n3453)
         );
  AOI21_X1 U4229 ( .B1(n4413), .B2(n3454), .A(n3453), .ZN(n4417) );
  NAND2_X1 U4230 ( .A1(n3455), .A2(n3613), .ZN(n4414) );
  AND3_X1 U4231 ( .A1(n4415), .A2(n4637), .A3(n4414), .ZN(n3459) );
  INV_X1 U4232 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3457) );
  INV_X1 U4233 ( .A(n3456), .ZN(n3634) );
  OAI22_X1 U4234 ( .A1(n4507), .A2(n3457), .B1(n3634), .B2(n4261), .ZN(n3458)
         );
  AOI211_X1 U4235 ( .C1(n4413), .C2(n4638), .A(n3459), .B(n3458), .ZN(n3460)
         );
  OAI21_X1 U4236 ( .B1(n4417), .B2(n2229), .A(n3460), .ZN(U3276) );
  INV_X1 U4237 ( .A(n3461), .ZN(n3481) );
  INV_X1 U4238 ( .A(n3462), .ZN(n3464) );
  NOR2_X1 U4239 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  OAI22_X1 U4240 ( .A1(n3562), .A2(n3733), .B1(n3732), .B2(n3474), .ZN(n3468)
         );
  XNOR2_X1 U4241 ( .A(n3468), .B(n3467), .ZN(n3551) );
  OR2_X1 U4242 ( .A1(n3562), .A2(n2906), .ZN(n3471) );
  NAND2_X1 U4243 ( .A1(n3469), .A2(n2908), .ZN(n3470) );
  XNOR2_X1 U4244 ( .A(n3551), .B(n3555), .ZN(n3472) );
  XNOR2_X1 U4245 ( .A(n3553), .B(n3472), .ZN(n3473) );
  NAND2_X1 U4246 ( .A1(n3473), .A2(n4498), .ZN(n3480) );
  OAI22_X1 U4247 ( .A1(n4491), .A2(n3474), .B1(n3531), .B2(n3867), .ZN(n3478)
         );
  NOR2_X1 U4248 ( .A1(STATE_REG_SCAN_IN), .A2(n4879), .ZN(n4554) );
  INV_X1 U4249 ( .A(n4554), .ZN(n3475) );
  OAI21_X1 U4250 ( .B1(n3863), .B2(n3476), .A(n3475), .ZN(n3477) );
  NOR2_X1 U4251 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  OAI211_X1 U4252 ( .C1(n4503), .C2(n3481), .A(n3480), .B(n3479), .ZN(U3233)
         );
  INV_X1 U4253 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3485) );
  OAI22_X1 U4254 ( .A1(n3562), .A2(n4406), .B1(n3561), .B2(n4405), .ZN(n3483)
         );
  AOI211_X1 U4255 ( .C1(n4681), .C2(n3484), .A(n3483), .B(n3482), .ZN(n3487)
         );
  MUX2_X1 U4256 ( .A(n3485), .B(n3487), .S(n4690), .Z(n3486) );
  OAI21_X1 U4257 ( .B1(n3490), .B2(n4466), .A(n3486), .ZN(U3491) );
  INV_X1 U4258 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3488) );
  MUX2_X1 U4259 ( .A(n3488), .B(n3487), .S(n4700), .Z(n3489) );
  OAI21_X1 U4260 ( .B1(n3490), .B2(n4412), .A(n3489), .ZN(U3530) );
  INV_X1 U4261 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3493) );
  AOI21_X1 U4262 ( .B1(n3492), .B2(n4681), .A(n3491), .ZN(n3495) );
  MUX2_X1 U4263 ( .A(n3493), .B(n3495), .S(n4690), .Z(n3494) );
  OAI21_X1 U4264 ( .B1(n3498), .B2(n4466), .A(n3494), .ZN(U3493) );
  INV_X1 U4265 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3496) );
  MUX2_X1 U4266 ( .A(n3496), .B(n3495), .S(n4700), .Z(n3497) );
  OAI21_X1 U4267 ( .B1(n4412), .B2(n3498), .A(n3497), .ZN(U3531) );
  XNOR2_X1 U4268 ( .A(n3499), .B(n3931), .ZN(n3570) );
  INV_X1 U4269 ( .A(n3570), .ZN(n3510) );
  NAND2_X1 U4270 ( .A1(n3500), .A2(n3878), .ZN(n3501) );
  XNOR2_X1 U4271 ( .A(n3501), .B(n3931), .ZN(n3502) );
  OAI22_X1 U4272 ( .A1(n3502), .A2(n4182), .B1(n4407), .B2(n4296), .ZN(n3569)
         );
  INV_X1 U4273 ( .A(n4415), .ZN(n3504) );
  INV_X1 U4274 ( .A(n3544), .ZN(n3503) );
  OAI21_X1 U4275 ( .B1(n3504), .B2(n3865), .A(n3503), .ZN(n3576) );
  NOR2_X1 U4276 ( .A1(n3576), .A2(n4339), .ZN(n3508) );
  AOI22_X1 U4277 ( .A1(n2229), .A2(REG2_REG_15__SCAN_IN), .B1(n3860), .B2(
        n4634), .ZN(n3506) );
  NAND2_X1 U4278 ( .A1(n4313), .A2(n4049), .ZN(n3505) );
  OAI211_X1 U4279 ( .C1(n4307), .C2(n3865), .A(n3506), .B(n3505), .ZN(n3507)
         );
  AOI211_X1 U4280 ( .C1(n3569), .C2(n4507), .A(n3508), .B(n3507), .ZN(n3509)
         );
  OAI21_X1 U4281 ( .B1(n3510), .B2(n4342), .A(n3509), .ZN(U3275) );
  INV_X1 U4282 ( .A(n3511), .ZN(n3536) );
  NAND2_X1 U4283 ( .A1(n3515), .A2(n2908), .ZN(n3513) );
  NAND2_X1 U4284 ( .A1(n3516), .A2(n3739), .ZN(n3512) );
  NAND2_X1 U4285 ( .A1(n3513), .A2(n3512), .ZN(n3514) );
  XNOR2_X1 U4286 ( .A(n3514), .B(n2947), .ZN(n3522) );
  NAND2_X1 U4287 ( .A1(n3515), .A2(n3741), .ZN(n3518) );
  NAND2_X1 U4288 ( .A1(n3516), .A2(n2908), .ZN(n3517) );
  NAND2_X1 U4289 ( .A1(n3518), .A2(n3517), .ZN(n3521) );
  NAND2_X1 U4290 ( .A1(n3522), .A2(n3521), .ZN(n3519) );
  OAI211_X1 U4291 ( .C1(n3552), .C2(n3551), .A(n3553), .B(n3519), .ZN(n3525)
         );
  INV_X1 U4292 ( .A(n3519), .ZN(n3556) );
  INV_X1 U4293 ( .A(n3551), .ZN(n3520) );
  NOR3_X1 U4294 ( .A1(n3556), .A2(n3520), .A3(n3555), .ZN(n3523) );
  NOR2_X1 U4295 ( .A1(n3522), .A2(n3521), .ZN(n3557) );
  NOR2_X1 U4296 ( .A1(n3523), .A2(n3557), .ZN(n3524) );
  NAND2_X1 U4297 ( .A1(n3525), .A2(n3524), .ZN(n3620) );
  OAI22_X1 U4298 ( .A1(n3628), .A2(n3733), .B1(n3732), .B2(n3529), .ZN(n3526)
         );
  XOR2_X1 U4299 ( .A(n2947), .B(n3526), .Z(n3621) );
  OAI22_X1 U4300 ( .A1(n3628), .A2(n2906), .B1(n3733), .B2(n3529), .ZN(n3624)
         );
  XNOR2_X1 U4301 ( .A(n3621), .B(n3624), .ZN(n3527) );
  XNOR2_X1 U4302 ( .A(n3620), .B(n3527), .ZN(n3528) );
  NAND2_X1 U4303 ( .A1(n3528), .A2(n4498), .ZN(n3535) );
  OAI22_X1 U4304 ( .A1(n4491), .A2(n3529), .B1(n3864), .B2(n3867), .ZN(n3533)
         );
  AND2_X1 U4305 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4573) );
  INV_X1 U4306 ( .A(n4573), .ZN(n3530) );
  OAI21_X1 U4307 ( .B1(n3863), .B2(n3531), .A(n3530), .ZN(n3532) );
  NOR2_X1 U4308 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  OAI211_X1 U4309 ( .C1(n4503), .C2(n3536), .A(n3535), .B(n3534), .ZN(U3231)
         );
  XNOR2_X1 U4310 ( .A(n3537), .B(n3942), .ZN(n3541) );
  NAND2_X1 U4311 ( .A1(n3653), .A2(n4327), .ZN(n3539) );
  NAND2_X1 U4312 ( .A1(n4486), .A2(n4241), .ZN(n3538) );
  OAI211_X1 U4313 ( .C1(n3845), .C2(n4296), .A(n3539), .B(n3538), .ZN(n3540)
         );
  AOI21_X1 U4314 ( .B1(n3541), .B2(n4324), .A(n3540), .ZN(n3588) );
  OAI21_X1 U4315 ( .B1(n3543), .B2(n3942), .A(n3542), .ZN(n3587) );
  OR2_X1 U4316 ( .A1(n3587), .A2(n4342), .ZN(n3549) );
  NOR2_X1 U4317 ( .A1(n3544), .A2(n4490), .ZN(n3545) );
  OR2_X1 U4318 ( .A1(n3579), .A2(n3545), .ZN(n3595) );
  INV_X1 U4319 ( .A(n3595), .ZN(n3547) );
  OAI22_X1 U4320 ( .A1(n4507), .A2(n4597), .B1(n4502), .B2(n4261), .ZN(n3546)
         );
  AOI21_X1 U4321 ( .B1(n3547), .B2(n4637), .A(n3546), .ZN(n3548) );
  OAI211_X1 U4322 ( .C1(n2229), .C2(n3588), .A(n3549), .B(n3548), .ZN(U3274)
         );
  INV_X1 U4323 ( .A(n3550), .ZN(n3567) );
  AOI21_X1 U4324 ( .B1(n3553), .B2(n3552), .A(n3551), .ZN(n3554) );
  AOI21_X1 U4325 ( .B1(n2433), .B2(n3555), .A(n3554), .ZN(n3559) );
  NOR2_X1 U4326 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  XNOR2_X1 U4327 ( .A(n3559), .B(n3558), .ZN(n3560) );
  NAND2_X1 U4328 ( .A1(n3560), .A2(n4498), .ZN(n3566) );
  OAI22_X1 U4329 ( .A1(n4491), .A2(n3561), .B1(n3628), .B2(n3867), .ZN(n3564)
         );
  NAND2_X1 U4330 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4559) );
  OAI21_X1 U4331 ( .B1(n3863), .B2(n3562), .A(n4559), .ZN(n3563) );
  NOR2_X1 U4332 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  OAI211_X1 U4333 ( .C1(n4503), .C2(n3567), .A(n3566), .B(n3565), .ZN(U3221)
         );
  INV_X1 U4334 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3571) );
  OAI22_X1 U4335 ( .A1(n3864), .A2(n4406), .B1(n3865), .B2(n4405), .ZN(n3568)
         );
  AOI211_X1 U4336 ( .C1(n3570), .C2(n4681), .A(n3569), .B(n3568), .ZN(n3573)
         );
  MUX2_X1 U4337 ( .A(n3571), .B(n3573), .S(n4700), .Z(n3572) );
  OAI21_X1 U4338 ( .B1(n4412), .B2(n3576), .A(n3572), .ZN(U3533) );
  INV_X1 U4339 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3574) );
  MUX2_X1 U4340 ( .A(n3574), .B(n3573), .S(n4690), .Z(n3575) );
  OAI21_X1 U4341 ( .B1(n3576), .B2(n4466), .A(n3575), .ZN(U3497) );
  NAND2_X1 U4342 ( .A1(n3604), .A2(n3601), .ZN(n3917) );
  XOR2_X1 U4343 ( .A(n3917), .B(n3577), .Z(n4410) );
  INV_X1 U4344 ( .A(n4410), .ZN(n3586) );
  XOR2_X1 U4345 ( .A(n3917), .B(n3603), .Z(n3578) );
  OAI22_X1 U4346 ( .A1(n3578), .A2(n4182), .B1(n4332), .B2(n4296), .ZN(n4409)
         );
  OAI21_X1 U4347 ( .B1(n3579), .B2(n4404), .A(n3599), .ZN(n4467) );
  NOR2_X1 U4348 ( .A1(n4467), .A2(n4339), .ZN(n3584) );
  AOI22_X1 U4349 ( .A1(n2229), .A2(REG2_REG_17__SCAN_IN), .B1(n3580), .B2(
        n4634), .ZN(n3582) );
  NAND2_X1 U4350 ( .A1(n4313), .A2(n4048), .ZN(n3581) );
  OAI211_X1 U4351 ( .C1(n4307), .C2(n4404), .A(n3582), .B(n3581), .ZN(n3583)
         );
  AOI211_X1 U4352 ( .C1(n4409), .C2(n4507), .A(n3584), .B(n3583), .ZN(n3585)
         );
  OAI21_X1 U4353 ( .B1(n3586), .B2(n4342), .A(n3585), .ZN(U3273) );
  OR2_X1 U4354 ( .A1(n3587), .A2(n4402), .ZN(n3589) );
  NAND2_X1 U4355 ( .A1(n3589), .A2(n3588), .ZN(n3592) );
  MUX2_X1 U4356 ( .A(REG0_REG_16__SCAN_IN), .B(n3592), .S(n4690), .Z(n3590) );
  INV_X1 U4357 ( .A(n3590), .ZN(n3591) );
  OAI21_X1 U4358 ( .B1(n3595), .B2(n4466), .A(n3591), .ZN(U3499) );
  MUX2_X1 U4359 ( .A(REG1_REG_16__SCAN_IN), .B(n3592), .S(n4700), .Z(n3593) );
  INV_X1 U4360 ( .A(n3593), .ZN(n3594) );
  OAI21_X1 U4361 ( .B1(n4412), .B2(n3595), .A(n3594), .ZN(U3534) );
  INV_X1 U4362 ( .A(n3597), .ZN(n3598) );
  AOI21_X1 U4363 ( .B1(n3923), .B2(n3596), .A(n3598), .ZN(n4403) );
  INV_X1 U4364 ( .A(n3599), .ZN(n3600) );
  OAI211_X1 U4365 ( .C1(n3600), .C2(n3844), .A(n4669), .B(n4333), .ZN(n4400)
         );
  INV_X1 U4366 ( .A(n3601), .ZN(n3602) );
  NAND2_X1 U4367 ( .A1(n4231), .A2(n3604), .ZN(n4321) );
  XNOR2_X1 U4368 ( .A(n4321), .B(n3923), .ZN(n3607) );
  AOI22_X1 U4369 ( .A1(n4312), .A2(n4328), .B1(n4327), .B2(n3668), .ZN(n3605)
         );
  OAI21_X1 U4370 ( .B1(n3845), .B2(n4406), .A(n3605), .ZN(n3606) );
  AOI21_X1 U4371 ( .B1(n3607), .B2(n4324), .A(n3606), .ZN(n4401) );
  OAI21_X1 U4372 ( .B1(n4473), .B2(n4400), .A(n4401), .ZN(n3610) );
  INV_X1 U4373 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4093) );
  INV_X1 U4374 ( .A(n3608), .ZN(n3850) );
  OAI22_X1 U4375 ( .A1(n4507), .A2(n4093), .B1(n3850), .B2(n4261), .ZN(n3609)
         );
  AOI21_X1 U4376 ( .B1(n3610), .B2(n4507), .A(n3609), .ZN(n3611) );
  OAI21_X1 U4377 ( .B1(n4403), .B2(n4342), .A(n3611), .ZN(U3272) );
  OAI22_X1 U4378 ( .A1(n3864), .A2(n3733), .B1(n3732), .B2(n3629), .ZN(n3612)
         );
  XNOR2_X1 U4379 ( .A(n3612), .B(n3742), .ZN(n3619) );
  INV_X1 U4380 ( .A(n3619), .ZN(n3617) );
  OR2_X1 U4381 ( .A1(n3864), .A2(n2906), .ZN(n3615) );
  NAND2_X1 U4382 ( .A1(n3613), .A2(n2908), .ZN(n3614) );
  NAND2_X1 U4383 ( .A1(n3615), .A2(n3614), .ZN(n3618) );
  INV_X1 U4384 ( .A(n3618), .ZN(n3616) );
  NAND2_X1 U4385 ( .A1(n3617), .A2(n3616), .ZN(n3644) );
  NAND2_X1 U4386 ( .A1(n3619), .A2(n3618), .ZN(n3642) );
  NAND2_X1 U4387 ( .A1(n3644), .A2(n3642), .ZN(n3626) );
  NAND2_X1 U4388 ( .A1(n3620), .A2(n3621), .ZN(n3625) );
  INV_X1 U4389 ( .A(n3620), .ZN(n3623) );
  INV_X1 U4390 ( .A(n3621), .ZN(n3622) );
  XOR2_X1 U4391 ( .A(n3626), .B(n3643), .Z(n3627) );
  NAND2_X1 U4392 ( .A1(n3627), .A2(n4498), .ZN(n3633) );
  OAI22_X1 U4393 ( .A1(n4491), .A2(n3629), .B1(n3628), .B2(n3863), .ZN(n3631)
         );
  NAND2_X1 U4394 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4579) );
  OAI21_X1 U4395 ( .B1(n3867), .B2(n3646), .A(n4579), .ZN(n3630) );
  NOR2_X1 U4396 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  OAI211_X1 U4397 ( .C1(n4503), .C2(n3634), .A(n3633), .B(n3632), .ZN(U3212)
         );
  INV_X1 U4398 ( .A(n3740), .ZN(n3747) );
  NAND2_X1 U4399 ( .A1(n4180), .A2(n4313), .ZN(n3636) );
  AOI22_X1 U4400 ( .A1(n3752), .A2(n4634), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2229), .ZN(n3635) );
  OAI211_X1 U4401 ( .C1(n4307), .C2(n3747), .A(n3636), .B(n3635), .ZN(n3639)
         );
  NOR2_X1 U4402 ( .A1(n3637), .A2(n2229), .ZN(n3638) );
  AOI211_X1 U4403 ( .C1(n4637), .C2(n2474), .A(n3639), .B(n3638), .ZN(n3640)
         );
  OAI21_X1 U4404 ( .B1(n3641), .B2(n4342), .A(n3640), .ZN(U3262) );
  OAI22_X1 U4405 ( .A1(n3646), .A2(n3733), .B1(n3865), .B2(n3732), .ZN(n3647)
         );
  XOR2_X1 U4406 ( .A(n2947), .B(n3647), .Z(n3651) );
  NAND2_X1 U4407 ( .A1(n4486), .A2(n3741), .ZN(n3650) );
  NAND2_X1 U4408 ( .A1(n3648), .A2(n2908), .ZN(n3649) );
  NAND2_X1 U4409 ( .A1(n3650), .A2(n3649), .ZN(n4495) );
  OAI22_X1 U4410 ( .A1(n4407), .A2(n3733), .B1(n4490), .B2(n3732), .ZN(n3652)
         );
  XNOR2_X1 U4411 ( .A(n3652), .B(n3742), .ZN(n3657) );
  OR2_X1 U4412 ( .A1(n4407), .A2(n2906), .ZN(n3655) );
  NAND2_X1 U4413 ( .A1(n3653), .A2(n2908), .ZN(n3654) );
  NAND2_X1 U4414 ( .A1(n3655), .A2(n3654), .ZN(n3656) );
  NOR2_X1 U4415 ( .A1(n3657), .A2(n3656), .ZN(n3658) );
  AOI21_X1 U4416 ( .B1(n3657), .B2(n3656), .A(n3658), .ZN(n4496) );
  OAI22_X1 U4417 ( .A1(n3845), .A2(n3733), .B1(n4404), .B2(n3732), .ZN(n3659)
         );
  XNOR2_X1 U4418 ( .A(n3659), .B(n3742), .ZN(n3662) );
  OR2_X1 U4419 ( .A1(n3845), .A2(n2906), .ZN(n3661) );
  OR2_X1 U4420 ( .A1(n4404), .A2(n3733), .ZN(n3660) );
  NAND2_X1 U4421 ( .A1(n3661), .A2(n3660), .ZN(n3663) );
  NAND2_X1 U4422 ( .A1(n3662), .A2(n3663), .ZN(n3799) );
  NAND2_X1 U4423 ( .A1(n3800), .A2(n3799), .ZN(n3666) );
  INV_X1 U4424 ( .A(n3662), .ZN(n3665) );
  INV_X1 U4425 ( .A(n3663), .ZN(n3664) );
  NAND2_X1 U4426 ( .A1(n3665), .A2(n3664), .ZN(n3798) );
  OAI22_X1 U4427 ( .A1(n4332), .A2(n3733), .B1(n3844), .B2(n3732), .ZN(n3667)
         );
  XNOR2_X1 U4428 ( .A(n3667), .B(n3742), .ZN(n3671) );
  OR2_X1 U4429 ( .A1(n4332), .A2(n2906), .ZN(n3670) );
  NAND2_X1 U4430 ( .A1(n3668), .A2(n2908), .ZN(n3669) );
  NAND2_X1 U4431 ( .A1(n3670), .A2(n3669), .ZN(n3672) );
  NAND2_X1 U4432 ( .A1(n3671), .A2(n3672), .ZN(n3841) );
  INV_X1 U4433 ( .A(n3671), .ZN(n3674) );
  INV_X1 U4434 ( .A(n3672), .ZN(n3673) );
  NAND2_X1 U4435 ( .A1(n3674), .A2(n3673), .ZN(n3840) );
  NAND2_X1 U4436 ( .A1(n4312), .A2(n2908), .ZN(n3676) );
  NAND2_X1 U4437 ( .A1(n4326), .A2(n3739), .ZN(n3675) );
  NAND2_X1 U4438 ( .A1(n3676), .A2(n3675), .ZN(n3677) );
  XNOR2_X1 U4439 ( .A(n3677), .B(n3742), .ZN(n3678) );
  AOI22_X1 U4440 ( .A1(n4312), .A2(n3741), .B1(n2908), .B2(n4326), .ZN(n3679)
         );
  XNOR2_X1 U4441 ( .A(n3678), .B(n3679), .ZN(n3769) );
  INV_X1 U4442 ( .A(n3678), .ZN(n3680) );
  NAND2_X1 U4443 ( .A1(n4329), .A2(n2908), .ZN(n3684) );
  NAND2_X1 U4444 ( .A1(n3686), .A2(n3739), .ZN(n3683) );
  NAND2_X1 U4445 ( .A1(n3684), .A2(n3683), .ZN(n3685) );
  XNOR2_X1 U4446 ( .A(n3685), .B(n3467), .ZN(n3695) );
  INV_X1 U4447 ( .A(n3695), .ZN(n3689) );
  AND2_X1 U4448 ( .A1(n3686), .A2(n2908), .ZN(n3687) );
  AOI21_X1 U4449 ( .B1(n4329), .B2(n3741), .A(n3687), .ZN(n3694) );
  INV_X1 U4450 ( .A(n3694), .ZN(n3688) );
  NAND2_X1 U4451 ( .A1(n3689), .A2(n3688), .ZN(n3820) );
  OAI22_X1 U4452 ( .A1(n4297), .A2(n3733), .B1(n4384), .B2(n3732), .ZN(n3690)
         );
  XNOR2_X1 U4453 ( .A(n3690), .B(n3742), .ZN(n3780) );
  OR2_X1 U4454 ( .A1(n4297), .A2(n2906), .ZN(n3693) );
  NAND2_X1 U4455 ( .A1(n3691), .A2(n2908), .ZN(n3692) );
  NAND2_X1 U4456 ( .A1(n3693), .A2(n3692), .ZN(n3779) );
  NAND2_X1 U4457 ( .A1(n3695), .A2(n3694), .ZN(n3819) );
  OAI21_X1 U4458 ( .B1(n3780), .B2(n3779), .A(n3819), .ZN(n3696) );
  INV_X1 U4459 ( .A(n3780), .ZN(n3698) );
  INV_X1 U4460 ( .A(n3779), .ZN(n3697) );
  NOR2_X1 U4461 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  AOI22_X1 U4462 ( .A1(n4280), .A2(n2908), .B1(n4258), .B2(n3739), .ZN(n3701)
         );
  XNOR2_X1 U4463 ( .A(n3701), .B(n3742), .ZN(n3703) );
  AOI22_X1 U4464 ( .A1(n4280), .A2(n3741), .B1(n4258), .B2(n2908), .ZN(n3704)
         );
  XNOR2_X1 U4465 ( .A(n3703), .B(n3704), .ZN(n3830) );
  INV_X1 U4466 ( .A(n3703), .ZN(n3706) );
  INV_X1 U4467 ( .A(n3704), .ZN(n3705) );
  NOR2_X1 U4468 ( .A1(n3706), .A2(n3705), .ZN(n3763) );
  NAND2_X1 U4469 ( .A1(n4267), .A2(n2908), .ZN(n3708) );
  OR2_X1 U4470 ( .A1(n4247), .A2(n3732), .ZN(n3707) );
  NAND2_X1 U4471 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  XNOR2_X1 U4472 ( .A(n3709), .B(n3467), .ZN(n3713) );
  NOR2_X1 U4473 ( .A1(n4247), .A2(n3733), .ZN(n3710) );
  AOI21_X1 U4474 ( .B1(n4267), .B2(n3741), .A(n3710), .ZN(n3712) );
  XNOR2_X1 U4475 ( .A(n3713), .B(n3712), .ZN(n3762) );
  NOR2_X1 U4476 ( .A1(n3763), .A2(n3762), .ZN(n3711) );
  NOR2_X1 U4477 ( .A1(n3713), .A2(n3712), .ZN(n3715) );
  OAI22_X1 U4478 ( .A1(n4244), .A2(n2906), .B1(n4368), .B2(n3733), .ZN(n3717)
         );
  OAI22_X1 U4479 ( .A1(n4244), .A2(n3733), .B1(n4368), .B2(n3732), .ZN(n3714)
         );
  XNOR2_X1 U4480 ( .A(n3714), .B(n3742), .ZN(n3812) );
  NAND2_X1 U4481 ( .A1(n3809), .A2(n3812), .ZN(n3719) );
  INV_X1 U4482 ( .A(n3715), .ZN(n3716) );
  NAND2_X1 U4483 ( .A1(n2466), .A2(n3716), .ZN(n3718) );
  NAND2_X1 U4484 ( .A1(n3718), .A2(n3717), .ZN(n3810) );
  NAND2_X1 U4485 ( .A1(n3719), .A2(n3810), .ZN(n3792) );
  NOR2_X1 U4486 ( .A1(n4200), .A2(n3732), .ZN(n3720) );
  AOI21_X1 U4487 ( .B1(n4215), .B2(n2908), .A(n3720), .ZN(n3721) );
  XNOR2_X1 U4488 ( .A(n3721), .B(n3742), .ZN(n3724) );
  NOR2_X1 U4489 ( .A1(n4200), .A2(n3733), .ZN(n3722) );
  AOI21_X1 U4490 ( .B1(n4215), .B2(n3741), .A(n3722), .ZN(n3723) );
  NAND2_X1 U4491 ( .A1(n3724), .A2(n3723), .ZN(n3790) );
  OR2_X1 U4492 ( .A1(n3724), .A2(n3723), .ZN(n3791) );
  NAND2_X1 U4493 ( .A1(n4197), .A2(n2908), .ZN(n3727) );
  OR2_X1 U4494 ( .A1(n4186), .A2(n3732), .ZN(n3726) );
  NAND2_X1 U4495 ( .A1(n3727), .A2(n3726), .ZN(n3728) );
  XNOR2_X1 U4496 ( .A(n3728), .B(n3467), .ZN(n3731) );
  NOR2_X1 U4497 ( .A1(n4186), .A2(n3733), .ZN(n3729) );
  AOI21_X1 U4498 ( .B1(n4197), .B2(n3741), .A(n3729), .ZN(n3730) );
  NOR2_X1 U4499 ( .A1(n3731), .A2(n3730), .ZN(n3851) );
  OAI22_X1 U4500 ( .A1(n3748), .A2(n3733), .B1(n3732), .B2(n4355), .ZN(n3734)
         );
  XNOR2_X1 U4501 ( .A(n3734), .B(n3742), .ZN(n3736) );
  OAI22_X1 U4502 ( .A1(n3748), .A2(n2906), .B1(n3733), .B2(n4355), .ZN(n3735)
         );
  XNOR2_X1 U4503 ( .A(n3736), .B(n3735), .ZN(n3755) );
  INV_X1 U4504 ( .A(n3735), .ZN(n3738) );
  INV_X1 U4505 ( .A(n3736), .ZN(n3737) );
  AOI22_X1 U4506 ( .A1(n4149), .A2(n2908), .B1(n3740), .B2(n3739), .ZN(n3745)
         );
  AOI22_X1 U4507 ( .A1(n4149), .A2(n3741), .B1(n3740), .B2(n2908), .ZN(n3743)
         );
  XNOR2_X1 U4508 ( .A(n3743), .B(n3742), .ZN(n3744) );
  XOR2_X1 U4509 ( .A(n3745), .B(n3744), .Z(n3746) );
  OAI22_X1 U4510 ( .A1(n4491), .A2(n3747), .B1(STATE_REG_SCAN_IN), .B2(n4780), 
        .ZN(n3751) );
  INV_X1 U4511 ( .A(n4044), .ZN(n3749) );
  OAI22_X1 U4512 ( .A1(n3749), .A2(n3867), .B1(n3748), .B2(n3863), .ZN(n3750)
         );
  AOI211_X1 U4513 ( .C1(n3752), .C2(n3834), .A(n3751), .B(n3750), .ZN(n3753)
         );
  OAI21_X1 U4514 ( .B1(n3754), .B2(n3858), .A(n3753), .ZN(U3217) );
  AOI22_X1 U4515 ( .A1(n4197), .A2(n4487), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3758) );
  NAND2_X1 U4516 ( .A1(n3756), .A2(n4162), .ZN(n3757) );
  OAI211_X1 U4517 ( .C1(n4160), .C2(n3867), .A(n3758), .B(n3757), .ZN(n3759)
         );
  AOI21_X1 U4518 ( .B1(n4165), .B2(n3834), .A(n3759), .ZN(n3760) );
  OAI21_X1 U4519 ( .B1(n3761), .B2(n3858), .A(n3760), .ZN(U3211) );
  OAI21_X1 U4520 ( .B1(n2234), .B2(n3763), .A(n3762), .ZN(n3764) );
  NAND3_X1 U4521 ( .A1(n2466), .A2(n3764), .A3(n4498), .ZN(n3768) );
  INV_X1 U4522 ( .A(n4280), .ZN(n3784) );
  NOR2_X1 U4523 ( .A1(n3784), .A2(n3863), .ZN(n3766) );
  OAI22_X1 U4524 ( .A1(n4244), .A2(n3867), .B1(n4491), .B2(n4247), .ZN(n3765)
         );
  AOI211_X1 U4525 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3766), .B(n3765), .ZN(n3767) );
  OAI211_X1 U4526 ( .C1(n4503), .C2(n4249), .A(n3768), .B(n3767), .ZN(U3213)
         );
  INV_X1 U4527 ( .A(n4337), .ZN(n3777) );
  XNOR2_X1 U4528 ( .A(n3770), .B(n3769), .ZN(n3771) );
  NAND2_X1 U4529 ( .A1(n3771), .A2(n4498), .ZN(n3776) );
  OAI22_X1 U4530 ( .A1(n4491), .A2(n4335), .B1(n4385), .B2(n3867), .ZN(n3774)
         );
  AND2_X1 U4531 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4131) );
  INV_X1 U4532 ( .A(n4131), .ZN(n3772) );
  OAI21_X1 U4533 ( .B1(n3863), .B2(n4332), .A(n3772), .ZN(n3773) );
  NOR2_X1 U4534 ( .A1(n3774), .A2(n3773), .ZN(n3775) );
  OAI211_X1 U4535 ( .C1(n4503), .C2(n3777), .A(n3776), .B(n3775), .ZN(U3216)
         );
  INV_X1 U4536 ( .A(n4284), .ZN(n3789) );
  INV_X1 U4537 ( .A(n3819), .ZN(n3778) );
  OAI21_X1 U4538 ( .B1(n3821), .B2(n3778), .A(n3820), .ZN(n3782) );
  XNOR2_X1 U4539 ( .A(n3780), .B(n3779), .ZN(n3781) );
  XNOR2_X1 U4540 ( .A(n3782), .B(n3781), .ZN(n3783) );
  NAND2_X1 U4541 ( .A1(n3783), .A2(n4498), .ZN(n3788) );
  OAI22_X1 U4542 ( .A1(n4491), .A2(n4384), .B1(n3784), .B2(n3867), .ZN(n3786)
         );
  OAI22_X1 U4543 ( .A1(n3863), .A2(n4385), .B1(STATE_REG_SCAN_IN), .B2(n4983), 
        .ZN(n3785) );
  NOR2_X1 U4544 ( .A1(n3786), .A2(n3785), .ZN(n3787) );
  OAI211_X1 U4545 ( .C1(n4503), .C2(n3789), .A(n3788), .B(n3787), .ZN(U3220)
         );
  NAND2_X1 U4546 ( .A1(n3791), .A2(n3790), .ZN(n3793) );
  XOR2_X1 U4547 ( .A(n3793), .B(n3792), .Z(n3797) );
  OAI22_X1 U4548 ( .A1(n4244), .A2(n3863), .B1(STATE_REG_SCAN_IN), .B2(n4955), 
        .ZN(n3795) );
  OAI22_X1 U4549 ( .A1(n5076), .A2(n3867), .B1(n4491), .B2(n4200), .ZN(n3794)
         );
  AOI211_X1 U4550 ( .C1(n4203), .C2(n3834), .A(n3795), .B(n3794), .ZN(n3796)
         );
  OAI21_X1 U4551 ( .B1(n3797), .B2(n3858), .A(n3796), .ZN(U3222) );
  NAND2_X1 U4552 ( .A1(n3799), .A2(n3798), .ZN(n3801) );
  XOR2_X1 U4553 ( .A(n3801), .B(n3800), .Z(n3802) );
  NAND2_X1 U4554 ( .A1(n3802), .A2(n4498), .ZN(n3807) );
  OAI22_X1 U4555 ( .A1(n4491), .A2(n4404), .B1(n4332), .B2(n3867), .ZN(n3805)
         );
  INV_X1 U4556 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U4557 ( .A1(STATE_REG_SCAN_IN), .A2(n4972), .ZN(n4611) );
  INV_X1 U4558 ( .A(n4611), .ZN(n3803) );
  OAI21_X1 U4559 ( .B1(n3863), .B2(n4407), .A(n3803), .ZN(n3804) );
  NOR2_X1 U4560 ( .A1(n3805), .A2(n3804), .ZN(n3806) );
  OAI211_X1 U4561 ( .C1(n4503), .C2(n3808), .A(n3807), .B(n3806), .ZN(U3225)
         );
  NAND2_X1 U4562 ( .A1(n3810), .A2(n3809), .ZN(n3811) );
  XOR2_X1 U4563 ( .A(n3812), .B(n3811), .Z(n3818) );
  INV_X1 U4564 ( .A(n4220), .ZN(n3816) );
  OAI22_X1 U4565 ( .A1(n4369), .A2(n3863), .B1(STATE_REG_SCAN_IN), .B2(n3813), 
        .ZN(n3815) );
  OAI22_X1 U4566 ( .A1(n4178), .A2(n3867), .B1(n4491), .B2(n4368), .ZN(n3814)
         );
  AOI211_X1 U4567 ( .C1(n3816), .C2(n3834), .A(n3815), .B(n3814), .ZN(n3817)
         );
  OAI21_X1 U4568 ( .B1(n3818), .B2(n3858), .A(n3817), .ZN(U3226) );
  INV_X1 U4569 ( .A(n4305), .ZN(n3829) );
  NAND2_X1 U4570 ( .A1(n3820), .A2(n3819), .ZN(n3822) );
  XOR2_X1 U4571 ( .A(n3822), .B(n3821), .Z(n3823) );
  NAND2_X1 U4572 ( .A1(n3823), .A2(n4498), .ZN(n3828) );
  OAI22_X1 U4573 ( .A1(n4491), .A2(n4391), .B1(n4297), .B2(n3867), .ZN(n3826)
         );
  INV_X1 U4574 ( .A(n4312), .ZN(n4392) );
  OAI22_X1 U4575 ( .A1(n3863), .A2(n4392), .B1(STATE_REG_SCAN_IN), .B2(n3824), 
        .ZN(n3825) );
  NOR2_X1 U4576 ( .A1(n3826), .A2(n3825), .ZN(n3827) );
  OAI211_X1 U4577 ( .C1(n4503), .C2(n3829), .A(n3828), .B(n3827), .ZN(U3230)
         );
  AOI21_X1 U4578 ( .B1(n3830), .B2(n2254), .A(n2234), .ZN(n3837) );
  INV_X1 U4579 ( .A(n4262), .ZN(n3835) );
  INV_X1 U4580 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3831) );
  OAI22_X1 U4581 ( .A1(n3863), .A2(n4297), .B1(STATE_REG_SCAN_IN), .B2(n3831), 
        .ZN(n3833) );
  OAI22_X1 U4582 ( .A1(n4491), .A2(n4270), .B1(n4369), .B2(n3867), .ZN(n3832)
         );
  AOI211_X1 U4583 ( .C1(n3835), .C2(n3834), .A(n3833), .B(n3832), .ZN(n3836)
         );
  OAI21_X1 U4584 ( .B1(n3837), .B2(n3858), .A(n3836), .ZN(U3232) );
  NOR2_X1 U4585 ( .A1(n3838), .A2(n2416), .ZN(n3843) );
  AOI21_X1 U4586 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n3842) );
  OAI21_X1 U4587 ( .B1(n3843), .B2(n3842), .A(n4498), .ZN(n3849) );
  OAI22_X1 U4588 ( .A1(n4491), .A2(n3844), .B1(n4392), .B2(n3867), .ZN(n3847)
         );
  INV_X1 U4589 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4904) );
  OAI22_X1 U4590 ( .A1(n3863), .A2(n3845), .B1(STATE_REG_SCAN_IN), .B2(n4904), 
        .ZN(n3846) );
  NOR2_X1 U4591 ( .A1(n3847), .A2(n3846), .ZN(n3848) );
  OAI211_X1 U4592 ( .C1(n4503), .C2(n3850), .A(n3849), .B(n3848), .ZN(U3235)
         );
  NOR2_X1 U4593 ( .A1(n3851), .A2(n2260), .ZN(n3852) );
  XNOR2_X1 U4594 ( .A(n3853), .B(n3852), .ZN(n3859) );
  NOR2_X1 U4595 ( .A1(n4503), .A2(n4185), .ZN(n3856) );
  AOI22_X1 U4596 ( .A1(n4215), .A2(n4487), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3854) );
  OAI21_X1 U4597 ( .B1(n4491), .B2(n4186), .A(n3854), .ZN(n3855) );
  AOI211_X1 U4598 ( .C1(n4180), .C2(n4485), .A(n3856), .B(n3855), .ZN(n3857)
         );
  OAI21_X1 U4599 ( .B1(n3859), .B2(n3858), .A(n3857), .ZN(U3237) );
  INV_X1 U4600 ( .A(n3860), .ZN(n3872) );
  NAND2_X1 U4601 ( .A1(n4493), .A2(n4494), .ZN(n3861) );
  XNOR2_X1 U4602 ( .A(n3861), .B(n4495), .ZN(n3862) );
  NAND2_X1 U4603 ( .A1(n3862), .A2(n4498), .ZN(n3871) );
  OAI22_X1 U4604 ( .A1(n4491), .A2(n3865), .B1(n3864), .B2(n3863), .ZN(n3869)
         );
  NOR2_X1 U4605 ( .A1(STATE_REG_SCAN_IN), .A2(n2678), .ZN(n4591) );
  INV_X1 U4606 ( .A(n4591), .ZN(n3866) );
  OAI21_X1 U4607 ( .B1(n3867), .B2(n4407), .A(n3866), .ZN(n3868) );
  NOR2_X1 U4608 ( .A1(n3869), .A2(n3868), .ZN(n3870) );
  OAI211_X1 U4609 ( .C1(n4503), .C2(n3872), .A(n3871), .B(n3870), .ZN(U3238)
         );
  NAND2_X1 U4610 ( .A1(n2546), .A2(DATAI_31_), .ZN(n4139) );
  INV_X1 U4611 ( .A(n4139), .ZN(n4142) );
  NAND2_X1 U4612 ( .A1(n2546), .A2(DATAI_30_), .ZN(n4351) );
  AND2_X1 U4613 ( .A1(n4043), .A2(n4351), .ZN(n3911) );
  INV_X1 U4614 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4143) );
  NAND2_X1 U4615 ( .A1(n3873), .A2(REG1_REG_31__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4616 ( .A1(n2766), .A2(REG0_REG_31__SCAN_IN), .ZN(n3874) );
  OAI211_X1 U4617 ( .C1(n3876), .C2(n4143), .A(n3875), .B(n3874), .ZN(n4042)
         );
  NOR2_X1 U4618 ( .A1(n4042), .A2(n4139), .ZN(n3910) );
  INV_X1 U4619 ( .A(n3877), .ZN(n3907) );
  AND2_X1 U4620 ( .A1(n3929), .A2(n3907), .ZN(n4015) );
  INV_X1 U4621 ( .A(n4015), .ZN(n3892) );
  NAND2_X1 U4622 ( .A1(n3878), .A2(n3881), .ZN(n3997) );
  NAND2_X1 U4623 ( .A1(n3880), .A2(n3879), .ZN(n3987) );
  NAND2_X1 U4624 ( .A1(n3987), .A2(n3881), .ZN(n3996) );
  OAI21_X1 U4625 ( .B1(n3882), .B2(n3997), .A(n3996), .ZN(n3884) );
  INV_X1 U4626 ( .A(n3883), .ZN(n3999) );
  AOI21_X1 U4627 ( .B1(n3884), .B2(n4002), .A(n3999), .ZN(n3887) );
  INV_X1 U4628 ( .A(n4233), .ZN(n3886) );
  OAI21_X1 U4629 ( .B1(n3887), .B2(n3886), .A(n3885), .ZN(n3888) );
  INV_X1 U4630 ( .A(n3888), .ZN(n3890) );
  OAI21_X1 U4631 ( .B1(n3890), .B2(n4009), .A(n3889), .ZN(n3891) );
  OAI221_X1 U4632 ( .B1(n3892), .B2(n4011), .C1(n3892), .C2(n3891), .A(n4019), 
        .ZN(n3894) );
  NAND2_X1 U4633 ( .A1(n4042), .A2(n4139), .ZN(n4023) );
  OAI21_X1 U4634 ( .B1(n4043), .B2(n4351), .A(n4023), .ZN(n3914) );
  INV_X1 U4635 ( .A(n3914), .ZN(n3893) );
  OAI21_X1 U4636 ( .B1(n4044), .B2(n4147), .A(n3893), .ZN(n3899) );
  OR4_X1 U4637 ( .A1(n3894), .A2(n3898), .A3(n3897), .A4(n3899), .ZN(n3904) );
  AOI21_X1 U4638 ( .B1(n4044), .B2(n4147), .A(n3895), .ZN(n3900) );
  NAND2_X1 U4639 ( .A1(n3900), .A2(n3896), .ZN(n4016) );
  INV_X1 U4640 ( .A(n4159), .ZN(n3902) );
  OR2_X1 U4641 ( .A1(n3898), .A2(n3897), .ZN(n3901) );
  AOI21_X1 U4642 ( .B1(n3901), .B2(n3900), .A(n3899), .ZN(n4020) );
  OAI21_X1 U4643 ( .B1(n4016), .B2(n3902), .A(n4020), .ZN(n3903) );
  INV_X1 U4644 ( .A(n4042), .ZN(n4141) );
  INV_X1 U4645 ( .A(n4351), .ZN(n4348) );
  AOI22_X1 U4646 ( .A1(n3904), .A2(n3903), .B1(n4141), .B2(n4348), .ZN(n3905)
         );
  AOI211_X1 U4647 ( .C1(n4142), .C2(n3911), .A(n3910), .B(n3905), .ZN(n4031)
         );
  NAND2_X1 U4648 ( .A1(n3907), .A2(n3906), .ZN(n4211) );
  AND2_X1 U4649 ( .A1(n3909), .A2(n3908), .ZN(n4303) );
  INV_X1 U4650 ( .A(n3910), .ZN(n3913) );
  INV_X1 U4651 ( .A(n3911), .ZN(n3912) );
  NAND2_X1 U4652 ( .A1(n3913), .A2(n3912), .ZN(n4024) );
  NOR2_X1 U4653 ( .A1(n3914), .A2(n4024), .ZN(n3915) );
  NAND2_X1 U4654 ( .A1(n3916), .A2(n3915), .ZN(n3918) );
  NOR4_X1 U4655 ( .A1(n4211), .A2(n4303), .A3(n3918), .A4(n3917), .ZN(n3928)
         );
  NOR4_X1 U4656 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3927)
         );
  NOR4_X1 U4657 ( .A1(n2724), .A2(n2785), .A3(n3925), .A4(n3924), .ZN(n3926)
         );
  NAND3_X1 U4658 ( .A1(n3928), .A2(n3927), .A3(n3926), .ZN(n3947) );
  XNOR2_X1 U4659 ( .A(n4312), .B(n4326), .ZN(n4323) );
  INV_X1 U4660 ( .A(n3929), .ZN(n3930) );
  OR2_X1 U4661 ( .A1(n3930), .A2(n4173), .ZN(n4192) );
  XNOR2_X1 U4662 ( .A(n4267), .B(n4247), .ZN(n4236) );
  NOR4_X1 U4663 ( .A1(n4192), .A2(n3932), .A3(n3931), .A4(n4236), .ZN(n3933)
         );
  NAND4_X1 U4664 ( .A1(n4159), .A2(n4323), .A3(n3934), .A4(n3933), .ZN(n3946)
         );
  NOR2_X1 U4665 ( .A1(n3936), .A2(n3935), .ZN(n4177) );
  INV_X1 U4666 ( .A(n3937), .ZN(n4234) );
  NOR4_X1 U4667 ( .A1(n4275), .A2(n3939), .A3(n2783), .A4(n3938), .ZN(n3944)
         );
  NOR4_X1 U4668 ( .A1(n4265), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3943)
         );
  NAND3_X1 U4669 ( .A1(n4177), .A2(n3944), .A3(n3943), .ZN(n3945) );
  OR4_X1 U4670 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3951) );
  OAI21_X1 U4671 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n4028) );
  INV_X1 U4672 ( .A(n3952), .ZN(n3956) );
  OAI211_X1 U4673 ( .C1(n3956), .C2(n3955), .A(n3954), .B(n3953), .ZN(n3959)
         );
  NAND3_X1 U4674 ( .A1(n3959), .A2(n3958), .A3(n3957), .ZN(n3962) );
  NAND3_X1 U4675 ( .A1(n3962), .A2(n3961), .A3(n3960), .ZN(n3965) );
  NAND3_X1 U4676 ( .A1(n3965), .A2(n3964), .A3(n3963), .ZN(n3968) );
  NAND4_X1 U4677 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3979), .ZN(n3971)
         );
  NAND3_X1 U4678 ( .A1(n3971), .A2(n3970), .A3(n3969), .ZN(n3978) );
  AND2_X1 U4679 ( .A1(n3973), .A2(n3972), .ZN(n3980) );
  INV_X1 U4680 ( .A(n3974), .ZN(n3977) );
  INV_X1 U4681 ( .A(n3975), .ZN(n3976) );
  AOI211_X1 U4682 ( .C1(n3978), .C2(n3980), .A(n3977), .B(n3976), .ZN(n3988)
         );
  INV_X1 U4683 ( .A(n3979), .ZN(n3983) );
  INV_X1 U4684 ( .A(n3980), .ZN(n3982) );
  NOR3_X1 U4685 ( .A1(n3983), .A2(n3982), .A3(n3981), .ZN(n3985) );
  INV_X1 U4686 ( .A(n3990), .ZN(n3984) );
  OAI21_X1 U4687 ( .B1(n3985), .B2(n3984), .A(n3996), .ZN(n3986) );
  OAI21_X1 U4688 ( .B1(n3988), .B2(n3987), .A(n3986), .ZN(n3994) );
  NAND2_X1 U4689 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  NAND4_X1 U4690 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n4001)
         );
  INV_X1 U4691 ( .A(n3995), .ZN(n3998) );
  OAI21_X1 U4692 ( .B1(n3998), .B2(n3997), .A(n3996), .ZN(n4000) );
  AOI21_X1 U4693 ( .B1(n4001), .B2(n4000), .A(n3999), .ZN(n4006) );
  INV_X1 U4694 ( .A(n4002), .ZN(n4005) );
  INV_X1 U4695 ( .A(n4003), .ZN(n4004) );
  OAI21_X1 U4696 ( .B1(n4006), .B2(n4005), .A(n4004), .ZN(n4008) );
  AOI211_X1 U4697 ( .C1(n4008), .C2(n4233), .A(n4007), .B(n4232), .ZN(n4010)
         );
  NOR2_X1 U4698 ( .A1(n4010), .A2(n4009), .ZN(n4013) );
  OAI21_X1 U4699 ( .B1(n4013), .B2(n4012), .A(n4011), .ZN(n4014) );
  NAND2_X1 U4700 ( .A1(n4015), .A2(n4014), .ZN(n4018) );
  AOI211_X1 U4701 ( .C1(n4019), .C2(n4018), .A(n4017), .B(n4016), .ZN(n4022)
         );
  INV_X1 U4702 ( .A(n4020), .ZN(n4021) );
  NOR2_X1 U4703 ( .A1(n4022), .A2(n4021), .ZN(n4025) );
  OAI21_X1 U4704 ( .B1(n4025), .B2(n4024), .A(n4023), .ZN(n4027) );
  MUX2_X1 U4705 ( .A(n4028), .B(n4027), .S(n4026), .Z(n4029) );
  OAI21_X1 U4706 ( .B1(n4031), .B2(n4030), .A(n4029), .ZN(n4032) );
  XNOR2_X1 U4707 ( .A(n4032), .B(n4133), .ZN(n4041) );
  INV_X1 U4708 ( .A(n4033), .ZN(n4038) );
  AOI21_X1 U4709 ( .B1(n4035), .B2(n4034), .A(n4967), .ZN(n4036) );
  OAI21_X1 U4710 ( .B1(n4038), .B2(n4037), .A(n4036), .ZN(n4039) );
  OAI21_X1 U4711 ( .B1(n4041), .B2(n4040), .A(n4039), .ZN(U3239) );
  MUX2_X1 U4712 ( .A(n4042), .B(DATAO_REG_31__SCAN_IN), .S(n4057), .Z(U3581)
         );
  MUX2_X1 U4713 ( .A(n4043), .B(DATAO_REG_30__SCAN_IN), .S(n4057), .Z(U3580)
         );
  MUX2_X1 U4714 ( .A(n4044), .B(DATAO_REG_29__SCAN_IN), .S(n4057), .Z(U3579)
         );
  MUX2_X1 U4715 ( .A(DATAO_REG_28__SCAN_IN), .B(n4149), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4716 ( .A(n4180), .B(DATAO_REG_27__SCAN_IN), .S(n4057), .Z(U3577)
         );
  MUX2_X1 U4717 ( .A(n4215), .B(DATAO_REG_25__SCAN_IN), .S(n4057), .Z(U3575)
         );
  MUX2_X1 U4718 ( .A(n4045), .B(DATAO_REG_24__SCAN_IN), .S(n4057), .Z(U3574)
         );
  MUX2_X1 U4719 ( .A(n4267), .B(DATAO_REG_23__SCAN_IN), .S(n4057), .Z(U3573)
         );
  MUX2_X1 U4720 ( .A(n4280), .B(DATAO_REG_22__SCAN_IN), .S(n4057), .Z(U3572)
         );
  MUX2_X1 U4721 ( .A(DATAO_REG_21__SCAN_IN), .B(n4046), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4722 ( .A(n4312), .B(DATAO_REG_19__SCAN_IN), .S(n4057), .Z(U3569)
         );
  MUX2_X1 U4723 ( .A(DATAO_REG_18__SCAN_IN), .B(n4047), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4724 ( .A(DATAO_REG_17__SCAN_IN), .B(n4484), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4725 ( .A(DATAO_REG_16__SCAN_IN), .B(n4048), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4726 ( .A(n4486), .B(DATAO_REG_15__SCAN_IN), .S(n4057), .Z(U3565)
         );
  MUX2_X1 U4727 ( .A(DATAO_REG_14__SCAN_IN), .B(n4049), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4728 ( .A(n4050), .B(DATAO_REG_10__SCAN_IN), .S(n4057), .Z(U3560)
         );
  MUX2_X1 U4729 ( .A(n4051), .B(DATAO_REG_9__SCAN_IN), .S(n4057), .Z(U3559) );
  MUX2_X1 U4730 ( .A(n4052), .B(DATAO_REG_6__SCAN_IN), .S(n4057), .Z(U3556) );
  MUX2_X1 U4731 ( .A(n4053), .B(DATAO_REG_5__SCAN_IN), .S(n4057), .Z(U3555) );
  MUX2_X1 U4732 ( .A(DATAO_REG_4__SCAN_IN), .B(n4054), .S(U4043), .Z(U3554) );
  MUX2_X1 U4733 ( .A(n2228), .B(DATAO_REG_3__SCAN_IN), .S(n4057), .Z(U3553) );
  MUX2_X1 U4734 ( .A(DATAO_REG_2__SCAN_IN), .B(n4056), .S(U4043), .Z(U3552) );
  MUX2_X1 U4735 ( .A(DATAO_REG_1__SCAN_IN), .B(n2547), .S(U4043), .Z(U3551) );
  MUX2_X1 U4736 ( .A(n4058), .B(DATAO_REG_0__SCAN_IN), .S(n4057), .Z(U3550) );
  NAND2_X1 U4737 ( .A1(n4059), .A2(n2230), .ZN(n4070) );
  AOI22_X1 U4738 ( .A1(n4612), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4069) );
  INV_X1 U4739 ( .A(n4060), .ZN(n4063) );
  OAI211_X1 U4740 ( .C1(n4063), .C2(n4062), .A(n4568), .B(n4061), .ZN(n4068)
         );
  OAI211_X1 U4741 ( .C1(n4066), .C2(n4065), .A(n4613), .B(n4064), .ZN(n4067)
         );
  NAND4_X1 U4742 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(U3241)
         );
  XOR2_X1 U4743 ( .A(REG1_REG_18__SCAN_IN), .B(n4474), .Z(n4123) );
  NOR2_X1 U4744 ( .A1(n4119), .A2(REG1_REG_17__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U4745 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4115), .ZN(n4086) );
  INV_X1 U4746 ( .A(n4115), .ZN(n4650) );
  AOI22_X1 U4747 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4115), .B1(n4650), .B2(
        n3571), .ZN(n4594) );
  NAND2_X1 U4748 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4111), .ZN(n4083) );
  INV_X1 U4749 ( .A(n4111), .ZN(n4653) );
  AOI22_X1 U4750 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4111), .B1(n4653), .B2(
        n3496), .ZN(n4576) );
  INV_X1 U4751 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U4752 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4097), .B1(n4655), .B2(
        n4698), .ZN(n4547) );
  NAND2_X1 U4753 ( .A1(n4098), .A2(REG1_REG_9__SCAN_IN), .ZN(n4078) );
  INV_X1 U4754 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4071) );
  INV_X1 U4755 ( .A(n4098), .ZN(n4657) );
  AOI22_X1 U4756 ( .A1(n4098), .A2(REG1_REG_9__SCAN_IN), .B1(n4071), .B2(n4657), .ZN(n4526) );
  INV_X1 U4757 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4074) );
  OAI21_X1 U4758 ( .B1(n4075), .B2(n4074), .A(n4073), .ZN(n4076) );
  NAND2_X1 U4759 ( .A1(n4514), .A2(n4076), .ZN(n4077) );
  NAND2_X1 U4760 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U4761 ( .A1(n4535), .A2(n4079), .ZN(n4080) );
  NAND2_X1 U4762 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U4763 ( .A1(n4080), .A2(n4541), .ZN(n4546) );
  NAND2_X1 U4764 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U4765 ( .A1(n4556), .A2(n4081), .ZN(n4082) );
  NAND2_X1 U4766 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4563), .ZN(n4562) );
  NAND2_X1 U4767 ( .A1(n4096), .A2(n4084), .ZN(n4085) );
  NAND2_X1 U4768 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U4769 ( .A1(n4085), .A2(n4584), .ZN(n4593) );
  NOR2_X1 U4770 ( .A1(n4116), .A2(n4087), .ZN(n4088) );
  INV_X1 U4771 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U4772 ( .A1(n4119), .A2(n4828), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4646), .ZN(n4614) );
  INV_X1 U4773 ( .A(n4474), .ZN(n4092) );
  NOR2_X1 U4774 ( .A1(STATE_REG_SCAN_IN), .A2(n4904), .ZN(n4090) );
  AOI21_X1 U4775 ( .B1(n4612), .B2(ADDR_REG_18__SCAN_IN), .A(n4090), .ZN(n4091) );
  OAI21_X1 U4776 ( .B1(n4619), .B2(n4092), .A(n4091), .ZN(n4122) );
  NOR2_X1 U4777 ( .A1(n4474), .A2(n4093), .ZN(n4094) );
  AOI21_X1 U4778 ( .B1(n4474), .B2(n4093), .A(n4094), .ZN(n4121) );
  NOR2_X1 U4779 ( .A1(n4119), .A2(REG2_REG_17__SCAN_IN), .ZN(n4095) );
  AOI21_X1 U4780 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4119), .A(n4095), .ZN(n4609) );
  INV_X1 U4781 ( .A(n4096), .ZN(n4651) );
  INV_X1 U4782 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4567) );
  NOR2_X1 U4783 ( .A1(n4567), .A2(n4653), .ZN(n4566) );
  NAND2_X1 U4784 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4097), .ZN(n4108) );
  INV_X1 U4785 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4952) );
  AOI22_X1 U4786 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4097), .B1(n4655), .B2(
        n4952), .ZN(n4550) );
  NAND2_X1 U4787 ( .A1(n4098), .A2(REG2_REG_9__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U4788 ( .A1(n4098), .A2(REG2_REG_9__SCAN_IN), .B1(n4902), .B2(n4657), .ZN(n4529) );
  INV_X1 U4789 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4101) );
  INV_X1 U4790 ( .A(n4099), .ZN(n4100) );
  NAND2_X1 U4791 ( .A1(n4514), .A2(n4103), .ZN(n4104) );
  NAND2_X1 U4792 ( .A1(n4529), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U4793 ( .A1(n4535), .A2(n4106), .ZN(n4107) );
  NAND2_X1 U4794 ( .A1(n4556), .A2(n4109), .ZN(n4110) );
  NOR2_X1 U4795 ( .A1(n4651), .A2(n4112), .ZN(n4113) );
  NAND2_X1 U4796 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4115), .ZN(n4114) );
  OAI21_X1 U4797 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4115), .A(n4114), .ZN(n4588) );
  INV_X1 U4798 ( .A(n4116), .ZN(n4648) );
  NAND2_X1 U4799 ( .A1(n4117), .A2(n4648), .ZN(n4118) );
  INV_X1 U4800 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4597) );
  NAND2_X1 U4801 ( .A1(n4609), .A2(n4607), .ZN(n4608) );
  AOI22_X1 U4802 ( .A1(n4124), .A2(n4123), .B1(n4474), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n4127) );
  INV_X1 U4803 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4125) );
  MUX2_X1 U4804 ( .A(n4125), .B(REG1_REG_19__SCAN_IN), .S(n4473), .Z(n4126) );
  XNOR2_X1 U4805 ( .A(n4127), .B(n4126), .ZN(n4137) );
  INV_X1 U4806 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4129) );
  MUX2_X1 U4807 ( .A(REG2_REG_19__SCAN_IN), .B(n4129), .S(n4473), .Z(n4130) );
  AOI21_X1 U4808 ( .B1(n4612), .B2(ADDR_REG_19__SCAN_IN), .A(n4131), .ZN(n4132) );
  OAI21_X1 U4809 ( .B1(n4619), .B2(n4133), .A(n4132), .ZN(n4134) );
  OAI21_X1 U4810 ( .B1(n4138), .B2(n4137), .A(n4136), .ZN(U3259) );
  XNOR2_X1 U4811 ( .A(n4346), .B(n4139), .ZN(n4422) );
  NOR2_X1 U4812 ( .A1(n4141), .A2(n4140), .ZN(n4349) );
  AOI21_X1 U4813 ( .B1(n4142), .B2(n4327), .A(n4349), .ZN(n4419) );
  MUX2_X1 U4814 ( .A(n4143), .B(n4419), .S(n4507), .Z(n4144) );
  OAI21_X1 U4815 ( .B1(n4422), .B2(n4339), .A(n4144), .ZN(U3260) );
  INV_X1 U4816 ( .A(n4145), .ZN(n4156) );
  INV_X1 U4817 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4146) );
  OAI22_X1 U4818 ( .A1(n4307), .A2(n4147), .B1(n4146), .B2(n4507), .ZN(n4148)
         );
  AOI21_X1 U4819 ( .B1(n4149), .B2(n4313), .A(n4148), .ZN(n4155) );
  OAI22_X1 U4820 ( .A1(n4151), .A2(n4339), .B1(n4150), .B2(n4261), .ZN(n4152)
         );
  OAI21_X1 U4821 ( .B1(n4153), .B2(n4152), .A(n4507), .ZN(n4154) );
  OAI211_X1 U4822 ( .C1(n4156), .C2(n4342), .A(n4155), .B(n4154), .ZN(U3354)
         );
  XNOR2_X1 U4823 ( .A(n4157), .B(n4159), .ZN(n4358) );
  INV_X1 U4824 ( .A(n4358), .ZN(n4171) );
  XOR2_X1 U4825 ( .A(n4159), .B(n4158), .Z(n4161) );
  OAI22_X1 U4826 ( .A1(n4161), .A2(n4182), .B1(n4160), .B2(n4296), .ZN(n4357)
         );
  NAND2_X1 U4827 ( .A1(n2233), .A2(n4162), .ZN(n4163) );
  NAND2_X1 U4828 ( .A1(n4164), .A2(n4163), .ZN(n4429) );
  NOR2_X1 U4829 ( .A1(n4429), .A2(n4339), .ZN(n4169) );
  AOI22_X1 U4830 ( .A1(n4165), .A2(n4634), .B1(REG2_REG_27__SCAN_IN), .B2(
        n2229), .ZN(n4167) );
  NAND2_X1 U4831 ( .A1(n4197), .A2(n4313), .ZN(n4166) );
  OAI211_X1 U4832 ( .C1(n4307), .C2(n4355), .A(n4167), .B(n4166), .ZN(n4168)
         );
  AOI211_X1 U4833 ( .C1(n4357), .C2(n4507), .A(n4169), .B(n4168), .ZN(n4170)
         );
  OAI21_X1 U4834 ( .B1(n4171), .B2(n4342), .A(n4170), .ZN(U3263) );
  XNOR2_X1 U4835 ( .A(n4172), .B(n4177), .ZN(n4362) );
  INV_X1 U4836 ( .A(n4362), .ZN(n4190) );
  INV_X1 U4837 ( .A(n4173), .ZN(n4174) );
  NAND2_X1 U4838 ( .A1(n4175), .A2(n4174), .ZN(n4176) );
  XOR2_X1 U4839 ( .A(n4177), .B(n4176), .Z(n4183) );
  OAI22_X1 U4840 ( .A1(n4178), .A2(n4406), .B1(n4186), .B2(n4405), .ZN(n4179)
         );
  AOI21_X1 U4841 ( .B1(n4180), .B2(n4328), .A(n4179), .ZN(n4181) );
  OAI21_X1 U4842 ( .B1(n4183), .B2(n4182), .A(n4181), .ZN(n4361) );
  OAI22_X1 U4843 ( .A1(n4185), .A2(n4261), .B1(n4184), .B2(n4507), .ZN(n4188)
         );
  OAI21_X1 U4844 ( .B1(n2330), .B2(n4186), .A(n2233), .ZN(n4433) );
  NOR2_X1 U4845 ( .A1(n4433), .A2(n4339), .ZN(n4187) );
  AOI211_X1 U4846 ( .C1(n4361), .C2(n4507), .A(n4188), .B(n4187), .ZN(n4189)
         );
  OAI21_X1 U4847 ( .B1(n4190), .B2(n4342), .A(n4189), .ZN(U3264) );
  XOR2_X1 U4848 ( .A(n4192), .B(n4191), .Z(n4365) );
  INV_X1 U4849 ( .A(n4365), .ZN(n4207) );
  INV_X1 U4850 ( .A(n4192), .ZN(n4193) );
  XNOR2_X1 U4851 ( .A(n4194), .B(n4193), .ZN(n4195) );
  NAND2_X1 U4852 ( .A1(n4195), .A2(n4324), .ZN(n4199) );
  OAI22_X1 U4853 ( .A1(n4244), .A2(n4406), .B1(n4200), .B2(n4405), .ZN(n4196)
         );
  AOI21_X1 U4854 ( .B1(n4197), .B2(n4328), .A(n4196), .ZN(n4198) );
  NAND2_X1 U4855 ( .A1(n4199), .A2(n4198), .ZN(n4364) );
  OR2_X1 U4856 ( .A1(n4218), .A2(n4200), .ZN(n4201) );
  NAND2_X1 U4857 ( .A1(n4202), .A2(n4201), .ZN(n4437) );
  AOI22_X1 U4858 ( .A1(n4203), .A2(n4634), .B1(n2229), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n4204) );
  OAI21_X1 U4859 ( .B1(n4437), .B2(n4339), .A(n4204), .ZN(n4205) );
  AOI21_X1 U4860 ( .B1(n4507), .B2(n4364), .A(n4205), .ZN(n4206) );
  OAI21_X1 U4861 ( .B1(n4207), .B2(n4342), .A(n4206), .ZN(U3265) );
  XOR2_X1 U4862 ( .A(n4211), .B(n4208), .Z(n4372) );
  INV_X1 U4863 ( .A(n4372), .ZN(n4227) );
  NAND2_X1 U4864 ( .A1(n4210), .A2(n4209), .ZN(n4213) );
  INV_X1 U4865 ( .A(n4211), .ZN(n4212) );
  XNOR2_X1 U4866 ( .A(n4213), .B(n4212), .ZN(n4214) );
  NAND2_X1 U4867 ( .A1(n4214), .A2(n4324), .ZN(n4217) );
  NAND2_X1 U4868 ( .A1(n4215), .A2(n4328), .ZN(n4216) );
  NAND2_X1 U4869 ( .A1(n4217), .A2(n4216), .ZN(n4371) );
  INV_X1 U4870 ( .A(n4218), .ZN(n4219) );
  OAI21_X1 U4871 ( .B1(n4245), .B2(n4368), .A(n4219), .ZN(n4441) );
  OAI22_X1 U4872 ( .A1(n4507), .A2(n4221), .B1(n4220), .B2(n4261), .ZN(n4223)
         );
  NOR2_X1 U4873 ( .A1(n4307), .A2(n4368), .ZN(n4222) );
  AOI211_X1 U4874 ( .C1(n4313), .C2(n4267), .A(n4223), .B(n4222), .ZN(n4224)
         );
  OAI21_X1 U4875 ( .B1(n4441), .B2(n4339), .A(n4224), .ZN(n4225) );
  AOI21_X1 U4876 ( .B1(n4507), .B2(n4371), .A(n4225), .ZN(n4226) );
  OAI21_X1 U4877 ( .B1(n4227), .B2(n4342), .A(n4226), .ZN(U3266) );
  XNOR2_X1 U4878 ( .A(n4228), .B(n4236), .ZN(n4376) );
  INV_X1 U4879 ( .A(n4376), .ZN(n4254) );
  INV_X1 U4880 ( .A(n4229), .ZN(n4230) );
  AOI21_X1 U4881 ( .B1(n4292), .B2(n4233), .A(n4232), .ZN(n4278) );
  INV_X1 U4882 ( .A(n4275), .ZN(n4277) );
  AOI21_X1 U4883 ( .B1(n4278), .B2(n4277), .A(n4234), .ZN(n4266) );
  OAI21_X1 U4884 ( .B1(n4266), .B2(n4265), .A(n4235), .ZN(n4238) );
  INV_X1 U4885 ( .A(n4236), .ZN(n4237) );
  XNOR2_X1 U4886 ( .A(n4238), .B(n4237), .ZN(n4239) );
  NAND2_X1 U4887 ( .A1(n4239), .A2(n4324), .ZN(n4243) );
  AOI22_X1 U4888 ( .A1(n4280), .A2(n4241), .B1(n4327), .B2(n4240), .ZN(n4242)
         );
  OAI211_X1 U4889 ( .C1(n4244), .C2(n4296), .A(n4243), .B(n4242), .ZN(n4375)
         );
  INV_X1 U4890 ( .A(n4260), .ZN(n4248) );
  INV_X1 U4891 ( .A(n4245), .ZN(n4246) );
  OAI21_X1 U4892 ( .B1(n4248), .B2(n4247), .A(n4246), .ZN(n4445) );
  NOR2_X1 U4893 ( .A1(n4445), .A2(n4339), .ZN(n4252) );
  OAI22_X1 U4894 ( .A1(n4507), .A2(n4250), .B1(n4249), .B2(n4261), .ZN(n4251)
         );
  AOI211_X1 U4895 ( .C1(n4375), .C2(n4507), .A(n4252), .B(n4251), .ZN(n4253)
         );
  OAI21_X1 U4896 ( .B1(n4254), .B2(n4342), .A(n4253), .ZN(U3267) );
  NOR2_X1 U4897 ( .A1(n4255), .A2(n4265), .ZN(n4256) );
  OR2_X1 U4898 ( .A1(n4257), .A2(n4256), .ZN(n4379) );
  NAND2_X1 U4899 ( .A1(n4283), .A2(n4258), .ZN(n4259) );
  NAND2_X1 U4900 ( .A1(n4260), .A2(n4259), .ZN(n4449) );
  INV_X1 U4901 ( .A(n4449), .ZN(n4264) );
  OAI22_X1 U4902 ( .A1(n4507), .A2(n4941), .B1(n4262), .B2(n4261), .ZN(n4263)
         );
  AOI21_X1 U4903 ( .B1(n4264), .B2(n4637), .A(n4263), .ZN(n4274) );
  XNOR2_X1 U4904 ( .A(n4266), .B(n4265), .ZN(n4272) );
  NAND2_X1 U4905 ( .A1(n4267), .A2(n4328), .ZN(n4269) );
  OR2_X1 U4906 ( .A1(n4297), .A2(n4406), .ZN(n4268) );
  OAI211_X1 U4907 ( .C1(n4405), .C2(n4270), .A(n4269), .B(n4268), .ZN(n4271)
         );
  AOI21_X1 U4908 ( .B1(n4272), .B2(n4324), .A(n4271), .ZN(n4380) );
  OR2_X1 U4909 ( .A1(n2229), .A2(n4380), .ZN(n4273) );
  OAI211_X1 U4910 ( .C1(n4379), .C2(n4342), .A(n4274), .B(n4273), .ZN(U3268)
         );
  XNOR2_X1 U4911 ( .A(n4276), .B(n4275), .ZN(n4388) );
  INV_X1 U4912 ( .A(n4388), .ZN(n4290) );
  XNOR2_X1 U4913 ( .A(n4278), .B(n4277), .ZN(n4279) );
  NAND2_X1 U4914 ( .A1(n4279), .A2(n4324), .ZN(n4282) );
  NAND2_X1 U4915 ( .A1(n4280), .A2(n4328), .ZN(n4281) );
  NAND2_X1 U4916 ( .A1(n4282), .A2(n4281), .ZN(n4387) );
  OAI21_X1 U4917 ( .B1(n4308), .B2(n4384), .A(n4283), .ZN(n4453) );
  NOR2_X1 U4918 ( .A1(n4453), .A2(n4339), .ZN(n4288) );
  AOI22_X1 U4919 ( .A1(n2229), .A2(REG2_REG_21__SCAN_IN), .B1(n4284), .B2(
        n4634), .ZN(n4286) );
  NAND2_X1 U4920 ( .A1(n4313), .A2(n4329), .ZN(n4285) );
  OAI211_X1 U4921 ( .C1(n4307), .C2(n4384), .A(n4286), .B(n4285), .ZN(n4287)
         );
  AOI211_X1 U4922 ( .C1(n4387), .C2(n4507), .A(n4288), .B(n4287), .ZN(n4289)
         );
  OAI21_X1 U4923 ( .B1(n4290), .B2(n4342), .A(n4289), .ZN(U3269) );
  NAND2_X1 U4924 ( .A1(n4292), .A2(n4291), .ZN(n4294) );
  INV_X1 U4925 ( .A(n4303), .ZN(n4293) );
  XNOR2_X1 U4926 ( .A(n4294), .B(n4293), .ZN(n4295) );
  NAND2_X1 U4927 ( .A1(n4295), .A2(n4324), .ZN(n4299) );
  OR2_X1 U4928 ( .A1(n4297), .A2(n4296), .ZN(n4298) );
  NAND2_X1 U4929 ( .A1(n4299), .A2(n4298), .ZN(n4394) );
  INV_X1 U4930 ( .A(n4394), .ZN(n4316) );
  AOI21_X1 U4931 ( .B1(n4317), .B2(n4301), .A(n4300), .ZN(n4302) );
  XOR2_X1 U4932 ( .A(n4303), .B(n4302), .Z(n4395) );
  NAND2_X1 U4933 ( .A1(n4395), .A2(n4304), .ZN(n4315) );
  AOI22_X1 U4934 ( .A1(n2229), .A2(REG2_REG_20__SCAN_IN), .B1(n4305), .B2(
        n4634), .ZN(n4306) );
  OAI21_X1 U4935 ( .B1(n4391), .B2(n4307), .A(n4306), .ZN(n4311) );
  INV_X1 U4936 ( .A(n4308), .ZN(n4309) );
  OAI21_X1 U4937 ( .B1(n4334), .B2(n4391), .A(n4309), .ZN(n4457) );
  NOR2_X1 U4938 ( .A1(n4457), .A2(n4339), .ZN(n4310) );
  AOI211_X1 U4939 ( .C1(n4313), .C2(n4312), .A(n4311), .B(n4310), .ZN(n4314)
         );
  OAI211_X1 U4940 ( .C1(n2229), .C2(n4316), .A(n4315), .B(n4314), .ZN(U3270)
         );
  XOR2_X1 U4941 ( .A(n4323), .B(n4317), .Z(n4398) );
  INV_X1 U4942 ( .A(n4398), .ZN(n4343) );
  INV_X1 U4943 ( .A(n4318), .ZN(n4320) );
  OAI21_X1 U4944 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4322) );
  XOR2_X1 U4945 ( .A(n4323), .B(n4322), .Z(n4325) );
  NAND2_X1 U4946 ( .A1(n4325), .A2(n4324), .ZN(n4331) );
  AOI22_X1 U4947 ( .A1(n4329), .A2(n4328), .B1(n4327), .B2(n4326), .ZN(n4330)
         );
  OAI211_X1 U4948 ( .C1(n4332), .C2(n4406), .A(n4331), .B(n4330), .ZN(n4397)
         );
  INV_X1 U4949 ( .A(n4333), .ZN(n4336) );
  OAI21_X1 U4950 ( .B1(n4336), .B2(n4335), .A(n2337), .ZN(n4461) );
  AOI22_X1 U4951 ( .A1(n2229), .A2(REG2_REG_19__SCAN_IN), .B1(n4337), .B2(
        n4634), .ZN(n4338) );
  OAI21_X1 U4952 ( .B1(n4461), .B2(n4339), .A(n4338), .ZN(n4340) );
  AOI21_X1 U4953 ( .B1(n4397), .B2(n4507), .A(n4340), .ZN(n4341) );
  OAI21_X1 U4954 ( .B1(n4343), .B2(n4342), .A(n4341), .ZN(U3271) );
  NOR2_X1 U4955 ( .A1(n4419), .A2(n4697), .ZN(n4344) );
  AOI21_X1 U4956 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4697), .A(n4344), .ZN(n4345) );
  OAI21_X1 U4957 ( .B1(n4422), .B2(n4412), .A(n4345), .ZN(U3549) );
  INV_X1 U4958 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4354) );
  AOI21_X1 U4959 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4505) );
  NAND2_X1 U4960 ( .A1(n4505), .A2(n2866), .ZN(n4353) );
  INV_X1 U4961 ( .A(n4349), .ZN(n4350) );
  OAI21_X1 U4962 ( .B1(n4351), .B2(n4405), .A(n4350), .ZN(n4504) );
  NAND2_X1 U4963 ( .A1(n4504), .A2(n4700), .ZN(n4352) );
  OAI211_X1 U4964 ( .C1(n4700), .C2(n4354), .A(n4353), .B(n4352), .ZN(U3548)
         );
  INV_X1 U4965 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4359) );
  OAI22_X1 U4966 ( .A1(n5076), .A2(n4406), .B1(n4355), .B2(n4405), .ZN(n4356)
         );
  AOI211_X1 U4967 ( .C1(n4358), .C2(n4681), .A(n4357), .B(n4356), .ZN(n4426)
         );
  MUX2_X1 U4968 ( .A(n4359), .B(n4426), .S(n4700), .Z(n4360) );
  OAI21_X1 U4969 ( .B1(n4412), .B2(n4429), .A(n4360), .ZN(U3545) );
  INV_X1 U4970 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4837) );
  AOI21_X1 U4971 ( .B1(n4362), .B2(n4681), .A(n4361), .ZN(n4430) );
  MUX2_X1 U4972 ( .A(n4837), .B(n4430), .S(n4700), .Z(n4363) );
  OAI21_X1 U4973 ( .B1(n4412), .B2(n4433), .A(n4363), .ZN(U3544) );
  INV_X1 U4974 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4366) );
  AOI21_X1 U4975 ( .B1(n4365), .B2(n4681), .A(n4364), .ZN(n4434) );
  MUX2_X1 U4976 ( .A(n4366), .B(n4434), .S(n4700), .Z(n4367) );
  OAI21_X1 U4977 ( .B1(n4412), .B2(n4437), .A(n4367), .ZN(U3543) );
  INV_X1 U4978 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4373) );
  OAI22_X1 U4979 ( .A1(n4369), .A2(n4406), .B1(n4368), .B2(n4405), .ZN(n4370)
         );
  AOI211_X1 U4980 ( .C1(n4372), .C2(n4681), .A(n4371), .B(n4370), .ZN(n4438)
         );
  MUX2_X1 U4981 ( .A(n4373), .B(n4438), .S(n4700), .Z(n4374) );
  OAI21_X1 U4982 ( .B1(n4412), .B2(n4441), .A(n4374), .ZN(U3542) );
  INV_X1 U4983 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4377) );
  AOI21_X1 U4984 ( .B1(n4376), .B2(n4681), .A(n4375), .ZN(n4442) );
  MUX2_X1 U4985 ( .A(n4377), .B(n4442), .S(n4700), .Z(n4378) );
  OAI21_X1 U4986 ( .B1(n4412), .B2(n4445), .A(n4378), .ZN(U3541) );
  OR2_X1 U4987 ( .A1(n4379), .A2(n4402), .ZN(n4381) );
  NAND2_X1 U4988 ( .A1(n4381), .A2(n4380), .ZN(n4446) );
  MUX2_X1 U4989 ( .A(n4446), .B(REG1_REG_22__SCAN_IN), .S(n4697), .Z(n4382) );
  INV_X1 U4990 ( .A(n4382), .ZN(n4383) );
  OAI21_X1 U4991 ( .B1(n4412), .B2(n4449), .A(n4383), .ZN(U3540) );
  INV_X1 U4992 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4389) );
  OAI22_X1 U4993 ( .A1(n4385), .A2(n4406), .B1(n4405), .B2(n4384), .ZN(n4386)
         );
  AOI211_X1 U4994 ( .C1(n4388), .C2(n4681), .A(n4387), .B(n4386), .ZN(n4450)
         );
  MUX2_X1 U4995 ( .A(n4389), .B(n4450), .S(n4700), .Z(n4390) );
  OAI21_X1 U4996 ( .B1(n4412), .B2(n4453), .A(n4390), .ZN(U3539) );
  INV_X1 U4997 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4891) );
  OAI22_X1 U4998 ( .A1(n4392), .A2(n4406), .B1(n4391), .B2(n4405), .ZN(n4393)
         );
  AOI211_X1 U4999 ( .C1(n4395), .C2(n4681), .A(n4394), .B(n4393), .ZN(n4454)
         );
  MUX2_X1 U5000 ( .A(n4891), .B(n4454), .S(n4700), .Z(n4396) );
  OAI21_X1 U5001 ( .B1(n4412), .B2(n4457), .A(n4396), .ZN(U3538) );
  AOI21_X1 U5002 ( .B1(n4398), .B2(n4681), .A(n4397), .ZN(n4458) );
  MUX2_X1 U5003 ( .A(n4125), .B(n4458), .S(n4700), .Z(n4399) );
  OAI21_X1 U5004 ( .B1(n4412), .B2(n4461), .A(n4399), .ZN(U3537) );
  OAI211_X1 U5005 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4462)
         );
  MUX2_X1 U5006 ( .A(REG1_REG_18__SCAN_IN), .B(n4462), .S(n4700), .Z(U3536) );
  OAI22_X1 U5007 ( .A1(n4407), .A2(n4406), .B1(n4405), .B2(n4404), .ZN(n4408)
         );
  AOI211_X1 U5008 ( .C1(n4410), .C2(n4681), .A(n4409), .B(n4408), .ZN(n4463)
         );
  MUX2_X1 U5009 ( .A(n4828), .B(n4463), .S(n4700), .Z(n4411) );
  OAI21_X1 U5010 ( .B1(n4412), .B2(n4467), .A(n4411), .ZN(U3535) );
  INV_X1 U5011 ( .A(n4413), .ZN(n4418) );
  NAND3_X1 U5012 ( .A1(n4415), .A2(n4669), .A3(n4414), .ZN(n4416) );
  OAI211_X1 U5013 ( .C1(n4418), .C2(n4664), .A(n4417), .B(n4416), .ZN(n4468)
         );
  MUX2_X1 U5014 ( .A(REG1_REG_14__SCAN_IN), .B(n4468), .S(n4700), .Z(U3532) );
  NOR2_X1 U5015 ( .A1(n4419), .A2(n4689), .ZN(n4420) );
  AOI21_X1 U5016 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4689), .A(n4420), .ZN(n4421) );
  OAI21_X1 U5017 ( .B1(n4422), .B2(n4466), .A(n4421), .ZN(U3517) );
  INV_X1 U5018 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4814) );
  NAND2_X1 U5019 ( .A1(n4505), .A2(n4423), .ZN(n4425) );
  NAND2_X1 U5020 ( .A1(n4504), .A2(n4690), .ZN(n4424) );
  OAI211_X1 U5021 ( .C1(n4690), .C2(n4814), .A(n4425), .B(n4424), .ZN(U3516)
         );
  INV_X1 U5022 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4427) );
  MUX2_X1 U5023 ( .A(n4427), .B(n4426), .S(n4690), .Z(n4428) );
  OAI21_X1 U5024 ( .B1(n4429), .B2(n4466), .A(n4428), .ZN(U3513) );
  INV_X1 U5025 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U5026 ( .A(n4431), .B(n4430), .S(n4690), .Z(n4432) );
  OAI21_X1 U5027 ( .B1(n4433), .B2(n4466), .A(n4432), .ZN(U3512) );
  INV_X1 U5028 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4435) );
  MUX2_X1 U5029 ( .A(n4435), .B(n4434), .S(n4690), .Z(n4436) );
  OAI21_X1 U5030 ( .B1(n4437), .B2(n4466), .A(n4436), .ZN(U3511) );
  INV_X1 U5031 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4439) );
  MUX2_X1 U5032 ( .A(n4439), .B(n4438), .S(n4690), .Z(n4440) );
  OAI21_X1 U5033 ( .B1(n4441), .B2(n4466), .A(n4440), .ZN(U3510) );
  INV_X1 U5034 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4443) );
  MUX2_X1 U5035 ( .A(n4443), .B(n4442), .S(n4690), .Z(n4444) );
  OAI21_X1 U5036 ( .B1(n4445), .B2(n4466), .A(n4444), .ZN(U3509) );
  MUX2_X1 U5037 ( .A(REG0_REG_22__SCAN_IN), .B(n4446), .S(n4690), .Z(n4447) );
  INV_X1 U5038 ( .A(n4447), .ZN(n4448) );
  OAI21_X1 U5039 ( .B1(n4449), .B2(n4466), .A(n4448), .ZN(U3508) );
  INV_X1 U5040 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4451) );
  MUX2_X1 U5041 ( .A(n4451), .B(n4450), .S(n4690), .Z(n4452) );
  OAI21_X1 U5042 ( .B1(n4453), .B2(n4466), .A(n4452), .ZN(U3507) );
  INV_X1 U5043 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4455) );
  MUX2_X1 U5044 ( .A(n4455), .B(n4454), .S(n4690), .Z(n4456) );
  OAI21_X1 U5045 ( .B1(n4457), .B2(n4466), .A(n4456), .ZN(U3506) );
  INV_X1 U5046 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4459) );
  MUX2_X1 U5047 ( .A(n4459), .B(n4458), .S(n4690), .Z(n4460) );
  OAI21_X1 U5048 ( .B1(n4461), .B2(n4466), .A(n4460), .ZN(U3505) );
  MUX2_X1 U5049 ( .A(REG0_REG_18__SCAN_IN), .B(n4462), .S(n4690), .Z(U3503) );
  INV_X1 U5050 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4464) );
  MUX2_X1 U5051 ( .A(n4464), .B(n4463), .S(n4690), .Z(n4465) );
  OAI21_X1 U5052 ( .B1(n4467), .B2(n4466), .A(n4465), .ZN(U3501) );
  MUX2_X1 U5053 ( .A(REG0_REG_14__SCAN_IN), .B(n4468), .S(n4690), .Z(U3495) );
  MUX2_X1 U5054 ( .A(n4469), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5055 ( .A(DATAI_27_), .B(n4470), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5056 ( .A(n4471), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5057 ( .A(DATAI_20_), .B(n4472), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5058 ( .A(n4473), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5059 ( .A(n4474), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5060 ( .A(DATAI_7_), .B(n4475), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5061 ( .A(n4476), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5062 ( .A(DATAI_4_), .B(n4477), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5063 ( .A(DATAI_3_), .B(n4478), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5064 ( .A(n4479), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5065 ( .A(n2230), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5066 ( .A(DATAI_28_), .ZN(n4481) );
  AOI22_X1 U5067 ( .A1(STATE_REG_SCAN_IN), .A2(n4482), .B1(n4481), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U5068 ( .A1(STATE_REG_SCAN_IN), .A2(n4483), .ZN(n4601) );
  AOI21_X1 U5069 ( .B1(n4485), .B2(n4484), .A(n4601), .ZN(n4489) );
  NAND2_X1 U5070 ( .A1(n4487), .A2(n4486), .ZN(n4488) );
  OAI211_X1 U5071 ( .C1(n4491), .C2(n4490), .A(n4489), .B(n4488), .ZN(n4492)
         );
  INV_X1 U5072 ( .A(n4492), .ZN(n4501) );
  OAI21_X1 U5073 ( .B1(n2457), .B2(n4495), .A(n4494), .ZN(n4497) );
  XNOR2_X1 U5074 ( .A(n4497), .B(n4496), .ZN(n4499) );
  NAND2_X1 U5075 ( .A1(n4499), .A2(n4498), .ZN(n4500) );
  OAI211_X1 U5076 ( .C1(n4503), .C2(n4502), .A(n4501), .B(n4500), .ZN(U3223)
         );
  AOI22_X1 U5077 ( .A1(n4505), .A2(n4637), .B1(n4507), .B2(n4504), .ZN(n4506)
         );
  OAI21_X1 U5078 ( .B1(n2882), .B2(n4507), .A(n4506), .ZN(U3261) );
  AOI21_X1 U5079 ( .B1(n3064), .B2(n4509), .A(n4508), .ZN(n4510) );
  XNOR2_X1 U5080 ( .A(n4510), .B(IR_REG_0__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5081 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4612), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4511) );
  OAI21_X1 U5082 ( .B1(n4513), .B2(n4512), .A(n4511), .ZN(U3240) );
  OAI211_X1 U5083 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4516), .A(n4568), .B(n4515), 
        .ZN(n4517) );
  NAND2_X1 U5084 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  AOI21_X1 U5085 ( .B1(n4612), .B2(ADDR_REG_8__SCAN_IN), .A(n4519), .ZN(n4523)
         );
  OAI211_X1 U5086 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4521), .A(n4613), .B(n4520), 
        .ZN(n4522) );
  OAI211_X1 U5087 ( .C1(n4619), .C2(n2355), .A(n4523), .B(n4522), .ZN(U3248)
         );
  OAI211_X1 U5088 ( .C1(n4526), .C2(n4525), .A(n4613), .B(n4524), .ZN(n4531)
         );
  OAI211_X1 U5089 ( .C1(n4529), .C2(n4528), .A(n4568), .B(n4527), .ZN(n4530)
         );
  OAI211_X1 U5090 ( .C1(n4619), .C2(n4657), .A(n4531), .B(n4530), .ZN(n4532)
         );
  AOI211_X1 U5091 ( .C1(n4612), .C2(ADDR_REG_9__SCAN_IN), .A(n4533), .B(n4532), 
        .ZN(n4534) );
  INV_X1 U5092 ( .A(n4534), .ZN(U3249) );
  OAI211_X1 U5093 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4537), .A(n4568), .B(n4536), .ZN(n4539) );
  NAND2_X1 U5094 ( .A1(n4539), .A2(n4538), .ZN(n4540) );
  AOI21_X1 U5095 ( .B1(n4612), .B2(ADDR_REG_10__SCAN_IN), .A(n4540), .ZN(n4544) );
  OAI211_X1 U5096 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4542), .A(n4613), .B(n4541), .ZN(n4543) );
  OAI211_X1 U5097 ( .C1(n4619), .C2(n2344), .A(n4544), .B(n4543), .ZN(U3250)
         );
  OAI211_X1 U5098 ( .C1(n4547), .C2(n4546), .A(n4613), .B(n4545), .ZN(n4552)
         );
  OAI211_X1 U5099 ( .C1(n4550), .C2(n4549), .A(n4568), .B(n4548), .ZN(n4551)
         );
  OAI211_X1 U5100 ( .C1(n4619), .C2(n4655), .A(n4552), .B(n4551), .ZN(n4553)
         );
  AOI211_X1 U5101 ( .C1(n4612), .C2(ADDR_REG_11__SCAN_IN), .A(n4554), .B(n4553), .ZN(n4555) );
  INV_X1 U5102 ( .A(n4555), .ZN(U3251) );
  OAI211_X1 U5103 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4558), .A(n4568), .B(n4557), .ZN(n4560) );
  NAND2_X1 U5104 ( .A1(n4560), .A2(n4559), .ZN(n4561) );
  AOI21_X1 U5105 ( .B1(n4612), .B2(ADDR_REG_12__SCAN_IN), .A(n4561), .ZN(n4565) );
  OAI211_X1 U5106 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4563), .A(n4613), .B(n4562), .ZN(n4564) );
  OAI211_X1 U5107 ( .C1(n4619), .C2(n2352), .A(n4565), .B(n4564), .ZN(U3252)
         );
  AOI21_X1 U5108 ( .B1(n4567), .B2(n4653), .A(n4566), .ZN(n4571) );
  OAI21_X1 U5109 ( .B1(n4571), .B2(n4570), .A(n4568), .ZN(n4569) );
  AOI21_X1 U5110 ( .B1(n4571), .B2(n4570), .A(n4569), .ZN(n4572) );
  AOI211_X1 U5111 ( .C1(n4612), .C2(ADDR_REG_13__SCAN_IN), .A(n4573), .B(n4572), .ZN(n4578) );
  OAI211_X1 U5112 ( .C1(n4576), .C2(n4575), .A(n4613), .B(n4574), .ZN(n4577)
         );
  OAI211_X1 U5113 ( .C1(n4619), .C2(n4653), .A(n4578), .B(n4577), .ZN(U3253)
         );
  INV_X1 U5114 ( .A(n4579), .ZN(n4583) );
  AOI211_X1 U5115 ( .C1(n3457), .C2(n4581), .A(n4580), .B(n4606), .ZN(n4582)
         );
  AOI211_X1 U5116 ( .C1(n4612), .C2(ADDR_REG_14__SCAN_IN), .A(n4583), .B(n4582), .ZN(n4587) );
  OAI211_X1 U5117 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4585), .A(n4613), .B(n4584), .ZN(n4586) );
  OAI211_X1 U5118 ( .C1(n4619), .C2(n4651), .A(n4587), .B(n4586), .ZN(U3254)
         );
  AOI211_X1 U5119 ( .C1(n4589), .C2(n4588), .A(n2249), .B(n4606), .ZN(n4590)
         );
  AOI211_X1 U5120 ( .C1(n4612), .C2(ADDR_REG_15__SCAN_IN), .A(n4591), .B(n4590), .ZN(n4596) );
  OAI211_X1 U5121 ( .C1(n4594), .C2(n4593), .A(n4613), .B(n4592), .ZN(n4595)
         );
  OAI211_X1 U5122 ( .C1(n4619), .C2(n4650), .A(n4596), .B(n4595), .ZN(U3255)
         );
  AOI221_X1 U5123 ( .B1(n4599), .B2(n4598), .C1(n4597), .C2(n4598), .A(n4606), 
        .ZN(n4600) );
  AOI211_X1 U5124 ( .C1(n4612), .C2(ADDR_REG_16__SCAN_IN), .A(n4601), .B(n4600), .ZN(n4605) );
  OAI221_X1 U5125 ( .B1(n4603), .B2(REG1_REG_16__SCAN_IN), .C1(n4603), .C2(
        n4602), .A(n4613), .ZN(n4604) );
  OAI211_X1 U5126 ( .C1(n4619), .C2(n4648), .A(n4605), .B(n4604), .ZN(U3256)
         );
  AOI221_X1 U5127 ( .B1(n4609), .B2(n4608), .C1(n4607), .C2(n4608), .A(n4606), 
        .ZN(n4610) );
  AOI211_X1 U5128 ( .C1(n4612), .C2(ADDR_REG_17__SCAN_IN), .A(n4611), .B(n4610), .ZN(n4618) );
  OAI221_X1 U5129 ( .B1(n4616), .B2(n4615), .C1(n4616), .C2(n4614), .A(n4613), 
        .ZN(n4617) );
  OAI211_X1 U5130 ( .C1(n4619), .C2(n4646), .A(n4618), .B(n4617), .ZN(U3257)
         );
  AOI22_X1 U5131 ( .A1(n4620), .A2(n4634), .B1(REG2_REG_10__SCAN_IN), .B2(
        n2229), .ZN(n4625) );
  INV_X1 U5132 ( .A(n4621), .ZN(n4622) );
  AOI22_X1 U5133 ( .A1(n4623), .A2(n4638), .B1(n4637), .B2(n4622), .ZN(n4624)
         );
  OAI211_X1 U5134 ( .C1(n2229), .C2(n4626), .A(n4625), .B(n4624), .ZN(U3280)
         );
  AOI22_X1 U5135 ( .A1(n4627), .A2(n4634), .B1(REG2_REG_8__SCAN_IN), .B2(n2229), .ZN(n4632) );
  INV_X1 U5136 ( .A(n4628), .ZN(n4629) );
  AOI22_X1 U5137 ( .A1(n4630), .A2(n4638), .B1(n4637), .B2(n4629), .ZN(n4631)
         );
  OAI211_X1 U5138 ( .C1(n2229), .C2(n4633), .A(n4632), .B(n4631), .ZN(U3282)
         );
  AOI22_X1 U5139 ( .A1(n4635), .A2(n4634), .B1(REG2_REG_6__SCAN_IN), .B2(n2229), .ZN(n4641) );
  AOI22_X1 U5140 ( .A1(n4639), .A2(n4638), .B1(n4637), .B2(n4636), .ZN(n4640)
         );
  OAI211_X1 U5141 ( .C1(n2229), .C2(n4642), .A(n4641), .B(n4640), .ZN(U3284)
         );
  INV_X1 U5142 ( .A(D_REG_31__SCAN_IN), .ZN(n4885) );
  NOR2_X1 U5143 ( .A1(n4644), .A2(n4885), .ZN(U3291) );
  AND2_X1 U5144 ( .A1(D_REG_30__SCAN_IN), .A2(n4643), .ZN(U3292) );
  INV_X1 U5145 ( .A(D_REG_29__SCAN_IN), .ZN(n4804) );
  NOR2_X1 U5146 ( .A1(n4644), .A2(n4804), .ZN(U3293) );
  INV_X1 U5147 ( .A(D_REG_28__SCAN_IN), .ZN(n4935) );
  NOR2_X1 U5148 ( .A1(n4644), .A2(n4935), .ZN(U3294) );
  AND2_X1 U5149 ( .A1(D_REG_27__SCAN_IN), .A2(n4643), .ZN(U3295) );
  AND2_X1 U5150 ( .A1(D_REG_26__SCAN_IN), .A2(n4643), .ZN(U3296) );
  INV_X1 U5151 ( .A(D_REG_25__SCAN_IN), .ZN(n4899) );
  NOR2_X1 U5152 ( .A1(n4644), .A2(n4899), .ZN(U3297) );
  INV_X1 U5153 ( .A(D_REG_24__SCAN_IN), .ZN(n4951) );
  NOR2_X1 U5154 ( .A1(n4644), .A2(n4951), .ZN(U3298) );
  AND2_X1 U5155 ( .A1(n4643), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  AND2_X1 U5156 ( .A1(D_REG_22__SCAN_IN), .A2(n4643), .ZN(U3300) );
  AND2_X1 U5157 ( .A1(D_REG_21__SCAN_IN), .A2(n4643), .ZN(U3301) );
  AND2_X1 U5158 ( .A1(D_REG_20__SCAN_IN), .A2(n4643), .ZN(U3302) );
  AND2_X1 U5159 ( .A1(D_REG_19__SCAN_IN), .A2(n4643), .ZN(U3303) );
  AND2_X1 U5160 ( .A1(D_REG_18__SCAN_IN), .A2(n4643), .ZN(U3304) );
  AND2_X1 U5161 ( .A1(D_REG_17__SCAN_IN), .A2(n4643), .ZN(U3305) );
  AND2_X1 U5162 ( .A1(D_REG_16__SCAN_IN), .A2(n4643), .ZN(U3306) );
  AND2_X1 U5163 ( .A1(D_REG_15__SCAN_IN), .A2(n4643), .ZN(U3307) );
  INV_X1 U5164 ( .A(D_REG_14__SCAN_IN), .ZN(n4958) );
  NOR2_X1 U5165 ( .A1(n4644), .A2(n4958), .ZN(U3308) );
  AND2_X1 U5166 ( .A1(D_REG_13__SCAN_IN), .A2(n4643), .ZN(U3309) );
  AND2_X1 U5167 ( .A1(D_REG_12__SCAN_IN), .A2(n4643), .ZN(U3310) );
  AND2_X1 U5168 ( .A1(n4643), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  INV_X1 U5169 ( .A(D_REG_10__SCAN_IN), .ZN(n4800) );
  NOR2_X1 U5170 ( .A1(n4644), .A2(n4800), .ZN(U3312) );
  INV_X1 U5171 ( .A(D_REG_9__SCAN_IN), .ZN(n4942) );
  NOR2_X1 U5172 ( .A1(n4644), .A2(n4942), .ZN(U3313) );
  AND2_X1 U5173 ( .A1(n4643), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  INV_X1 U5174 ( .A(D_REG_7__SCAN_IN), .ZN(n4917) );
  NOR2_X1 U5175 ( .A1(n4644), .A2(n4917), .ZN(U3315) );
  INV_X1 U5176 ( .A(D_REG_6__SCAN_IN), .ZN(n4793) );
  NOR2_X1 U5177 ( .A1(n4644), .A2(n4793), .ZN(U3316) );
  AND2_X1 U5178 ( .A1(D_REG_5__SCAN_IN), .A2(n4643), .ZN(U3317) );
  INV_X1 U5179 ( .A(D_REG_4__SCAN_IN), .ZN(n4794) );
  NOR2_X1 U5180 ( .A1(n4644), .A2(n4794), .ZN(U3318) );
  AND2_X1 U5181 ( .A1(D_REG_3__SCAN_IN), .A2(n4643), .ZN(U3319) );
  INV_X1 U5182 ( .A(D_REG_2__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U5183 ( .A1(n4644), .A2(n4795), .ZN(U3320) );
  INV_X1 U5184 ( .A(DATAI_23_), .ZN(n4954) );
  AOI21_X1 U5185 ( .B1(U3149), .B2(n4954), .A(n4645), .ZN(U3329) );
  AOI22_X1 U5186 ( .A1(STATE_REG_SCAN_IN), .A2(n4646), .B1(n2711), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5187 ( .A(DATAI_16_), .ZN(n4647) );
  AOI22_X1 U5188 ( .A1(STATE_REG_SCAN_IN), .A2(n4648), .B1(n4647), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5189 ( .A(DATAI_15_), .ZN(n4649) );
  AOI22_X1 U5190 ( .A1(STATE_REG_SCAN_IN), .A2(n4650), .B1(n4649), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5191 ( .A(DATAI_14_), .ZN(n4767) );
  AOI22_X1 U5192 ( .A1(STATE_REG_SCAN_IN), .A2(n4651), .B1(n4767), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5193 ( .A(DATAI_13_), .ZN(n4652) );
  AOI22_X1 U5194 ( .A1(STATE_REG_SCAN_IN), .A2(n4653), .B1(n4652), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5195 ( .A(DATAI_12_), .ZN(n4980) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n2352), .B1(n4980), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5197 ( .A(DATAI_11_), .ZN(n4654) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4655), .B1(n4654), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5199 ( .A(DATAI_10_), .ZN(n4985) );
  AOI22_X1 U5200 ( .A1(STATE_REG_SCAN_IN), .A2(n2344), .B1(n4985), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5201 ( .A(DATAI_9_), .ZN(n4656) );
  AOI22_X1 U5202 ( .A1(STATE_REG_SCAN_IN), .A2(n4657), .B1(n4656), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5203 ( .A(DATAI_8_), .ZN(n4658) );
  AOI22_X1 U5204 ( .A1(STATE_REG_SCAN_IN), .A2(n2355), .B1(n4658), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5205 ( .A(DATAI_0_), .ZN(n4659) );
  AOI22_X1 U5206 ( .A1(STATE_REG_SCAN_IN), .A2(n3065), .B1(n4659), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5207 ( .C1(n4688), .C2(n4662), .A(n4661), .B(n4660), .ZN(n4691)
         );
  INV_X1 U5208 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U5209 ( .A1(n4690), .A2(n4691), .B1(n4803), .B2(n4689), .ZN(U3467)
         );
  OAI22_X1 U5210 ( .A1(n4665), .A2(n4664), .B1(n4683), .B2(n4663), .ZN(n4666)
         );
  NOR2_X1 U5211 ( .A1(n4667), .A2(n4666), .ZN(n4692) );
  INV_X1 U5212 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U5213 ( .A1(n4690), .A2(n4692), .B1(n4973), .B2(n4689), .ZN(U3469)
         );
  AND3_X1 U5214 ( .A1(n4670), .A2(n4669), .A3(n4668), .ZN(n4672) );
  AOI211_X1 U5215 ( .C1(n4688), .C2(n4673), .A(n4672), .B(n4671), .ZN(n4693)
         );
  INV_X1 U5216 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4806) );
  AOI22_X1 U5217 ( .A1(n4690), .A2(n4693), .B1(n4806), .B2(n4689), .ZN(U3471)
         );
  INV_X1 U5218 ( .A(n4674), .ZN(n4676) );
  AOI211_X1 U5219 ( .C1(n4677), .C2(n4688), .A(n4676), .B(n4675), .ZN(n4695)
         );
  INV_X1 U5220 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5221 ( .A1(n4690), .A2(n4695), .B1(n4678), .B2(n4689), .ZN(U3475)
         );
  AOI211_X1 U5222 ( .C1(n4682), .C2(n4681), .A(n4680), .B(n4679), .ZN(n4696)
         );
  INV_X1 U5223 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U5224 ( .A1(n4690), .A2(n4696), .B1(n4965), .B2(n4689), .ZN(U3481)
         );
  NOR2_X1 U5225 ( .A1(n4684), .A2(n4683), .ZN(n4686) );
  AOI211_X1 U5226 ( .C1(n4688), .C2(n4687), .A(n4686), .B(n4685), .ZN(n4699)
         );
  INV_X1 U5227 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U5228 ( .A1(n4690), .A2(n4699), .B1(n4901), .B2(n4689), .ZN(U3489)
         );
  AOI22_X1 U5229 ( .A1(n4700), .A2(n4691), .B1(n3064), .B2(n4697), .ZN(U3518)
         );
  AOI22_X1 U5230 ( .A1(n4700), .A2(n4692), .B1(n3031), .B2(n4697), .ZN(U3519)
         );
  AOI22_X1 U5231 ( .A1(n4700), .A2(n4693), .B1(n4905), .B2(n4697), .ZN(U3520)
         );
  AOI22_X1 U5232 ( .A1(n4700), .A2(n4695), .B1(n4694), .B2(n4697), .ZN(U3522)
         );
  AOI22_X1 U5233 ( .A1(n4700), .A2(n4696), .B1(n4074), .B2(n4697), .ZN(U3525)
         );
  AOI22_X1 U5234 ( .A1(n4700), .A2(n4699), .B1(n4698), .B2(n4697), .ZN(U3529)
         );
  AOI22_X1 U5235 ( .A1(DATAI_18_), .A2(keyinput237), .B1(DATAI_13_), .B2(
        keyinput238), .ZN(n4701) );
  OAI221_X1 U5236 ( .B1(DATAI_18_), .B2(keyinput237), .C1(DATAI_13_), .C2(
        keyinput238), .A(n4701), .ZN(n4708) );
  AOI22_X1 U5237 ( .A1(DATAI_6_), .A2(keyinput181), .B1(DATAI_10_), .B2(
        keyinput141), .ZN(n4702) );
  OAI221_X1 U5238 ( .B1(DATAI_6_), .B2(keyinput181), .C1(DATAI_10_), .C2(
        keyinput141), .A(n4702), .ZN(n4707) );
  AOI22_X1 U5239 ( .A1(DATAI_4_), .A2(keyinput223), .B1(DATAI_5_), .B2(
        keyinput166), .ZN(n4703) );
  OAI221_X1 U5240 ( .B1(DATAI_4_), .B2(keyinput223), .C1(DATAI_5_), .C2(
        keyinput166), .A(n4703), .ZN(n4706) );
  AOI22_X1 U5241 ( .A1(DATAI_0_), .A2(keyinput232), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput184), .ZN(n4704) );
  OAI221_X1 U5242 ( .B1(DATAI_0_), .B2(keyinput232), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput184), .A(n4704), .ZN(n4705) );
  NOR4_X1 U5243 ( .A1(n4708), .A2(n4707), .A3(n4706), .A4(n4705), .ZN(n4736)
         );
  AOI22_X1 U5244 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput250), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput169), .ZN(n4709) );
  OAI221_X1 U5245 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput250), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput169), .A(n4709), .ZN(n4716) );
  AOI22_X1 U5246 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput185), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput161), .ZN(n4710) );
  OAI221_X1 U5247 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput185), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput161), .A(n4710), .ZN(n4715) );
  AOI22_X1 U5248 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput239), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput230), .ZN(n4711) );
  OAI221_X1 U5249 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput239), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput230), .A(n4711), .ZN(n4714) );
  AOI22_X1 U5250 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput198), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput211), .ZN(n4712) );
  OAI221_X1 U5251 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput198), .C1(
        IR_REG_23__SCAN_IN), .C2(keyinput211), .A(n4712), .ZN(n4713) );
  NOR4_X1 U5252 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4735)
         );
  AOI22_X1 U5253 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput196), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput152), .ZN(n4717) );
  OAI221_X1 U5254 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput196), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput152), .A(n4717), .ZN(n4724) );
  AOI22_X1 U5255 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput248), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput236), .ZN(n4718) );
  OAI221_X1 U5256 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput248), .C1(
        D_REG_11__SCAN_IN), .C2(keyinput236), .A(n4718), .ZN(n4723) );
  AOI22_X1 U5257 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput154), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput129), .ZN(n4719) );
  OAI221_X1 U5258 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput154), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput129), .A(n4719), .ZN(n4722) );
  AOI22_X1 U5259 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput179), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput224), .ZN(n4720) );
  OAI221_X1 U5260 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput179), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput224), .A(n4720), .ZN(n4721) );
  NOR4_X1 U5261 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4734)
         );
  AOI22_X1 U5262 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput165), .B1(
        REG0_REG_3__SCAN_IN), .B2(keyinput142), .ZN(n4725) );
  OAI221_X1 U5263 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput165), .C1(
        REG0_REG_3__SCAN_IN), .C2(keyinput142), .A(n4725), .ZN(n4732) );
  AOI22_X1 U5264 ( .A1(REG0_REG_5__SCAN_IN), .A2(keyinput255), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput205), .ZN(n4726) );
  OAI221_X1 U5265 ( .B1(REG0_REG_5__SCAN_IN), .B2(keyinput255), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput205), .A(n4726), .ZN(n4731) );
  AOI22_X1 U5266 ( .A1(REG0_REG_12__SCAN_IN), .A2(keyinput134), .B1(
        REG0_REG_19__SCAN_IN), .B2(keyinput151), .ZN(n4727) );
  OAI221_X1 U5267 ( .B1(REG0_REG_12__SCAN_IN), .B2(keyinput134), .C1(
        REG0_REG_19__SCAN_IN), .C2(keyinput151), .A(n4727), .ZN(n4730) );
  AOI22_X1 U5268 ( .A1(REG0_REG_22__SCAN_IN), .A2(keyinput158), .B1(
        REG0_REG_26__SCAN_IN), .B2(keyinput157), .ZN(n4728) );
  OAI221_X1 U5269 ( .B1(REG0_REG_22__SCAN_IN), .B2(keyinput158), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput157), .A(n4728), .ZN(n4729) );
  NOR4_X1 U5270 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4733)
         );
  NAND4_X1 U5271 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .ZN(n4874)
         );
  AOI22_X1 U5272 ( .A1(REG1_REG_1__SCAN_IN), .A2(keyinput242), .B1(
        REG1_REG_6__SCAN_IN), .B2(keyinput150), .ZN(n4737) );
  OAI221_X1 U5273 ( .B1(REG1_REG_1__SCAN_IN), .B2(keyinput242), .C1(
        REG1_REG_6__SCAN_IN), .C2(keyinput150), .A(n4737), .ZN(n4744) );
  AOI22_X1 U5274 ( .A1(REG1_REG_11__SCAN_IN), .A2(keyinput137), .B1(
        REG1_REG_22__SCAN_IN), .B2(keyinput226), .ZN(n4738) );
  OAI221_X1 U5275 ( .B1(REG1_REG_11__SCAN_IN), .B2(keyinput137), .C1(
        REG1_REG_22__SCAN_IN), .C2(keyinput226), .A(n4738), .ZN(n4743) );
  AOI22_X1 U5276 ( .A1(REG2_REG_6__SCAN_IN), .A2(keyinput225), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput219), .ZN(n4739) );
  OAI221_X1 U5277 ( .B1(REG2_REG_6__SCAN_IN), .B2(keyinput225), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput219), .A(n4739), .ZN(n4742) );
  AOI22_X1 U5278 ( .A1(REG2_REG_15__SCAN_IN), .A2(keyinput138), .B1(
        REG2_REG_10__SCAN_IN), .B2(keyinput227), .ZN(n4740) );
  OAI221_X1 U5279 ( .B1(REG2_REG_15__SCAN_IN), .B2(keyinput138), .C1(
        REG2_REG_10__SCAN_IN), .C2(keyinput227), .A(n4740), .ZN(n4741) );
  NOR4_X1 U5280 ( .A1(n4744), .A2(n4743), .A3(n4742), .A4(n4741), .ZN(n4775)
         );
  AOI22_X1 U5281 ( .A1(REG2_REG_11__SCAN_IN), .A2(keyinput178), .B1(
        REG2_REG_21__SCAN_IN), .B2(keyinput253), .ZN(n4745) );
  OAI221_X1 U5282 ( .B1(REG2_REG_11__SCAN_IN), .B2(keyinput178), .C1(
        REG2_REG_21__SCAN_IN), .C2(keyinput253), .A(n4745), .ZN(n4752) );
  AOI22_X1 U5283 ( .A1(REG2_REG_30__SCAN_IN), .A2(keyinput228), .B1(
        REG2_REG_27__SCAN_IN), .B2(keyinput200), .ZN(n4746) );
  OAI221_X1 U5284 ( .B1(REG2_REG_30__SCAN_IN), .B2(keyinput228), .C1(
        REG2_REG_27__SCAN_IN), .C2(keyinput200), .A(n4746), .ZN(n4751) );
  AOI22_X1 U5285 ( .A1(ADDR_REG_8__SCAN_IN), .A2(keyinput175), .B1(
        ADDR_REG_12__SCAN_IN), .B2(keyinput144), .ZN(n4747) );
  OAI221_X1 U5286 ( .B1(ADDR_REG_8__SCAN_IN), .B2(keyinput175), .C1(
        ADDR_REG_12__SCAN_IN), .C2(keyinput144), .A(n4747), .ZN(n4750) );
  AOI22_X1 U5287 ( .A1(DATAO_REG_10__SCAN_IN), .A2(keyinput131), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput143), .ZN(n4748) );
  OAI221_X1 U5288 ( .B1(DATAO_REG_10__SCAN_IN), .B2(keyinput131), .C1(
        DATAO_REG_8__SCAN_IN), .C2(keyinput143), .A(n4748), .ZN(n4749) );
  NOR4_X1 U5289 ( .A1(n4752), .A2(n4751), .A3(n4750), .A4(n4749), .ZN(n4774)
         );
  AOI22_X1 U5290 ( .A1(DATAO_REG_13__SCAN_IN), .A2(keyinput203), .B1(
        DATAO_REG_11__SCAN_IN), .B2(keyinput172), .ZN(n4753) );
  OAI221_X1 U5291 ( .B1(DATAO_REG_13__SCAN_IN), .B2(keyinput203), .C1(
        DATAO_REG_11__SCAN_IN), .C2(keyinput172), .A(n4753), .ZN(n4760) );
  AOI22_X1 U5292 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput201), .B1(
        B_REG_SCAN_IN), .B2(keyinput130), .ZN(n4754) );
  OAI221_X1 U5293 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput201), .C1(
        B_REG_SCAN_IN), .C2(keyinput130), .A(n4754), .ZN(n4759) );
  AOI22_X1 U5294 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput163), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput139), .ZN(n4755) );
  OAI221_X1 U5295 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput163), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput139), .A(n4755), .ZN(n4758) );
  INV_X1 U5296 ( .A(DATAI_30_), .ZN(n4889) );
  AOI22_X1 U5297 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput197), .B1(n4889), 
        .B2(keyinput156), .ZN(n4756) );
  OAI221_X1 U5298 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput197), .C1(n4889), 
        .C2(keyinput156), .A(n4756), .ZN(n4757) );
  NOR4_X1 U5299 ( .A1(n4760), .A2(n4759), .A3(n4758), .A4(n4757), .ZN(n4773)
         );
  AOI22_X1 U5300 ( .A1(n4762), .A2(keyinput170), .B1(keyinput162), .B2(n4954), 
        .ZN(n4761) );
  OAI221_X1 U5301 ( .B1(n4762), .B2(keyinput170), .C1(n4954), .C2(keyinput162), 
        .A(n4761), .ZN(n4771) );
  INV_X1 U5302 ( .A(DATAI_22_), .ZN(n4949) );
  AOI22_X1 U5303 ( .A1(n4949), .A2(keyinput191), .B1(keyinput243), .B2(n4916), 
        .ZN(n4763) );
  OAI221_X1 U5304 ( .B1(n4949), .B2(keyinput191), .C1(n4916), .C2(keyinput243), 
        .A(n4763), .ZN(n4770) );
  INV_X1 U5305 ( .A(DATAI_20_), .ZN(n4765) );
  INV_X1 U5306 ( .A(DATAI_19_), .ZN(n4914) );
  AOI22_X1 U5307 ( .A1(n4765), .A2(keyinput213), .B1(keyinput192), .B2(n4914), 
        .ZN(n4764) );
  OAI221_X1 U5308 ( .B1(n4765), .B2(keyinput213), .C1(n4914), .C2(keyinput192), 
        .A(n4764), .ZN(n4769) );
  AOI22_X1 U5309 ( .A1(n4767), .A2(keyinput190), .B1(keyinput149), .B2(n4980), 
        .ZN(n4766) );
  OAI221_X1 U5310 ( .B1(n4767), .B2(keyinput190), .C1(n4980), .C2(keyinput149), 
        .A(n4766), .ZN(n4768) );
  NOR4_X1 U5311 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4772)
         );
  NAND4_X1 U5312 ( .A1(n4775), .A2(n4774), .A3(n4773), .A4(n4772), .ZN(n4873)
         );
  INV_X1 U5313 ( .A(DATAI_7_), .ZN(n4888) );
  AOI22_X1 U5314 ( .A1(n4888), .A2(keyinput148), .B1(keyinput145), .B2(n2367), 
        .ZN(n4776) );
  OAI221_X1 U5315 ( .B1(n4888), .B2(keyinput148), .C1(n2367), .C2(keyinput145), 
        .A(n4776), .ZN(n4785) );
  INV_X1 U5316 ( .A(DATAI_3_), .ZN(n4979) );
  AOI22_X1 U5317 ( .A1(n4979), .A2(keyinput133), .B1(n2560), .B2(keyinput135), 
        .ZN(n4777) );
  OAI221_X1 U5318 ( .B1(n4979), .B2(keyinput133), .C1(n2560), .C2(keyinput135), 
        .A(n4777), .ZN(n4784) );
  INV_X1 U5319 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4780) );
  INV_X1 U5320 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5321 ( .A1(n4780), .A2(keyinput160), .B1(keyinput217), .B2(n4779), 
        .ZN(n4778) );
  OAI221_X1 U5322 ( .B1(n4780), .B2(keyinput160), .C1(n4779), .C2(keyinput217), 
        .A(n4778), .ZN(n4783) );
  AOI22_X1 U5323 ( .A1(n4972), .A2(keyinput153), .B1(keyinput136), .B2(n3074), 
        .ZN(n4781) );
  OAI221_X1 U5324 ( .B1(n4972), .B2(keyinput153), .C1(n3074), .C2(keyinput136), 
        .A(n4781), .ZN(n4782) );
  NOR4_X1 U5325 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4824)
         );
  XOR2_X1 U5326 ( .A(IR_REG_9__SCAN_IN), .B(keyinput221), .Z(n4788) );
  XOR2_X1 U5327 ( .A(IR_REG_13__SCAN_IN), .B(keyinput189), .Z(n4787) );
  XNOR2_X1 U5328 ( .A(keyinput215), .B(n2774), .ZN(n4786) );
  NOR3_X1 U5329 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(n4791) );
  XOR2_X1 U5330 ( .A(n2617), .B(keyinput206), .Z(n4790) );
  XNOR2_X1 U5331 ( .A(IR_REG_26__SCAN_IN), .B(keyinput240), .ZN(n4789) );
  NAND3_X1 U5332 ( .A1(n4791), .A2(n4790), .A3(n4789), .ZN(n4798) );
  AOI22_X1 U5333 ( .A1(n4794), .A2(keyinput254), .B1(keyinput188), .B2(n4793), 
        .ZN(n4792) );
  OAI221_X1 U5334 ( .B1(n4794), .B2(keyinput254), .C1(n4793), .C2(keyinput188), 
        .A(n4792), .ZN(n4797) );
  XNOR2_X1 U5335 ( .A(n4795), .B(keyinput244), .ZN(n4796) );
  NOR3_X1 U5336 ( .A1(n4798), .A2(n4797), .A3(n4796), .ZN(n4823) );
  AOI22_X1 U5337 ( .A1(n4800), .A2(keyinput194), .B1(keyinput246), .B2(n4917), 
        .ZN(n4799) );
  OAI221_X1 U5338 ( .B1(n4800), .B2(keyinput194), .C1(n4917), .C2(keyinput246), 
        .A(n4799), .ZN(n4810) );
  AOI22_X1 U5339 ( .A1(n4935), .A2(keyinput202), .B1(n4885), .B2(keyinput245), 
        .ZN(n4801) );
  OAI221_X1 U5340 ( .B1(n4935), .B2(keyinput202), .C1(n4885), .C2(keyinput245), 
        .A(n4801), .ZN(n4809) );
  AOI22_X1 U5341 ( .A1(n4804), .A2(keyinput207), .B1(keyinput249), .B2(n4803), 
        .ZN(n4802) );
  OAI221_X1 U5342 ( .B1(n4804), .B2(keyinput207), .C1(n4803), .C2(keyinput249), 
        .A(n4802), .ZN(n4808) );
  AOI22_X1 U5343 ( .A1(n4806), .A2(keyinput233), .B1(n4970), .B2(keyinput177), 
        .ZN(n4805) );
  OAI221_X1 U5344 ( .B1(n4806), .B2(keyinput233), .C1(n4970), .C2(keyinput177), 
        .A(n4805), .ZN(n4807) );
  NOR4_X1 U5345 ( .A1(n4810), .A2(n4809), .A3(n4808), .A4(n4807), .ZN(n4822)
         );
  AOI22_X1 U5346 ( .A1(n4965), .A2(keyinput155), .B1(keyinput216), .B2(n4901), 
        .ZN(n4811) );
  OAI221_X1 U5347 ( .B1(n4965), .B2(keyinput155), .C1(n4901), .C2(keyinput216), 
        .A(n4811), .ZN(n4820) );
  AOI22_X1 U5348 ( .A1(n3574), .A2(keyinput252), .B1(n4427), .B2(keyinput168), 
        .ZN(n4812) );
  OAI221_X1 U5349 ( .B1(n3574), .B2(keyinput252), .C1(n4427), .C2(keyinput168), 
        .A(n4812), .ZN(n4819) );
  AOI22_X1 U5350 ( .A1(n4814), .A2(keyinput220), .B1(n4905), .B2(keyinput204), 
        .ZN(n4813) );
  OAI221_X1 U5351 ( .B1(n4814), .B2(keyinput220), .C1(n4905), .C2(keyinput204), 
        .A(n4813), .ZN(n4818) );
  AOI22_X1 U5352 ( .A1(n4074), .A2(keyinput212), .B1(n4816), .B2(keyinput132), 
        .ZN(n4815) );
  OAI221_X1 U5353 ( .B1(n4074), .B2(keyinput212), .C1(n4816), .C2(keyinput132), 
        .A(n4815), .ZN(n4817) );
  NOR4_X1 U5354 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4821)
         );
  NAND4_X1 U5355 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .ZN(n4872)
         );
  INV_X1 U5356 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4919) );
  INV_X1 U5357 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5358 ( .A1(n4919), .A2(keyinput235), .B1(n4826), .B2(keyinput209), 
        .ZN(n4825) );
  OAI221_X1 U5359 ( .B1(n4919), .B2(keyinput235), .C1(n4826), .C2(keyinput209), 
        .A(n4825), .ZN(n4834) );
  INV_X1 U5360 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4920) );
  AOI22_X1 U5361 ( .A1(n4920), .A2(keyinput234), .B1(n4828), .B2(keyinput214), 
        .ZN(n4827) );
  OAI221_X1 U5362 ( .B1(n4920), .B2(keyinput234), .C1(n4828), .C2(keyinput214), 
        .A(n4827), .ZN(n4833) );
  AOI22_X1 U5363 ( .A1(n4891), .A2(keyinput164), .B1(n4389), .B2(keyinput140), 
        .ZN(n4829) );
  OAI221_X1 U5364 ( .B1(n4891), .B2(keyinput164), .C1(n4389), .C2(keyinput140), 
        .A(n4829), .ZN(n4832) );
  AOI22_X1 U5365 ( .A1(n4377), .A2(keyinput159), .B1(n4366), .B2(keyinput247), 
        .ZN(n4830) );
  OAI221_X1 U5366 ( .B1(n4377), .B2(keyinput159), .C1(n4366), .C2(keyinput247), 
        .A(n4830), .ZN(n4831) );
  NOR4_X1 U5367 ( .A1(n4834), .A2(n4833), .A3(n4832), .A4(n4831), .ZN(n4870)
         );
  INV_X1 U5368 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5369 ( .A1(n4837), .A2(keyinput222), .B1(keyinput193), .B2(n4836), 
        .ZN(n4835) );
  OAI221_X1 U5370 ( .B1(n4837), .B2(keyinput222), .C1(n4836), .C2(keyinput193), 
        .A(n4835), .ZN(n4844) );
  AOI22_X1 U5371 ( .A1(n2536), .A2(keyinput176), .B1(n4944), .B2(keyinput210), 
        .ZN(n4838) );
  OAI221_X1 U5372 ( .B1(n2536), .B2(keyinput176), .C1(n4944), .C2(keyinput210), 
        .A(n4838), .ZN(n4843) );
  AOI22_X1 U5373 ( .A1(n4101), .A2(keyinput147), .B1(n4902), .B2(keyinput208), 
        .ZN(n4839) );
  OAI221_X1 U5374 ( .B1(n4101), .B2(keyinput147), .C1(n4902), .C2(keyinput208), 
        .A(n4839), .ZN(n4842) );
  AOI22_X1 U5375 ( .A1(n4093), .A2(keyinput171), .B1(n4250), .B2(keyinput218), 
        .ZN(n4840) );
  OAI221_X1 U5376 ( .B1(n4093), .B2(keyinput171), .C1(n4250), .C2(keyinput218), 
        .A(n4840), .ZN(n4841) );
  NOR4_X1 U5377 ( .A1(n4844), .A2(n4843), .A3(n4842), .A4(n4841), .ZN(n4869)
         );
  INV_X1 U5378 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U5379 ( .A1(n4941), .A2(keyinput186), .B1(keyinput183), .B2(n4221), 
        .ZN(n4845) );
  OAI221_X1 U5380 ( .B1(n4941), .B2(keyinput186), .C1(n4221), .C2(keyinput183), 
        .A(n4845), .ZN(n4856) );
  AOI22_X1 U5381 ( .A1(n4146), .A2(keyinput128), .B1(keyinput199), .B2(n4143), 
        .ZN(n4846) );
  OAI221_X1 U5382 ( .B1(n4146), .B2(keyinput128), .C1(n4143), .C2(keyinput199), 
        .A(n4846), .ZN(n4855) );
  INV_X1 U5383 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4849) );
  INV_X1 U5384 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4848) );
  AOI22_X1 U5385 ( .A1(n4849), .A2(keyinput173), .B1(keyinput231), .B2(n4848), 
        .ZN(n4847) );
  OAI221_X1 U5386 ( .B1(n4849), .B2(keyinput173), .C1(n4848), .C2(keyinput231), 
        .A(n4847), .ZN(n4854) );
  INV_X1 U5387 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U5388 ( .A1(n4852), .A2(keyinput187), .B1(keyinput182), .B2(n4851), 
        .ZN(n4850) );
  OAI221_X1 U5389 ( .B1(n4852), .B2(keyinput187), .C1(n4851), .C2(keyinput182), 
        .A(n4850), .ZN(n4853) );
  NOR4_X1 U5390 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n4868)
         );
  INV_X1 U5391 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4858) );
  AOI22_X1 U5392 ( .A1(n4968), .A2(keyinput146), .B1(keyinput167), .B2(n4858), 
        .ZN(n4857) );
  OAI221_X1 U5393 ( .B1(n4968), .B2(keyinput146), .C1(n4858), .C2(keyinput167), 
        .A(n4857), .ZN(n4866) );
  AOI22_X1 U5394 ( .A1(n4860), .A2(keyinput251), .B1(n2678), .B2(keyinput229), 
        .ZN(n4859) );
  OAI221_X1 U5395 ( .B1(n4860), .B2(keyinput251), .C1(n2678), .C2(keyinput229), 
        .A(n4859), .ZN(n4865) );
  AOI22_X1 U5396 ( .A1(n4879), .A2(keyinput241), .B1(n4904), .B2(keyinput180), 
        .ZN(n4861) );
  OAI221_X1 U5397 ( .B1(n4879), .B2(keyinput241), .C1(n4904), .C2(keyinput180), 
        .A(n4861), .ZN(n4864) );
  AOI22_X1 U5398 ( .A1(n4942), .A2(keyinput195), .B1(keyinput174), .B2(n4955), 
        .ZN(n4862) );
  OAI221_X1 U5399 ( .B1(n4942), .B2(keyinput195), .C1(n4955), .C2(keyinput174), 
        .A(n4862), .ZN(n4863) );
  NOR4_X1 U5400 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n4867)
         );
  NAND4_X1 U5401 ( .A1(n4870), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(n4871)
         );
  NOR4_X1 U5402 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(n5075)
         );
  AOI22_X1 U5403 ( .A1(REG1_REG_11__SCAN_IN), .A2(keyinput9), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput1), .ZN(n4875) );
  OAI221_X1 U5404 ( .B1(REG1_REG_11__SCAN_IN), .B2(keyinput9), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput1), .A(n4875), .ZN(n4883) );
  AOI22_X1 U5405 ( .A1(REG2_REG_0__SCAN_IN), .A2(keyinput65), .B1(
        IR_REG_13__SCAN_IN), .B2(keyinput61), .ZN(n4876) );
  OAI221_X1 U5406 ( .B1(REG2_REG_0__SCAN_IN), .B2(keyinput65), .C1(
        IR_REG_13__SCAN_IN), .C2(keyinput61), .A(n4876), .ZN(n4882) );
  AOI22_X1 U5407 ( .A1(ADDR_REG_16__SCAN_IN), .A2(keyinput45), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput57), .ZN(n4877) );
  OAI221_X1 U5408 ( .B1(ADDR_REG_16__SCAN_IN), .B2(keyinput45), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput57), .A(n4877), .ZN(n4881) );
  AOI22_X1 U5409 ( .A1(n4879), .A2(keyinput113), .B1(n2678), .B2(keyinput101), 
        .ZN(n4878) );
  OAI221_X1 U5410 ( .B1(n4879), .B2(keyinput113), .C1(n2678), .C2(keyinput101), 
        .A(n4878), .ZN(n4880) );
  NOR4_X1 U5411 ( .A1(n4883), .A2(n4882), .A3(n4881), .A4(n4880), .ZN(n4931)
         );
  INV_X1 U5412 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U5413 ( .A1(n4886), .A2(keyinput125), .B1(n4885), .B2(keyinput117), 
        .ZN(n4884) );
  OAI221_X1 U5414 ( .B1(n4886), .B2(keyinput125), .C1(n4885), .C2(keyinput117), 
        .A(n4884), .ZN(n4897) );
  AOI22_X1 U5415 ( .A1(n4889), .A2(keyinput28), .B1(n4888), .B2(keyinput20), 
        .ZN(n4887) );
  OAI221_X1 U5416 ( .B1(n4889), .B2(keyinput28), .C1(n4888), .C2(keyinput20), 
        .A(n4887), .ZN(n4896) );
  AOI22_X1 U5417 ( .A1(n4891), .A2(keyinput36), .B1(n2491), .B2(keyinput24), 
        .ZN(n4890) );
  OAI221_X1 U5418 ( .B1(n4891), .B2(keyinput36), .C1(n2491), .C2(keyinput24), 
        .A(n4890), .ZN(n4895) );
  AOI22_X1 U5419 ( .A1(n4427), .A2(keyinput40), .B1(keyinput44), .B2(n4893), 
        .ZN(n4892) );
  OAI221_X1 U5420 ( .B1(n4427), .B2(keyinput40), .C1(n4893), .C2(keyinput44), 
        .A(n4892), .ZN(n4894) );
  NOR4_X1 U5421 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4930)
         );
  AOI22_X1 U5422 ( .A1(n2882), .A2(keyinput100), .B1(n4899), .B2(keyinput96), 
        .ZN(n4898) );
  OAI221_X1 U5423 ( .B1(n2882), .B2(keyinput100), .C1(n4899), .C2(keyinput96), 
        .A(n4898), .ZN(n4911) );
  AOI22_X1 U5424 ( .A1(n4902), .A2(keyinput80), .B1(keyinput88), .B2(n4901), 
        .ZN(n4900) );
  OAI221_X1 U5425 ( .B1(n4902), .B2(keyinput80), .C1(n4901), .C2(keyinput88), 
        .A(n4900), .ZN(n4910) );
  AOI22_X1 U5426 ( .A1(n2536), .A2(keyinput48), .B1(n4904), .B2(keyinput52), 
        .ZN(n4903) );
  OAI221_X1 U5427 ( .B1(n2536), .B2(keyinput48), .C1(n4904), .C2(keyinput52), 
        .A(n4903), .ZN(n4909) );
  XOR2_X1 U5428 ( .A(n4905), .B(keyinput76), .Z(n4907) );
  XNOR2_X1 U5429 ( .A(IR_REG_24__SCAN_IN), .B(keyinput68), .ZN(n4906) );
  NAND2_X1 U5430 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  NOR4_X1 U5431 ( .A1(n4911), .A2(n4910), .A3(n4909), .A4(n4908), .ZN(n4929)
         );
  INV_X1 U5432 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4913) );
  AOI22_X1 U5433 ( .A1(n4914), .A2(keyinput64), .B1(keyinput127), .B2(n4913), 
        .ZN(n4912) );
  OAI221_X1 U5434 ( .B1(n4914), .B2(keyinput64), .C1(n4913), .C2(keyinput127), 
        .A(n4912), .ZN(n4927) );
  AOI22_X1 U5435 ( .A1(n4917), .A2(keyinput118), .B1(keyinput115), .B2(n4916), 
        .ZN(n4915) );
  OAI221_X1 U5436 ( .B1(n4917), .B2(keyinput118), .C1(n4916), .C2(keyinput115), 
        .A(n4915), .ZN(n4926) );
  AOI22_X1 U5437 ( .A1(n4920), .A2(keyinput106), .B1(n4919), .B2(keyinput107), 
        .ZN(n4918) );
  OAI221_X1 U5438 ( .B1(n4920), .B2(keyinput106), .C1(n4919), .C2(keyinput107), 
        .A(n4918), .ZN(n4925) );
  INV_X1 U5439 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4923) );
  INV_X1 U5440 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4922) );
  AOI22_X1 U5441 ( .A1(n4923), .A2(keyinput98), .B1(keyinput99), .B2(n4922), 
        .ZN(n4921) );
  OAI221_X1 U5442 ( .B1(n4923), .B2(keyinput98), .C1(n4922), .C2(keyinput99), 
        .A(n4921), .ZN(n4924) );
  NOR4_X1 U5443 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n4928)
         );
  NAND4_X1 U5444 ( .A1(n4931), .A2(n4930), .A3(n4929), .A4(n4928), .ZN(n5074)
         );
  AOI22_X1 U5445 ( .A1(n4934), .A2(keyinput75), .B1(n4933), .B2(keyinput70), 
        .ZN(n4932) );
  OAI221_X1 U5446 ( .B1(n4934), .B2(keyinput75), .C1(n4933), .C2(keyinput70), 
        .A(n4932), .ZN(n4939) );
  XNOR2_X1 U5447 ( .A(n4935), .B(keyinput74), .ZN(n4938) );
  XNOR2_X1 U5448 ( .A(n4936), .B(keyinput83), .ZN(n4937) );
  OR3_X1 U5449 ( .A1(n4939), .A2(n4938), .A3(n4937), .ZN(n4947) );
  AOI22_X1 U5450 ( .A1(n4942), .A2(keyinput67), .B1(keyinput58), .B2(n4941), 
        .ZN(n4940) );
  OAI221_X1 U5451 ( .B1(n4942), .B2(keyinput67), .C1(n4941), .C2(keyinput58), 
        .A(n4940), .ZN(n4946) );
  AOI22_X1 U5452 ( .A1(n4944), .A2(keyinput82), .B1(n2774), .B2(keyinput87), 
        .ZN(n4943) );
  OAI221_X1 U5453 ( .B1(n4944), .B2(keyinput82), .C1(n2774), .C2(keyinput87), 
        .A(n4943), .ZN(n4945) );
  NOR3_X1 U5454 ( .A1(n4947), .A2(n4946), .A3(n4945), .ZN(n4997) );
  AOI22_X1 U5455 ( .A1(n4949), .A2(keyinput63), .B1(keyinput55), .B2(n4221), 
        .ZN(n4948) );
  OAI221_X1 U5456 ( .B1(n4949), .B2(keyinput63), .C1(n4221), .C2(keyinput55), 
        .A(n4948), .ZN(n4962) );
  AOI22_X1 U5457 ( .A1(n4952), .A2(keyinput50), .B1(n4951), .B2(keyinput51), 
        .ZN(n4950) );
  OAI221_X1 U5458 ( .B1(n4952), .B2(keyinput50), .C1(n4951), .C2(keyinput51), 
        .A(n4950), .ZN(n4961) );
  AOI22_X1 U5459 ( .A1(n4955), .A2(keyinput46), .B1(keyinput34), .B2(n4954), 
        .ZN(n4953) );
  OAI221_X1 U5460 ( .B1(n4955), .B2(keyinput46), .C1(n4954), .C2(keyinput34), 
        .A(n4953), .ZN(n4960) );
  INV_X1 U5461 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U5462 ( .A1(n4958), .A2(keyinput26), .B1(keyinput30), .B2(n4957), 
        .ZN(n4956) );
  OAI221_X1 U5463 ( .B1(n4958), .B2(keyinput26), .C1(n4957), .C2(keyinput30), 
        .A(n4956), .ZN(n4959) );
  NOR4_X1 U5464 ( .A1(n4962), .A2(n4961), .A3(n4960), .A4(n4959), .ZN(n4996)
         );
  INV_X1 U5465 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U5466 ( .A1(n4965), .A2(keyinput27), .B1(keyinput14), .B2(n4964), 
        .ZN(n4963) );
  OAI221_X1 U5467 ( .B1(n4965), .B2(keyinput27), .C1(n4964), .C2(keyinput14), 
        .A(n4963), .ZN(n4977) );
  AOI22_X1 U5468 ( .A1(n4968), .A2(keyinput18), .B1(n4967), .B2(keyinput2), 
        .ZN(n4966) );
  OAI221_X1 U5469 ( .B1(n4968), .B2(keyinput18), .C1(n4967), .C2(keyinput2), 
        .A(n4966), .ZN(n4976) );
  AOI22_X1 U5470 ( .A1(n2560), .A2(keyinput7), .B1(keyinput49), .B2(n4970), 
        .ZN(n4969) );
  OAI221_X1 U5471 ( .B1(n2560), .B2(keyinput7), .C1(n4970), .C2(keyinput49), 
        .A(n4969), .ZN(n4975) );
  AOI22_X1 U5472 ( .A1(n4973), .A2(keyinput37), .B1(n4972), .B2(keyinput25), 
        .ZN(n4971) );
  OAI221_X1 U5473 ( .B1(n4973), .B2(keyinput37), .C1(n4972), .C2(keyinput25), 
        .A(n4971), .ZN(n4974) );
  NOR4_X1 U5474 ( .A1(n4977), .A2(n4976), .A3(n4975), .A4(n4974), .ZN(n4995)
         );
  AOI22_X1 U5475 ( .A1(n4980), .A2(keyinput21), .B1(keyinput5), .B2(n4979), 
        .ZN(n4978) );
  OAI221_X1 U5476 ( .B1(n4980), .B2(keyinput21), .C1(n4979), .C2(keyinput5), 
        .A(n4978), .ZN(n4993) );
  INV_X1 U5477 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4982) );
  AOI22_X1 U5478 ( .A1(n4983), .A2(keyinput33), .B1(n4982), .B2(keyinput73), 
        .ZN(n4981) );
  OAI221_X1 U5479 ( .B1(n4983), .B2(keyinput33), .C1(n4982), .C2(keyinput73), 
        .A(n4981), .ZN(n4992) );
  INV_X1 U5480 ( .A(DATAI_6_), .ZN(n4986) );
  AOI22_X1 U5481 ( .A1(n4986), .A2(keyinput53), .B1(n4985), .B2(keyinput13), 
        .ZN(n4984) );
  OAI221_X1 U5482 ( .B1(n4986), .B2(keyinput53), .C1(n4985), .C2(keyinput13), 
        .A(n4984), .ZN(n4991) );
  XOR2_X1 U5483 ( .A(n4987), .B(keyinput69), .Z(n4989) );
  XNOR2_X1 U5484 ( .A(IR_REG_9__SCAN_IN), .B(keyinput93), .ZN(n4988) );
  NAND2_X1 U5485 ( .A1(n4989), .A2(n4988), .ZN(n4990) );
  NOR4_X1 U5486 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n4994)
         );
  NAND4_X1 U5487 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), .ZN(n5073)
         );
  OAI22_X1 U5488 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput56), .B1(
        REG3_REG_0__SCAN_IN), .B2(keyinput8), .ZN(n4998) );
  AOI221_X1 U5489 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput56), .C1(keyinput8), 
        .C2(REG3_REG_0__SCAN_IN), .A(n4998), .ZN(n5005) );
  OAI22_X1 U5490 ( .A1(REG2_REG_27__SCAN_IN), .A2(keyinput72), .B1(keyinput17), 
        .B2(DATAI_1_), .ZN(n4999) );
  AOI221_X1 U5491 ( .B1(REG2_REG_27__SCAN_IN), .B2(keyinput72), .C1(DATAI_1_), 
        .C2(keyinput17), .A(n4999), .ZN(n5004) );
  OAI22_X1 U5492 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput60), .B1(keyinput4), 
        .B2(REG1_REG_10__SCAN_IN), .ZN(n5000) );
  AOI221_X1 U5493 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput60), .C1(
        REG1_REG_10__SCAN_IN), .C2(keyinput4), .A(n5000), .ZN(n5003) );
  OAI22_X1 U5494 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput32), .B1(
        ADDR_REG_12__SCAN_IN), .B2(keyinput16), .ZN(n5001) );
  AOI221_X1 U5495 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput32), .C1(keyinput16), .C2(ADDR_REG_12__SCAN_IN), .A(n5001), .ZN(n5002) );
  NAND4_X1 U5496 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n5033)
         );
  OAI22_X1 U5497 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput108), .B1(DATAI_0_), 
        .B2(keyinput104), .ZN(n5006) );
  AOI221_X1 U5498 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput108), .C1(keyinput104), 
        .C2(DATAI_0_), .A(n5006), .ZN(n5013) );
  OAI22_X1 U5499 ( .A1(REG1_REG_7__SCAN_IN), .A2(keyinput84), .B1(keyinput103), 
        .B2(ADDR_REG_15__SCAN_IN), .ZN(n5007) );
  AOI221_X1 U5500 ( .B1(REG1_REG_7__SCAN_IN), .B2(keyinput84), .C1(
        ADDR_REG_15__SCAN_IN), .C2(keyinput103), .A(n5007), .ZN(n5012) );
  OAI22_X1 U5501 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput120), .B1(keyinput92), 
        .B2(REG0_REG_30__SCAN_IN), .ZN(n5008) );
  AOI221_X1 U5502 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput120), .C1(
        REG0_REG_30__SCAN_IN), .C2(keyinput92), .A(n5008), .ZN(n5011) );
  OAI22_X1 U5503 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput116), .B1(keyinput124), 
        .B2(REG0_REG_15__SCAN_IN), .ZN(n5009) );
  AOI221_X1 U5504 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput116), .C1(
        REG0_REG_15__SCAN_IN), .C2(keyinput124), .A(n5009), .ZN(n5010) );
  NAND4_X1 U5505 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n5032)
         );
  OAI22_X1 U5506 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput121), .B1(keyinput109), .B2(DATAI_18_), .ZN(n5014) );
  AOI221_X1 U5507 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput121), .C1(DATAI_18_), 
        .C2(keyinput109), .A(n5014), .ZN(n5021) );
  OAI22_X1 U5508 ( .A1(REG1_REG_16__SCAN_IN), .A2(keyinput81), .B1(keyinput77), 
        .B2(REG0_REG_6__SCAN_IN), .ZN(n5015) );
  AOI221_X1 U5509 ( .B1(REG1_REG_16__SCAN_IN), .B2(keyinput81), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput77), .A(n5015), .ZN(n5020) );
  OAI22_X1 U5510 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput41), .B1(keyinput29), 
        .B2(REG0_REG_26__SCAN_IN), .ZN(n5016) );
  AOI221_X1 U5511 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput41), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput29), .A(n5016), .ZN(n5019) );
  OAI22_X1 U5512 ( .A1(REG2_REG_6__SCAN_IN), .A2(keyinput97), .B1(
        REG0_REG_2__SCAN_IN), .B2(keyinput105), .ZN(n5017) );
  AOI221_X1 U5513 ( .B1(REG2_REG_6__SCAN_IN), .B2(keyinput97), .C1(keyinput105), .C2(REG0_REG_2__SCAN_IN), .A(n5017), .ZN(n5018) );
  NAND4_X1 U5514 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n5031)
         );
  OAI22_X1 U5515 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput11), .B1(
        REG0_REG_19__SCAN_IN), .B2(keyinput23), .ZN(n5022) );
  AOI221_X1 U5516 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput11), .C1(keyinput23), 
        .C2(REG0_REG_19__SCAN_IN), .A(n5022), .ZN(n5029) );
  OAI22_X1 U5517 ( .A1(REG1_REG_21__SCAN_IN), .A2(keyinput12), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput15), .ZN(n5023) );
  AOI221_X1 U5518 ( .B1(REG1_REG_21__SCAN_IN), .B2(keyinput12), .C1(keyinput15), .C2(DATAO_REG_8__SCAN_IN), .A(n5023), .ZN(n5028) );
  OAI22_X1 U5519 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput89), .B1(keyinput85), 
        .B2(DATAI_20_), .ZN(n5024) );
  AOI221_X1 U5520 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput89), .C1(DATAI_20_), 
        .C2(keyinput85), .A(n5024), .ZN(n5027) );
  OAI22_X1 U5521 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput19), .B1(
        DATAO_REG_10__SCAN_IN), .B2(keyinput3), .ZN(n5025) );
  AOI221_X1 U5522 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput19), .C1(keyinput3), 
        .C2(DATAO_REG_10__SCAN_IN), .A(n5025), .ZN(n5026) );
  NAND4_X1 U5523 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n5030)
         );
  NOR4_X1 U5524 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5071)
         );
  OAI22_X1 U5525 ( .A1(DATAI_14_), .A2(keyinput62), .B1(DATAO_REG_7__SCAN_IN), 
        .B2(keyinput54), .ZN(n5034) );
  AOI221_X1 U5526 ( .B1(DATAI_14_), .B2(keyinput62), .C1(keyinput54), .C2(
        DATAO_REG_7__SCAN_IN), .A(n5034), .ZN(n5041) );
  OAI22_X1 U5527 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput78), .B1(
        D_REG_10__SCAN_IN), .B2(keyinput66), .ZN(n5035) );
  AOI221_X1 U5528 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput78), .C1(keyinput66), 
        .C2(D_REG_10__SCAN_IN), .A(n5035), .ZN(n5040) );
  OAI22_X1 U5529 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput22), .B1(
        REG2_REG_15__SCAN_IN), .B2(keyinput10), .ZN(n5036) );
  AOI221_X1 U5530 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput22), .C1(keyinput10), 
        .C2(REG2_REG_15__SCAN_IN), .A(n5036), .ZN(n5039) );
  OAI22_X1 U5531 ( .A1(DATAI_29_), .A2(keyinput42), .B1(DATAI_5_), .B2(
        keyinput38), .ZN(n5037) );
  AOI221_X1 U5532 ( .B1(DATAI_29_), .B2(keyinput42), .C1(keyinput38), .C2(
        DATAI_5_), .A(n5037), .ZN(n5038) );
  NAND4_X1 U5533 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n5069)
         );
  OAI22_X1 U5534 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput126), .B1(keyinput122), 
        .B2(REG3_REG_10__SCAN_IN), .ZN(n5042) );
  AOI221_X1 U5535 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput126), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput122), .A(n5042), .ZN(n5049) );
  OAI22_X1 U5536 ( .A1(DATAI_13_), .A2(keyinput110), .B1(keyinput114), .B2(
        REG1_REG_1__SCAN_IN), .ZN(n5043) );
  AOI221_X1 U5537 ( .B1(DATAI_13_), .B2(keyinput110), .C1(REG1_REG_1__SCAN_IN), 
        .C2(keyinput114), .A(n5043), .ZN(n5048) );
  OAI22_X1 U5538 ( .A1(REG2_REG_23__SCAN_IN), .A2(keyinput90), .B1(
        REG1_REG_17__SCAN_IN), .B2(keyinput86), .ZN(n5044) );
  AOI221_X1 U5539 ( .B1(REG2_REG_23__SCAN_IN), .B2(keyinput90), .C1(keyinput86), .C2(REG1_REG_17__SCAN_IN), .A(n5044), .ZN(n5047) );
  OAI22_X1 U5540 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput102), .B1(
        REG1_REG_26__SCAN_IN), .B2(keyinput94), .ZN(n5045) );
  AOI221_X1 U5541 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput102), .C1(keyinput94), 
        .C2(REG1_REG_26__SCAN_IN), .A(n5045), .ZN(n5046) );
  NAND4_X1 U5542 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n5068)
         );
  OAI22_X1 U5543 ( .A1(REG2_REG_29__SCAN_IN), .A2(keyinput0), .B1(keyinput123), 
        .B2(DATAO_REG_20__SCAN_IN), .ZN(n5050) );
  AOI221_X1 U5544 ( .B1(REG2_REG_29__SCAN_IN), .B2(keyinput0), .C1(
        DATAO_REG_20__SCAN_IN), .C2(keyinput123), .A(n5050), .ZN(n5057) );
  OAI22_X1 U5545 ( .A1(REG1_REG_25__SCAN_IN), .A2(keyinput119), .B1(keyinput39), .B2(DATAO_REG_26__SCAN_IN), .ZN(n5051) );
  AOI221_X1 U5546 ( .B1(REG1_REG_25__SCAN_IN), .B2(keyinput119), .C1(
        DATAO_REG_26__SCAN_IN), .C2(keyinput39), .A(n5051), .ZN(n5056) );
  OAI22_X1 U5547 ( .A1(REG1_REG_29__SCAN_IN), .A2(keyinput91), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput111), .ZN(n5052) );
  AOI221_X1 U5548 ( .B1(REG1_REG_29__SCAN_IN), .B2(keyinput91), .C1(
        keyinput111), .C2(IR_REG_0__SCAN_IN), .A(n5052), .ZN(n5055) );
  OAI22_X1 U5549 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput112), .B1(DATAI_4_), 
        .B2(keyinput95), .ZN(n5053) );
  AOI221_X1 U5550 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput112), .C1(keyinput95), 
        .C2(DATAI_4_), .A(n5053), .ZN(n5054) );
  NAND4_X1 U5551 ( .A1(n5057), .A2(n5056), .A3(n5055), .A4(n5054), .ZN(n5067)
         );
  OAI22_X1 U5552 ( .A1(REG2_REG_31__SCAN_IN), .A2(keyinput71), .B1(keyinput47), 
        .B2(ADDR_REG_8__SCAN_IN), .ZN(n5058) );
  AOI221_X1 U5553 ( .B1(REG2_REG_31__SCAN_IN), .B2(keyinput71), .C1(
        ADDR_REG_8__SCAN_IN), .C2(keyinput47), .A(n5058), .ZN(n5065) );
  OAI22_X1 U5554 ( .A1(REG0_REG_12__SCAN_IN), .A2(keyinput6), .B1(
        ADDR_REG_4__SCAN_IN), .B2(keyinput59), .ZN(n5059) );
  AOI221_X1 U5555 ( .B1(REG0_REG_12__SCAN_IN), .B2(keyinput6), .C1(keyinput59), 
        .C2(ADDR_REG_4__SCAN_IN), .A(n5059), .ZN(n5064) );
  OAI22_X1 U5556 ( .A1(REG1_REG_23__SCAN_IN), .A2(keyinput31), .B1(
        REG2_REG_18__SCAN_IN), .B2(keyinput43), .ZN(n5060) );
  AOI221_X1 U5557 ( .B1(REG1_REG_23__SCAN_IN), .B2(keyinput31), .C1(keyinput43), .C2(REG2_REG_18__SCAN_IN), .A(n5060), .ZN(n5063) );
  OAI22_X1 U5558 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput79), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput35), .ZN(n5061) );
  AOI221_X1 U5559 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput79), .C1(keyinput35), 
        .C2(D_REG_8__SCAN_IN), .A(n5061), .ZN(n5062) );
  NAND4_X1 U5560 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n5066)
         );
  NOR4_X1 U5561 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n5070)
         );
  NAND2_X1 U5562 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  NOR4_X1 U5563 ( .A1(n5075), .A2(n5074), .A3(n5073), .A4(n5072), .ZN(n5079)
         );
  NAND2_X1 U5564 ( .A1(n5076), .A2(U4043), .ZN(n5077) );
  OAI21_X1 U5565 ( .B1(U4043), .B2(DATAO_REG_26__SCAN_IN), .A(n5077), .ZN(
        n5078) );
  XNOR2_X1 U5566 ( .A(n5079), .B(n5078), .ZN(U3576) );
  CLKBUF_X1 U2471 ( .A(n2750), .Z(n2827) );
  CLKBUF_X2 U2474 ( .A(n2550), .Z(n2766) );
  CLKBUF_X1 U2476 ( .A(n4055), .Z(n2228) );
endmodule

