

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10965, n10966, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246;

  NAND2_X1 U11072 ( .A1(n15672), .A2(n11080), .ZN(n15618) );
  NAND2_X1 U11073 ( .A1(n16470), .A2(n11422), .ZN(n16414) );
  OR2_X1 U11074 ( .A1(n16265), .A2(n11322), .ZN(n11324) );
  INV_X2 U11075 ( .A(n20269), .ZN(n20458) );
  NOR2_X1 U11076 ( .A1(n18176), .A2(n20814), .ZN(n18175) );
  INV_X1 U11077 ( .A(n20738), .ZN(n20063) );
  INV_X1 U11078 ( .A(n13390), .ZN(n13273) );
  CLKBUF_X2 U11079 ( .A(n15077), .Z(n10971) );
  INV_X2 U11080 ( .A(n12366), .ZN(n12345) );
  CLKBUF_X2 U11081 ( .A(n15091), .Z(n10970) );
  CLKBUF_X2 U11082 ( .A(n11603), .Z(n12295) );
  NOR2_X1 U11084 ( .A1(n13815), .A2(n14089), .ZN(n14113) );
  CLKBUF_X2 U11086 ( .A(n15077), .Z(n10972) );
  INV_X4 U11087 ( .A(n11019), .ZN(n17740) );
  AND2_X1 U11088 ( .A1(n10989), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12726) );
  NOR2_X2 U11089 ( .A1(n14093), .A2(n21946), .ZN(n13839) );
  NAND2_X1 U11090 ( .A1(n12989), .A2(n12544), .ZN(n13188) );
  AND2_X1 U11091 ( .A1(n15284), .A2(n14293), .ZN(n15415) );
  NOR2_X1 U11092 ( .A1(n20727), .A2(n15041), .ZN(n15066) );
  CLKBUF_X2 U11093 ( .A(n11596), .Z(n12139) );
  AND2_X1 U11094 ( .A1(n16098), .A2(n11537), .ZN(n11687) );
  AND2_X1 U11095 ( .A1(n16098), .A2(n13958), .ZN(n11707) );
  AND2_X1 U11096 ( .A1(n13840), .A2(n16097), .ZN(n11709) );
  AND2_X1 U11097 ( .A1(n13818), .A2(n11543), .ZN(n11665) );
  AND2_X1 U11098 ( .A1(n13818), .A2(n11542), .ZN(n11686) );
  INV_X4 U11099 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12450) );
  CLKBUF_X2 U11100 ( .A(n11591), .Z(n12293) );
  AND2_X1 U11101 ( .A1(n13833), .A2(n11532), .ZN(n11591) );
  CLKBUF_X1 U11103 ( .A(n15588), .Z(n10968) );
  INV_X1 U11104 ( .A(n20714), .ZN(n15040) );
  INV_X1 U11105 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21165) );
  INV_X1 U11106 ( .A(n13785), .ZN(n13878) );
  OR2_X1 U11107 ( .A1(n13580), .A2(n11215), .ZN(n13583) );
  NAND2_X1 U11109 ( .A1(n11127), .A2(n11036), .ZN(n16462) );
  AND2_X1 U11110 ( .A1(n12614), .A2(n12613), .ZN(n19138) );
  CLKBUF_X3 U11111 ( .A(n15066), .Z(n17700) );
  NAND3_X1 U11112 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20721) );
  NAND2_X1 U11113 ( .A1(n11385), .A2(n13579), .ZN(n13580) );
  XNOR2_X1 U11114 ( .A(n14442), .B(n21715), .ZN(n13827) );
  NAND2_X1 U11115 ( .A1(n11868), .A2(n11858), .ZN(n13508) );
  INV_X1 U11116 ( .A(n11645), .ZN(n21667) );
  NOR2_X1 U11117 ( .A1(n16267), .A2(n16266), .ZN(n16265) );
  XNOR2_X1 U11118 ( .A(n13177), .B(n13176), .ZN(n16104) );
  AND2_X1 U11119 ( .A1(n11414), .A2(n11150), .ZN(n11149) );
  INV_X1 U11121 ( .A(n18020), .ZN(n17976) );
  INV_X1 U11122 ( .A(n21068), .ZN(n21142) );
  NOR2_X1 U11123 ( .A1(n18175), .A2(n17808), .ZN(n18163) );
  INV_X2 U11124 ( .A(n15588), .ZN(n15607) );
  INV_X1 U11125 ( .A(n10973), .ZN(n13182) );
  NAND2_X1 U11126 ( .A1(n14033), .A2(n14032), .ZN(n14129) );
  AND2_X1 U11128 ( .A1(n12605), .A2(n12600), .ZN(n18349) );
  NAND2_X1 U11129 ( .A1(n16627), .A2(n11289), .ZN(n16577) );
  AND2_X1 U11130 ( .A1(n21111), .A2(n20063), .ZN(n21182) );
  INV_X1 U11131 ( .A(n18003), .ZN(n18050) );
  INV_X1 U11132 ( .A(n18195), .ZN(n18221) );
  NAND2_X1 U11133 ( .A1(n18021), .A2(n18003), .ZN(n18215) );
  NAND2_X1 U11134 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20713) );
  AOI211_X1 U11135 ( .C1(n17788), .C2(n17785), .A(n15270), .B(n20743), .ZN(
        n21195) );
  INV_X1 U11136 ( .A(n18215), .ZN(n18205) );
  INV_X4 U11137 ( .A(n12935), .ZN(n12969) );
  OR2_X2 U11138 ( .A1(n12590), .A2(n12589), .ZN(n13084) );
  AND2_X1 U11139 ( .A1(n11539), .A2(n16098), .ZN(n11603) );
  INV_X2 U11140 ( .A(n15470), .ZN(n10965) );
  OAI211_X2 U11141 ( .C1(n13444), .C2(n13447), .A(n13445), .B(n15502), .ZN(
        n12981) );
  MUX2_X2 U11142 ( .A(n12472), .B(n12471), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19437) );
  INV_X2 U11143 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10966) );
  AND2_X1 U11144 ( .A1(n13840), .A2(n16098), .ZN(n11702) );
  NAND2_X2 U11145 ( .A1(n11256), .A2(n11255), .ZN(n17587) );
  AND2_X1 U11146 ( .A1(n21946), .A2(n14364), .ZN(n15588) );
  BUF_X4 U11147 ( .A(n15091), .Z(n10969) );
  NOR2_X1 U11148 ( .A1(n15041), .A2(n15039), .ZN(n15091) );
  AND2_X4 U11149 ( .A1(n11458), .A2(n10966), .ZN(n12502) );
  AND2_X2 U11150 ( .A1(n12415), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11458) );
  AOI211_X2 U11151 ( .C1(n16671), .C2(n17273), .A(n16416), .B(n16415), .ZN(
        n16417) );
  NOR2_X1 U11152 ( .A1(n15041), .A2(n15040), .ZN(n15077) );
  INV_X1 U11154 ( .A(n12460), .ZN(n12967) );
  AND2_X4 U11156 ( .A1(n14293), .A2(n10966), .ZN(n12503) );
  INV_X2 U11157 ( .A(n11024), .ZN(n17687) );
  NAND2_X1 U11158 ( .A1(n15513), .A2(n11503), .ZN(n18569) );
  OR2_X1 U11159 ( .A1(n16164), .A2(n16163), .ZN(n16647) );
  OR3_X1 U11160 ( .A1(n21031), .A2(n18037), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17987) );
  NAND2_X1 U11161 ( .A1(n18064), .A2(n17950), .ZN(n18011) );
  INV_X1 U11162 ( .A(n18125), .ZN(n18106) );
  NAND3_X1 U11164 ( .A1(n11026), .A2(n11528), .A3(n11002), .ZN(n12693) );
  INV_X4 U11165 ( .A(n18226), .ZN(n18214) );
  AND2_X2 U11166 ( .A1(n14220), .A2(n11084), .ZN(n16380) );
  NAND2_X1 U11167 ( .A1(n20063), .A2(n21224), .ZN(n18226) );
  AND2_X1 U11168 ( .A1(n11164), .A2(n11163), .ZN(n21162) );
  AND2_X1 U11169 ( .A1(n12598), .A2(n12609), .ZN(n19190) );
  BUF_X1 U11170 ( .A(n13945), .Z(n18624) );
  NOR2_X1 U11172 ( .A1(n14617), .A2(n14470), .ZN(n14834) );
  OAI21_X2 U11173 ( .B1(n20498), .B2(n20497), .A(n20496), .ZN(n20670) );
  NOR2_X1 U11174 ( .A1(n13256), .A2(n13255), .ZN(n14469) );
  AOI21_X1 U11175 ( .B1(n13986), .B2(n11514), .A(n13251), .ZN(n13256) );
  NOR2_X1 U11176 ( .A1(n12809), .A2(n12780), .ZN(n12784) );
  INV_X1 U11177 ( .A(n12586), .ZN(n13171) );
  OR2_X1 U11178 ( .A1(n12547), .A2(n13761), .ZN(n12586) );
  AND3_X1 U11179 ( .A1(n11287), .A2(n13191), .A3(n11286), .ZN(n12556) );
  NAND2_X1 U11180 ( .A1(n14347), .A2(n19594), .ZN(n12547) );
  INV_X2 U11181 ( .A(n20495), .ZN(n20055) );
  NAND2_X1 U11182 ( .A1(n10981), .A2(n12461), .ZN(n13975) );
  INV_X2 U11183 ( .A(n11630), .ZN(n11656) );
  NAND2_X2 U11184 ( .A1(n12458), .A2(n12457), .ZN(n12519) );
  CLKBUF_X2 U11185 ( .A(n19780), .Z(n21230) );
  INV_X1 U11186 ( .A(n10992), .ZN(n10994) );
  CLKBUF_X2 U11187 ( .A(n11686), .Z(n12292) );
  CLKBUF_X1 U11188 ( .A(n12633), .Z(n15283) );
  CLKBUF_X1 U11189 ( .A(n12502), .Z(n15471) );
  INV_X1 U11190 ( .A(n15051), .ZN(n10992) );
  BUF_X4 U11191 ( .A(n15089), .Z(n10976) );
  INV_X2 U11192 ( .A(n12431), .ZN(n10996) );
  INV_X4 U11194 ( .A(n12431), .ZN(n15462) );
  INV_X4 U11195 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11243) );
  INV_X2 U11196 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12415) );
  NOR2_X1 U11197 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20714) );
  INV_X4 U11198 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20712) );
  INV_X2 U11199 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U11200 ( .A1(n11147), .A2(n16516), .ZN(n11146) );
  XNOR2_X1 U11201 ( .A(n16437), .B(n16436), .ZN(n16692) );
  OR2_X1 U11202 ( .A1(n15877), .A2(n11086), .ZN(n11379) );
  NAND2_X1 U11203 ( .A1(n11238), .A2(n11462), .ZN(n16437) );
  AND2_X1 U11204 ( .A1(n11461), .A2(n11459), .ZN(n16421) );
  NOR2_X1 U11205 ( .A1(n11426), .A2(n16710), .ZN(n16453) );
  NAND2_X1 U11206 ( .A1(n16445), .A2(n11462), .ZN(n11461) );
  OR2_X2 U11207 ( .A1(n16499), .A2(n16494), .ZN(n16492) );
  NAND2_X1 U11208 ( .A1(n11324), .A2(n11328), .ZN(n15461) );
  NAND2_X1 U11209 ( .A1(n11417), .A2(n11419), .ZN(n16499) );
  NAND2_X1 U11210 ( .A1(n19944), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13579) );
  NOR2_X1 U11211 ( .A1(n17253), .A2(n13578), .ZN(n19946) );
  NAND2_X1 U11212 ( .A1(n11186), .A2(n11377), .ZN(n17253) );
  XNOR2_X1 U11213 ( .A(n15437), .B(n11512), .ZN(n16267) );
  AND2_X1 U11214 ( .A1(n13458), .A2(n13457), .ZN(n11515) );
  AND2_X1 U11215 ( .A1(n16475), .A2(n16476), .ZN(n16588) );
  OAI21_X1 U11216 ( .B1(n11378), .B2(n11376), .A(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11375) );
  AOI21_X1 U11217 ( .B1(n11413), .B2(n13065), .A(n18597), .ZN(n11412) );
  AND2_X1 U11218 ( .A1(n11204), .A2(n11202), .ZN(n18009) );
  AND2_X1 U11219 ( .A1(n16299), .A2(n11085), .ZN(n16273) );
  NOR2_X1 U11220 ( .A1(n19919), .A2(n11039), .ZN(n11377) );
  NAND2_X1 U11221 ( .A1(n11223), .A2(n18373), .ZN(n12848) );
  NOR2_X1 U11222 ( .A1(n11018), .A2(n16304), .ZN(n16303) );
  INV_X1 U11223 ( .A(n18011), .ZN(n17981) );
  NAND2_X1 U11224 ( .A1(n19883), .A2(n16043), .ZN(n15902) );
  AND2_X1 U11225 ( .A1(n19883), .A2(n21255), .ZN(n15966) );
  OR2_X1 U11226 ( .A1(n15679), .A2(n15551), .ZN(n15657) );
  OR2_X2 U11227 ( .A1(n16335), .A2(n16189), .ZN(n11020) );
  NAND2_X1 U11228 ( .A1(n17952), .A2(n17836), .ZN(n17891) );
  INV_X2 U11229 ( .A(n19894), .ZN(n19945) );
  NAND2_X1 U11230 ( .A1(n18057), .A2(n21034), .ZN(n17952) );
  NAND2_X1 U11231 ( .A1(n11116), .A2(n11115), .ZN(n13070) );
  INV_X2 U11232 ( .A(n13560), .ZN(n19894) );
  NAND2_X1 U11233 ( .A1(n18058), .A2(n21101), .ZN(n18057) );
  NAND2_X1 U11234 ( .A1(n14688), .A2(n14687), .ZN(n14864) );
  AND2_X1 U11235 ( .A1(n11110), .A2(n12846), .ZN(n13071) );
  AND2_X1 U11236 ( .A1(n12930), .A2(n12929), .ZN(n12931) );
  NAND2_X1 U11237 ( .A1(n16766), .A2(n11097), .ZN(n16221) );
  NOR2_X1 U11238 ( .A1(n14649), .A2(n14648), .ZN(n14688) );
  NAND2_X1 U11239 ( .A1(n12739), .A2(n12738), .ZN(n12741) );
  NAND2_X1 U11240 ( .A1(n14459), .A2(n11079), .ZN(n14649) );
  AND2_X1 U11241 ( .A1(n13530), .A2(n13786), .ZN(n13550) );
  OR2_X1 U11242 ( .A1(n12724), .A2(n12723), .ZN(n12739) );
  OR2_X1 U11243 ( .A1(n14263), .A2(n14264), .ZN(n14416) );
  AND3_X1 U11244 ( .A1(n12655), .A2(n12645), .A3(n12646), .ZN(n11026) );
  OR2_X1 U11245 ( .A1(n14224), .A2(n14223), .ZN(n14263) );
  NAND2_X1 U11246 ( .A1(n11433), .A2(n11435), .ZN(n21752) );
  NAND2_X1 U11247 ( .A1(n14017), .A2(n14016), .ZN(n14353) );
  AND2_X1 U11248 ( .A1(n12603), .A2(n18624), .ZN(n19121) );
  AND2_X1 U11249 ( .A1(n12603), .A2(n12609), .ZN(n19160) );
  NAND2_X1 U11250 ( .A1(n11784), .A2(n11783), .ZN(n11856) );
  NAND2_X1 U11251 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18145), .ZN(
        n17820) );
  AND2_X1 U11252 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  OR2_X2 U11253 ( .A1(n21227), .A2(n14359), .ZN(n14663) );
  CLKBUF_X1 U11254 ( .A(n13827), .Z(n21753) );
  NAND2_X1 U11255 ( .A1(n13949), .A2(n13948), .ZN(n14015) );
  NOR2_X1 U11256 ( .A1(n16129), .A2(n16128), .ZN(n16130) );
  INV_X1 U11257 ( .A(n21179), .ZN(n21019) );
  NAND2_X1 U11258 ( .A1(n20738), .A2(n21111), .ZN(n21179) );
  NOR2_X2 U11259 ( .A1(n21085), .A2(n21184), .ZN(n21111) );
  NAND2_X1 U11260 ( .A1(n11846), .A2(n11845), .ZN(n13484) );
  NAND2_X1 U11261 ( .A1(n12599), .A2(n12608), .ZN(n16241) );
  NOR2_X1 U11262 ( .A1(n11496), .A2(n11495), .ZN(n11494) );
  OR2_X2 U11263 ( .A1(n13660), .A2(n14364), .ZN(n13884) );
  XNOR2_X1 U11264 ( .A(n13772), .B(n13950), .ZN(n13766) );
  NAND2_X1 U11265 ( .A1(n11845), .A2(n11720), .ZN(n11834) );
  NAND2_X1 U11266 ( .A1(n12871), .A2(n12872), .ZN(n12878) );
  NOR2_X2 U11267 ( .A1(n16352), .A2(n19591), .ZN(n14780) );
  NOR2_X2 U11268 ( .A1(n14748), .A2(n19591), .ZN(n14749) );
  NOR2_X2 U11269 ( .A1(n14754), .A2(n19591), .ZN(n14755) );
  INV_X1 U11270 ( .A(n12594), .ZN(n12606) );
  NOR2_X2 U11271 ( .A1(n16365), .A2(n19591), .ZN(n14600) );
  AND2_X2 U11272 ( .A1(n12381), .A2(n12380), .ZN(n15546) );
  INV_X2 U11273 ( .A(n16284), .ZN(n14161) );
  INV_X1 U11274 ( .A(n18349), .ZN(n18587) );
  NOR2_X1 U11275 ( .A1(n13085), .A2(n11499), .ZN(n11498) );
  NAND2_X1 U11276 ( .A1(n11155), .A2(n11154), .ZN(n12580) );
  NAND2_X1 U11277 ( .A1(n20696), .A2(n20012), .ZN(n16991) );
  OR2_X1 U11278 ( .A1(n12593), .A2(n12592), .ZN(n12600) );
  NAND3_X1 U11279 ( .A1(n11120), .A2(n12565), .A3(n12566), .ZN(n12592) );
  OAI221_X2 U11280 ( .B1(n20692), .B2(n20690), .C1(n20692), .C2(n20689), .A(
        n17783), .ZN(n21068) );
  OR2_X1 U11281 ( .A1(n13256), .A2(n13252), .ZN(n14473) );
  NAND2_X1 U11282 ( .A1(n12576), .A2(n11157), .ZN(n11156) );
  NOR2_X1 U11283 ( .A1(n12849), .A2(n11244), .ZN(n12857) );
  AND2_X1 U11284 ( .A1(n11122), .A2(n11083), .ZN(n12534) );
  OAI211_X1 U11285 ( .C1(n17020), .C2(n11664), .A(n13813), .B(n11663), .ZN(
        n11727) );
  AND2_X1 U11286 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  OAI211_X2 U11287 ( .C1(n11493), .C2(n18340), .A(n12554), .B(n11492), .ZN(
        n12582) );
  INV_X2 U11288 ( .A(n13099), .ZN(n13161) );
  AND2_X1 U11289 ( .A1(n12575), .A2(n11032), .ZN(n11157) );
  INV_X2 U11290 ( .A(n13171), .ZN(n13169) );
  NAND2_X1 U11291 ( .A1(n12791), .A2(n12790), .ZN(n12809) );
  INV_X2 U11292 ( .A(n13099), .ZN(n10978) );
  AND2_X1 U11293 ( .A1(n12803), .A2(n12802), .ZN(n12791) );
  OR2_X1 U11294 ( .A1(n10988), .A2(n12577), .ZN(n11032) );
  NOR2_X1 U11295 ( .A1(n12586), .A2(n12548), .ZN(n12549) );
  CLKBUF_X1 U11296 ( .A(n13628), .Z(n15538) );
  AND2_X1 U11297 ( .A1(n13968), .A2(n13967), .ZN(n13247) );
  NOR2_X1 U11298 ( .A1(n15253), .A2(n11274), .ZN(n15243) );
  OAI21_X1 U11299 ( .B1(n15269), .B2(n11047), .A(n15242), .ZN(n15253) );
  NAND2_X1 U11300 ( .A1(n12561), .A2(n11287), .ZN(n11493) );
  NAND2_X1 U11301 ( .A1(n11471), .A2(n13238), .ZN(n13967) );
  MUX2_X1 U11302 ( .A(n12545), .B(n13186), .S(n19437), .Z(n12561) );
  AND2_X1 U11303 ( .A1(n11254), .A2(n17794), .ZN(n17797) );
  NAND2_X1 U11304 ( .A1(n11636), .A2(n11635), .ZN(n11653) );
  NAND2_X1 U11305 ( .A1(n11241), .A2(n11242), .ZN(n12803) );
  INV_X1 U11306 ( .A(n12545), .ZN(n13191) );
  NAND2_X1 U11307 ( .A1(n11640), .A2(n14164), .ZN(n16089) );
  NAND2_X1 U11308 ( .A1(n13224), .A2(n13228), .ZN(n13417) );
  AOI21_X1 U11309 ( .B1(n11639), .B2(n21946), .A(n11631), .ZN(n11636) );
  NAND2_X1 U11310 ( .A1(n11273), .A2(n11272), .ZN(n12545) );
  INV_X1 U11311 ( .A(n13013), .ZN(n14347) );
  NOR2_X1 U11312 ( .A1(n20550), .A2(n20669), .ZN(n17796) );
  AND2_X2 U11313 ( .A1(n21859), .A2(n11645), .ZN(n14114) );
  NAND2_X1 U11314 ( .A1(n12523), .A2(n12520), .ZN(n13013) );
  INV_X1 U11315 ( .A(n13197), .ZN(n12567) );
  NAND3_X2 U11316 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(n20592) );
  NAND2_X1 U11317 ( .A1(n12691), .A2(n12690), .ZN(n13248) );
  INV_X1 U11318 ( .A(n13975), .ZN(n13974) );
  INV_X1 U11319 ( .A(n20736), .ZN(n20558) );
  INV_X1 U11320 ( .A(n12998), .ZN(n12525) );
  OR2_X1 U11321 ( .A1(n12667), .A2(n12666), .ZN(n13233) );
  NAND2_X1 U11322 ( .A1(n12530), .A2(n13181), .ZN(n13197) );
  NAND3_X1 U11323 ( .A1(n15063), .A2(n15062), .A3(n15061), .ZN(n20495) );
  AND2_X1 U11324 ( .A1(n14112), .A2(n22037), .ZN(n12335) );
  NOR2_X1 U11325 ( .A1(n11630), .A2(n11847), .ZN(n11994) );
  OR2_X1 U11326 ( .A1(n12679), .A2(n12678), .ZN(n13243) );
  AND3_X1 U11327 ( .A1(n11040), .A2(n11279), .A3(n11277), .ZN(n20736) );
  OR2_X1 U11328 ( .A1(n12705), .A2(n12704), .ZN(n13229) );
  NAND2_X1 U11329 ( .A1(n11160), .A2(n11159), .ZN(n20557) );
  OR2_X1 U11330 ( .A1(n12642), .A2(n12641), .ZN(n13260) );
  OR2_X1 U11331 ( .A1(n12845), .A2(n12844), .ZN(n13264) );
  INV_X2 U11332 ( .A(U212), .ZN(n10979) );
  NOR2_X1 U11333 ( .A1(n11632), .A2(n11630), .ZN(n13472) );
  INV_X2 U11334 ( .A(n12516), .ZN(n18335) );
  INV_X1 U11335 ( .A(n11632), .ZN(n14112) );
  INV_X1 U11336 ( .A(n14093), .ZN(n11633) );
  OR2_X2 U11337 ( .A1(n11560), .A2(n11559), .ZN(n21946) );
  OR2_X1 U11338 ( .A1(n11549), .A2(n11548), .ZN(n14093) );
  NOR2_X1 U11339 ( .A1(n11357), .A2(n11356), .ZN(n11360) );
  OR2_X2 U11340 ( .A1(n11580), .A2(n11579), .ZN(n14164) );
  NAND2_X2 U11341 ( .A1(U214), .A2(n19958), .ZN(n19999) );
  NAND2_X1 U11342 ( .A1(n12493), .A2(n12492), .ZN(n12516) );
  AND4_X1 U11343 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12758) );
  AND4_X1 U11344 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11626) );
  AND3_X1 U11345 ( .A1(n12430), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12429), .ZN(n12434) );
  AND4_X1 U11346 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12441) );
  CLKBUF_X3 U11347 ( .A(n11596), .Z(n12300) );
  AND2_X2 U11348 ( .A1(n15462), .A2(n12450), .ZN(n12656) );
  INV_X2 U11349 ( .A(n10992), .ZN(n10993) );
  BUF_X2 U11350 ( .A(n15066), .Z(n17742) );
  INV_X4 U11352 ( .A(n17518), .ZN(n17701) );
  BUF_X2 U11353 ( .A(n15076), .Z(n17765) );
  AND2_X2 U11355 ( .A1(n11540), .A2(n13958), .ZN(n11772) );
  INV_X1 U11356 ( .A(n11024), .ZN(n17464) );
  OR2_X1 U11357 ( .A1(n15254), .A2(n15041), .ZN(n17518) );
  INV_X2 U11358 ( .A(n19711), .ZN(n19763) );
  OR2_X1 U11359 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20721), .ZN(
        n11511) );
  NAND2_X1 U11360 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21165), .ZN(
        n15039) );
  NAND2_X1 U11361 ( .A1(n20712), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15038) );
  AND2_X1 U11362 ( .A1(n11541), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11538) );
  NOR2_X1 U11363 ( .A1(n11531), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11539) );
  AND2_X1 U11364 ( .A1(n16093), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11540) );
  AND2_X2 U11365 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14293) );
  OR2_X1 U11366 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20054) );
  AND2_X2 U11367 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16097) );
  AND2_X1 U11368 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13958) );
  NOR2_X2 U11369 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16098) );
  AND2_X1 U11370 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13833) );
  INV_X1 U11371 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16093) );
  AND2_X1 U11372 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11543) );
  INV_X2 U11373 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11847) );
  NOR2_X2 U11374 ( .A1(n20919), .A2(n20924), .ZN(n21084) );
  INV_X4 U11375 ( .A(n17587), .ZN(n17735) );
  INV_X1 U11376 ( .A(n12516), .ZN(n10980) );
  NOR2_X1 U11377 ( .A1(n15040), .A2(n15038), .ZN(n15089) );
  INV_X1 U11378 ( .A(n12459), .ZN(n10981) );
  INV_X1 U11379 ( .A(n12459), .ZN(n12460) );
  NAND3_X2 U11380 ( .A1(n12542), .A2(n13188), .A3(n12541), .ZN(n13180) );
  AND2_X4 U11381 ( .A1(n15475), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12743) );
  AND2_X1 U11382 ( .A1(n14293), .A2(n10966), .ZN(n10982) );
  AND2_X2 U11383 ( .A1(n14293), .A2(n10966), .ZN(n10983) );
  INV_X1 U11384 ( .A(n11021), .ZN(n10984) );
  OR2_X1 U11385 ( .A1(n20054), .A2(n15254), .ZN(n11021) );
  AND2_X1 U11387 ( .A1(n11458), .A2(n10966), .ZN(n10986) );
  NOR2_X2 U11388 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12636) );
  INV_X2 U11389 ( .A(n15470), .ZN(n10987) );
  OR2_X1 U11390 ( .A1(n12547), .A2(n13761), .ZN(n10988) );
  NAND2_X2 U11391 ( .A1(n12543), .A2(n12570), .ZN(n12574) );
  AND2_X4 U11392 ( .A1(n14293), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10989) );
  NOR2_X1 U11393 ( .A1(n20713), .A2(n15039), .ZN(n15208) );
  INV_X4 U11394 ( .A(n15941), .ZN(n19883) );
  INV_X4 U11395 ( .A(n11511), .ZN(n17737) );
  XNOR2_X1 U11396 ( .A(n12597), .B(n12596), .ZN(n13945) );
  AND2_X1 U11397 ( .A1(n11264), .A2(n11263), .ZN(n12594) );
  INV_X1 U11398 ( .A(n20592), .ZN(n10990) );
  OAI211_X1 U11399 ( .C1(n12527), .C2(n12515), .A(n12514), .B(n18334), .ZN(
        n13192) );
  INV_X1 U11400 ( .A(n15283), .ZN(n10991) );
  NOR4_X1 U11401 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A4(n20732), .ZN(n15051) );
  NAND2_X1 U11402 ( .A1(n21679), .A2(n11740), .ZN(n13964) );
  AND2_X1 U11403 ( .A1(n10998), .A2(n12519), .ZN(n13224) );
  AND2_X4 U11404 ( .A1(n11538), .A2(n11537), .ZN(n11596) );
  NAND2_X1 U11405 ( .A1(n11153), .A2(n13055), .ZN(n13058) );
  AND2_X1 U11406 ( .A1(n13818), .A2(n11542), .ZN(n10995) );
  NOR2_X1 U11407 ( .A1(n12619), .A2(n12610), .ZN(n19264) );
  INV_X1 U11408 ( .A(n16470), .ZN(n11426) );
  NAND2_X1 U11409 ( .A1(n16470), .A2(n11423), .ZN(n16424) );
  NAND2_X2 U11410 ( .A1(n11408), .A2(n12529), .ZN(n14332) );
  AOI22_X1 U11411 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14626), .B1(n14625), 
        .B2(n18340), .ZN(n18557) );
  AND4_X2 U11412 ( .A1(n13181), .A2(n19437), .A3(n14750), .A4(n12519), .ZN(
        n12523) );
  NOR2_X2 U11413 ( .A1(n14510), .A2(n14509), .ZN(n14547) );
  XNOR2_X2 U11414 ( .A(n13052), .B(n13053), .ZN(n14615) );
  NAND2_X2 U11415 ( .A1(n14534), .A2(n13051), .ZN(n13052) );
  NOR2_X2 U11416 ( .A1(n14420), .A2(n14419), .ZN(n14461) );
  AND2_X2 U11417 ( .A1(n14685), .A2(n11334), .ZN(n15014) );
  NOR2_X4 U11418 ( .A1(n14654), .A2(n14653), .ZN(n14685) );
  INV_X1 U11419 ( .A(n12460), .ZN(n10998) );
  NAND2_X1 U11420 ( .A1(n11407), .A2(n11406), .ZN(n12459) );
  NOR2_X1 U11421 ( .A1(n12460), .A2(n12519), .ZN(n11272) );
  INV_X1 U11422 ( .A(n12495), .ZN(n11273) );
  INV_X1 U11423 ( .A(n12741), .ZN(n11116) );
  INV_X1 U11424 ( .A(n12740), .ZN(n11115) );
  AOI21_X1 U11425 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19154), .A(
        n12778), .ZN(n12995) );
  NOR2_X1 U11426 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  INV_X1 U11427 ( .A(n12775), .ZN(n12777) );
  NAND2_X1 U11428 ( .A1(n12461), .A2(n12459), .ZN(n12538) );
  AOI21_X1 U11429 ( .B1(n20269), .B2(n20343), .A(n20358), .ZN(n11297) );
  OR2_X1 U11430 ( .A1(n12377), .A2(n12376), .ZN(n12381) );
  NAND2_X1 U11431 ( .A1(n13485), .A2(n11834), .ZN(n11836) );
  CLKBUF_X1 U11432 ( .A(n15079), .Z(n17759) );
  NAND2_X1 U11433 ( .A1(n11646), .A2(n14114), .ZN(n11655) );
  NAND2_X1 U11434 ( .A1(n19203), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U11435 ( .A1(n12582), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12535) );
  CLKBUF_X1 U11436 ( .A(n11757), .Z(n12301) );
  OR2_X1 U11437 ( .A1(n11715), .A2(n11714), .ZN(n13497) );
  NOR2_X1 U11438 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11532) );
  NOR2_X1 U11439 ( .A1(n20535), .A2(n17755), .ZN(n17753) );
  NOR2_X2 U11440 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12323) );
  OR2_X1 U11441 ( .A1(n14164), .A2(n11847), .ZN(n12317) );
  INV_X1 U11442 ( .A(n11375), .ZN(n11374) );
  INV_X1 U11443 ( .A(n13498), .ZN(n13486) );
  NAND3_X1 U11444 ( .A1(n11523), .A2(n12445), .A3(n12444), .ZN(n11406) );
  NOR2_X1 U11445 ( .A1(n11485), .A2(n11486), .ZN(n11484) );
  INV_X1 U11446 ( .A(n15509), .ZN(n11485) );
  NOR2_X1 U11447 ( .A1(n11346), .A2(n16306), .ZN(n11344) );
  NAND2_X1 U11448 ( .A1(n16296), .A2(n16288), .ZN(n11346) );
  AND2_X1 U11449 ( .A1(n16765), .A2(n16361), .ZN(n11489) );
  AND2_X1 U11450 ( .A1(n11066), .A2(n11475), .ZN(n11474) );
  INV_X1 U11451 ( .A(n14800), .ZN(n11475) );
  AND2_X1 U11452 ( .A1(n12516), .A2(n19262), .ZN(n13228) );
  NAND2_X1 U11453 ( .A1(n11490), .A2(n11491), .ZN(n12461) );
  NAND2_X1 U11454 ( .A1(n11463), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11462) );
  INV_X1 U11455 ( .A(n16443), .ZN(n11463) );
  NAND2_X1 U11456 ( .A1(n11118), .A2(n12571), .ZN(n12593) );
  NOR2_X1 U11457 ( .A1(n11270), .A2(n12957), .ZN(n11269) );
  INV_X1 U11458 ( .A(n13417), .ZN(n13410) );
  INV_X1 U11459 ( .A(n19437), .ZN(n12530) );
  NAND2_X1 U11460 ( .A1(n20592), .A2(n15245), .ZN(n17782) );
  AOI21_X1 U11461 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21176), .A(
        n15135), .ZN(n15257) );
  NOR2_X1 U11462 ( .A1(n20495), .A2(n10990), .ZN(n15246) );
  INV_X1 U11463 ( .A(n21183), .ZN(n17788) );
  NAND2_X1 U11464 ( .A1(n12390), .A2(n21229), .ZN(n13779) );
  AND2_X1 U11465 ( .A1(n11847), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12326) );
  NOR2_X2 U11466 ( .A1(n15618), .A2(n15605), .ZN(n15604) );
  INV_X1 U11467 ( .A(n16026), .ZN(n11361) );
  OR2_X1 U11468 ( .A1(n19946), .A2(n19945), .ZN(n11385) );
  NAND2_X1 U11469 ( .A1(n14869), .A2(n11025), .ZN(n19884) );
  OAI21_X1 U11470 ( .B1(n11836), .B2(n11212), .A(n11766), .ZN(n11434) );
  NAND2_X1 U11471 ( .A1(n11214), .A2(n11213), .ZN(n11766) );
  NOR2_X1 U11472 ( .A1(n21687), .A2(n21686), .ZN(n21821) );
  AND2_X1 U11473 ( .A1(n13078), .A2(n13079), .ZN(n17292) );
  NOR2_X1 U11474 ( .A1(n13058), .A2(n11288), .ZN(n11413) );
  INV_X1 U11475 ( .A(n13061), .ZN(n11288) );
  NAND2_X1 U11476 ( .A1(n13066), .A2(n13057), .ZN(n11151) );
  AND2_X1 U11477 ( .A1(n13030), .A2(n12525), .ZN(n12999) );
  NOR2_X1 U11478 ( .A1(n17320), .A2(n17305), .ZN(n19223) );
  INV_X1 U11479 ( .A(n12532), .ZN(n15487) );
  NAND2_X1 U11480 ( .A1(n20342), .A2(n20269), .ZN(n11295) );
  NAND2_X1 U11481 ( .A1(n20736), .A2(n20557), .ZN(n20506) );
  INV_X1 U11482 ( .A(n20670), .ZN(n20505) );
  INV_X1 U11483 ( .A(n16991), .ZN(n20497) );
  NAND3_X1 U11484 ( .A1(n21198), .A2(n21178), .A3(n21221), .ZN(n20498) );
  AOI22_X1 U11485 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15049) );
  AOI211_X1 U11486 ( .C1(n10993), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n15047), .B(n15046), .ZN(n15048) );
  AOI22_X1 U11487 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15050) );
  INV_X1 U11488 ( .A(n21182), .ZN(n21026) );
  OR2_X1 U11489 ( .A1(n19901), .A2(n15936), .ZN(n11177) );
  NAND2_X1 U11490 ( .A1(n14333), .A2(n18345), .ZN(n18664) );
  NOR3_X1 U11491 ( .A1(n20632), .A2(n20592), .A3(n11276), .ZN(n20593) );
  NAND2_X1 U11492 ( .A1(n20592), .A2(n20670), .ZN(n20658) );
  AND4_X1 U11493 ( .A1(n11647), .A2(n11655), .A3(n14108), .A4(n13805), .ZN(
        n11650) );
  INV_X1 U11494 ( .A(n12832), .ZN(n11114) );
  NOR2_X1 U11495 ( .A1(n12711), .A2(n15448), .ZN(n11113) );
  AND2_X1 U11496 ( .A1(n11856), .A2(n11867), .ZN(n11219) );
  OR2_X1 U11497 ( .A1(n11679), .A2(n11678), .ZN(n13551) );
  NAND2_X1 U11498 ( .A1(n21667), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11750) );
  OR2_X1 U11499 ( .A1(n11764), .A2(n11763), .ZN(n13496) );
  NAND2_X1 U11500 ( .A1(n11166), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11723) );
  NAND2_X1 U11501 ( .A1(n11724), .A2(n11170), .ZN(n11166) );
  INV_X1 U11502 ( .A(n11651), .ZN(n11170) );
  NAND2_X1 U11503 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11612) );
  NOR2_X1 U11504 ( .A1(n16093), .A2(n11213), .ZN(n11169) );
  NAND2_X1 U11505 ( .A1(n11651), .A2(n11169), .ZN(n11167) );
  NAND2_X1 U11506 ( .A1(n11323), .A2(n11331), .ZN(n11322) );
  OR2_X1 U11507 ( .A1(n15443), .A2(n11332), .ZN(n11331) );
  INV_X1 U11508 ( .A(n11527), .ZN(n11323) );
  INV_X1 U11509 ( .A(n16262), .ZN(n11332) );
  NOR2_X1 U11510 ( .A1(n11333), .A2(n16262), .ZN(n11330) );
  AND2_X1 U11511 ( .A1(n12912), .A2(n11230), .ZN(n11229) );
  NAND2_X1 U11512 ( .A1(n11234), .A2(n11231), .ZN(n11230) );
  AND2_X1 U11513 ( .A1(n11073), .A2(n13229), .ZN(n11469) );
  NAND2_X1 U11514 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11140) );
  AOI22_X1 U11515 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19160), .B1(
        n19121), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U11516 ( .A1(n11137), .A2(n11134), .ZN(n11133) );
  NAND2_X1 U11517 ( .A1(n19190), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U11518 ( .A1(n19250), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11141) );
  NAND2_X1 U11519 ( .A1(n14741), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11138) );
  NAND2_X1 U11520 ( .A1(n19236), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U11521 ( .A1(n12552), .A2(n12553), .ZN(n11264) );
  NOR2_X1 U11522 ( .A1(n14031), .A2(n19480), .ZN(n14023) );
  NAND2_X1 U11523 ( .A1(n12773), .A2(n12772), .ZN(n12775) );
  NAND2_X1 U11524 ( .A1(n11751), .A2(n11750), .ZN(n12379) );
  INV_X1 U11525 ( .A(n22037), .ZN(n12343) );
  AND2_X1 U11526 ( .A1(n11630), .A2(n14164), .ZN(n12397) );
  AND2_X1 U11527 ( .A1(n11456), .A2(n15633), .ZN(n11455) );
  AND2_X1 U11528 ( .A1(n15646), .A2(n15659), .ZN(n11456) );
  NOR2_X1 U11529 ( .A1(n15763), .A2(n11453), .ZN(n11452) );
  INV_X1 U11530 ( .A(n11094), .ZN(n11453) );
  OR2_X1 U11531 ( .A1(n11447), .A2(n11103), .ZN(n11446) );
  NOR2_X1 U11532 ( .A1(n11449), .A2(n11448), .ZN(n11447) );
  NOR2_X1 U11533 ( .A1(n14661), .A2(n14962), .ZN(n11448) );
  INV_X1 U11534 ( .A(n13541), .ZN(n11364) );
  NAND2_X1 U11535 ( .A1(n11217), .A2(n13537), .ZN(n13540) );
  OR2_X1 U11536 ( .A1(n14245), .A2(n11368), .ZN(n11172) );
  OR2_X1 U11537 ( .A1(n19871), .A2(n11370), .ZN(n11368) );
  INV_X1 U11538 ( .A(n11366), .ZN(n11365) );
  OAI21_X1 U11539 ( .B1(n19871), .B2(n11367), .A(n11050), .ZN(n11366) );
  NAND2_X1 U11540 ( .A1(n11369), .A2(n13521), .ZN(n11367) );
  NOR2_X1 U11541 ( .A1(n14191), .A2(n14233), .ZN(n14232) );
  NAND2_X1 U11542 ( .A1(n11836), .A2(n11431), .ZN(n11430) );
  NOR2_X1 U11543 ( .A1(n11765), .A2(n11432), .ZN(n11431) );
  INV_X1 U11544 ( .A(n12323), .ZN(n12315) );
  AND2_X1 U11545 ( .A1(n11092), .A2(n11395), .ZN(n11394) );
  INV_X1 U11546 ( .A(n15648), .ZN(n11395) );
  NAND2_X1 U11547 ( .A1(n11391), .A2(n15756), .ZN(n11390) );
  INV_X1 U11548 ( .A(n15767), .ZN(n11391) );
  INV_X1 U11549 ( .A(n15698), .ZN(n11392) );
  NAND2_X1 U11550 ( .A1(n15964), .A2(n11377), .ZN(n11373) );
  OR2_X1 U11551 ( .A1(n13575), .A2(n19894), .ZN(n11378) );
  INV_X1 U11552 ( .A(n13562), .ZN(n11185) );
  NAND2_X1 U11553 ( .A1(n11400), .A2(n14994), .ZN(n11399) );
  INV_X1 U11554 ( .A(n14947), .ZN(n11400) );
  NAND2_X1 U11555 ( .A1(n11188), .A2(n13786), .ZN(n13491) );
  INV_X1 U11556 ( .A(n12397), .ZN(n14089) );
  AND2_X1 U11557 ( .A1(n14112), .A2(n13551), .ZN(n13548) );
  OR2_X1 U11558 ( .A1(n11693), .A2(n11692), .ZN(n13498) );
  NAND2_X1 U11559 ( .A1(n14112), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11751) );
  NAND2_X1 U11560 ( .A1(n11211), .A2(n11210), .ZN(n11209) );
  NAND2_X1 U11561 ( .A1(n11734), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11210) );
  NAND2_X1 U11562 ( .A1(n11765), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11211) );
  AND2_X1 U11563 ( .A1(n11656), .A2(n22037), .ZN(n11642) );
  NAND4_X1 U11564 ( .A1(n13839), .A2(n21859), .A3(n12343), .A4(n21667), .ZN(
        n13815) );
  OR2_X1 U11565 ( .A1(n11590), .A2(n11589), .ZN(n11632) );
  AND2_X1 U11566 ( .A1(n21743), .A2(n11744), .ZN(n21668) );
  AND3_X2 U11567 ( .A1(n13488), .A2(n15798), .A3(n13472), .ZN(n14115) );
  AND2_X1 U11568 ( .A1(n12913), .A2(n12903), .ZN(n11253) );
  AND2_X1 U11569 ( .A1(n10974), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U11570 ( .A1(n11245), .A2(n12854), .ZN(n11244) );
  INV_X1 U11571 ( .A(n11247), .ZN(n11245) );
  NOR2_X1 U11572 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15284) );
  INV_X1 U11573 ( .A(n14863), .ZN(n11336) );
  INV_X1 U11574 ( .A(n14084), .ZN(n11477) );
  INV_X1 U11575 ( .A(n14507), .ZN(n11502) );
  AND2_X1 U11576 ( .A1(n11465), .A2(n11235), .ZN(n11234) );
  NAND2_X1 U11577 ( .A1(n12867), .A2(n11236), .ZN(n11235) );
  NOR2_X1 U11578 ( .A1(n16601), .A2(n11466), .ZN(n11465) );
  INV_X1 U11579 ( .A(n16634), .ZN(n11236) );
  INV_X1 U11580 ( .A(n14040), .ZN(n11497) );
  AND2_X1 U11581 ( .A1(n13075), .A2(n13079), .ZN(n11418) );
  AND3_X1 U11582 ( .A1(n13378), .A2(n13377), .A3(n13376), .ZN(n14466) );
  INV_X1 U11583 ( .A(n14035), .ZN(n11499) );
  NAND2_X1 U11584 ( .A1(n13013), .A2(n12524), .ZN(n13420) );
  NOR2_X1 U11585 ( .A1(n12538), .A2(n19594), .ZN(n12539) );
  NAND2_X1 U11586 ( .A1(n13757), .A2(n19262), .ZN(n14019) );
  NAND2_X1 U11587 ( .A1(n15439), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14013) );
  NAND2_X1 U11588 ( .A1(n12511), .A2(n12512), .ZN(n12527) );
  INV_X1 U11589 ( .A(n12988), .ZN(n13007) );
  AND2_X1 U11590 ( .A1(n18340), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14022) );
  NOR2_X1 U11591 ( .A1(n11312), .A2(n11315), .ZN(n11311) );
  INV_X1 U11592 ( .A(n11313), .ZN(n11312) );
  AND3_X1 U11593 ( .A1(n11201), .A2(n11030), .A3(n11200), .ZN(n17984) );
  INV_X1 U11594 ( .A(n17982), .ZN(n11200) );
  NAND2_X1 U11595 ( .A1(n18009), .A2(n17983), .ZN(n11201) );
  NAND2_X1 U11596 ( .A1(n17891), .A2(n11203), .ZN(n17955) );
  AND2_X1 U11597 ( .A1(n20927), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11203) );
  NOR2_X1 U11598 ( .A1(n18101), .A2(n20755), .ZN(n17830) );
  AND2_X1 U11599 ( .A1(n11198), .A2(n21034), .ZN(n17831) );
  OR2_X1 U11600 ( .A1(n17828), .A2(n11199), .ZN(n11198) );
  NAND2_X1 U11601 ( .A1(n18072), .A2(n11104), .ZN(n11199) );
  OR2_X1 U11602 ( .A1(n18127), .A2(n18099), .ZN(n17853) );
  NAND2_X1 U11603 ( .A1(n17753), .A2(n17789), .ZN(n17752) );
  NAND2_X1 U11604 ( .A1(n18151), .A2(n17779), .ZN(n17852) );
  NAND2_X1 U11605 ( .A1(n18172), .A2(n17775), .ZN(n17777) );
  NAND2_X1 U11606 ( .A1(n18202), .A2(n17772), .ZN(n17773) );
  OR2_X1 U11607 ( .A1(n16992), .A2(n11158), .ZN(n20692) );
  NAND2_X1 U11608 ( .A1(n20012), .A2(n17784), .ZN(n11158) );
  NOR2_X1 U11609 ( .A1(n20692), .A2(n20717), .ZN(n20720) );
  OR2_X1 U11610 ( .A1(n16089), .A2(n11648), .ZN(n13874) );
  NOR2_X1 U11611 ( .A1(n11438), .A2(n11437), .ZN(n11436) );
  INV_X1 U11612 ( .A(n11439), .ZN(n11438) );
  INV_X1 U11613 ( .A(n15774), .ZN(n11437) );
  NAND2_X1 U11614 ( .A1(n15546), .A2(n13627), .ZN(n13660) );
  AND2_X1 U11615 ( .A1(n15545), .A2(n14250), .ZN(n13627) );
  AND2_X1 U11616 ( .A1(n15671), .A2(n12205), .ZN(n15672) );
  NAND2_X1 U11617 ( .A1(n12181), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12222) );
  AND2_X1 U11618 ( .A1(n12116), .A2(n12115), .ZN(n15697) );
  AND2_X1 U11619 ( .A1(n12084), .A2(n11452), .ZN(n15765) );
  AND2_X1 U11620 ( .A1(n11888), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11890) );
  AND2_X1 U11621 ( .A1(n11172), .A2(n11365), .ZN(n13539) );
  NAND2_X1 U11622 ( .A1(n13539), .A2(n13538), .ZN(n14580) );
  OAI21_X1 U11623 ( .B1(n13584), .B2(n16025), .A(n19945), .ZN(n15868) );
  NAND2_X1 U11624 ( .A1(n15867), .A2(n15868), .ZN(n15877) );
  NAND2_X1 U11625 ( .A1(n13580), .A2(n15902), .ZN(n11183) );
  NAND2_X1 U11626 ( .A1(n11183), .A2(n11181), .ZN(n11180) );
  NAND2_X1 U11627 ( .A1(n15885), .A2(n16042), .ZN(n11181) );
  INV_X1 U11628 ( .A(n15885), .ZN(n11215) );
  NOR2_X1 U11629 ( .A1(n11023), .A2(n15686), .ZN(n15688) );
  NAND2_X1 U11630 ( .A1(n19894), .A2(n21404), .ZN(n11216) );
  INV_X1 U11631 ( .A(n13560), .ZN(n15941) );
  NAND2_X1 U11632 ( .A1(n13556), .A2(n13555), .ZN(n14869) );
  INV_X1 U11633 ( .A(n14871), .ZN(n13556) );
  AOI21_X1 U11634 ( .B1(n14100), .B2(n14099), .A(n21561), .ZN(n14118) );
  NAND2_X1 U11635 ( .A1(n11732), .A2(n11731), .ZN(n11740) );
  NAND2_X1 U11636 ( .A1(n11729), .A2(n11730), .ZN(n21679) );
  NOR2_X1 U11637 ( .A1(n11653), .A2(n11637), .ZN(n13628) );
  AND2_X1 U11638 ( .A1(n13508), .A2(n21658), .ZN(n21702) );
  BUF_X1 U11639 ( .A(n11632), .Z(n21991) );
  NOR2_X1 U11640 ( .A1(n21775), .A2(n22129), .ZN(n21835) );
  AOI21_X1 U11641 ( .B1(n21810), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22129), 
        .ZN(n21848) );
  NOR2_X2 U11642 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21852) );
  NAND2_X1 U11643 ( .A1(n11213), .A2(n21666), .ZN(n22129) );
  AND2_X1 U11644 ( .A1(n12547), .A2(n14332), .ZN(n14337) );
  INV_X1 U11645 ( .A(n12874), .ZN(n12871) );
  AND2_X1 U11646 ( .A1(n10975), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12860) );
  OR2_X1 U11647 ( .A1(n14338), .A2(n18661), .ZN(n13612) );
  INV_X1 U11648 ( .A(n14512), .ZN(n14509) );
  NOR2_X1 U11649 ( .A1(n11063), .A2(n11339), .ZN(n11338) );
  INV_X1 U11650 ( .A(n14261), .ZN(n11339) );
  AND2_X1 U11651 ( .A1(n11285), .A2(n13191), .ZN(n14279) );
  NOR2_X1 U11652 ( .A1(n12544), .A2(n13197), .ZN(n11285) );
  INV_X1 U11653 ( .A(n11020), .ZN(n11481) );
  NOR2_X1 U11654 ( .A1(n16172), .A2(n13413), .ZN(n11483) );
  INV_X1 U11655 ( .A(n16265), .ZN(n11326) );
  NAND2_X1 U11656 ( .A1(n11345), .A2(n11344), .ZN(n11343) );
  INV_X1 U11657 ( .A(n16283), .ZN(n11345) );
  INV_X1 U11658 ( .A(n16223), .ZN(n11487) );
  AND3_X1 U11659 ( .A1(n13364), .A2(n13363), .A3(n13362), .ZN(n14410) );
  AND2_X1 U11660 ( .A1(n12531), .A2(n12567), .ZN(n13190) );
  AND2_X1 U11661 ( .A1(n13929), .A2(n13928), .ZN(n17337) );
  AOI21_X1 U11662 ( .B1(n12867), .B2(n16609), .A(n11049), .ZN(n11468) );
  NAND2_X1 U11663 ( .A1(n16637), .A2(n16634), .ZN(n16608) );
  AND4_X1 U11664 ( .A1(n12747), .A2(n12746), .A3(n12745), .A4(n12744), .ZN(
        n12759) );
  NOR2_X2 U11665 ( .A1(n16414), .A2(n13452), .ZN(n15507) );
  AND2_X1 U11666 ( .A1(n11267), .A2(n12962), .ZN(n11265) );
  NAND2_X1 U11667 ( .A1(n11269), .A2(n12959), .ZN(n11268) );
  INV_X1 U11668 ( .A(n16275), .ZN(n11507) );
  NAND2_X1 U11669 ( .A1(n16299), .A2(n11065), .ZN(n16274) );
  NAND2_X1 U11670 ( .A1(n16466), .A2(n11457), .ZN(n11127) );
  NAND2_X1 U11671 ( .A1(n16467), .A2(n16733), .ZN(n11457) );
  NOR2_X1 U11672 ( .A1(n13056), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11152) );
  NAND2_X1 U11673 ( .A1(n11048), .A2(n11153), .ZN(n13067) );
  NAND2_X1 U11674 ( .A1(n11500), .A2(n11498), .ZN(n14039) );
  NAND2_X1 U11675 ( .A1(n12597), .A2(n12596), .ZN(n12581) );
  INV_X1 U11676 ( .A(n16755), .ZN(n16807) );
  NAND2_X1 U11677 ( .A1(n13766), .A2(n13765), .ZN(n13953) );
  XNOR2_X1 U11678 ( .A(n14015), .B(n14013), .ZN(n13955) );
  AND2_X1 U11679 ( .A1(n19162), .A2(n17309), .ZN(n19257) );
  OR2_X1 U11680 ( .A1(n19162), .A2(n17309), .ZN(n19124) );
  NAND2_X1 U11681 ( .A1(n18653), .A2(n18340), .ZN(n14594) );
  INV_X1 U11682 ( .A(n19281), .ZN(n19591) );
  AND2_X1 U11683 ( .A1(n14277), .A2(n14276), .ZN(n16957) );
  AOI21_X1 U11684 ( .B1(n18326), .B2(n21619), .A(n18322), .ZN(n20739) );
  AND2_X1 U11685 ( .A1(n11294), .A2(n20269), .ZN(n20378) );
  NAND2_X1 U11686 ( .A1(n11297), .A2(n20377), .ZN(n11296) );
  INV_X1 U11687 ( .A(n11311), .ZN(n11308) );
  AND2_X1 U11688 ( .A1(n17972), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18053) );
  AND2_X1 U11689 ( .A1(n17992), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17972) );
  NOR2_X1 U11690 ( .A1(n11317), .A2(n11318), .ZN(n11316) );
  NAND2_X1 U11691 ( .A1(n18203), .A2(n18204), .ZN(n18202) );
  NOR2_X1 U11692 ( .A1(n15096), .A2(n11280), .ZN(n11279) );
  AOI21_X1 U11693 ( .B1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n17700), .A(
        n11278), .ZN(n11277) );
  OAI211_X1 U11694 ( .C1(n15141), .C2(n15140), .A(n15257), .B(n15258), .ZN(
        n21183) );
  INV_X1 U11695 ( .A(n15128), .ZN(n20748) );
  INV_X1 U11696 ( .A(n15105), .ZN(n11159) );
  NOR2_X1 U11697 ( .A1(n15104), .A2(n11161), .ZN(n11160) );
  AOI21_X1 U11698 ( .B1(n15613), .B2(P1_REIP_REG_31__SCAN_IN), .A(n11404), 
        .ZN(n11403) );
  OAI21_X1 U11699 ( .B1(n15601), .B2(P1_REIP_REG_31__SCAN_IN), .A(n15600), 
        .ZN(n11404) );
  AND2_X1 U11700 ( .A1(n14663), .A2(n14380), .ZN(n21530) );
  AND2_X1 U11701 ( .A1(n14374), .A2(n14369), .ZN(n21490) );
  AND2_X1 U11702 ( .A1(n13793), .A2(n12393), .ZN(n12395) );
  AND2_X1 U11703 ( .A1(n11382), .A2(n19949), .ZN(n11380) );
  XNOR2_X1 U11704 ( .A(n15604), .B(n12328), .ZN(n15549) );
  NAND2_X1 U11705 ( .A1(n19927), .A2(n15937), .ZN(n11178) );
  NAND2_X1 U11706 ( .A1(n21546), .A2(n13476), .ZN(n19901) );
  AND2_X1 U11707 ( .A1(n19901), .A2(n14009), .ZN(n19927) );
  XNOR2_X1 U11708 ( .A(n15598), .B(n11405), .ZN(n15993) );
  INV_X1 U11709 ( .A(n15599), .ZN(n11405) );
  XNOR2_X1 U11710 ( .A(n15935), .B(n15568), .ZN(n21393) );
  INV_X1 U11711 ( .A(n19939), .ZN(n15933) );
  INV_X1 U11712 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21823) );
  NAND2_X1 U11713 ( .A1(n11837), .A2(n11836), .ZN(n21687) );
  INV_X1 U11714 ( .A(n22185), .ZN(n22188) );
  AND3_X1 U11715 ( .A1(n16962), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18345) );
  NAND2_X1 U11716 ( .A1(n18664), .A2(n13433), .ZN(n17268) );
  NAND2_X1 U11717 ( .A1(n17268), .A2(n17000), .ZN(n17296) );
  OR2_X1 U11718 ( .A1(n16155), .A2(n15514), .ZN(n11503) );
  OR2_X1 U11719 ( .A1(n16715), .A2(n13205), .ZN(n16691) );
  INV_X1 U11720 ( .A(n16696), .ZN(n11227) );
  NAND2_X1 U11721 ( .A1(n11151), .A2(n11031), .ZN(n11410) );
  INV_X1 U11722 ( .A(n18607), .ZN(n18625) );
  NAND2_X1 U11723 ( .A1(n13951), .A2(n13774), .ZN(n17305) );
  INV_X1 U11724 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19262) );
  INV_X1 U11725 ( .A(n17309), .ZN(n19491) );
  AND2_X1 U11726 ( .A1(n13767), .A2(n13953), .ZN(n17320) );
  OR2_X1 U11727 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  XNOR2_X1 U11728 ( .A(n14352), .B(n14353), .ZN(n19162) );
  AND2_X1 U11729 ( .A1(n20482), .A2(n20481), .ZN(n11305) );
  AND2_X1 U11730 ( .A1(n11298), .A2(n20269), .ZN(n20357) );
  AND2_X1 U11731 ( .A1(n20621), .A2(n11017), .ZN(n20605) );
  NOR2_X1 U11732 ( .A1(n20569), .A2(n20570), .ZN(n20633) );
  AOI22_X1 U11733 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U11734 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15075) );
  AOI211_X1 U11735 ( .C1(n10977), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n15072), .B(n15071), .ZN(n15073) );
  INV_X1 U11736 ( .A(n20637), .ZN(n20638) );
  NOR2_X1 U11737 ( .A1(n20651), .A2(n20650), .ZN(n20649) );
  NOR2_X1 U11738 ( .A1(n20657), .A2(n20655), .ZN(n20556) );
  NOR2_X1 U11739 ( .A1(n17676), .A2(n17675), .ZN(n21021) );
  NOR2_X1 U11740 ( .A1(n20506), .A2(n20505), .ZN(n20631) );
  NOR2_X1 U11741 ( .A1(n20505), .A2(n20499), .ZN(n20667) );
  INV_X1 U11742 ( .A(n20592), .ZN(n20671) );
  NAND2_X1 U11743 ( .A1(n20670), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n20665) );
  INV_X1 U11744 ( .A(n20631), .ZN(n20673) );
  AND2_X1 U11745 ( .A1(n11262), .A2(n11261), .ZN(n20998) );
  NAND2_X1 U11746 ( .A1(n20984), .A2(n21065), .ZN(n11261) );
  NAND2_X1 U11747 ( .A1(n20983), .A2(n21182), .ZN(n11262) );
  NOR3_X1 U11748 ( .A1(n20994), .A2(n21092), .A3(n11258), .ZN(n11257) );
  NAND2_X1 U11749 ( .A1(n11260), .A2(n11259), .ZN(n11258) );
  INV_X1 U11750 ( .A(n21030), .ZN(n11259) );
  OR2_X1 U11751 ( .A1(n21076), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11260) );
  XNOR2_X1 U11752 ( .A(n18047), .B(n21004), .ZN(n20993) );
  NAND2_X1 U11753 ( .A1(n11194), .A2(n11193), .ZN(n11192) );
  NOR2_X1 U11754 ( .A1(n21029), .A2(n21030), .ZN(n11193) );
  INV_X1 U11755 ( .A(n21028), .ZN(n11194) );
  NOR2_X2 U11756 ( .A1(n21021), .A2(n20846), .ZN(n21152) );
  INV_X1 U11757 ( .A(n21152), .ZN(n21133) );
  NOR2_X1 U11758 ( .A1(n12867), .A2(n16586), .ZN(n11231) );
  AND2_X1 U11759 ( .A1(n11234), .A2(n11233), .ZN(n11232) );
  INV_X1 U11760 ( .A(n12619), .ZN(n11137) );
  OAI21_X1 U11761 ( .B1(n12611), .B2(n19480), .A(n11135), .ZN(n11134) );
  NAND2_X1 U11762 ( .A1(n11136), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11135) );
  INV_X1 U11763 ( .A(n12610), .ZN(n11136) );
  NAND2_X1 U11764 ( .A1(n14750), .A2(n12532), .ZN(n12495) );
  AND2_X1 U11765 ( .A1(n19274), .A2(n16959), .ZN(n12795) );
  XNOR2_X1 U11766 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12985) );
  CLKBUF_X2 U11767 ( .A(n11687), .Z(n12302) );
  NOR2_X1 U11768 ( .A1(n14661), .A2(n11450), .ZN(n11449) );
  CLKBUF_X2 U11769 ( .A(n11709), .Z(n12294) );
  CLKBUF_X2 U11770 ( .A(n11680), .Z(n12303) );
  CLKBUF_X2 U11771 ( .A(n11707), .Z(n12291) );
  CLKBUF_X2 U11772 ( .A(n11702), .Z(n12304) );
  OR2_X1 U11773 ( .A1(n11820), .A2(n11819), .ZN(n13535) );
  OR2_X1 U11774 ( .A1(n11807), .A2(n11806), .ZN(n13532) );
  OR2_X1 U11775 ( .A1(n11795), .A2(n11794), .ZN(n13523) );
  CLKBUF_X2 U11776 ( .A(n11665), .Z(n12146) );
  NOR2_X1 U11777 ( .A1(n11660), .A2(n11659), .ZN(n11661) );
  NAND2_X1 U11778 ( .A1(n14106), .A2(n11530), .ZN(n11659) );
  AND2_X1 U11779 ( .A1(n11633), .A2(n21946), .ZN(n13488) );
  AND2_X1 U11780 ( .A1(n12544), .A2(n13007), .ZN(n13027) );
  OR2_X1 U11781 ( .A1(n12736), .A2(n12735), .ZN(n12781) );
  INV_X1 U11782 ( .A(n11468), .ZN(n11466) );
  OR2_X1 U11783 ( .A1(n12556), .A2(n16959), .ZN(n11119) );
  NAND2_X1 U11784 ( .A1(n11321), .A2(n11075), .ZN(n12558) );
  NAND2_X1 U11785 ( .A1(n12556), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U11786 ( .A1(n12567), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11145) );
  INV_X1 U11787 ( .A(n14466), .ZN(n11478) );
  NOR2_X1 U11788 ( .A1(n11114), .A2(n11113), .ZN(n11112) );
  INV_X1 U11789 ( .A(n12833), .ZN(n11111) );
  NAND2_X1 U11790 ( .A1(n12562), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11492) );
  NOR2_X1 U11791 ( .A1(n15436), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13219) );
  NOR2_X1 U11792 ( .A1(n12689), .A2(n12688), .ZN(n12690) );
  NAND2_X1 U11793 ( .A1(n12517), .A2(n12545), .ZN(n12560) );
  NAND2_X1 U11794 ( .A1(n10981), .A2(n12532), .ZN(n12521) );
  NAND2_X1 U11795 ( .A1(n12521), .A2(n12538), .ZN(n13017) );
  OAI211_X1 U11796 ( .C1(n13017), .C2(n13016), .A(n12462), .B(n12519), .ZN(
        n13186) );
  NAND2_X1 U11797 ( .A1(n13975), .A2(n13016), .ZN(n12462) );
  AOI21_X1 U11798 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21169), .A(
        n15129), .ZN(n15139) );
  AND2_X1 U11799 ( .A1(n17804), .A2(n17805), .ZN(n17792) );
  AND2_X1 U11800 ( .A1(n20544), .A2(n17796), .ZN(n17756) );
  AND2_X1 U11801 ( .A1(n15607), .A2(n13785), .ZN(n14193) );
  NAND2_X1 U11802 ( .A1(n13881), .A2(n11386), .ZN(n14053) );
  OAI211_X1 U11803 ( .C1(n13878), .C2(P1_EBX_REG_1__SCAN_IN), .A(n15607), .B(
        n13880), .ZN(n11386) );
  NAND2_X1 U11804 ( .A1(n12374), .A2(n12373), .ZN(n12387) );
  OR2_X1 U11805 ( .A1(n12372), .A2(n12371), .ZN(n12374) );
  NOR2_X1 U11806 ( .A1(n11442), .A2(n11440), .ZN(n11439) );
  INV_X1 U11807 ( .A(n11441), .ZN(n11440) );
  INV_X1 U11808 ( .A(n15725), .ZN(n11442) );
  OR2_X1 U11809 ( .A1(n16089), .A2(n11213), .ZN(n12320) );
  NOR2_X1 U11810 ( .A1(n15787), .A2(n15033), .ZN(n11441) );
  NAND2_X1 U11811 ( .A1(n11978), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U11812 ( .A1(n11443), .A2(n11449), .ZN(n14937) );
  XNOR2_X1 U11813 ( .A(n13530), .B(n11823), .ZN(n13542) );
  AND2_X1 U11814 ( .A1(n11428), .A2(n14169), .ZN(n11429) );
  INV_X1 U11815 ( .A(n14183), .ZN(n11428) );
  INV_X1 U11816 ( .A(n14193), .ZN(n15590) );
  OR2_X1 U11817 ( .A1(n11782), .A2(n11781), .ZN(n13515) );
  NAND3_X1 U11818 ( .A1(n21991), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n11645), 
        .ZN(n12366) );
  AND2_X1 U11819 ( .A1(n11613), .A2(n11612), .ZN(n11359) );
  NOR2_X1 U11820 ( .A1(n11034), .A2(n11003), .ZN(n11358) );
  OAI211_X1 U11821 ( .C1(n11724), .C2(n11168), .A(n11722), .B(n11167), .ZN(
        n11726) );
  INV_X1 U11822 ( .A(n11169), .ZN(n11168) );
  INV_X1 U11823 ( .A(n13484), .ZN(n21686) );
  OAI21_X1 U11824 ( .B1(n21556), .B2(n16083), .A(n16096), .ZN(n21666) );
  AND2_X1 U11825 ( .A1(n10974), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12898) );
  OR2_X1 U11826 ( .A1(n12883), .A2(n12881), .ZN(n12900) );
  NAND2_X1 U11827 ( .A1(n12893), .A2(n12894), .ZN(n12883) );
  AND2_X1 U11828 ( .A1(n10974), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12881) );
  AND2_X1 U11829 ( .A1(n12885), .A2(n12886), .ZN(n12893) );
  NOR2_X1 U11830 ( .A1(n12891), .A2(n12889), .ZN(n12885) );
  NAND2_X1 U11831 ( .A1(n11240), .A2(n12877), .ZN(n12891) );
  INV_X1 U11832 ( .A(n12878), .ZN(n11240) );
  AND2_X1 U11833 ( .A1(n10974), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12889) );
  NAND2_X1 U11834 ( .A1(n10974), .A2(n12771), .ZN(n11241) );
  NOR2_X1 U11835 ( .A1(n11330), .A2(n11329), .ZN(n11328) );
  INV_X1 U11836 ( .A(n16256), .ZN(n11329) );
  INV_X1 U11837 ( .A(n16726), .ZN(n11488) );
  NOR2_X1 U11838 ( .A1(n11480), .A2(n14410), .ZN(n11479) );
  INV_X1 U11839 ( .A(n14219), .ZN(n11480) );
  INV_X1 U11840 ( .A(n14083), .ZN(n11476) );
  INV_X1 U11841 ( .A(n15439), .ZN(n14031) );
  INV_X1 U11842 ( .A(n12989), .ZN(n12531) );
  NAND2_X1 U11843 ( .A1(n16125), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16127) );
  NAND2_X1 U11844 ( .A1(n13072), .A2(n13071), .ZN(n13077) );
  NAND2_X1 U11845 ( .A1(n11271), .A2(n12959), .ZN(n11267) );
  AND2_X1 U11846 ( .A1(n11424), .A2(n16660), .ZN(n11423) );
  INV_X1 U11847 ( .A(n11425), .ZN(n11424) );
  AND2_X1 U11848 ( .A1(n12944), .A2(n11460), .ZN(n11459) );
  INV_X1 U11849 ( .A(n16201), .ZN(n11508) );
  NAND2_X1 U11850 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11425) );
  AND2_X1 U11851 ( .A1(n16289), .A2(n11510), .ZN(n11509) );
  INV_X1 U11852 ( .A(n16220), .ZN(n11510) );
  INV_X1 U11853 ( .A(n14930), .ZN(n11506) );
  INV_X1 U11854 ( .A(n14865), .ZN(n11505) );
  NAND2_X1 U11855 ( .A1(n11015), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U11856 ( .A1(n13057), .A2(n12935), .ZN(n11223) );
  OR2_X1 U11857 ( .A1(n13042), .A2(n13248), .ZN(n12692) );
  NOR2_X1 U11858 ( .A1(n11132), .A2(n11131), .ZN(n11130) );
  OR2_X1 U11859 ( .A1(n15527), .A2(n13049), .ZN(n13050) );
  INV_X1 U11860 ( .A(n11264), .ZN(n11123) );
  INV_X1 U11861 ( .A(n12544), .ZN(n11287) );
  NAND2_X2 U11862 ( .A1(n10980), .A2(n19594), .ZN(n12544) );
  NAND2_X1 U11863 ( .A1(n13760), .A2(n13759), .ZN(n13772) );
  NAND2_X1 U11864 ( .A1(n15439), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13950) );
  NAND2_X1 U11865 ( .A1(n12617), .A2(n12609), .ZN(n12830) );
  AND2_X1 U11866 ( .A1(n11470), .A2(n14021), .ZN(n12617) );
  AND2_X1 U11867 ( .A1(n13995), .A2(n18587), .ZN(n11470) );
  AOI21_X1 U11868 ( .B1(n12502), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12424), .ZN(n12427) );
  AND2_X1 U11869 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12424) );
  INV_X1 U11870 ( .A(n12538), .ZN(n12520) );
  INV_X1 U11871 ( .A(n15254), .ZN(n11255) );
  INV_X1 U11872 ( .A(n15038), .ZN(n11256) );
  NOR2_X1 U11873 ( .A1(n20067), .A2(n11314), .ZN(n11313) );
  NOR2_X1 U11874 ( .A1(n20134), .A2(n11302), .ZN(n11301) );
  XNOR2_X1 U11875 ( .A(n20669), .B(n20550), .ZN(n17758) );
  NOR2_X1 U11876 ( .A1(n17846), .A2(n20892), .ZN(n18076) );
  NAND2_X1 U11877 ( .A1(n18126), .A2(n17827), .ZN(n17828) );
  NAND2_X1 U11878 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17853), .ZN(
        n20863) );
  INV_X1 U11879 ( .A(n15097), .ZN(n11278) );
  INV_X1 U11880 ( .A(n15098), .ZN(n11280) );
  OR2_X1 U11881 ( .A1(n20736), .A2(n20557), .ZN(n15260) );
  INV_X1 U11882 ( .A(n20506), .ZN(n20678) );
  NAND2_X1 U11883 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15254) );
  NAND2_X1 U11884 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11162) );
  INV_X1 U11885 ( .A(n12392), .ZN(n11165) );
  NAND2_X1 U11886 ( .A1(n15688), .A2(n11394), .ZN(n15650) );
  NOR2_X1 U11887 ( .A1(n15793), .A2(n15726), .ZN(n15780) );
  NOR3_X1 U11888 ( .A1(n14948), .A2(n11058), .A3(n14947), .ZN(n14995) );
  NOR2_X1 U11889 ( .A1(n14241), .A2(n14240), .ZN(n14438) );
  AND2_X1 U11890 ( .A1(n14062), .A2(n14061), .ZN(n14214) );
  AND2_X1 U11891 ( .A1(n12343), .A2(n14164), .ZN(n15798) );
  NAND2_X1 U11892 ( .A1(n14045), .A2(n11855), .ZN(n14170) );
  NAND2_X1 U11893 ( .A1(n21859), .A2(n21667), .ZN(n12392) );
  AOI21_X1 U11894 ( .B1(n13884), .B2(n14251), .A(n21587), .ZN(n19767) );
  INV_X1 U11895 ( .A(n12317), .ZN(n12327) );
  AND2_X1 U11896 ( .A1(n12264), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12265) );
  NOR2_X1 U11897 ( .A1(n12222), .A2(n15915), .ZN(n12223) );
  NAND2_X1 U11898 ( .A1(n12223), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12263) );
  AND2_X1 U11899 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12180), .ZN(
        n12181) );
  OR2_X1 U11900 ( .A1(n12186), .A2(n12185), .ZN(n15685) );
  NOR2_X1 U11901 ( .A1(n12130), .A2(n15936), .ZN(n12131) );
  NAND2_X1 U11902 ( .A1(n12131), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12179) );
  AND2_X1 U11903 ( .A1(n11072), .A2(n15752), .ZN(n11451) );
  AND2_X1 U11904 ( .A1(n12084), .A2(n11072), .ZN(n15753) );
  NOR2_X1 U11905 ( .A1(n12098), .A2(n15944), .ZN(n12099) );
  NAND2_X1 U11906 ( .A1(n12099), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U11907 ( .A1(n12084), .A2(n11094), .ZN(n15764) );
  NOR2_X1 U11908 ( .A1(n12064), .A2(n15957), .ZN(n12065) );
  NAND2_X1 U11909 ( .A1(n12065), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12098) );
  AND2_X1 U11910 ( .A1(n12014), .A2(n11439), .ZN(n15775) );
  NOR2_X1 U11911 ( .A1(n12031), .A2(n12030), .ZN(n12032) );
  INV_X1 U11912 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U11913 ( .A1(n12032), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U11914 ( .A1(n11997), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12031) );
  NAND2_X1 U11915 ( .A1(n12014), .A2(n12013), .ZN(n15788) );
  NOR2_X1 U11916 ( .A1(n11982), .A2(n15970), .ZN(n11997) );
  NOR2_X1 U11917 ( .A1(n11446), .A2(n11445), .ZN(n11444) );
  INV_X1 U11918 ( .A(n14988), .ZN(n11445) );
  AND2_X1 U11919 ( .A1(n11937), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U11920 ( .A1(n11938), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11977) );
  NOR2_X1 U11921 ( .A1(n11922), .A2(n14552), .ZN(n11937) );
  INV_X1 U11922 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14552) );
  NAND2_X1 U11923 ( .A1(n11171), .A2(n11221), .ZN(n14871) );
  AOI21_X1 U11924 ( .B1(n19879), .B2(n11364), .A(n11043), .ZN(n11221) );
  AND3_X1 U11925 ( .A1(n11907), .A2(n11906), .A3(n11905), .ZN(n14483) );
  AND2_X1 U11926 ( .A1(n11890), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11908) );
  AOI21_X1 U11927 ( .B1(n13531), .B2(n11994), .A(n11892), .ZN(n14233) );
  AND2_X1 U11928 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11824), .ZN(
        n11874) );
  AND2_X1 U11929 ( .A1(n15546), .A2(n14102), .ZN(n17035) );
  OAI21_X1 U11930 ( .B1(n11433), .B2(n11432), .A(n11042), .ZN(n11833) );
  OAI21_X1 U11931 ( .B1(n21687), .B2(n11432), .A(n11840), .ZN(n13871) );
  AOI21_X1 U11932 ( .B1(n13484), .B2(n11656), .A(n11847), .ZN(n14005) );
  INV_X1 U11933 ( .A(n15580), .ZN(n15596) );
  NAND2_X1 U11934 ( .A1(n15688), .A2(n11096), .ZN(n15637) );
  INV_X1 U11935 ( .A(n15635), .ZN(n11393) );
  NOR2_X1 U11936 ( .A1(n15637), .A2(n15622), .ZN(n15621) );
  NAND2_X1 U11937 ( .A1(n15688), .A2(n11092), .ZN(n15663) );
  AND2_X1 U11938 ( .A1(n15688), .A2(n15674), .ZN(n15676) );
  AND2_X1 U11939 ( .A1(n15579), .A2(n15578), .ZN(n15686) );
  OR2_X1 U11940 ( .A1(n11390), .A2(n15749), .ZN(n11389) );
  INV_X1 U11941 ( .A(n21378), .ZN(n11372) );
  NOR3_X1 U11942 ( .A1(n15768), .A2(n11392), .A3(n15767), .ZN(n15757) );
  NOR2_X1 U11943 ( .A1(n15768), .A2(n15767), .ZN(n15769) );
  NOR2_X1 U11944 ( .A1(n15932), .A2(n11077), .ZN(n19937) );
  NAND2_X1 U11945 ( .A1(n11373), .A2(n11374), .ZN(n15932) );
  NAND2_X1 U11946 ( .A1(n11173), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n19939) );
  INV_X1 U11947 ( .A(n19937), .ZN(n11173) );
  OR2_X1 U11948 ( .A1(n15778), .A2(n15714), .ZN(n15768) );
  NAND2_X1 U11949 ( .A1(n11184), .A2(n11006), .ZN(n11186) );
  OR2_X1 U11950 ( .A1(n14869), .A2(n11185), .ZN(n11184) );
  OR2_X1 U11951 ( .A1(n15791), .A2(n15790), .ZN(n15793) );
  NAND2_X1 U11952 ( .A1(n11398), .A2(n11397), .ZN(n11396) );
  INV_X1 U11953 ( .A(n11399), .ZN(n11398) );
  NOR2_X1 U11954 ( .A1(n11058), .A2(n15035), .ZN(n11397) );
  NOR2_X1 U11955 ( .A1(n14948), .A2(n14947), .ZN(n15028) );
  OR2_X1 U11956 ( .A1(n14542), .A2(n14543), .ZN(n14948) );
  AND2_X1 U11957 ( .A1(n14438), .A2(n14437), .ZN(n14490) );
  NAND2_X1 U11958 ( .A1(n11388), .A2(n11387), .ZN(n14241) );
  NOR2_X1 U11959 ( .A1(n14197), .A2(n14198), .ZN(n11387) );
  INV_X1 U11960 ( .A(n14212), .ZN(n11388) );
  NAND2_X1 U11961 ( .A1(n14214), .A2(n14213), .ZN(n14212) );
  XNOR2_X1 U11962 ( .A(n14008), .B(n13492), .ZN(n13940) );
  NOR2_X1 U11963 ( .A1(n14110), .A2(n21242), .ZN(n21327) );
  OAI21_X1 U11964 ( .B1(n13484), .B2(n13510), .A(n13483), .ZN(n14006) );
  NAND2_X1 U11965 ( .A1(n14006), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14008) );
  AND2_X1 U11966 ( .A1(n15607), .A2(n14056), .ZN(n15580) );
  OAI21_X1 U11967 ( .B1(n21699), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11698), 
        .ZN(n11841) );
  OAI21_X1 U11968 ( .B1(n11696), .B2(n11213), .A(n11695), .ZN(n11697) );
  NAND2_X1 U11969 ( .A1(n11746), .A2(n11745), .ZN(n11747) );
  NAND2_X1 U11970 ( .A1(n11207), .A2(n11206), .ZN(n11857) );
  AND2_X1 U11971 ( .A1(n11208), .A2(n11834), .ZN(n11206) );
  AOI21_X1 U11972 ( .B1(n13964), .B2(n11734), .A(n11209), .ZN(n11208) );
  NAND2_X1 U11973 ( .A1(n11785), .A2(n11856), .ZN(n11868) );
  XNOR2_X1 U11974 ( .A(n11728), .B(n11727), .ZN(n21699) );
  INV_X1 U11975 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13830) );
  NOR2_X1 U11976 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13818) );
  OR2_X2 U11977 ( .A1(n11570), .A2(n11569), .ZN(n22037) );
  INV_X1 U11978 ( .A(n21741), .ZN(n21789) );
  INV_X2 U11979 ( .A(n14364), .ZN(n21859) );
  AND2_X1 U11980 ( .A1(n21549), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12394) );
  NAND2_X1 U11981 ( .A1(n15546), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16096) );
  INV_X1 U11982 ( .A(n12394), .ZN(n17053) );
  NOR2_X1 U11983 ( .A1(n21549), .A2(n11847), .ZN(n16083) );
  NAND2_X1 U11984 ( .A1(n11246), .A2(n12851), .ZN(n12976) );
  INV_X1 U11985 ( .A(n12849), .ZN(n11246) );
  OR2_X1 U11986 ( .A1(n12966), .A2(n12965), .ZN(n12973) );
  OR2_X1 U11987 ( .A1(n12954), .A2(n12953), .ZN(n12966) );
  AND2_X1 U11988 ( .A1(n12947), .A2(n12946), .ZN(n12948) );
  NAND2_X1 U11989 ( .A1(n12948), .A2(n12949), .ZN(n12954) );
  NOR2_X1 U11990 ( .A1(n11250), .A2(n11249), .ZN(n11248) );
  INV_X1 U11991 ( .A(n12939), .ZN(n11250) );
  NAND2_X1 U11992 ( .A1(n12931), .A2(n12932), .ZN(n12938) );
  AND2_X1 U11993 ( .A1(n11253), .A2(n11252), .ZN(n11251) );
  INV_X1 U11994 ( .A(n11102), .ZN(n11252) );
  INV_X1 U11995 ( .A(n16114), .ZN(n13435) );
  AND2_X1 U11996 ( .A1(n16110), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16113) );
  NAND2_X1 U11997 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16113), .ZN(
        n16114) );
  NOR2_X1 U11998 ( .A1(n14714), .A2(n14713), .ZN(n16110) );
  NAND2_X1 U11999 ( .A1(n12859), .A2(n12858), .ZN(n12874) );
  INV_X1 U12000 ( .A(n12860), .ZN(n12858) );
  NAND2_X1 U12001 ( .A1(n12853), .A2(n12851), .ZN(n11247) );
  INV_X1 U12002 ( .A(n11341), .ZN(n11340) );
  INV_X1 U12003 ( .A(n14229), .ZN(n14227) );
  NAND2_X1 U12004 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14128) );
  INV_X1 U12005 ( .A(n11484), .ZN(n11482) );
  AND2_X1 U12006 ( .A1(n16162), .A2(n16161), .ZN(n16164) );
  XNOR2_X1 U12007 ( .A(n16278), .B(n15429), .ZN(n16272) );
  AND2_X1 U12008 ( .A1(n13399), .A2(n13398), .ZN(n16203) );
  NOR2_X2 U12009 ( .A1(n16221), .A2(n16203), .ZN(n16333) );
  NAND2_X1 U12010 ( .A1(n16280), .A2(n16279), .ZN(n16278) );
  INV_X1 U12011 ( .A(n11344), .ZN(n11342) );
  NAND2_X1 U12012 ( .A1(n16766), .A2(n11489), .ZN(n16725) );
  NAND2_X1 U12013 ( .A1(n16766), .A2(n11090), .ZN(n16723) );
  AND2_X1 U12014 ( .A1(n13387), .A2(n13386), .ZN(n16370) );
  AND2_X1 U12015 ( .A1(n11001), .A2(n11335), .ZN(n11334) );
  INV_X1 U12016 ( .A(n14984), .ZN(n11335) );
  NAND2_X1 U12017 ( .A1(n14220), .A2(n11479), .ZN(n14465) );
  NAND2_X1 U12018 ( .A1(n14220), .A2(n14219), .ZN(n14411) );
  NAND2_X1 U12019 ( .A1(n11474), .A2(n11473), .ZN(n11472) );
  INV_X1 U12020 ( .A(n16892), .ZN(n11473) );
  NAND2_X1 U12021 ( .A1(n11476), .A2(n11066), .ZN(n14801) );
  AND3_X1 U12022 ( .A1(n13232), .A2(n13231), .A3(n13230), .ZN(n14617) );
  NAND2_X1 U12023 ( .A1(n14030), .A2(n14029), .ZN(n14033) );
  NOR2_X1 U12024 ( .A1(n14031), .A2(n14895), .ZN(n14032) );
  XNOR2_X1 U12025 ( .A(n13247), .B(n13241), .ZN(n13981) );
  XOR2_X1 U12026 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13436), .Z(
        n14625) );
  AND2_X1 U12027 ( .A1(n16130), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16133) );
  OR2_X1 U12028 ( .A1(n16127), .A2(n18548), .ZN(n16129) );
  NAND2_X1 U12029 ( .A1(n11239), .A2(n11460), .ZN(n11238) );
  INV_X1 U12030 ( .A(n16445), .ZN(n11239) );
  OR2_X1 U12031 ( .A1(n16120), .A2(n18514), .ZN(n16122) );
  NAND2_X1 U12032 ( .A1(n16117), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16116) );
  INV_X1 U12033 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16511) );
  NOR2_X1 U12034 ( .A1(n16831), .A2(n16839), .ZN(n11293) );
  OR2_X1 U12035 ( .A1(n14712), .A2(n18425), .ZN(n14714) );
  INV_X1 U12036 ( .A(n14545), .ZN(n11501) );
  NAND2_X1 U12037 ( .A1(n14710), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14712) );
  NAND2_X1 U12038 ( .A1(n14459), .A2(n14458), .ZN(n14506) );
  NAND2_X1 U12039 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n14706), .ZN(
        n14705) );
  NAND2_X1 U12040 ( .A1(n17293), .A2(n17292), .ZN(n17291) );
  NAND2_X1 U12041 ( .A1(n11500), .A2(n11494), .ZN(n14156) );
  NAND2_X1 U12042 ( .A1(n11497), .A2(n14158), .ZN(n11495) );
  INV_X1 U12043 ( .A(n11498), .ZN(n11496) );
  AND2_X1 U12044 ( .A1(n11500), .A2(n11100), .ZN(n14157) );
  NOR2_X1 U12045 ( .A1(n14846), .A2(n14701), .ZN(n14704) );
  NAND2_X1 U12046 ( .A1(n12592), .A2(n12593), .ZN(n12605) );
  NOR2_X2 U12047 ( .A1(n16170), .A2(n16156), .ZN(n16155) );
  NOR2_X1 U12048 ( .A1(n16169), .A2(n12935), .ZN(n16399) );
  AND2_X1 U12049 ( .A1(n11423), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11422) );
  AND2_X1 U12050 ( .A1(n12960), .A2(n16675), .ZN(n16434) );
  OR2_X1 U12051 ( .A1(n12960), .A2(n16675), .ZN(n16433) );
  NAND2_X1 U12052 ( .A1(n16299), .A2(n11509), .ZN(n16218) );
  NAND2_X1 U12053 ( .A1(n16299), .A2(n16289), .ZN(n16291) );
  NAND2_X1 U12054 ( .A1(n12927), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11128) );
  NAND2_X1 U12055 ( .A1(n12917), .A2(n16486), .ZN(n11129) );
  AND2_X1 U12056 ( .A1(n16766), .A2(n16765), .ZN(n16768) );
  INV_X1 U12057 ( .A(n11420), .ZN(n11419) );
  NAND2_X1 U12058 ( .A1(n16640), .A2(n11418), .ZN(n11417) );
  OAI21_X1 U12059 ( .B1(n17292), .B2(n11421), .A(n13208), .ZN(n11420) );
  NOR3_X1 U12060 ( .A1(n14864), .A2(n14930), .A3(n14865), .ZN(n14971) );
  NOR2_X1 U12061 ( .A1(n11290), .A2(n16853), .ZN(n11289) );
  NOR2_X1 U12062 ( .A1(n11291), .A2(n11290), .ZN(n16576) );
  NAND2_X1 U12063 ( .A1(n16627), .A2(n11015), .ZN(n16596) );
  NOR2_X1 U12064 ( .A1(n11291), .A2(n16905), .ZN(n16606) );
  AND3_X1 U12065 ( .A1(n13287), .A2(n13286), .A3(n13285), .ZN(n14084) );
  NOR2_X1 U12066 ( .A1(n14083), .A2(n14084), .ZN(n14085) );
  NAND2_X1 U12067 ( .A1(n11225), .A2(n12818), .ZN(n11125) );
  NAND2_X1 U12068 ( .A1(n11411), .A2(n13065), .ZN(n16944) );
  OR2_X1 U12069 ( .A1(n13059), .A2(n11413), .ZN(n11411) );
  AND2_X1 U12070 ( .A1(n11151), .A2(n13058), .ZN(n13059) );
  NOR2_X1 U12071 ( .A1(n13180), .A2(n13197), .ZN(n14280) );
  OR2_X1 U12072 ( .A1(n13423), .A2(n13199), .ZN(n16755) );
  INV_X1 U12073 ( .A(n13772), .ZN(n13951) );
  AOI21_X1 U12074 ( .B1(n16241), .B2(n14022), .A(n13764), .ZN(n13765) );
  INV_X2 U12075 ( .A(n18557), .ZN(n18535) );
  NAND2_X1 U12076 ( .A1(n19162), .A2(n19491), .ZN(n17321) );
  INV_X1 U12077 ( .A(n19185), .ZN(n19184) );
  NAND2_X1 U12078 ( .A1(n17320), .A2(n17305), .ZN(n19182) );
  NAND2_X1 U12079 ( .A1(n12598), .A2(n18624), .ZN(n14774) );
  AND2_X1 U12080 ( .A1(n17320), .A2(n19195), .ZN(n19256) );
  INV_X1 U12081 ( .A(n14781), .ZN(n19593) );
  NAND2_X1 U12082 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19281), .ZN(n14781) );
  INV_X1 U12083 ( .A(n14783), .ZN(n19597) );
  INV_X1 U12084 ( .A(n14782), .ZN(n19598) );
  NAND3_X1 U12085 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15486), .A3(n19231), 
        .ZN(n14783) );
  NAND3_X1 U12086 ( .A1(n13649), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19231), 
        .ZN(n14782) );
  INV_X1 U12087 ( .A(n19119), .ZN(n19242) );
  INV_X1 U12088 ( .A(n19124), .ZN(n19120) );
  AND2_X1 U12089 ( .A1(n13011), .A2(n17302), .ZN(n18645) );
  NAND2_X1 U12090 ( .A1(n18340), .A2(n16962), .ZN(n18637) );
  OR2_X1 U12091 ( .A1(n17782), .A2(n20557), .ZN(n11274) );
  INV_X1 U12092 ( .A(n20741), .ZN(n21178) );
  OR2_X1 U12093 ( .A1(n20342), .A2(n20343), .ZN(n11298) );
  INV_X1 U12094 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20305) );
  NOR2_X1 U12095 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20160), .ZN(n20187) );
  AOI211_X1 U12096 ( .C1(n15066), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n15060), .B(n15059), .ZN(n15061) );
  NOR2_X1 U12097 ( .A1(n20013), .A2(n16990), .ZN(n18279) );
  NAND2_X1 U12098 ( .A1(n20738), .A2(n15243), .ZN(n20012) );
  NAND2_X1 U12099 ( .A1(n18053), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18022) );
  AND2_X1 U12100 ( .A1(n17922), .A2(n11013), .ZN(n17992) );
  INV_X1 U12101 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17921) );
  NOR2_X2 U12102 ( .A1(n17893), .A2(n17921), .ZN(n17922) );
  NAND2_X1 U12103 ( .A1(n18059), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17823) );
  NOR2_X1 U12104 ( .A1(n17848), .A2(n20265), .ZN(n18059) );
  NAND4_X1 U12105 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A4(n18067), .ZN(n17848) );
  NOR2_X1 U12106 ( .A1(n18093), .A2(n20217), .ZN(n18067) );
  INV_X1 U12107 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20217) );
  NOR2_X1 U12108 ( .A1(n18116), .A2(n18095), .ZN(n20200) );
  INV_X1 U12109 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18095) );
  NAND3_X1 U12110 ( .A1(n11299), .A2(n20200), .A3(n11301), .ZN(n18093) );
  INV_X1 U12111 ( .A(n20863), .ZN(n20750) );
  NOR2_X1 U12112 ( .A1(n20103), .A2(n11300), .ZN(n18148) );
  INV_X1 U12113 ( .A(n11301), .ZN(n11300) );
  INV_X1 U12114 ( .A(n18177), .ZN(n18181) );
  XNOR2_X1 U12115 ( .A(n17758), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18204) );
  AND2_X1 U12116 ( .A1(n11033), .A2(n21037), .ZN(n17991) );
  NAND2_X1 U12117 ( .A1(n17991), .A2(n18099), .ZN(n17990) );
  INV_X1 U12118 ( .A(n17959), .ZN(n11204) );
  NOR2_X1 U12119 ( .A1(n17955), .A2(n21054), .ZN(n11202) );
  NAND2_X1 U12120 ( .A1(n11350), .A2(n17952), .ZN(n17960) );
  AND2_X1 U12121 ( .A1(n17953), .A2(n11082), .ZN(n11350) );
  NOR2_X1 U12122 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17960), .ZN(
        n17959) );
  AND2_X1 U12123 ( .A1(n11349), .A2(n11197), .ZN(n18058) );
  NAND2_X1 U12124 ( .A1(n17829), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11349) );
  NOR2_X1 U12125 ( .A1(n17831), .A2(n11069), .ZN(n11197) );
  NAND2_X1 U12126 ( .A1(n18076), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20919) );
  NOR2_X1 U12127 ( .A1(n20924), .A2(n20917), .ZN(n20915) );
  INV_X1 U12128 ( .A(n21138), .ZN(n20893) );
  NAND2_X1 U12129 ( .A1(n18140), .A2(n17781), .ZN(n18127) );
  NAND2_X1 U12130 ( .A1(n18127), .A2(n18128), .ZN(n18126) );
  XNOR2_X1 U12131 ( .A(n17852), .B(n11205), .ZN(n18141) );
  INV_X1 U12132 ( .A(n17780), .ZN(n11205) );
  NAND2_X1 U12133 ( .A1(n18166), .A2(n17778), .ZN(n18152) );
  NAND2_X1 U12134 ( .A1(n18152), .A2(n18153), .ZN(n18151) );
  XNOR2_X1 U12135 ( .A(n17777), .B(n11348), .ZN(n18167) );
  INV_X1 U12136 ( .A(n17776), .ZN(n11348) );
  NAND2_X1 U12137 ( .A1(n18167), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18166) );
  NAND2_X1 U12138 ( .A1(n18191), .A2(n17774), .ZN(n18173) );
  NAND2_X1 U12139 ( .A1(n18173), .A2(n18174), .ZN(n18172) );
  NAND2_X1 U12140 ( .A1(n17785), .A2(n20006), .ZN(n21090) );
  INV_X1 U12141 ( .A(n20713), .ZN(n20704) );
  INV_X1 U12142 ( .A(n20719), .ZN(n11282) );
  INV_X1 U12143 ( .A(n20720), .ZN(n20688) );
  NAND2_X1 U12144 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20732), .ZN(
        n20727) );
  INV_X1 U12145 ( .A(n20696), .ZN(n20681) );
  NOR2_X2 U12146 ( .A1(n15117), .A2(n15116), .ZN(n20746) );
  NAND2_X1 U12147 ( .A1(n21182), .A2(n17788), .ZN(n11163) );
  NAND2_X1 U12148 ( .A1(n21019), .A2(n21180), .ZN(n11164) );
  INV_X1 U12149 ( .A(n21218), .ZN(n21221) );
  NAND2_X2 U12150 ( .A1(n12407), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21662)
         );
  NAND2_X1 U12151 ( .A1(n13656), .A2(n13660), .ZN(n21227) );
  AND2_X1 U12152 ( .A1(n15647), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15629) );
  NOR2_X1 U12153 ( .A1(n21453), .A2(n15708), .ZN(n21475) );
  INV_X1 U12154 ( .A(n21529), .ZN(n21505) );
  INV_X1 U12155 ( .A(n14663), .ZN(n15550) );
  INV_X1 U12156 ( .A(n21485), .ZN(n15720) );
  INV_X1 U12157 ( .A(n21530), .ZN(n21519) );
  INV_X1 U12158 ( .A(n15796), .ZN(n19866) );
  INV_X1 U12159 ( .A(n19870), .ZN(n15794) );
  AND2_X1 U12160 ( .A1(n13876), .A2(n13875), .ZN(n19870) );
  AND2_X1 U12161 ( .A1(n13785), .A2(n14250), .ZN(n13875) );
  INV_X1 U12162 ( .A(n19865), .ZN(n15785) );
  INV_X1 U12163 ( .A(n19866), .ZN(n15783) );
  AND2_X1 U12164 ( .A1(n15852), .A2(n14166), .ZN(n21653) );
  INV_X1 U12165 ( .A(n21653), .ZN(n15866) );
  NAND2_X1 U12166 ( .A1(n15864), .A2(n14167), .ZN(n15863) );
  NOR2_X2 U12167 ( .A1(n13660), .A2(n14088), .ZN(n13934) );
  NOR2_X1 U12168 ( .A1(n13478), .A2(n15873), .ZN(n13479) );
  AOI21_X1 U12169 ( .B1(n15620), .B2(n15617), .A(n15619), .ZN(n15883) );
  OAI21_X1 U12170 ( .B1(n15646), .B2(n15644), .A(n15645), .ZN(n15901) );
  AOI21_X1 U12171 ( .B1(n15661), .B2(n15660), .A(n15644), .ZN(n15908) );
  NAND2_X1 U12172 ( .A1(n21390), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n11176) );
  INV_X1 U12173 ( .A(n21512), .ZN(n21646) );
  INV_X1 U12174 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15944) );
  INV_X1 U12175 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15957) );
  NAND2_X1 U12176 ( .A1(n14580), .A2(n13541), .ZN(n19878) );
  NAND2_X1 U12177 ( .A1(n11371), .A2(n13521), .ZN(n19872) );
  NAND2_X1 U12178 ( .A1(n14245), .A2(n14244), .ZN(n11371) );
  NAND2_X1 U12179 ( .A1(n13591), .A2(n13590), .ZN(n11384) );
  AOI21_X1 U12180 ( .B1(n11009), .B2(n13585), .A(n11383), .ZN(n11382) );
  INV_X1 U12181 ( .A(n13592), .ZN(n11383) );
  XNOR2_X1 U12182 ( .A(n15877), .B(n11218), .ZN(n16016) );
  INV_X1 U12183 ( .A(n15878), .ZN(n11218) );
  INV_X1 U12184 ( .A(n11179), .ZN(n15888) );
  OAI211_X1 U12185 ( .C1(n11183), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11182), .B(n11180), .ZN(n11179) );
  INV_X1 U12186 ( .A(n15886), .ZN(n11182) );
  NAND2_X1 U12187 ( .A1(n15903), .A2(n13584), .ZN(n11362) );
  OR2_X1 U12188 ( .A1(n13580), .A2(n11216), .ZN(n15920) );
  XNOR2_X1 U12189 ( .A(n13580), .B(n11068), .ZN(n21400) );
  OR2_X1 U12190 ( .A1(n13480), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21401) );
  NAND2_X1 U12191 ( .A1(n14869), .A2(n13559), .ZN(n14901) );
  NOR2_X1 U12192 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21415), .ZN(
        n14174) );
  AND2_X1 U12193 ( .A1(n14118), .A2(n14117), .ZN(n21409) );
  AND2_X1 U12194 ( .A1(n14118), .A2(n14105), .ZN(n21411) );
  INV_X1 U12195 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21824) );
  NAND2_X1 U12196 ( .A1(n11836), .A2(n11212), .ZN(n11435) );
  AND2_X1 U12197 ( .A1(n15538), .A2(n14364), .ZN(n17021) );
  NOR2_X1 U12198 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16094) );
  INV_X1 U12199 ( .A(n21710), .ZN(n22157) );
  OAI21_X1 U12200 ( .B1(n22162), .B2(n21721), .A(n21835), .ZN(n22164) );
  AND2_X1 U12201 ( .A1(n21742), .A2(n21821), .ZN(n22181) );
  OAI211_X1 U12202 ( .C1(n22186), .C2(n21805), .A(n21780), .B(n21761), .ZN(
        n22189) );
  OAI21_X1 U12203 ( .B1(n21788), .B2(n21787), .A(n21848), .ZN(n22207) );
  OAI211_X1 U12204 ( .C1(n22211), .C2(n21805), .A(n21835), .B(n21804), .ZN(
        n22214) );
  AOI22_X1 U12205 ( .A1(n21803), .A2(n21800), .B1(n21799), .B2(n21798), .ZN(
        n22218) );
  OAI211_X1 U12206 ( .C1(n22226), .C2(n21836), .A(n21835), .B(n21834), .ZN(
        n22229) );
  NOR2_X1 U12207 ( .A1(n22129), .A2(n21661), .ZN(n21845) );
  NOR2_X1 U12208 ( .A1(n22129), .A2(n21857), .ZN(n21895) );
  NOR2_X1 U12209 ( .A1(n22129), .A2(n21900), .ZN(n21939) );
  INV_X1 U12210 ( .A(n21968), .ZN(n21984) );
  NOR2_X1 U12211 ( .A1(n22129), .A2(n21944), .ZN(n21983) );
  INV_X1 U12212 ( .A(n22014), .ZN(n22030) );
  NOR2_X1 U12213 ( .A1(n22129), .A2(n21989), .ZN(n22029) );
  INV_X1 U12214 ( .A(n22062), .ZN(n22078) );
  NOR2_X1 U12215 ( .A1(n22129), .A2(n22035), .ZN(n22077) );
  NOR2_X1 U12216 ( .A1(n22129), .A2(n22083), .ZN(n22123) );
  AND2_X1 U12217 ( .A1(n21822), .A2(n21741), .ZN(n22238) );
  NOR2_X1 U12218 ( .A1(n22129), .A2(n22128), .ZN(n22235) );
  NAND2_X1 U12219 ( .A1(n12394), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21561) );
  INV_X1 U12220 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21549) );
  INV_X1 U12221 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21585) );
  INV_X1 U12222 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19796) );
  NOR2_X1 U12223 ( .A1(n13612), .A2(n12547), .ZN(n14635) );
  INV_X1 U12224 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18565) );
  INV_X1 U12225 ( .A(n18509), .ZN(n18572) );
  NAND2_X1 U12226 ( .A1(n18341), .A2(n14631), .ZN(n18576) );
  OR3_X1 U12227 ( .A1(n14641), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n21594), 
        .ZN(n18511) );
  INV_X1 U12228 ( .A(n18643), .ZN(n18558) );
  OR2_X1 U12229 ( .A1(n13374), .A2(n13373), .ZN(n14686) );
  OR2_X1 U12230 ( .A1(n13361), .A2(n13360), .ZN(n14656) );
  OR2_X1 U12231 ( .A1(n13348), .A2(n13347), .ZN(n14548) );
  CLKBUF_X1 U12232 ( .A(n14654), .Z(n14652) );
  OR2_X1 U12233 ( .A1(n13335), .A2(n13334), .ZN(n14512) );
  OR2_X1 U12234 ( .A1(n13322), .A2(n13321), .ZN(n14462) );
  CLKBUF_X1 U12235 ( .A(n14510), .Z(n14508) );
  OR2_X1 U12236 ( .A1(n13309), .A2(n13308), .ZN(n14422) );
  OR2_X1 U12237 ( .A1(n13297), .A2(n13296), .ZN(n14261) );
  CLKBUF_X1 U12238 ( .A(n14420), .Z(n14418) );
  NOR2_X1 U12239 ( .A1(n14128), .A2(n19296), .ZN(n11341) );
  INV_X1 U12240 ( .A(n16302), .ZN(n16307) );
  AND2_X1 U12241 ( .A1(n13769), .A2(n18345), .ZN(n16284) );
  OR2_X1 U12242 ( .A1(n14161), .A2(n13976), .ZN(n16302) );
  XNOR2_X1 U12243 ( .A(n13419), .B(n13418), .ZN(n19110) );
  NAND2_X1 U12244 ( .A1(n11481), .A2(n11091), .ZN(n13419) );
  NAND2_X1 U12245 ( .A1(n11326), .A2(n11325), .ZN(n16260) );
  NOR2_X1 U12246 ( .A1(n11527), .A2(n11333), .ZN(n11325) );
  AND2_X1 U12247 ( .A1(n15489), .A2(n15485), .ZN(n19583) );
  AND2_X1 U12248 ( .A1(n15489), .A2(n15488), .ZN(n19582) );
  AND2_X1 U12249 ( .A1(n15489), .A2(n10974), .ZN(n19581) );
  NAND2_X1 U12250 ( .A1(n13975), .A2(n15489), .ZN(n14684) );
  NAND2_X1 U12251 ( .A1(n13973), .A2(n13972), .ZN(n19496) );
  INV_X1 U12252 ( .A(n19342), .ZN(n19586) );
  INV_X1 U12253 ( .A(n16373), .ZN(n19585) );
  INV_X1 U12254 ( .A(n19496), .ZN(n19579) );
  NAND2_X1 U12256 ( .A1(n16152), .A2(n17273), .ZN(n13464) );
  INV_X1 U12257 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16457) );
  NAND2_X1 U12258 ( .A1(n11467), .A2(n11468), .ZN(n16600) );
  NAND2_X1 U12259 ( .A1(n16608), .A2(n12867), .ZN(n11467) );
  INV_X1 U12260 ( .A(n17294), .ZN(n17270) );
  INV_X1 U12261 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17269) );
  INV_X1 U12262 ( .A(n17296), .ZN(n17273) );
  INV_X1 U12263 ( .A(n17268), .ZN(n17286) );
  INV_X1 U12264 ( .A(n18614), .ZN(n18627) );
  INV_X1 U12265 ( .A(n11415), .ZN(n11414) );
  NAND2_X1 U12266 ( .A1(n13067), .A2(n11416), .ZN(n14833) );
  AND2_X1 U12267 ( .A1(n11500), .A2(n13084), .ZN(n14036) );
  INV_X1 U12268 ( .A(n18427), .ZN(n18600) );
  OR2_X1 U12269 ( .A1(n13423), .A2(n13184), .ZN(n18615) );
  INV_X1 U12270 ( .A(n16241), .ZN(n13995) );
  OR2_X1 U12271 ( .A1(n13423), .A2(n13422), .ZN(n18603) );
  INV_X1 U12272 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19274) );
  INV_X1 U12273 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19272) );
  INV_X1 U12274 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19172) );
  INV_X1 U12275 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19154) );
  OR2_X1 U12276 ( .A1(n17321), .A2(n17320), .ZN(n19212) );
  CLKBUF_X1 U12277 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n16959) );
  NOR2_X1 U12278 ( .A1(n14591), .A2(n19262), .ZN(n18653) );
  INV_X1 U12279 ( .A(n17305), .ZN(n19195) );
  OR2_X1 U12280 ( .A1(n13955), .A2(n13954), .ZN(n13956) );
  AOI21_X1 U12281 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17001), .A(n16958), .ZN(
        n18579) );
  INV_X1 U12282 ( .A(n19676), .ZN(n19678) );
  OAI22_X1 U12283 ( .A1(n19239), .A2(n19235), .B1(n19234), .B2(n19233), .ZN(
        n19673) );
  OR2_X1 U12284 ( .A1(n17321), .A2(n19182), .ZN(n19564) );
  INV_X1 U12285 ( .A(n19641), .ZN(n19553) );
  NOR2_X1 U12286 ( .A1(n19185), .A2(n19143), .ZN(n19625) );
  INV_X1 U12287 ( .A(n19534), .ZN(n19538) );
  AOI22_X1 U12288 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19597), .ZN(n19387) );
  INV_X1 U12289 ( .A(n19697), .ZN(n19700) );
  AOI22_X1 U12290 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19597), .ZN(n19470) );
  INV_X1 U12291 ( .A(n19473), .ZN(n19475) );
  INV_X1 U12292 ( .A(n19430), .ZN(n19432) );
  NAND2_X1 U12293 ( .A1(n19120), .A2(n19256), .ZN(n19614) );
  AOI22_X1 U12294 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19597), .ZN(n19331) );
  INV_X1 U12295 ( .A(n19271), .ZN(n19293) );
  INV_X1 U12296 ( .A(n19690), .ZN(n19704) );
  INV_X1 U12297 ( .A(n19642), .ZN(n19698) );
  AOI22_X1 U12298 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19597), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19598), .ZN(n19697) );
  INV_X1 U12299 ( .A(n19578), .ZN(n19569) );
  INV_X1 U12300 ( .A(n19531), .ZN(n19536) );
  AND2_X1 U12301 ( .A1(n13001), .A2(n19593), .ZN(n19535) );
  AOI22_X1 U12302 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_18__SCAN_IN), .B2(n19597), .ZN(n19534) );
  INV_X1 U12303 ( .A(n19470), .ZN(n19477) );
  INV_X1 U12304 ( .A(n19452), .ZN(n19474) );
  AOI22_X1 U12305 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19597), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19598), .ZN(n19473) );
  AOI22_X1 U12306 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19597), .ZN(n19430) );
  INV_X1 U12307 ( .A(n19435), .ZN(n19427) );
  INV_X1 U12308 ( .A(n19384), .ZN(n19392) );
  INV_X1 U12309 ( .A(n19387), .ZN(n19389) );
  AOI22_X1 U12310 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19597), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19598), .ZN(n19334) );
  INV_X1 U12311 ( .A(n19331), .ZN(n19336) );
  AOI22_X1 U12312 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19597), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19598), .ZN(n19271) );
  INV_X1 U12313 ( .A(n19602), .ZN(n19705) );
  NAND2_X1 U12314 ( .A1(n19120), .A2(n19242), .ZN(n19544) );
  INV_X1 U12315 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17375) );
  OR2_X1 U12316 ( .A1(n21177), .A2(n20013), .ZN(n20059) );
  NOR2_X1 U12317 ( .A1(n15243), .A2(n15262), .ZN(n21158) );
  NAND2_X1 U12318 ( .A1(n21221), .A2(n21178), .ZN(n20013) );
  INV_X1 U12319 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20057) );
  NOR2_X1 U12320 ( .A1(n17823), .A2(n20305), .ZN(n20312) );
  NOR2_X1 U12321 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20303), .ZN(n20315) );
  NOR2_X1 U12322 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20213), .ZN(n20234) );
  INV_X1 U12323 ( .A(n20490), .ZN(n20407) );
  INV_X1 U12324 ( .A(n20486), .ZN(n20451) );
  NAND4_X1 U12325 ( .A1(n21129), .A2(n20059), .A3(n21205), .A4(n21216), .ZN(
        n20490) );
  INV_X1 U12326 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17420) );
  NOR2_X1 U12327 ( .A1(n20125), .A2(n17411), .ZN(n17422) );
  INV_X1 U12328 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17725) );
  INV_X1 U12329 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17712) );
  INV_X1 U12330 ( .A(n17655), .ZN(n17657) );
  NAND2_X1 U12331 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(P3_EAX_REG_25__SCAN_IN), 
        .ZN(n11275) );
  NAND2_X1 U12332 ( .A1(n11281), .A2(n10999), .ZN(n20569) );
  NOR2_X1 U12333 ( .A1(n20577), .A2(n20582), .ZN(n20576) );
  NAND4_X1 U12334 ( .A1(n20556), .A2(P3_EAX_REG_13__SCAN_IN), .A3(
        P3_EAX_REG_12__SCAN_IN), .A4(n20555), .ZN(n20651) );
  NOR2_X1 U12335 ( .A1(n20554), .A2(n20524), .ZN(n20518) );
  NAND4_X1 U12336 ( .A1(n20662), .A2(P3_EAX_REG_4__SCAN_IN), .A3(
        P3_EAX_REG_5__SCAN_IN), .A4(n20503), .ZN(n20657) );
  NOR2_X1 U12337 ( .A1(n17686), .A2(n17685), .ZN(n20535) );
  NOR2_X1 U12338 ( .A1(n20546), .A2(n20547), .ZN(n20539) );
  INV_X1 U12339 ( .A(n17790), .ZN(n20669) );
  NOR2_X1 U12340 ( .A1(n20665), .A2(n20664), .ZN(n20662) );
  NOR2_X2 U12341 ( .A1(n21196), .A2(n20013), .ZN(n20046) );
  NOR2_X2 U12342 ( .A1(n20012), .A2(n20498), .ZN(n20051) );
  CLKBUF_X1 U12343 ( .A(n20043), .Z(n20050) );
  NAND2_X1 U12344 ( .A1(n11308), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U12345 ( .A1(n18053), .A2(n11093), .ZN(n11309) );
  OR2_X1 U12346 ( .A1(n18053), .A2(n20485), .ZN(n11310) );
  OAI211_X1 U12347 ( .C1(n18049), .C2(n18048), .A(n18054), .B(n11105), .ZN(
        n11355) );
  OR2_X1 U12348 ( .A1(n18051), .A2(n18050), .ZN(n11353) );
  NAND2_X1 U12349 ( .A1(n17990), .A2(n21037), .ZN(n17985) );
  NAND2_X1 U12350 ( .A1(n17922), .A2(n11000), .ZN(n18006) );
  NAND2_X1 U12351 ( .A1(n17922), .A2(n11008), .ZN(n17936) );
  INV_X1 U12352 ( .A(n18064), .ZN(n17870) );
  NAND3_X1 U12353 ( .A1(n21574), .A2(n18221), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18003) );
  NOR2_X2 U12354 ( .A1(n21021), .A2(n18225), .ZN(n18122) );
  INV_X1 U12355 ( .A(n18122), .ZN(n18139) );
  NAND2_X1 U12356 ( .A1(n11299), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18157) );
  INV_X1 U12357 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20134) );
  INV_X1 U12358 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20067) );
  INV_X1 U12359 ( .A(n21038), .ZN(n11190) );
  NOR2_X1 U12360 ( .A1(n21179), .A2(n20749), .ZN(n21065) );
  AOI21_X1 U12361 ( .B1(n20874), .B2(n20912), .A(n21092), .ZN(n21150) );
  INV_X1 U12362 ( .A(n21111), .ZN(n21059) );
  NOR2_X1 U12363 ( .A1(n21092), .A2(n21026), .ZN(n20955) );
  NAND2_X1 U12364 ( .A1(n21136), .A2(n21019), .ZN(n20846) );
  INV_X1 U12365 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21176) );
  INV_X1 U12366 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20732) );
  NOR2_X1 U12367 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20057), .ZN(n21201) );
  NAND2_X1 U12368 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21621), .ZN(n18324) );
  INV_X1 U12369 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22244) );
  OR2_X1 U12370 ( .A1(n13649), .A2(n13608), .ZN(n19958) );
  CLKBUF_X1 U12371 ( .A(n18690), .Z(n19008) );
  AOI21_X1 U12372 ( .B1(n15993), .B2(n21490), .A(n11402), .ZN(n15602) );
  INV_X1 U12373 ( .A(n11403), .ZN(n11402) );
  AOI21_X1 U12374 ( .B1(n21393), .B2(n19949), .A(n11174), .ZN(n15938) );
  NAND2_X1 U12375 ( .A1(n11178), .A2(n11175), .ZN(n11174) );
  AND2_X1 U12376 ( .A1(n11177), .A2(n11176), .ZN(n11175) );
  NAND2_X1 U12377 ( .A1(n11004), .A2(n11146), .ZN(n16802) );
  OAI211_X1 U12378 ( .C1(n18607), .C2(n18569), .A(n15520), .B(n15521), .ZN(
        n15522) );
  NAND2_X1 U12379 ( .A1(n11227), .A2(n18623), .ZN(n11226) );
  NOR3_X1 U12380 ( .A1(n20480), .A2(n11305), .A3(n11304), .ZN(n11303) );
  OR2_X1 U12381 ( .A1(n20474), .A2(n11099), .ZN(n11306) );
  NAND2_X1 U12382 ( .A1(n20483), .A2(n11067), .ZN(n11304) );
  INV_X1 U12383 ( .A(n20605), .ZN(n20610) );
  NOR2_X1 U12384 ( .A1(n20632), .A2(n20592), .ZN(n20626) );
  INV_X1 U12385 ( .A(n20665), .ZN(n20675) );
  OAI21_X1 U12386 ( .B1(n20993), .B2(n18139), .A(n11351), .ZN(P3_U2801) );
  AND2_X1 U12387 ( .A1(n11354), .A2(n11352), .ZN(n11351) );
  NAND2_X1 U12388 ( .A1(n11353), .A2(n20446), .ZN(n11352) );
  INV_X1 U12389 ( .A(n11355), .ZN(n11354) );
  AOI21_X1 U12390 ( .B1(n20998), .B2(n11257), .A(n21004), .ZN(n20985) );
  NOR2_X1 U12391 ( .A1(n11029), .A2(n11190), .ZN(n11189) );
  AOI21_X1 U12392 ( .B1(n11196), .B2(n11195), .A(n11192), .ZN(n11191) );
  OR2_X1 U12393 ( .A1(n19958), .A2(n19993), .ZN(U212) );
  AND4_X1 U12394 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n11106), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n10999) );
  NOR2_X1 U12395 ( .A1(n15039), .A2(n15038), .ZN(n15065) );
  AND2_X1 U12396 ( .A1(n11011), .A2(n11316), .ZN(n11000) );
  AND2_X1 U12397 ( .A1(n11010), .A2(n14929), .ZN(n11001) );
  INV_X1 U12398 ( .A(n12574), .ZN(n13174) );
  NOR2_X1 U12399 ( .A1(n20054), .A2(n20727), .ZN(n15076) );
  NAND2_X1 U12400 ( .A1(n14685), .A2(n11001), .ZN(n14983) );
  NAND2_X1 U12401 ( .A1(n14685), .A2(n14686), .ZN(n14862) );
  AND2_X1 U12402 ( .A1(n12648), .A2(n12647), .ZN(n11002) );
  AND2_X1 U12403 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11003) );
  AND2_X1 U12404 ( .A1(n16517), .A2(n11108), .ZN(n11004) );
  OR2_X1 U12405 ( .A1(n16305), .A2(n11342), .ZN(n11005) );
  INV_X1 U12406 ( .A(n11377), .ZN(n11376) );
  AND2_X1 U12407 ( .A1(n11378), .A2(n11041), .ZN(n11006) );
  NAND2_X1 U12408 ( .A1(n11187), .A2(n11734), .ZN(n13485) );
  INV_X1 U12409 ( .A(n13485), .ZN(n11188) );
  INV_X1 U12410 ( .A(n16527), .ZN(n11147) );
  AND3_X1 U12411 ( .A1(n11222), .A2(n12693), .A3(n11073), .ZN(n11007) );
  INV_X1 U12412 ( .A(n13056), .ZN(n13062) );
  NAND2_X1 U12413 ( .A1(n11749), .A2(n14442), .ZN(n13802) );
  NAND2_X1 U12414 ( .A1(n13083), .A2(n13086), .ZN(n11500) );
  INV_X1 U12415 ( .A(n11994), .ZN(n11432) );
  AND2_X1 U12416 ( .A1(n11429), .A2(n14170), .ZN(n14182) );
  NAND2_X1 U12417 ( .A1(n14459), .A2(n11064), .ZN(n14504) );
  AND2_X1 U12418 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11008) );
  AND2_X1 U12419 ( .A1(n13587), .A2(n13586), .ZN(n11009) );
  AND2_X1 U12420 ( .A1(n11336), .A2(n14686), .ZN(n11010) );
  AND2_X1 U12421 ( .A1(n11008), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11011) );
  OR3_X1 U12422 ( .A1(n14948), .A2(n11399), .A3(n11058), .ZN(n11012) );
  AND2_X1 U12423 ( .A1(n11000), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11013) );
  AND2_X1 U12424 ( .A1(n11479), .A2(n11478), .ZN(n11014) );
  AND2_X1 U12425 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11015) );
  AND2_X1 U12426 ( .A1(n11293), .A2(n11107), .ZN(n11016) );
  AND3_X1 U12427 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(P3_EAX_REG_28__SCAN_IN), 
        .A3(P3_EAX_REG_27__SCAN_IN), .ZN(n11017) );
  AND2_X2 U12428 ( .A1(n15284), .A2(n11458), .ZN(n12673) );
  NAND3_X1 U12429 ( .A1(n11310), .A2(n11309), .A3(n11307), .ZN(n20269) );
  OR3_X1 U12430 ( .A1(n14864), .A2(n11504), .A3(n15016), .ZN(n11018) );
  OR2_X1 U12431 ( .A1(n20054), .A2(n15040), .ZN(n11019) );
  OR3_X1 U12432 ( .A1(n20632), .A2(n20592), .A3(n11275), .ZN(n11022) );
  AND2_X1 U12433 ( .A1(n10982), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12835) );
  OR3_X1 U12434 ( .A1(n15768), .A2(n11389), .A3(n11392), .ZN(n11023) );
  NAND2_X1 U12435 ( .A1(n12594), .A2(n12605), .ZN(n12599) );
  OR2_X1 U12436 ( .A1(n20732), .A2(n20721), .ZN(n11024) );
  NOR2_X1 U12437 ( .A1(n14538), .A2(n14661), .ZN(n14660) );
  AND2_X1 U12438 ( .A1(n13561), .A2(n13559), .ZN(n11025) );
  OAI21_X1 U12439 ( .B1(n16265), .B2(n11527), .A(n11333), .ZN(n11327) );
  AND2_X1 U12440 ( .A1(n15672), .A2(n15659), .ZN(n15644) );
  NAND2_X1 U12441 ( .A1(n12931), .A2(n11248), .ZN(n11027) );
  AND4_X1 U12442 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11028) );
  NOR3_X1 U12443 ( .A1(n21037), .A2(n21133), .A3(n21036), .ZN(n11029) );
  OR2_X1 U12444 ( .A1(n18099), .A2(n17959), .ZN(n11030) );
  AND2_X1 U12445 ( .A1(n13058), .A2(n13065), .ZN(n11031) );
  OR2_X1 U12446 ( .A1(n17984), .A2(n21031), .ZN(n11033) );
  AND2_X1 U12447 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11034) );
  NOR2_X1 U12448 ( .A1(n16188), .A2(n16171), .ZN(n13160) );
  AND2_X1 U12449 ( .A1(n16628), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16627) );
  INV_X1 U12450 ( .A(n16627), .ZN(n11291) );
  AND3_X1 U12451 ( .A1(n12478), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12477), .ZN(n11035) );
  OR2_X1 U12452 ( .A1(n16467), .A2(n16733), .ZN(n11036) );
  NOR2_X1 U12453 ( .A1(n20620), .A2(n20614), .ZN(n11037) );
  AND2_X1 U12454 ( .A1(n11319), .A2(n14028), .ZN(n14352) );
  NOR2_X1 U12455 ( .A1(n12549), .A2(n12550), .ZN(n11038) );
  INV_X1 U12456 ( .A(n13521), .ZN(n11370) );
  AND2_X1 U12457 ( .A1(n19894), .A2(n13563), .ZN(n11039) );
  NOR2_X1 U12458 ( .A1(n15748), .A2(n15685), .ZN(n15671) );
  NAND2_X1 U12459 ( .A1(n12581), .A2(n12580), .ZN(n13083) );
  AND4_X1 U12460 ( .A1(n15095), .A2(n15094), .A3(n15093), .A4(n15092), .ZN(
        n11040) );
  NAND2_X1 U12461 ( .A1(n16443), .A2(n11464), .ZN(n11460) );
  OR2_X1 U12462 ( .A1(n11025), .A2(n11185), .ZN(n11041) );
  AND2_X1 U12463 ( .A1(n11430), .A2(n11832), .ZN(n11042) );
  NAND2_X1 U12464 ( .A1(n17291), .A2(n13079), .ZN(n16628) );
  AND2_X1 U12465 ( .A1(n13547), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U12466 ( .A1(n12902), .A2(n12903), .ZN(n11044) );
  AND4_X1 U12467 ( .A1(n16488), .A2(n16484), .A3(n16479), .A4(n16478), .ZN(
        n11045) );
  OAI21_X1 U12468 ( .B1(n16637), .B2(n11237), .A(n11234), .ZN(n16475) );
  AND4_X1 U12469 ( .A1(n11112), .A2(n12825), .A3(n12826), .A4(n12831), .ZN(
        n11046) );
  NAND2_X1 U12470 ( .A1(n15260), .A2(n20691), .ZN(n11047) );
  AND2_X1 U12471 ( .A1(n13056), .A2(n13055), .ZN(n11048) );
  NAND2_X1 U12472 ( .A1(n16611), .A2(n16621), .ZN(n11049) );
  OR2_X1 U12473 ( .A1(n13529), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U12474 ( .A1(n19884), .A2(n13562), .ZN(n15950) );
  INV_X1 U12475 ( .A(n11723), .ZN(n11741) );
  AND3_X1 U12476 ( .A1(n12616), .A2(n11139), .A3(n11138), .ZN(n11051) );
  AND3_X1 U12477 ( .A1(n12416), .A2(n12417), .A3(n12450), .ZN(n11052) );
  AND3_X1 U12478 ( .A1(n12421), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12420), .ZN(n11053) );
  AND3_X1 U12479 ( .A1(n11614), .A2(n11619), .A3(n11625), .ZN(n11054) );
  NAND2_X1 U12480 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12848), .ZN(
        n11055) );
  INV_X1 U12481 ( .A(n13079), .ZN(n11421) );
  OR2_X1 U12482 ( .A1(n13077), .A2(n13076), .ZN(n13079) );
  AND2_X1 U12483 ( .A1(n11620), .A2(n11624), .ZN(n11056) );
  AND2_X1 U12484 ( .A1(n11374), .A2(n11372), .ZN(n11057) );
  OR2_X1 U12485 ( .A1(n14953), .A2(n15027), .ZN(n11058) );
  AND2_X1 U12486 ( .A1(n17922), .A2(n11011), .ZN(n11059) );
  INV_X1 U12487 ( .A(n12556), .ZN(n13099) );
  INV_X1 U12488 ( .A(n11765), .ZN(n11212) );
  AND2_X1 U12489 ( .A1(n12014), .A2(n11441), .ZN(n11060) );
  NOR2_X2 U12490 ( .A1(n21021), .A2(n17752), .ZN(n18099) );
  INV_X1 U12491 ( .A(n18099), .ZN(n21034) );
  AND2_X1 U12492 ( .A1(n14685), .A2(n11010), .ZN(n11061) );
  AND2_X1 U12493 ( .A1(n14220), .A2(n11014), .ZN(n11062) );
  OR2_X1 U12494 ( .A1(n14227), .A2(n11340), .ZN(n11063) );
  AND2_X1 U12495 ( .A1(n11502), .A2(n14458), .ZN(n11064) );
  AND2_X1 U12496 ( .A1(n11509), .A2(n11508), .ZN(n11065) );
  INV_X1 U12497 ( .A(n13802), .ZN(n11214) );
  NOR2_X1 U12498 ( .A1(n14538), .A2(n11446), .ZN(n14938) );
  NOR2_X1 U12499 ( .A1(n14431), .A2(n14483), .ZN(n14482) );
  NAND2_X1 U12500 ( .A1(n12533), .A2(n12547), .ZN(n13178) );
  AND2_X1 U12501 ( .A1(n14076), .A2(n11477), .ZN(n11066) );
  OR2_X1 U12502 ( .A1(n20484), .A2(n20485), .ZN(n11067) );
  XOR2_X1 U12503 ( .A(n19945), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n11068) );
  AND2_X1 U12504 ( .A1(n18099), .A2(n21109), .ZN(n11069) );
  NAND2_X1 U12505 ( .A1(n11476), .A2(n11474), .ZN(n11070) );
  NOR3_X1 U12506 ( .A1(n16305), .A2(n16306), .A3(n11347), .ZN(n16287) );
  NOR2_X1 U12507 ( .A1(n16305), .A2(n16306), .ZN(n16294) );
  OR3_X1 U12508 ( .A1(n15768), .A2(n11392), .A3(n11390), .ZN(n11071) );
  AND2_X1 U12509 ( .A1(n15697), .A2(n11452), .ZN(n11072) );
  AND2_X1 U12510 ( .A1(n12692), .A2(n12644), .ZN(n11073) );
  NAND2_X1 U12511 ( .A1(n20649), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20640) );
  INV_X1 U12512 ( .A(n20640), .ZN(n11281) );
  INV_X1 U12513 ( .A(n12867), .ZN(n11237) );
  OR2_X1 U12514 ( .A1(n14864), .A2(n11504), .ZN(n11074) );
  AND2_X1 U12515 ( .A1(n18637), .A2(n12557), .ZN(n11075) );
  OR2_X1 U12516 ( .A1(n12849), .A2(n11247), .ZN(n11076) );
  INV_X1 U12517 ( .A(n17975), .ZN(n18021) );
  NOR2_X1 U12518 ( .A1(n18222), .A2(n18195), .ZN(n17975) );
  OR2_X1 U12519 ( .A1(n15941), .A2(n21361), .ZN(n11077) );
  AND2_X1 U12520 ( .A1(n11641), .A2(n14164), .ZN(n11078) );
  AND2_X1 U12521 ( .A1(n11064), .A2(n11501), .ZN(n11079) );
  AND2_X1 U12522 ( .A1(n11455), .A2(n11454), .ZN(n11080) );
  INV_X1 U12523 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17933) );
  OR2_X1 U12524 ( .A1(n14864), .A2(n14865), .ZN(n11081) );
  INV_X1 U12525 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18340) );
  OR2_X1 U12526 ( .A1(n17954), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11082) );
  OR2_X1 U12527 ( .A1(n18637), .A2(n19272), .ZN(n11083) );
  AND2_X1 U12528 ( .A1(n11014), .A2(n16822), .ZN(n11084) );
  AND2_X1 U12529 ( .A1(n11065), .A2(n11507), .ZN(n11085) );
  OR2_X1 U12530 ( .A1(n11384), .A2(n13585), .ZN(n11086) );
  NOR2_X1 U12531 ( .A1(n21699), .A2(n11729), .ZN(n11087) );
  INV_X1 U12532 ( .A(n18608), .ZN(n18623) );
  NOR2_X1 U12533 ( .A1(n14129), .A2(n14128), .ZN(n14226) );
  AND2_X1 U12534 ( .A1(n18053), .A2(n11313), .ZN(n11088) );
  INV_X1 U12535 ( .A(n15443), .ZN(n11333) );
  NOR2_X1 U12536 ( .A1(n14129), .A2(n11063), .ZN(n14260) );
  AND2_X1 U12537 ( .A1(n11295), .A2(n11297), .ZN(n11089) );
  AND2_X1 U12538 ( .A1(n11489), .A2(n11488), .ZN(n11090) );
  AND2_X1 U12539 ( .A1(n11484), .A2(n11483), .ZN(n11091) );
  NAND2_X1 U12540 ( .A1(n17035), .A2(n14250), .ZN(n21546) );
  INV_X1 U12541 ( .A(n21546), .ZN(n19949) );
  AND2_X1 U12542 ( .A1(n15674), .A2(n15664), .ZN(n11092) );
  NAND2_X1 U12543 ( .A1(n13266), .A2(n13265), .ZN(n14078) );
  NAND3_X1 U12544 ( .A1(n15050), .A2(n15049), .A3(n15048), .ZN(n20738) );
  INV_X1 U12545 ( .A(n12932), .ZN(n11249) );
  INV_X1 U12546 ( .A(n16586), .ZN(n11233) );
  AND2_X1 U12547 ( .A1(n11311), .A2(n20485), .ZN(n11093) );
  AND2_X1 U12548 ( .A1(n12083), .A2(n12082), .ZN(n11094) );
  AND2_X1 U12549 ( .A1(n12161), .A2(n12160), .ZN(n11095) );
  AND2_X1 U12550 ( .A1(n11394), .A2(n11393), .ZN(n11096) );
  AND2_X1 U12551 ( .A1(n11090), .A2(n11487), .ZN(n11097) );
  NOR2_X1 U12552 ( .A1(n14948), .A2(n11396), .ZN(n11401) );
  AND2_X1 U12553 ( .A1(n11337), .A2(n11341), .ZN(n11098) );
  INV_X1 U12554 ( .A(n16296), .ZN(n11347) );
  OR2_X1 U12555 ( .A1(n20473), .A2(n20475), .ZN(n11099) );
  AND2_X1 U12556 ( .A1(n11498), .A2(n11497), .ZN(n11100) );
  AND2_X1 U12557 ( .A1(n11248), .A2(n12943), .ZN(n11101) );
  AND2_X1 U12558 ( .A1(n10974), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U12559 ( .A1(n15021), .A2(n14940), .ZN(n11103) );
  OR2_X1 U12560 ( .A1(n19011), .A2(n18714), .ZN(n18965) );
  INV_X1 U12561 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11318) );
  INV_X1 U12562 ( .A(n14934), .ZN(n11450) );
  AND2_X1 U12563 ( .A1(n20924), .A2(n20903), .ZN(n11104) );
  INV_X1 U12564 ( .A(n16161), .ZN(n11486) );
  AND2_X1 U12565 ( .A1(n13471), .A2(n21852), .ZN(n19948) );
  OR2_X1 U12566 ( .A1(n21129), .A2(n20457), .ZN(n11105) );
  INV_X1 U12567 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11427) );
  AND2_X1 U12568 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n11106) );
  INV_X1 U12569 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11315) );
  INV_X1 U12570 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11314) );
  INV_X1 U12571 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n11276) );
  AND2_X1 U12572 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11107) );
  OR2_X1 U12573 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11108) );
  INV_X1 U12574 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11302) );
  AND2_X1 U12575 ( .A1(n11016), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11109) );
  XNOR2_X2 U12576 ( .A(n13070), .B(n13071), .ZN(n13057) );
  NAND4_X1 U12577 ( .A1(n11046), .A2(n12823), .A3(n12824), .A4(n11111), .ZN(
        n11110) );
  NAND3_X1 U12578 ( .A1(n12693), .A2(n11222), .A3(n11469), .ZN(n12740) );
  AND2_X2 U12579 ( .A1(n11121), .A2(n11117), .ZN(n12597) );
  NAND3_X1 U12580 ( .A1(n11263), .A2(n12592), .A3(n12593), .ZN(n11117) );
  OAI21_X1 U12581 ( .B1(n12582), .B2(n12568), .A(n11119), .ZN(n11118) );
  NAND2_X1 U12582 ( .A1(n12574), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U12583 ( .A1(n11123), .A2(n11263), .ZN(n11121) );
  NAND4_X1 U12584 ( .A1(n11038), .A2(n12534), .A3(n12535), .A4(n12551), .ZN(
        n11263) );
  NAND2_X1 U12585 ( .A1(n12574), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U12586 ( .A1(n13178), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11122) );
  AND2_X2 U12587 ( .A1(n11055), .A2(n11124), .ZN(n16637) );
  NAND2_X1 U12588 ( .A1(n16942), .A2(n16943), .ZN(n11124) );
  XNOR2_X1 U12589 ( .A(n12848), .B(n18597), .ZN(n16943) );
  AND2_X2 U12590 ( .A1(n11126), .A2(n11125), .ZN(n16942) );
  NAND2_X1 U12591 ( .A1(n11224), .A2(n14831), .ZN(n11126) );
  NOR2_X2 U12592 ( .A1(n16421), .A2(n16395), .ZN(n16398) );
  NAND3_X1 U12593 ( .A1(n11129), .A2(n11128), .A3(n11045), .ZN(n16466) );
  NAND4_X1 U12594 ( .A1(n12531), .A2(n13224), .A3(n12532), .A4(n12567), .ZN(
        n11409) );
  NAND3_X1 U12595 ( .A1(n11130), .A2(n11051), .A3(n12626), .ZN(n11222) );
  NAND3_X1 U12596 ( .A1(n11141), .A2(n11133), .A3(n11142), .ZN(n11131) );
  NAND4_X1 U12597 ( .A1(n11140), .A2(n11143), .A3(n11144), .A4(n12604), .ZN(
        n11132) );
  NOR2_X2 U12598 ( .A1(n12619), .A2(n12611), .ZN(n14881) );
  NOR2_X2 U12599 ( .A1(n12621), .A2(n12611), .ZN(n19236) );
  NOR2_X2 U12600 ( .A1(n12621), .A2(n12618), .ZN(n14602) );
  NOR2_X2 U12601 ( .A1(n12619), .A2(n12620), .ZN(n19250) );
  NAND2_X1 U12602 ( .A1(n14778), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11144) );
  OR2_X2 U12603 ( .A1(n13180), .A2(n11145), .ZN(n12570) );
  NAND3_X1 U12604 ( .A1(n11004), .A2(n11146), .A3(n18623), .ZN(n11148) );
  NAND2_X1 U12605 ( .A1(n11148), .A2(n16801), .ZN(P2_U3028) );
  NAND2_X2 U12606 ( .A1(n11149), .A2(n13067), .ZN(n13066) );
  NAND2_X1 U12607 ( .A1(n14615), .A2(n14838), .ZN(n11153) );
  NAND2_X1 U12608 ( .A1(n11152), .A2(n14615), .ZN(n11150) );
  INV_X1 U12609 ( .A(n11156), .ZN(n11154) );
  INV_X1 U12610 ( .A(n12578), .ZN(n11155) );
  NAND2_X1 U12611 ( .A1(n12578), .A2(n11156), .ZN(n12579) );
  NOR2_X4 U12612 ( .A1(n16577), .A2(n16854), .ZN(n16551) );
  INV_X2 U12613 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20680) );
  NAND2_X2 U12614 ( .A1(n20720), .A2(n11282), .ZN(n20696) );
  NAND3_X1 U12615 ( .A1(n15106), .A2(n15107), .A3(n11162), .ZN(n11161) );
  AND2_X2 U12616 ( .A1(n18106), .A2(n21083), .ZN(n18064) );
  NOR2_X2 U12617 ( .A1(n21162), .A2(n21218), .ZN(n21224) );
  AND2_X2 U12618 ( .A1(n21177), .A2(n17784), .ZN(n21138) );
  NOR2_X2 U12619 ( .A1(n16991), .A2(n16992), .ZN(n21177) );
  NAND2_X1 U12620 ( .A1(n11653), .A2(n11165), .ZN(n13813) );
  OAI22_X1 U12621 ( .A1(n15546), .A2(n11165), .B1(n15545), .B2(n15544), .ZN(
        n19953) );
  NAND2_X1 U12622 ( .A1(n14372), .A2(n11165), .ZN(n14361) );
  AND2_X2 U12623 ( .A1(n11638), .A2(n12382), .ZN(n11724) );
  NAND3_X1 U12624 ( .A1(n11172), .A2(n11365), .A3(n11363), .ZN(n11171) );
  INV_X1 U12625 ( .A(n13539), .ZN(n14582) );
  NAND3_X1 U12626 ( .A1(n21679), .A2(n11213), .A3(n11740), .ZN(n11187) );
  INV_X1 U12627 ( .A(n21037), .ZN(n18045) );
  OAI21_X1 U12628 ( .B1(n21039), .B2(n11191), .A(n11189), .ZN(P3_U2834) );
  INV_X1 U12629 ( .A(n21020), .ZN(n11195) );
  OAI21_X1 U12630 ( .B1(n21033), .B2(n21021), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U12631 ( .A1(n21018), .A2(n21019), .ZN(n21033) );
  NAND2_X1 U12632 ( .A1(n13802), .A2(n11765), .ZN(n11207) );
  INV_X1 U12633 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n11213) );
  NAND2_X4 U12634 ( .A1(n11360), .A2(n11626), .ZN(n14364) );
  NAND3_X1 U12635 ( .A1(n13530), .A2(n13531), .A3(n13786), .ZN(n11217) );
  OR2_X2 U12636 ( .A1(n11887), .A2(n11886), .ZN(n13530) );
  AND2_X2 U12637 ( .A1(n16097), .A2(n13958), .ZN(n11708) );
  NAND2_X1 U12638 ( .A1(n11785), .A2(n11219), .ZN(n11879) );
  INV_X1 U12639 ( .A(n11879), .ZN(n11810) );
  OAI21_X1 U12640 ( .B1(n13538), .B2(n11364), .A(n19879), .ZN(n11220) );
  INV_X1 U12641 ( .A(n11220), .ZN(n11363) );
  NAND2_X1 U12642 ( .A1(n11222), .A2(n12644), .ZN(n11284) );
  NAND2_X1 U12643 ( .A1(n14830), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11224) );
  INV_X1 U12644 ( .A(n14830), .ZN(n11225) );
  NAND2_X1 U12645 ( .A1(n16695), .A2(n11226), .ZN(P2_U3021) );
  NAND2_X1 U12646 ( .A1(n16637), .A2(n11232), .ZN(n11228) );
  NAND2_X1 U12647 ( .A1(n11229), .A2(n11228), .ZN(n12918) );
  NAND2_X2 U12648 ( .A1(n12636), .A2(n10966), .ZN(n15470) );
  NAND2_X1 U12649 ( .A1(n13243), .A2(n13182), .ZN(n11242) );
  NAND3_X2 U12650 ( .A1(n12415), .A2(n11243), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12431) );
  NAND2_X1 U12651 ( .A1(n12931), .A2(n11101), .ZN(n12945) );
  NAND2_X1 U12652 ( .A1(n12902), .A2(n11253), .ZN(n12916) );
  NAND2_X1 U12653 ( .A1(n12902), .A2(n11251), .ZN(n12928) );
  NOR2_X2 U12654 ( .A1(n18130), .A2(n17822), .ZN(n17846) );
  NOR2_X2 U12656 ( .A1(n18188), .A2(n17803), .ZN(n17806) );
  INV_X1 U12657 ( .A(n17794), .ZN(n17795) );
  NOR2_X1 U12658 ( .A1(n18201), .A2(n18200), .ZN(n18199) );
  XNOR2_X1 U12659 ( .A(n17797), .B(n20789), .ZN(n18201) );
  NAND2_X1 U12660 ( .A1(n17796), .A2(n17798), .ZN(n11254) );
  AND2_X2 U12661 ( .A1(n12693), .A2(n12692), .ZN(n11283) );
  INV_X1 U12662 ( .A(n11461), .ZN(n11266) );
  OAI21_X2 U12663 ( .B1(n11268), .B2(n11266), .A(n11265), .ZN(n15504) );
  INV_X1 U12664 ( .A(n11459), .ZN(n11270) );
  INV_X1 U12665 ( .A(n12956), .ZN(n11271) );
  INV_X1 U12666 ( .A(n20593), .ZN(n20625) );
  NAND2_X1 U12667 ( .A1(n20621), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n20620) );
  NAND2_X1 U12668 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  XNOR2_X2 U12669 ( .A(n11284), .B(n11283), .ZN(n14533) );
  NOR2_X1 U12670 ( .A1(n13197), .A2(n18340), .ZN(n11286) );
  NAND2_X1 U12671 ( .A1(n16551), .A2(n11109), .ZN(n11292) );
  NAND2_X1 U12672 ( .A1(n16551), .A2(n11016), .ZN(n16517) );
  AND2_X1 U12673 ( .A1(n16551), .A2(n11293), .ZN(n16527) );
  NAND2_X1 U12674 ( .A1(n16551), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16820) );
  NAND2_X1 U12675 ( .A1(n11292), .A2(n16763), .ZN(n16500) );
  OR2_X1 U12676 ( .A1(n20342), .A2(n11296), .ZN(n11294) );
  INV_X1 U12677 ( .A(n11298), .ZN(n20356) );
  INV_X1 U12678 ( .A(n20103), .ZN(n11299) );
  NAND2_X1 U12679 ( .A1(n11306), .A2(n11303), .ZN(P3_U2640) );
  NOR2_X1 U12680 ( .A1(n20459), .A2(n20458), .ZN(n20474) );
  INV_X1 U12681 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11317) );
  AND2_X4 U12682 ( .A1(n12635), .A2(n10966), .ZN(n12501) );
  AND2_X2 U12683 ( .A1(n11243), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12635) );
  NAND2_X1 U12684 ( .A1(n14353), .A2(n14352), .ZN(n14030) );
  NAND2_X1 U12685 ( .A1(n11320), .A2(n14026), .ZN(n11319) );
  NAND2_X1 U12686 ( .A1(n14021), .A2(n14022), .ZN(n11320) );
  INV_X1 U12687 ( .A(n14129), .ZN(n11337) );
  NAND2_X1 U12688 ( .A1(n11337), .A2(n11338), .ZN(n14420) );
  OAI22_X2 U12689 ( .A1(n16305), .A2(n11343), .B1(n18335), .B2(n15424), .ZN(
        n16280) );
  OAI21_X2 U12690 ( .B1(n11723), .B2(n11541), .A(n11652), .ZN(n11728) );
  NAND3_X1 U12691 ( .A1(n11056), .A2(n11621), .A3(n11623), .ZN(n11356) );
  NAND4_X1 U12692 ( .A1(n11359), .A2(n11054), .A3(n11358), .A4(n11622), .ZN(
        n11357) );
  NAND3_X1 U12693 ( .A1(n15903), .A2(n13584), .A3(n11361), .ZN(n15867) );
  XNOR2_X1 U12694 ( .A(n11362), .B(n15898), .ZN(n16030) );
  INV_X1 U12695 ( .A(n14244), .ZN(n11369) );
  NAND2_X1 U12696 ( .A1(n11373), .A2(n11057), .ZN(n13576) );
  NAND3_X1 U12697 ( .A1(n11379), .A2(n11380), .A3(n11381), .ZN(n13593) );
  NAND2_X1 U12698 ( .A1(n15877), .A2(n11009), .ZN(n11381) );
  NAND3_X1 U12699 ( .A1(n11381), .A2(n11382), .A3(n11379), .ZN(n15996) );
  NAND2_X1 U12700 ( .A1(n13579), .A2(n19945), .ZN(n15911) );
  INV_X1 U12701 ( .A(n11401), .ZN(n15791) );
  NAND2_X1 U12702 ( .A1(n12441), .A2(n12450), .ZN(n11407) );
  NAND2_X1 U12703 ( .A1(n11409), .A2(n14332), .ZN(n12537) );
  INV_X1 U12704 ( .A(n12527), .ZN(n11408) );
  NAND2_X1 U12705 ( .A1(n11410), .A2(n11412), .ZN(n16945) );
  NAND2_X1 U12706 ( .A1(n13058), .A2(n13062), .ZN(n11416) );
  OAI21_X1 U12707 ( .B1(n13055), .B2(n13056), .A(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11415) );
  NAND2_X1 U12708 ( .A1(n16640), .A2(n13075), .ZN(n17293) );
  NOR2_X2 U12709 ( .A1(n11426), .A2(n11425), .ZN(n16441) );
  NOR2_X2 U12710 ( .A1(n11427), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13840) );
  NAND3_X1 U12711 ( .A1(n14192), .A2(n11429), .A3(n14170), .ZN(n14191) );
  NAND2_X1 U12712 ( .A1(n14170), .A2(n14169), .ZN(n14168) );
  OAI21_X1 U12713 ( .B1(n11836), .B2(n11766), .A(n11434), .ZN(n11433) );
  NAND2_X1 U12714 ( .A1(n12014), .A2(n11436), .ZN(n15777) );
  INV_X1 U12715 ( .A(n14538), .ZN(n11443) );
  NAND2_X1 U12716 ( .A1(n11443), .A2(n11444), .ZN(n14987) );
  NAND2_X1 U12717 ( .A1(n12084), .A2(n11451), .ZN(n15755) );
  NAND2_X1 U12718 ( .A1(n15672), .A2(n11455), .ZN(n15617) );
  AND2_X1 U12719 ( .A1(n15672), .A2(n11456), .ZN(n15632) );
  INV_X1 U12720 ( .A(n15620), .ZN(n11454) );
  AND3_X4 U12721 ( .A1(n12415), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15466) );
  INV_X1 U12722 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11464) );
  NAND2_X1 U12723 ( .A1(n12535), .A2(n12534), .ZN(n12553) );
  NAND2_X1 U12724 ( .A1(n11038), .A2(n12551), .ZN(n12552) );
  AND2_X1 U12725 ( .A1(n14021), .A2(n18587), .ZN(n12614) );
  XNOR2_X2 U12726 ( .A(n13083), .B(n13086), .ZN(n14021) );
  INV_X2 U12727 ( .A(n12461), .ZN(n12532) );
  OR2_X1 U12728 ( .A1(n13417), .A2(n12555), .ZN(n11471) );
  AND2_X2 U12729 ( .A1(n13228), .A2(n13182), .ZN(n13375) );
  MUX2_X1 U12730 ( .A(n12770), .B(n12769), .S(n13182), .Z(n12802) );
  MUX2_X1 U12731 ( .A(n12978), .B(n12977), .S(n13182), .Z(n16141) );
  NOR2_X2 U12732 ( .A1(n14083), .A2(n11472), .ZN(n16893) );
  NOR2_X1 U12733 ( .A1(n11020), .A2(n16172), .ZN(n16162) );
  OR3_X1 U12734 ( .A1(n11020), .A2(n11482), .A3(n16172), .ZN(n15511) );
  NAND3_X1 U12735 ( .A1(n11052), .A2(n12418), .A3(n12419), .ZN(n11490) );
  NAND3_X1 U12736 ( .A1(n11053), .A2(n12422), .A3(n12423), .ZN(n11491) );
  NAND2_X1 U12737 ( .A1(n12582), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12573) );
  NAND3_X1 U12738 ( .A1(n11506), .A2(n11505), .A3(n14970), .ZN(n11504) );
  NAND2_X1 U12739 ( .A1(n15864), .A2(n12397), .ZN(n12409) );
  NAND2_X1 U12740 ( .A1(n12335), .A2(n21667), .ZN(n11637) );
  NOR2_X2 U12741 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U12742 ( .A1(n12162), .A2(n11095), .ZN(n15748) );
  NAND2_X1 U12743 ( .A1(n18335), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13761) );
  NOR2_X1 U12744 ( .A1(n12547), .A2(n18335), .ZN(n12536) );
  NAND2_X1 U12745 ( .A1(n16152), .A2(n18625), .ZN(n13458) );
  NAND2_X1 U12746 ( .A1(n11078), .A2(n11516), .ZN(n13788) );
  AOI211_X2 U12747 ( .C1(n16650), .C2(n16653), .A(n16649), .B(n16648), .ZN(
        n16651) );
  AND2_X2 U12748 ( .A1(n11539), .A2(n11540), .ZN(n11752) );
  NOR2_X1 U12749 ( .A1(n13466), .A2(n13465), .ZN(n13470) );
  NAND2_X1 U12750 ( .A1(n11740), .A2(n11739), .ZN(n11748) );
  INV_X1 U12751 ( .A(n14432), .ZN(n11893) );
  INV_X1 U12752 ( .A(n14987), .ZN(n12014) );
  INV_X1 U12753 ( .A(n14048), .ZN(n11854) );
  OR2_X2 U12754 ( .A1(n14021), .A2(n18624), .ZN(n12619) );
  AND2_X1 U12755 ( .A1(n14021), .A2(n12595), .ZN(n12598) );
  AOI21_X1 U12756 ( .B1(n15605), .B2(n15618), .A(n15604), .ZN(n15875) );
  INV_X1 U12757 ( .A(n15755), .ZN(n12162) );
  AOI21_X2 U12758 ( .B1(n16462), .B2(n16458), .A(n16459), .ZN(n16445) );
  NAND2_X1 U12759 ( .A1(n13170), .A2(n13450), .ZN(n13177) );
  INV_X1 U12760 ( .A(n15671), .ZN(n15684) );
  NAND2_X1 U12761 ( .A1(n15549), .A2(n12396), .ZN(n12414) );
  NOR2_X1 U12762 ( .A1(n13508), .A2(n21752), .ZN(n21770) );
  AND2_X1 U12763 ( .A1(n21752), .A2(n14066), .ZN(n21742) );
  AND2_X1 U12764 ( .A1(n11856), .A2(n21752), .ZN(n21822) );
  AND2_X1 U12765 ( .A1(n15434), .A2(n15439), .ZN(n11512) );
  OR2_X1 U12766 ( .A1(n13459), .A2(n18608), .ZN(n11513) );
  INV_X1 U12767 ( .A(n15864), .ZN(n21649) );
  AOI21_X2 U12768 ( .B1(n13779), .B2(n12395), .A(n21561), .ZN(n15864) );
  INV_X1 U12769 ( .A(n21649), .ZN(n15852) );
  OR2_X1 U12770 ( .A1(n13247), .A2(n13246), .ZN(n11514) );
  INV_X1 U12771 ( .A(n13219), .ZN(n13391) );
  INV_X1 U12772 ( .A(n13218), .ZN(n13390) );
  AND2_X1 U12773 ( .A1(n14165), .A2(n14112), .ZN(n11516) );
  OR2_X1 U12774 ( .A1(n19276), .A2(n18637), .ZN(n18488) );
  OR2_X1 U12775 ( .A1(n15596), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11517) );
  INV_X1 U12776 ( .A(n13649), .ZN(n15486) );
  OR2_X1 U12777 ( .A1(n15596), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11518) );
  INV_X2 U12778 ( .A(n18965), .ZN(n19012) );
  INV_X1 U12779 ( .A(n19830), .ZN(n19838) );
  AND3_X1 U12780 ( .A1(n12474), .A2(n12450), .A3(n12473), .ZN(n11519) );
  NAND2_X1 U12781 ( .A1(n12789), .A2(n18362), .ZN(n14830) );
  INV_X2 U12782 ( .A(n17658), .ZN(n17654) );
  AND3_X1 U12783 ( .A1(n12489), .A2(n12488), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11520) );
  OR2_X1 U12784 ( .A1(n15596), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11521) );
  INV_X1 U12785 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18581) );
  OR2_X1 U12786 ( .A1(n15596), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11522) );
  AND3_X1 U12787 ( .A1(n12443), .A2(n12442), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11523) );
  AND3_X1 U12788 ( .A1(n12426), .A2(n12425), .A3(n12450), .ZN(n11524) );
  NOR2_X1 U12789 ( .A1(n21773), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11525) );
  OR2_X1 U12790 ( .A1(n16278), .A2(n15432), .ZN(n11526) );
  AND2_X1 U12791 ( .A1(n15437), .A2(n11512), .ZN(n11527) );
  AND3_X1 U12792 ( .A1(n12654), .A2(n12653), .A3(n12652), .ZN(n11528) );
  AND4_X1 U12793 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11529) );
  AND2_X2 U12794 ( .A1(n11537), .A2(n16097), .ZN(n11758) );
  AND2_X2 U12795 ( .A1(n11539), .A2(n16097), .ZN(n11681) );
  AND2_X1 U12796 ( .A1(n11658), .A2(n13805), .ZN(n11530) );
  INV_X1 U12797 ( .A(n13488), .ZN(n11648) );
  INV_X1 U12798 ( .A(n19138), .ZN(n12820) );
  AOI22_X1 U12799 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19190), .B1(
        n19160), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U12800 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12615), .B1(
        n19138), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12616) );
  INV_X1 U12801 ( .A(n12334), .ZN(n12342) );
  NAND2_X1 U12802 ( .A1(n12332), .A2(n12331), .ZN(n12361) );
  INV_X1 U12803 ( .A(n13420), .ZN(n12526) );
  INV_X1 U12804 ( .A(n14750), .ZN(n12494) );
  AND2_X1 U12805 ( .A1(n17062), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12371) );
  OR2_X1 U12806 ( .A1(n12174), .A2(n12173), .ZN(n12197) );
  AOI22_X1 U12807 ( .A1(n12556), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U12808 ( .A1(n12526), .A2(n12525), .ZN(n12554) );
  NAND2_X1 U12809 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14443), .ZN(
        n12373) );
  NAND2_X1 U12810 ( .A1(n12345), .A2(n13786), .ZN(n12375) );
  AND2_X1 U12811 ( .A1(n13548), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13549) );
  INV_X1 U12812 ( .A(n11697), .ZN(n11698) );
  INV_X1 U12813 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11531) );
  AND4_X1 U12814 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12756) );
  XNOR2_X1 U12815 ( .A(n12450), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12776) );
  OR2_X1 U12816 ( .A1(n12322), .A2(n15881), .ZN(n13478) );
  INV_X1 U12817 ( .A(n12179), .ZN(n12180) );
  INV_X1 U12818 ( .A(n11977), .ZN(n11978) );
  INV_X1 U12819 ( .A(n14583), .ZN(n13538) );
  OR2_X1 U12820 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  NAND2_X1 U12821 ( .A1(n13827), .A2(n11213), .ZN(n11784) );
  NOR2_X1 U12822 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17003), .ZN(
        n12994) );
  INV_X1 U12823 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14713) );
  INV_X1 U12824 ( .A(n13264), .ZN(n12847) );
  INV_X1 U12825 ( .A(n14422), .ZN(n14419) );
  AND2_X1 U12826 ( .A1(n13385), .A2(n13384), .ZN(n16790) );
  NOR2_X1 U12827 ( .A1(n16396), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12957) );
  AND2_X1 U12828 ( .A1(n13084), .A2(n12591), .ZN(n13086) );
  AND2_X1 U12829 ( .A1(n13044), .A2(n13243), .ZN(n13042) );
  INV_X1 U12830 ( .A(n12628), .ZN(n14278) );
  NOR2_X1 U12831 ( .A1(n20680), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n15256) );
  INV_X1 U12832 ( .A(n20734), .ZN(n15249) );
  NAND2_X1 U12833 ( .A1(n14663), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14362) );
  AND2_X1 U12834 ( .A1(n14363), .A2(n21829), .ZN(n14373) );
  OR2_X1 U12835 ( .A1(n12382), .A2(n13629), .ZN(n13654) );
  NAND2_X1 U12836 ( .A1(n12265), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12322) );
  INV_X1 U12837 ( .A(n12320), .ZN(n12286) );
  NAND2_X1 U12838 ( .A1(n11874), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11880) );
  NAND2_X1 U12839 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  OR2_X1 U12840 ( .A1(n13574), .A2(n15951), .ZN(n19919) );
  INV_X1 U12841 ( .A(n13510), .ZN(n13786) );
  NAND2_X1 U12842 ( .A1(n11841), .A2(n11842), .ZN(n11845) );
  NAND2_X1 U12843 ( .A1(n11771), .A2(n11770), .ZN(n21715) );
  NAND2_X1 U12844 ( .A1(n12516), .A2(n18334), .ZN(n12989) );
  AOI221_X1 U12845 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12995), 
        .C1(n18581), .C2(n12995), .A(n12994), .ZN(n13030) );
  INV_X1 U12846 ( .A(n14656), .ZN(n14653) );
  NAND2_X1 U12847 ( .A1(n18349), .A2(n14022), .ZN(n13760) );
  AND2_X1 U12848 ( .A1(n13405), .A2(n13404), .ZN(n16172) );
  AND2_X1 U12849 ( .A1(n13762), .A2(n15487), .ZN(n15439) );
  AND3_X1 U12850 ( .A1(n13312), .A2(n13311), .A3(n13310), .ZN(n14800) );
  NAND2_X1 U12851 ( .A1(n16133), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16132) );
  OR2_X1 U12852 ( .A1(n16122), .A2(n16121), .ZN(n16124) );
  INV_X1 U12853 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14698) );
  NOR2_X1 U12854 ( .A1(n15519), .A2(n15518), .ZN(n15520) );
  AND3_X1 U12855 ( .A1(n16544), .A2(n16528), .A3(n16532), .ZN(n16481) );
  AND2_X1 U12856 ( .A1(n14819), .A2(n12876), .ZN(n16586) );
  INV_X1 U12857 ( .A(n14774), .ZN(n14778) );
  INV_X1 U12858 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16962) );
  OAI21_X1 U12859 ( .B1(n15247), .B2(n21158), .A(n21196), .ZN(n16992) );
  INV_X1 U12860 ( .A(n17835), .ZN(n17913) );
  OAI21_X1 U12861 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n20741) );
  NAND2_X1 U12862 ( .A1(n11908), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11922) );
  NOR2_X1 U12863 ( .A1(n11880), .A2(n19877), .ZN(n11888) );
  NOR2_X1 U12864 ( .A1(n14362), .A2(n21667), .ZN(n14374) );
  NAND2_X1 U12865 ( .A1(n15852), .A2(n15798), .ZN(n21636) );
  INV_X1 U12866 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15915) );
  INV_X1 U12867 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15936) );
  INV_X1 U12868 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15970) );
  NOR2_X1 U12869 ( .A1(n13789), .A2(n13806), .ZN(n14102) );
  AND2_X1 U12870 ( .A1(n15567), .A2(n15566), .ZN(n15767) );
  AND2_X1 U12871 ( .A1(n14952), .A2(n14951), .ZN(n15027) );
  INV_X1 U12872 ( .A(n14900), .ZN(n13561) );
  AND2_X1 U12873 ( .A1(n14118), .A2(n15535), .ZN(n21325) );
  NAND2_X1 U12874 ( .A1(n22037), .A2(n14364), .ZN(n13510) );
  AND2_X1 U12875 ( .A1(n21239), .A2(n21238), .ZN(n21328) );
  INV_X1 U12876 ( .A(n21325), .ZN(n21367) );
  AND2_X1 U12877 ( .A1(n21841), .A2(n11768), .ZN(n21754) );
  INV_X1 U12878 ( .A(n21702), .ZN(n21711) );
  INV_X1 U12879 ( .A(n11856), .ZN(n14066) );
  NOR2_X1 U12880 ( .A1(n21799), .A2(n22129), .ZN(n21780) );
  INV_X1 U12881 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21810) );
  NAND3_X1 U12882 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n11213), .A3(n21666), 
        .ZN(n22132) );
  NAND2_X1 U12883 ( .A1(n13797), .A2(n13796), .ZN(n17044) );
  NOR2_X1 U12884 ( .A1(n13180), .A2(n13183), .ZN(n14327) );
  INV_X1 U12885 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18514) );
  AND2_X1 U12886 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n13435), .ZN(
        n16117) );
  INV_X1 U12887 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18425) );
  AND2_X1 U12888 ( .A1(n14707), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14709) );
  INV_X1 U12889 ( .A(n18528), .ZN(n18562) );
  NAND2_X1 U12890 ( .A1(n18562), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18564) );
  NAND2_X1 U12891 ( .A1(n15461), .A2(n15460), .ZN(n16248) );
  OR2_X1 U12892 ( .A1(n15438), .A2(n15442), .ZN(n16255) );
  INV_X1 U12893 ( .A(n15432), .ZN(n15429) );
  AND3_X1 U12894 ( .A1(n13325), .A2(n13324), .A3(n13323), .ZN(n16892) );
  NAND2_X1 U12895 ( .A1(n19594), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12998) );
  INV_X1 U12896 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18548) );
  NOR2_X1 U12897 ( .A1(n14705), .A2(n14698), .ZN(n14707) );
  INV_X1 U12898 ( .A(n13456), .ZN(n13457) );
  INV_X1 U12899 ( .A(n18603), .ZN(n18628) );
  AND2_X1 U12900 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19243) );
  AND2_X1 U12901 ( .A1(n19281), .A2(n19282), .ZN(n19231) );
  OR2_X1 U12902 ( .A1(n19162), .A2(n19491), .ZN(n19185) );
  NAND2_X1 U12903 ( .A1(n14594), .A2(n14593), .ZN(n19281) );
  NAND2_X1 U12904 ( .A1(n19263), .A2(n19262), .ZN(n19276) );
  NOR2_X1 U12905 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20328), .ZN(n20344) );
  NOR2_X1 U12906 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20239), .ZN(n20258) );
  NOR2_X1 U12907 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20188), .ZN(n20207) );
  INV_X1 U12908 ( .A(n20173), .ZN(n20192) );
  OR3_X1 U12909 ( .A1(n20738), .A2(n20495), .A3(n20494), .ZN(n20496) );
  INV_X1 U12910 ( .A(n20877), .ZN(n20876) );
  INV_X1 U12911 ( .A(n21021), .ZN(n20749) );
  INV_X1 U12912 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21169) );
  NOR3_X1 U12913 ( .A1(n17782), .A2(n20737), .A3(n20691), .ZN(n17785) );
  AND2_X1 U12914 ( .A1(n15629), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15614) );
  NOR2_X1 U12915 ( .A1(n15657), .A2(n17139), .ZN(n15647) );
  NOR2_X1 U12916 ( .A1(n21533), .A2(n21534), .ZN(n15690) );
  INV_X1 U12917 ( .A(n21475), .ZN(n21473) );
  AND2_X1 U12918 ( .A1(n14663), .A2(n14360), .ZN(n21525) );
  NOR2_X1 U12919 ( .A1(n19955), .A2(n15550), .ZN(n21495) );
  AND2_X1 U12920 ( .A1(n14374), .A2(n14366), .ZN(n21529) );
  AND2_X1 U12921 ( .A1(n14190), .A2(n14189), .ZN(n14198) );
  AND2_X1 U12922 ( .A1(n19870), .A2(n22131), .ZN(n19865) );
  NOR2_X2 U12923 ( .A1(n12409), .A2(n21662), .ZN(n21652) );
  INV_X1 U12924 ( .A(n19915), .ZN(n21664) );
  INV_X1 U12925 ( .A(n19901), .ZN(n19943) );
  INV_X1 U12926 ( .A(n21561), .ZN(n14250) );
  AND3_X1 U12927 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n21308), .ZN(n21240) );
  NOR2_X1 U12928 ( .A1(n21328), .A2(n14174), .ZN(n21310) );
  INV_X1 U12929 ( .A(n21239), .ZN(n21415) );
  INV_X1 U12930 ( .A(n21786), .ZN(n21701) );
  AND2_X1 U12931 ( .A1(n21702), .A2(n21793), .ZN(n22143) );
  AND2_X1 U12932 ( .A1(n21687), .A2(n21686), .ZN(n21816) );
  NOR2_X2 U12933 ( .A1(n21711), .A2(n21688), .ZN(n22156) );
  NOR2_X2 U12934 ( .A1(n21711), .A2(n21789), .ZN(n22163) );
  AND2_X1 U12935 ( .A1(n21742), .A2(n21816), .ZN(n22174) );
  NOR2_X1 U12936 ( .A1(n21687), .A2(n13484), .ZN(n21741) );
  AND2_X1 U12937 ( .A1(n21770), .A2(n21816), .ZN(n22199) );
  AND2_X1 U12938 ( .A1(n21783), .A2(n21832), .ZN(n21776) );
  NOR2_X2 U12939 ( .A1(n21790), .A2(n21789), .ZN(n22213) );
  AND2_X1 U12940 ( .A1(n21687), .A2(n13484), .ZN(n21793) );
  NOR2_X2 U12941 ( .A1(n21818), .A2(n21817), .ZN(n22228) );
  NAND2_X1 U12942 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21229) );
  AND2_X1 U12943 ( .A1(n21580), .A2(n11628), .ZN(n13777) );
  NOR2_X1 U12944 ( .A1(n13000), .A2(n12999), .ZN(n14591) );
  NAND2_X1 U12945 ( .A1(n16118), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16120) );
  INV_X1 U12946 ( .A(n18576), .ZN(n18531) );
  INV_X1 U12947 ( .A(n18488), .ZN(n18427) );
  AND2_X1 U12948 ( .A1(n14709), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14710) );
  INV_X1 U12949 ( .A(n18564), .ZN(n18529) );
  INV_X1 U12950 ( .A(n18511), .ZN(n18570) );
  OR2_X1 U12951 ( .A1(n15421), .A2(n15420), .ZN(n16288) );
  OR2_X1 U12952 ( .A1(n13284), .A2(n13283), .ZN(n14229) );
  OR2_X1 U12953 ( .A1(n15013), .A2(n15012), .ZN(n15015) );
  NAND2_X1 U12954 ( .A1(n13971), .A2(n18345), .ZN(n13973) );
  NOR2_X1 U12955 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17303), .ZN(n17358) );
  INV_X1 U12956 ( .A(n14633), .ZN(n13743) );
  NAND2_X1 U12957 ( .A1(n13464), .A2(n13463), .ZN(n13465) );
  NAND2_X1 U12958 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n14704), .ZN(
        n14703) );
  AND2_X1 U12959 ( .A1(n17268), .A2(n13751), .ZN(n17260) );
  INV_X1 U12960 ( .A(n17295), .ZN(n17274) );
  INV_X1 U12961 ( .A(n16466), .ZN(n16469) );
  NAND2_X1 U12962 ( .A1(n13040), .A2(n18345), .ZN(n13423) );
  OR2_X1 U12963 ( .A1(n13423), .A2(n13179), .ZN(n18607) );
  INV_X1 U12964 ( .A(n19276), .ZN(n19282) );
  OAI21_X1 U12965 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n19703) );
  NOR2_X2 U12966 ( .A1(n19279), .A2(n19182), .ZN(n19701) );
  OAI21_X1 U12967 ( .B1(n19268), .B2(n19276), .A(n19267), .ZN(n19687) );
  AND2_X1 U12968 ( .A1(n19257), .A2(n19242), .ZN(n19686) );
  OAI21_X1 U12969 ( .B1(n19239), .B2(n19238), .A(n19237), .ZN(n19672) );
  INV_X1 U12970 ( .A(n19564), .ZN(n19671) );
  INV_X1 U12971 ( .A(n19669), .ZN(n19659) );
  INV_X1 U12972 ( .A(n19649), .ZN(n19636) );
  OAI21_X1 U12973 ( .B1(n19179), .B2(n19178), .A(n19177), .ZN(n19631) );
  INV_X1 U12974 ( .A(n19628), .ZN(n19630) );
  OAI21_X1 U12975 ( .B1(n19157), .B2(n19156), .A(n19155), .ZN(n19618) );
  OAI21_X1 U12976 ( .B1(n14777), .B2(n14776), .A(n14775), .ZN(n19611) );
  INV_X1 U12977 ( .A(n19334), .ZN(n19337) );
  NOR2_X1 U12978 ( .A1(n10974), .A2(n14781), .ZN(n19388) );
  INV_X1 U12979 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19263) );
  INV_X1 U12980 ( .A(n18655), .ZN(n21594) );
  AND2_X1 U12981 ( .A1(n21612), .A2(n21598), .ZN(n17382) );
  INV_X1 U12982 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n16997) );
  NOR2_X1 U12983 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20380), .ZN(n20398) );
  NOR2_X1 U12984 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20355), .ZN(n20371) );
  NAND2_X1 U12985 ( .A1(n20061), .A2(n20062), .ZN(n20419) );
  OR2_X1 U12986 ( .A1(n20286), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n20303) );
  NOR2_X1 U12987 ( .A1(n20059), .A2(n20055), .ZN(n20062) );
  NOR3_X1 U12988 ( .A1(n20419), .A2(n20871), .A3(n20215), .ZN(n20253) );
  INV_X1 U12989 ( .A(n20419), .ZN(n20404) );
  INV_X1 U12990 ( .A(n20487), .ZN(n20472) );
  NOR2_X2 U12991 ( .A1(n21208), .A2(n20407), .ZN(n20432) );
  AND2_X1 U12992 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17502), .ZN(n17478) );
  INV_X1 U12993 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20146) );
  NOR3_X1 U12994 ( .A1(n20592), .A2(n20640), .A3(n20568), .ZN(n20586) );
  NOR2_X1 U12995 ( .A1(n20051), .A2(n20046), .ZN(n20043) );
  INV_X1 U12996 ( .A(n17846), .ZN(n20859) );
  AOI21_X2 U12997 ( .B1(n20004), .B2(n20057), .A(n21224), .ZN(n18195) );
  INV_X1 U12998 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18104) );
  INV_X1 U12999 ( .A(n21090), .ZN(n21184) );
  INV_X1 U13000 ( .A(n21118), .ZN(n21049) );
  NAND2_X1 U13001 ( .A1(n20057), .A2(n18693), .ZN(n19011) );
  INV_X1 U13002 ( .A(n18908), .ZN(n19094) );
  INV_X1 U13003 ( .A(n19078), .ZN(n19086) );
  INV_X1 U13004 ( .A(n19067), .ZN(n19081) );
  INV_X1 U13005 ( .A(n19050), .ZN(n19063) );
  INV_X1 U13006 ( .A(n19044), .ZN(n19058) );
  INV_X1 U13007 ( .A(n18923), .ZN(n18914) );
  INV_X1 U13008 ( .A(n18957), .ZN(n18959) );
  NOR2_X1 U13009 ( .A1(n20685), .A2(n21075), .ZN(n17662) );
  INV_X1 U13010 ( .A(n18324), .ZN(n18322) );
  NOR2_X1 U13011 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13608), .ZN(n18690)
         );
  INV_X1 U13012 ( .A(n13660), .ZN(n13664) );
  INV_X1 U13013 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21829) );
  INV_X1 U13014 ( .A(n21517), .ZN(n21544) );
  INV_X1 U13015 ( .A(n21490), .ZN(n21535) );
  INV_X1 U13016 ( .A(n21525), .ZN(n21537) );
  AND2_X1 U13017 ( .A1(n21537), .A2(n14361), .ZN(n14519) );
  NAND2_X1 U13018 ( .A1(n19870), .A2(n14164), .ZN(n15796) );
  OR2_X1 U13019 ( .A1(n12409), .A2(n21663), .ZN(n21657) );
  INV_X1 U13020 ( .A(n14908), .ZN(n14560) );
  AND2_X1 U13021 ( .A1(n13864), .A2(n13863), .ZN(n21900) );
  NAND2_X1 U13022 ( .A1(n19767), .A2(n11645), .ZN(n14578) );
  INV_X1 U13023 ( .A(n19767), .ZN(n19794) );
  INV_X1 U13024 ( .A(n13922), .ZN(n13938) );
  INV_X1 U13025 ( .A(n19927), .ZN(n19952) );
  OAI21_X1 U13026 ( .B1(n15022), .B2(n14940), .A(n14939), .ZN(n15975) );
  INV_X1 U13027 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19877) );
  INV_X1 U13028 ( .A(n21409), .ZN(n21389) );
  INV_X1 U13029 ( .A(n21411), .ZN(n21335) );
  INV_X1 U13030 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21825) );
  INV_X1 U13031 ( .A(n16984), .ZN(n16982) );
  AOI22_X1 U13032 ( .A1(n21673), .A2(n21670), .B1(n21775), .B2(n21714), .ZN(
        n22140) );
  NAND2_X1 U13033 ( .A1(n21702), .A2(n21816), .ZN(n22149) );
  AOI22_X1 U13034 ( .A1(n21693), .A2(n21695), .B1(n11525), .B2(n21775), .ZN(
        n22154) );
  INV_X1 U13035 ( .A(n21705), .ZN(n22160) );
  NAND2_X1 U13036 ( .A1(n21742), .A2(n21793), .ZN(n22172) );
  AOI22_X1 U13037 ( .A1(n21737), .A2(n21734), .B1(n21799), .B2(n11525), .ZN(
        n22178) );
  NAND2_X1 U13038 ( .A1(n21742), .A2(n21741), .ZN(n22185) );
  NAND2_X1 U13039 ( .A1(n21770), .A2(n21793), .ZN(n22197) );
  AOI22_X1 U13040 ( .A1(n21778), .A2(n21776), .B1(n21775), .B2(n21774), .ZN(
        n22204) );
  NAND2_X1 U13041 ( .A1(n21770), .A2(n21821), .ZN(n22210) );
  INV_X1 U13042 ( .A(n21895), .ZN(n21887) );
  INV_X1 U13043 ( .A(n22123), .ZN(n22115) );
  NAND2_X1 U13044 ( .A1(n21822), .A2(n21793), .ZN(n22224) );
  NAND2_X1 U13045 ( .A1(n21822), .A2(n21821), .ZN(n22242) );
  INV_X1 U13046 ( .A(n21564), .ZN(n21566) );
  OR2_X1 U13047 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n13777), .ZN(n21587) );
  INV_X1 U13048 ( .A(n19836), .ZN(n19834) );
  NOR2_X1 U13049 ( .A1(n13612), .A2(n14337), .ZN(n18341) );
  INV_X1 U13050 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21569) );
  NAND2_X1 U13051 ( .A1(n15511), .A2(n15510), .ZN(n18577) );
  OR3_X1 U13052 ( .A1(n14641), .A2(n16247), .A3(n14638), .ZN(n18509) );
  NAND2_X1 U13053 ( .A1(n14017), .A2(n13956), .ZN(n17309) );
  NOR2_X1 U13054 ( .A1(n19586), .A2(n19585), .ZN(n19348) );
  NAND2_X1 U13055 ( .A1(n19496), .A2(n13974), .ZN(n19342) );
  NAND2_X1 U13056 ( .A1(n17337), .A2(n12525), .ZN(n14154) );
  INV_X1 U13057 ( .A(n17337), .ZN(n17371) );
  OAI21_X1 U13058 ( .B1(n13616), .B2(n21594), .A(n14633), .ZN(n13631) );
  NAND2_X1 U13059 ( .A1(n14635), .A2(n15436), .ZN(n14633) );
  NAND2_X1 U13060 ( .A1(n13468), .A2(n17274), .ZN(n13469) );
  OR2_X1 U13061 ( .A1(n18664), .A2(n18335), .ZN(n17294) );
  OR2_X1 U13062 ( .A1(n18664), .A2(n15436), .ZN(n17295) );
  INV_X1 U13063 ( .A(n17260), .ZN(n17301) );
  OR2_X1 U13064 ( .A1(n13423), .A2(n13082), .ZN(n18608) );
  OR2_X1 U13065 ( .A1(n13423), .A2(n14325), .ZN(n18614) );
  AND2_X1 U13066 ( .A1(n18615), .A2(n16755), .ZN(n18593) );
  INV_X1 U13067 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15371) );
  AOI21_X1 U13068 ( .B1(n14884), .B2(n14885), .A(n19591), .ZN(n19709) );
  NAND2_X1 U13069 ( .A1(n19257), .A2(n19256), .ZN(n19696) );
  INV_X1 U13070 ( .A(n19686), .ZN(n19683) );
  NAND2_X1 U13071 ( .A1(n19257), .A2(n19223), .ZN(n19676) );
  OR2_X1 U13072 ( .A1(n17321), .A2(n14605), .ZN(n19669) );
  INV_X1 U13073 ( .A(n19666), .ZN(n19524) );
  AOI22_X1 U13074 ( .A1(n14740), .A2(n14739), .B1(n14738), .B2(n14737), .ZN(
        n19663) );
  NAND2_X1 U13075 ( .A1(n19196), .A2(n19195), .ZN(n19655) );
  NAND2_X1 U13076 ( .A1(n19184), .A2(n19183), .ZN(n19649) );
  NAND2_X1 U13077 ( .A1(n19184), .A2(n19256), .ZN(n19641) );
  NAND2_X1 U13078 ( .A1(n19184), .A2(n19242), .ZN(n19628) );
  AOI22_X1 U13079 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19597), .ZN(n19531) );
  INV_X1 U13080 ( .A(n19625), .ZN(n19621) );
  AOI22_X1 U13081 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19597), .ZN(n19690) );
  AOI22_X1 U13082 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19597), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19598), .ZN(n19435) );
  AOI22_X1 U13083 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19597), .ZN(n19572) );
  NAND2_X1 U13084 ( .A1(n19120), .A2(n19223), .ZN(n19602) );
  INV_X1 U13085 ( .A(n21572), .ZN(n16999) );
  AOI21_X1 U13086 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n16996), .A(n17382), 
        .ZN(n21604) );
  OR2_X1 U13087 ( .A1(n16997), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n17390) );
  INV_X1 U13088 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21574) );
  INV_X1 U13089 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20417) );
  INV_X1 U13090 ( .A(n20432), .ZN(n20484) );
  INV_X1 U13091 ( .A(n17564), .ZN(n17577) );
  INV_X1 U13092 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17414) );
  INV_X1 U13093 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17739) );
  INV_X1 U13094 ( .A(n20658), .ZN(n20663) );
  AND3_X1 U13095 ( .A1(n17710), .A2(n17709), .A3(n17708), .ZN(n20550) );
  INV_X1 U13096 ( .A(n20667), .ZN(n20676) );
  NAND2_X1 U13097 ( .A1(n18279), .A2(n20495), .ZN(n18304) );
  INV_X1 U13098 ( .A(n18279), .ZN(n18278) );
  INV_X1 U13099 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20664) );
  INV_X1 U13100 ( .A(n20051), .ZN(n20048) );
  INV_X1 U13101 ( .A(n20046), .ZN(n20053) );
  INV_X1 U13102 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21109) );
  INV_X1 U13103 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21149) );
  INV_X1 U13104 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n20924) );
  INV_X1 U13105 ( .A(n21136), .ZN(n21092) );
  NAND2_X1 U13106 ( .A1(n21129), .A2(n21092), .ZN(n21118) );
  INV_X1 U13107 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21174) );
  OAI211_X1 U13108 ( .C1(n21195), .C2(n21218), .A(n15271), .B(n16978), .ZN(
        n20730) );
  INV_X1 U13109 ( .A(n19104), .ZN(n19091) );
  INV_X1 U13110 ( .A(n19074), .ZN(n18989) );
  INV_X1 U13111 ( .A(n19052), .ZN(n18980) );
  INV_X1 U13112 ( .A(n19003), .ZN(n19001) );
  NAND2_X1 U13113 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21201), .ZN(n21218) );
  INV_X1 U13114 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21208) );
  INV_X1 U13115 ( .A(n16987), .ZN(n21577) );
  INV_X1 U13116 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20122) );
  INV_X1 U13117 ( .A(n21662), .ZN(n21663) );
  AND2_X2 U13118 ( .A1(n11538), .A2(n13840), .ZN(n11757) );
  AND2_X2 U13119 ( .A1(n11538), .A2(n13958), .ZN(n11680) );
  AOI22_X1 U13120 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11680), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U13121 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U13122 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U13123 ( .A1(n11687), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U13124 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11549) );
  AOI22_X1 U13125 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U13126 ( .A1(n11603), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U13127 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11545) );
  NOR2_X1 U13128 ( .A1(n11541), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11542) );
  AOI22_X1 U13129 ( .A1(n11686), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U13130 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  AOI22_X1 U13131 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11603), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U13132 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U13133 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11687), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11552) );
  BUF_X1 U13134 ( .A(n11708), .Z(n11550) );
  AOI22_X1 U13135 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11551) );
  NAND4_X1 U13136 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(
        n11560) );
  AOI22_X1 U13137 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U13138 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11686), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U13139 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U13140 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11555) );
  NAND4_X1 U13141 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11559) );
  AOI22_X1 U13142 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U13143 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U13144 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11687), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U13145 ( .A1(n11686), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11561) );
  NAND4_X1 U13146 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11570) );
  AOI22_X1 U13147 ( .A1(n11603), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U13148 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U13149 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U13150 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11565) );
  NAND4_X1 U13151 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11569) );
  AOI22_X1 U13152 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11603), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U13153 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U13154 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11687), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U13155 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11571) );
  NAND4_X1 U13156 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11580) );
  AOI22_X1 U13157 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U13158 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11686), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U13159 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U13160 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U13161 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11579) );
  AOI22_X1 U13162 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U13163 ( .A1(n11603), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11687), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U13164 ( .A1(n11686), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U13165 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U13166 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AOI22_X1 U13167 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U13168 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U13169 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13170 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U13171 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  AOI22_X1 U13172 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13173 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U13174 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11687), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U13175 ( .A1(n11758), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U13176 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11602) );
  AOI22_X1 U13177 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11603), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U13178 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U13179 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10995), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U13180 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U13181 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11601) );
  OR2_X2 U13182 ( .A1(n11602), .A2(n11601), .ZN(n11630) );
  AOI22_X1 U13183 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11603), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U13184 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13185 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11687), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U13186 ( .A1(n11680), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U13187 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U13188 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11686), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U13189 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U13190 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11591), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11608) );
  NAND2_X2 U13191 ( .A1(n11028), .A2(n11529), .ZN(n11645) );
  AND2_X2 U13192 ( .A1(n14115), .A2(n11645), .ZN(n15545) );
  NAND2_X1 U13193 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U13194 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11613) );
  NAND2_X1 U13195 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U13196 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U13197 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11616) );
  NAND2_X1 U13198 ( .A1(n11686), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U13199 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U13200 ( .A1(n11603), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U13201 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U13202 ( .A1(n11758), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11619) );
  NAND2_X1 U13203 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11625) );
  NAND2_X1 U13204 ( .A1(n11687), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11624) );
  NAND2_X1 U13205 ( .A1(n11591), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11623) );
  NAND2_X1 U13206 ( .A1(n21585), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21580) );
  INV_X1 U13207 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11627) );
  NAND2_X1 U13208 ( .A1(n11627), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U13209 ( .A1(n21859), .A2(n13777), .ZN(n11629) );
  AOI21_X1 U13210 ( .B1(n15545), .B2(n11629), .A(n14113), .ZN(n11638) );
  NAND2_X1 U13211 ( .A1(n11642), .A2(n21991), .ZN(n11639) );
  INV_X1 U13212 ( .A(n13472), .ZN(n11643) );
  NAND2_X1 U13213 ( .A1(n11643), .A2(n14164), .ZN(n11631) );
  NAND2_X1 U13214 ( .A1(n11630), .A2(n22037), .ZN(n11634) );
  NAND2_X1 U13216 ( .A1(n13628), .A2(n21859), .ZN(n12382) );
  INV_X1 U13217 ( .A(n11639), .ZN(n11640) );
  NAND2_X1 U13218 ( .A1(n12343), .A2(n11630), .ZN(n11641) );
  INV_X1 U13219 ( .A(n11642), .ZN(n14165) );
  NAND2_X1 U13220 ( .A1(n16089), .A2(n13788), .ZN(n11647) );
  INV_X1 U13221 ( .A(n12335), .ZN(n13806) );
  NAND2_X1 U13222 ( .A1(n11643), .A2(n13806), .ZN(n11644) );
  NAND2_X1 U13223 ( .A1(n11644), .A2(n14164), .ZN(n11646) );
  NAND2_X1 U13224 ( .A1(n12335), .A2(n15588), .ZN(n14108) );
  NAND2_X1 U13225 ( .A1(n21667), .A2(n14364), .ZN(n13805) );
  NAND2_X1 U13226 ( .A1(n11653), .A2(n21667), .ZN(n11649) );
  NAND3_X1 U13227 ( .A1(n11650), .A2(n11649), .A3(n13488), .ZN(n11651) );
  NAND2_X1 U13228 ( .A1(n16094), .A2(n11213), .ZN(n13480) );
  MUX2_X1 U13229 ( .A(n13480), .B(n12394), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11652) );
  INV_X1 U13230 ( .A(n16089), .ZN(n17020) );
  NAND2_X1 U13231 ( .A1(n13788), .A2(n14364), .ZN(n11664) );
  AND2_X1 U13232 ( .A1(n12392), .A2(n15607), .ZN(n13659) );
  NAND2_X1 U13233 ( .A1(n14165), .A2(n21946), .ZN(n11654) );
  NAND2_X1 U13234 ( .A1(n13659), .A2(n11654), .ZN(n11662) );
  INV_X1 U13235 ( .A(n11655), .ZN(n11660) );
  NAND2_X1 U13236 ( .A1(n13839), .A2(n11656), .ZN(n14106) );
  NAND2_X1 U13237 ( .A1(n16094), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11657) );
  AOI21_X1 U13238 ( .B1(n14093), .B2(n11645), .A(n11657), .ZN(n11658) );
  AOI22_X1 U13239 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11671) );
  BUF_X1 U13240 ( .A(n11752), .Z(n11666) );
  AOI22_X1 U13241 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U13242 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11686), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11669) );
  BUF_X1 U13243 ( .A(n11758), .Z(n11667) );
  AOI22_X1 U13244 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11668) );
  NAND4_X1 U13245 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n11679) );
  AOI22_X1 U13246 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11677) );
  BUF_X1 U13247 ( .A(n11772), .Z(n11672) );
  AOI22_X1 U13248 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11676) );
  INV_X1 U13249 ( .A(n11681), .ZN(n13838) );
  AOI22_X1 U13250 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11675) );
  BUF_X1 U13251 ( .A(n11708), .Z(n11673) );
  AOI22_X1 U13252 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11674) );
  NAND4_X1 U13253 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11678) );
  AOI22_X1 U13254 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n12303), .B1(
        n12304), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11685) );
  INV_X2 U13255 ( .A(n13838), .ZN(n12271) );
  AOI22_X1 U13256 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12271), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U13257 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U13258 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U13259 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11693) );
  AOI22_X1 U13260 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12295), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U13261 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U13262 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11686), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U13263 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12302), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11688) );
  NAND4_X1 U13264 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11692) );
  NAND2_X1 U13265 ( .A1(n13548), .A2(n13486), .ZN(n11696) );
  INV_X1 U13266 ( .A(n11751), .ZN(n11733) );
  INV_X1 U13267 ( .A(n13551), .ZN(n11694) );
  NAND3_X1 U13268 ( .A1(n11733), .A2(n11694), .A3(n13498), .ZN(n11695) );
  INV_X1 U13269 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11701) );
  AOI21_X1 U13270 ( .B1(n21667), .B2(n13498), .A(n11213), .ZN(n11700) );
  INV_X1 U13271 ( .A(n13548), .ZN(n11699) );
  OAI211_X1 U13272 ( .C1(n12366), .C2(n11701), .A(n11700), .B(n11699), .ZN(
        n11842) );
  INV_X1 U13273 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11718) );
  INV_X1 U13274 ( .A(n11750), .ZN(n11716) );
  AOI22_X1 U13275 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U13276 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U13277 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11686), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U13278 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11703) );
  NAND4_X1 U13279 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11715) );
  AOI22_X1 U13280 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U13281 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U13282 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U13283 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U13284 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11714) );
  NAND2_X1 U13285 ( .A1(n11716), .A2(n13497), .ZN(n11717) );
  OAI211_X1 U13286 ( .C1(n12366), .C2(n11718), .A(n11717), .B(n11751), .ZN(
        n11719) );
  INV_X1 U13287 ( .A(n11719), .ZN(n11720) );
  NAND2_X1 U13288 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11743) );
  OAI21_X1 U13289 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11743), .ZN(n21773) );
  NAND2_X1 U13290 ( .A1(n17053), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11736) );
  OAI21_X1 U13291 ( .B1(n13480), .B2(n21773), .A(n11736), .ZN(n11721) );
  INV_X1 U13292 ( .A(n11721), .ZN(n11722) );
  INV_X1 U13293 ( .A(n11724), .ZN(n11725) );
  AND2_X2 U13294 ( .A1(n11725), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11735) );
  XNOR2_X1 U13295 ( .A(n11726), .B(n11735), .ZN(n11729) );
  NAND2_X1 U13296 ( .A1(n11728), .A2(n11727), .ZN(n11730) );
  INV_X1 U13297 ( .A(n11729), .ZN(n11732) );
  INV_X1 U13298 ( .A(n11730), .ZN(n11731) );
  NAND2_X1 U13299 ( .A1(n11733), .A2(n13497), .ZN(n11734) );
  INV_X1 U13300 ( .A(n11735), .ZN(n11738) );
  AND2_X1 U13301 ( .A1(n11736), .A2(n16093), .ZN(n11737) );
  NAND2_X1 U13302 ( .A1(n11741), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11746) );
  INV_X1 U13303 ( .A(n11743), .ZN(n11742) );
  NAND2_X1 U13304 ( .A1(n11742), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21743) );
  NAND2_X1 U13305 ( .A1(n11743), .A2(n21824), .ZN(n11744) );
  INV_X1 U13306 ( .A(n13480), .ZN(n11769) );
  AOI22_X1 U13307 ( .A1(n21668), .A2(n11769), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17053), .ZN(n11745) );
  OR2_X2 U13308 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  NAND2_X2 U13309 ( .A1(n11748), .A2(n11747), .ZN(n14442) );
  AOI22_X1 U13310 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U13311 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U13312 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U13313 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11753) );
  NAND4_X1 U13314 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11764) );
  AOI22_X1 U13315 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U13316 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U13317 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U13318 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11759) );
  NAND4_X1 U13319 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11763) );
  AOI22_X1 U13320 ( .A1(n12379), .A2(n13496), .B1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12345), .ZN(n11765) );
  INV_X1 U13321 ( .A(n11857), .ZN(n11785) );
  NAND2_X1 U13322 ( .A1(n11741), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11771) );
  INV_X1 U13323 ( .A(n21743), .ZN(n11767) );
  NAND2_X1 U13324 ( .A1(n11767), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21841) );
  NAND2_X1 U13325 ( .A1(n21743), .A2(n21825), .ZN(n11768) );
  AOI22_X1 U13326 ( .A1(n21754), .A2(n11769), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17053), .ZN(n11770) );
  AOI22_X1 U13327 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U13328 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U13329 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U13330 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11773) );
  NAND4_X1 U13331 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11782) );
  AOI22_X1 U13332 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U13333 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U13334 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U13335 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11777) );
  NAND4_X1 U13336 ( .A1(n11780), .A2(n11779), .A3(n11778), .A4(n11777), .ZN(
        n11781) );
  AOI22_X1 U13337 ( .A1(n12379), .A2(n13515), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12345), .ZN(n11783) );
  AOI22_X1 U13338 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U13339 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U13340 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U13341 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U13342 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11795) );
  AOI22_X1 U13343 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U13344 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U13345 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U13346 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11790) );
  NAND4_X1 U13347 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11794) );
  NAND2_X1 U13348 ( .A1(n12379), .A2(n13523), .ZN(n11797) );
  NAND2_X1 U13349 ( .A1(n12345), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U13350 ( .A1(n11797), .A2(n11796), .ZN(n11867) );
  AOI22_X1 U13351 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13352 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U13353 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U13354 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11798) );
  NAND4_X1 U13355 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11807) );
  AOI22_X1 U13356 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U13357 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U13358 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U13359 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11802) );
  NAND4_X1 U13360 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11806) );
  NAND2_X1 U13361 ( .A1(n12379), .A2(n13532), .ZN(n11809) );
  NAND2_X1 U13362 ( .A1(n12345), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U13363 ( .A1(n11809), .A2(n11808), .ZN(n11878) );
  NAND2_X1 U13364 ( .A1(n11810), .A2(n11878), .ZN(n11887) );
  AOI22_X1 U13365 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U13366 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U13367 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U13368 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11811) );
  NAND4_X1 U13369 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11820) );
  AOI22_X1 U13370 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U13371 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U13372 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U13373 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11815) );
  NAND4_X1 U13374 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11819) );
  AOI22_X1 U13375 ( .A1(n12379), .A2(n13535), .B1(n12345), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11886) );
  NAND2_X1 U13376 ( .A1(n12379), .A2(n13551), .ZN(n11822) );
  NAND2_X1 U13377 ( .A1(n12345), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U13378 ( .A1(n11822), .A2(n11821), .ZN(n11823) );
  INV_X1 U13379 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11828) );
  NAND2_X1 U13380 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11859) );
  INV_X1 U13381 ( .A(n11859), .ZN(n11824) );
  NOR2_X1 U13382 ( .A1(n11890), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11825) );
  OR2_X1 U13383 ( .A1(n11908), .A2(n11825), .ZN(n21435) );
  NAND2_X1 U13384 ( .A1(n21435), .A2(n12323), .ZN(n11827) );
  NAND2_X1 U13385 ( .A1(n12326), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11826) );
  OAI211_X1 U13386 ( .C1(n12317), .C2(n11828), .A(n11827), .B(n11826), .ZN(
        n11829) );
  AOI21_X1 U13387 ( .B1(n13542), .B2(n11994), .A(n11829), .ZN(n14432) );
  AND2_X1 U13388 ( .A1(n12397), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11869) );
  XNOR2_X1 U13389 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14404) );
  AOI21_X1 U13390 ( .B1(n12323), .B2(n14404), .A(n12326), .ZN(n11830) );
  OAI21_X1 U13391 ( .B1(n12317), .B2(n19771), .A(n11830), .ZN(n11831) );
  AOI21_X1 U13392 ( .B1(n11869), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11831), .ZN(n11832) );
  NAND2_X1 U13393 ( .A1(n12326), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U13394 ( .A1(n11833), .A2(n11855), .ZN(n14048) );
  INV_X1 U13395 ( .A(n11834), .ZN(n11835) );
  NAND2_X1 U13396 ( .A1(n11835), .A2(n11188), .ZN(n11837) );
  INV_X1 U13397 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11838) );
  INV_X1 U13398 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14390) );
  OAI22_X1 U13399 ( .A1(n12317), .A2(n11838), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14390), .ZN(n11839) );
  AOI21_X1 U13400 ( .B1(n11869), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11839), .ZN(n11840) );
  INV_X1 U13401 ( .A(n11841), .ZN(n11844) );
  INV_X1 U13402 ( .A(n11842), .ZN(n11843) );
  NAND2_X1 U13403 ( .A1(n11844), .A2(n11843), .ZN(n11846) );
  INV_X1 U13404 ( .A(n21699), .ZN(n16086) );
  NAND2_X1 U13405 ( .A1(n16086), .A2(n11994), .ZN(n11851) );
  INV_X1 U13406 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n11848) );
  INV_X1 U13407 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14517) );
  OAI22_X1 U13408 ( .A1(n12317), .A2(n11848), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14517), .ZN(n11849) );
  AOI21_X1 U13409 ( .B1(n11869), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11849), .ZN(n11850) );
  NAND2_X1 U13410 ( .A1(n11851), .A2(n11850), .ZN(n14004) );
  NAND2_X1 U13411 ( .A1(n14005), .A2(n14004), .ZN(n14003) );
  OR2_X1 U13412 ( .A1(n14004), .A2(n12315), .ZN(n11852) );
  NAND2_X1 U13413 ( .A1(n14003), .A2(n11852), .ZN(n13872) );
  NAND2_X1 U13414 ( .A1(n13871), .A2(n13872), .ZN(n14047) );
  INV_X1 U13415 ( .A(n14047), .ZN(n11853) );
  NAND2_X1 U13416 ( .A1(n11854), .A2(n11853), .ZN(n14045) );
  NAND2_X1 U13417 ( .A1(n14066), .A2(n11857), .ZN(n11858) );
  INV_X1 U13418 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11864) );
  INV_X1 U13419 ( .A(n11874), .ZN(n11862) );
  INV_X1 U13420 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U13421 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  NAND2_X1 U13422 ( .A1(n11862), .A2(n11861), .ZN(n14381) );
  AOI22_X1 U13423 ( .A1(n14381), .A2(n12323), .B1(n12326), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11863) );
  OAI21_X1 U13424 ( .B1(n12317), .B2(n11864), .A(n11863), .ZN(n11865) );
  AOI21_X1 U13425 ( .B1(n11869), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11865), .ZN(n11866) );
  OAI21_X1 U13426 ( .B1(n13508), .B2(n11432), .A(n11866), .ZN(n14169) );
  XNOR2_X1 U13427 ( .A(n11868), .B(n11867), .ZN(n13514) );
  INV_X1 U13428 ( .A(n11869), .ZN(n11872) );
  INV_X1 U13429 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U13430 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11871) );
  NAND2_X1 U13431 ( .A1(n12327), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11870) );
  OAI211_X1 U13432 ( .C1(n11872), .C2(n14443), .A(n11871), .B(n11870), .ZN(
        n11873) );
  NAND2_X1 U13433 ( .A1(n11873), .A2(n12315), .ZN(n11876) );
  OAI21_X1 U13434 ( .B1(n11874), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11880), .ZN(n14451) );
  NAND2_X1 U13435 ( .A1(n14451), .A2(n12323), .ZN(n11875) );
  NAND2_X1 U13436 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  AOI21_X1 U13437 ( .B1(n13514), .B2(n11994), .A(n11877), .ZN(n14183) );
  XNOR2_X1 U13438 ( .A(n11879), .B(n11878), .ZN(n13522) );
  NAND2_X1 U13439 ( .A1(n13522), .A2(n11994), .ZN(n11885) );
  INV_X1 U13440 ( .A(n12326), .ZN(n12046) );
  AND2_X1 U13441 ( .A1(n11880), .A2(n19877), .ZN(n11881) );
  OR2_X1 U13442 ( .A1(n11881), .A2(n11888), .ZN(n19873) );
  NAND2_X1 U13443 ( .A1(n19873), .A2(n12323), .ZN(n11882) );
  OAI21_X1 U13444 ( .B1(n19877), .B2(n12046), .A(n11882), .ZN(n11883) );
  AOI21_X1 U13445 ( .B1(n12327), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11883), .ZN(
        n11884) );
  NAND2_X1 U13446 ( .A1(n11885), .A2(n11884), .ZN(n14192) );
  NAND2_X1 U13447 ( .A1(n11887), .A2(n11886), .ZN(n13531) );
  INV_X1 U13448 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19778) );
  NOR2_X1 U13449 ( .A1(n11888), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11889) );
  OR2_X1 U13450 ( .A1(n11890), .A2(n11889), .ZN(n21432) );
  AOI22_X1 U13451 ( .A1(n21432), .A2(n12323), .B1(n12326), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11891) );
  OAI21_X1 U13452 ( .B1(n12317), .B2(n19778), .A(n11891), .ZN(n11892) );
  NAND2_X1 U13453 ( .A1(n11893), .A2(n14232), .ZN(n14431) );
  INV_X1 U13454 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14502) );
  INV_X1 U13455 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14873) );
  OAI22_X1 U13456 ( .A1(n12317), .A2(n14502), .B1(n12046), .B2(n14873), .ZN(
        n11894) );
  INV_X1 U13457 ( .A(n11894), .ZN(n11907) );
  XNOR2_X1 U13458 ( .A(n11908), .B(n14873), .ZN(n14875) );
  OR2_X1 U13459 ( .A1(n14875), .A2(n12315), .ZN(n11906) );
  AOI22_X1 U13460 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U13461 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U13462 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U13463 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11895) );
  NAND4_X1 U13464 ( .A1(n11898), .A2(n11897), .A3(n11896), .A4(n11895), .ZN(
        n11904) );
  AOI22_X1 U13465 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12303), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U13466 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U13467 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U13468 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11899) );
  NAND4_X1 U13469 ( .A1(n11902), .A2(n11901), .A3(n11900), .A4(n11899), .ZN(
        n11903) );
  OAI21_X1 U13470 ( .B1(n11904), .B2(n11903), .A(n11994), .ZN(n11905) );
  XOR2_X1 U13471 ( .A(n14552), .B(n11922), .Z(n14904) );
  AOI22_X1 U13472 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U13473 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U13474 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U13475 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11909) );
  NAND4_X1 U13476 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11918) );
  AOI22_X1 U13477 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U13478 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U13479 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U13480 ( .A1(n11673), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U13481 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11917) );
  OR2_X1 U13482 ( .A1(n11918), .A2(n11917), .ZN(n11919) );
  AOI22_X1 U13483 ( .A1(n11994), .A2(n11919), .B1(n12326), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11921) );
  NAND2_X1 U13484 ( .A1(n12327), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11920) );
  OAI211_X1 U13485 ( .C1(n14904), .C2(n12315), .A(n11921), .B(n11920), .ZN(
        n14539) );
  NAND2_X1 U13486 ( .A1(n14482), .A2(n14539), .ZN(n14538) );
  XNOR2_X1 U13487 ( .A(n11937), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19889) );
  AOI22_X1 U13488 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U13489 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U13490 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U13491 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U13492 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11932) );
  AOI22_X1 U13493 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U13494 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U13495 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U13496 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U13497 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  NOR2_X1 U13498 ( .A1(n11932), .A2(n11931), .ZN(n11935) );
  NAND2_X1 U13499 ( .A1(n12327), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U13500 ( .A1(n12326), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11933) );
  OAI211_X1 U13501 ( .C1(n11432), .C2(n11935), .A(n11934), .B(n11933), .ZN(
        n11936) );
  AOI21_X1 U13502 ( .B1(n19889), .B2(n12323), .A(n11936), .ZN(n14661) );
  OAI21_X1 U13503 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11938), .A(
        n11977), .ZN(n21446) );
  AOI22_X1 U13504 ( .A1(n12323), .A2(n21446), .B1(n12326), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11939) );
  OAI21_X1 U13505 ( .B1(n12317), .B2(n19788), .A(n11939), .ZN(n14934) );
  AOI22_X1 U13506 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U13507 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U13508 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U13509 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U13510 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11949) );
  AOI22_X1 U13511 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U13512 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U13513 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U13514 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11944) );
  NAND4_X1 U13515 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11948) );
  OR2_X1 U13516 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  NAND2_X1 U13517 ( .A1(n11994), .A2(n11950), .ZN(n14962) );
  INV_X1 U13518 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U13519 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U13520 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U13521 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U13522 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U13523 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11960) );
  AOI22_X1 U13524 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13525 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13526 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U13527 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11955) );
  NAND4_X1 U13528 ( .A1(n11958), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11959) );
  OR2_X1 U13529 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  NAND2_X1 U13530 ( .A1(n11994), .A2(n11961), .ZN(n11965) );
  XNOR2_X1 U13531 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11977), .ZN(
        n21457) );
  INV_X1 U13532 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11962) );
  OAI22_X1 U13533 ( .A1(n21457), .A2(n12315), .B1(n12046), .B2(n11962), .ZN(
        n11963) );
  INV_X1 U13534 ( .A(n11963), .ZN(n11964) );
  OAI211_X1 U13535 ( .C1(n12317), .C2(n15026), .A(n11965), .B(n11964), .ZN(
        n15021) );
  INV_X1 U13536 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15001) );
  AOI22_X1 U13537 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U13538 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13539 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U13540 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11966) );
  NAND4_X1 U13541 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11975) );
  AOI22_X1 U13542 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U13543 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U13544 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U13545 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11970) );
  NAND4_X1 U13546 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n11974) );
  OR2_X1 U13547 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  NAND2_X1 U13548 ( .A1(n11994), .A2(n11976), .ZN(n11981) );
  INV_X1 U13549 ( .A(n11982), .ZN(n11979) );
  XNOR2_X1 U13550 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11979), .ZN(
        n14941) );
  AOI22_X1 U13551 ( .A1(n12323), .A2(n14941), .B1(n12326), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11980) );
  OAI211_X1 U13552 ( .C1(n12317), .C2(n15001), .A(n11981), .B(n11980), .ZN(
        n14940) );
  XOR2_X1 U13553 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11997), .Z(
        n21467) );
  AOI22_X1 U13554 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U13555 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U13556 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U13557 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11983) );
  NAND4_X1 U13558 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n11992) );
  AOI22_X1 U13559 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U13560 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U13561 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U13562 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U13563 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11991) );
  OR2_X1 U13564 ( .A1(n11992), .A2(n11991), .ZN(n11993) );
  AOI22_X1 U13565 ( .A1(n11994), .A2(n11993), .B1(n12326), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U13566 ( .A1(n12327), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11995) );
  OAI211_X1 U13567 ( .C1(n21467), .C2(n12315), .A(n11996), .B(n11995), .ZN(
        n14988) );
  XNOR2_X1 U13568 ( .A(n12031), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21478) );
  INV_X1 U13569 ( .A(n21478), .ZN(n12012) );
  AOI22_X1 U13570 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U13571 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U13572 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U13573 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U13574 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12007) );
  AOI22_X1 U13575 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U13576 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U13577 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U13578 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U13579 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  NOR2_X1 U13580 ( .A1(n12007), .A2(n12006), .ZN(n12010) );
  NAND2_X1 U13581 ( .A1(n12327), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12009) );
  NAND2_X1 U13582 ( .A1(n12326), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12008) );
  OAI211_X1 U13583 ( .C1(n11432), .C2(n12010), .A(n12009), .B(n12008), .ZN(
        n12011) );
  AOI21_X1 U13584 ( .B1(n12012), .B2(n12323), .A(n12011), .ZN(n15033) );
  INV_X1 U13585 ( .A(n15033), .ZN(n12013) );
  AOI22_X1 U13586 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U13587 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12303), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U13588 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U13589 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U13590 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12024) );
  AOI22_X1 U13591 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12301), .B1(
        n12304), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U13592 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U13593 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U13594 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U13595 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n12023) );
  NOR2_X1 U13596 ( .A1(n12024), .A2(n12023), .ZN(n12029) );
  INV_X1 U13597 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U13598 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12025) );
  OAI211_X1 U13599 ( .C1(n12317), .C2(n12026), .A(n12315), .B(n12025), .ZN(
        n12027) );
  INV_X1 U13600 ( .A(n12027), .ZN(n12028) );
  OAI21_X1 U13601 ( .B1(n12320), .B2(n12029), .A(n12028), .ZN(n12034) );
  OAI21_X1 U13602 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12032), .A(
        n12064), .ZN(n21487) );
  OR2_X1 U13603 ( .A1(n12315), .A2(n21487), .ZN(n12033) );
  NAND2_X1 U13604 ( .A1(n12034), .A2(n12033), .ZN(n15787) );
  AOI22_X1 U13605 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U13606 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U13607 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U13608 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U13609 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12044) );
  AOI22_X1 U13610 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U13611 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U13612 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U13613 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U13614 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12043) );
  NOR2_X1 U13615 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  OR2_X1 U13616 ( .A1(n12320), .A2(n12045), .ZN(n12049) );
  XNOR2_X1 U13617 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12064), .ZN(
        n15959) );
  OAI22_X1 U13618 ( .A1(n15959), .A2(n12315), .B1(n12046), .B2(n15957), .ZN(
        n12047) );
  AOI21_X1 U13619 ( .B1(n12327), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12047), .ZN(
        n12048) );
  NAND2_X1 U13620 ( .A1(n12049), .A2(n12048), .ZN(n15725) );
  AOI22_X1 U13621 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U13622 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U13623 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13624 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12050) );
  NAND4_X1 U13625 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12059) );
  AOI22_X1 U13626 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U13627 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U13628 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U13629 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12054) );
  NAND4_X1 U13630 ( .A1(n12057), .A2(n12056), .A3(n12055), .A4(n12054), .ZN(
        n12058) );
  NOR2_X1 U13631 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  OR2_X1 U13632 ( .A1(n12320), .A2(n12060), .ZN(n12068) );
  INV_X1 U13633 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12062) );
  NAND2_X1 U13634 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12061) );
  OAI211_X1 U13635 ( .C1(n12317), .C2(n12062), .A(n12315), .B(n12061), .ZN(
        n12063) );
  INV_X1 U13636 ( .A(n12063), .ZN(n12067) );
  OAI21_X1 U13637 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12065), .A(
        n12098), .ZN(n21497) );
  NOR2_X1 U13638 ( .A1(n21497), .A2(n12315), .ZN(n12066) );
  AOI21_X1 U13639 ( .B1(n12068), .B2(n12067), .A(n12066), .ZN(n15774) );
  INV_X2 U13640 ( .A(n15777), .ZN(n12084) );
  AOI22_X1 U13641 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U13642 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U13643 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U13644 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12069) );
  NAND4_X1 U13645 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12078) );
  AOI22_X1 U13646 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U13647 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U13648 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U13649 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12073) );
  NAND4_X1 U13650 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12077) );
  NOR2_X1 U13651 ( .A1(n12078), .A2(n12077), .ZN(n12081) );
  OAI21_X1 U13652 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15944), .A(n12315), 
        .ZN(n12079) );
  AOI21_X1 U13653 ( .B1(n12327), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12079), .ZN(
        n12080) );
  OAI21_X1 U13654 ( .B1(n12320), .B2(n12081), .A(n12080), .ZN(n12083) );
  XNOR2_X1 U13655 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12098), .ZN(
        n15946) );
  NAND2_X1 U13656 ( .A1(n12323), .A2(n15946), .ZN(n12082) );
  AOI22_X1 U13657 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U13658 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U13659 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U13660 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U13661 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12094) );
  AOI22_X1 U13662 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U13663 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U13664 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U13665 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U13666 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12093) );
  NOR2_X1 U13667 ( .A1(n12094), .A2(n12093), .ZN(n12097) );
  OAI21_X1 U13668 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21829), .A(
        n11847), .ZN(n12096) );
  NAND2_X1 U13669 ( .A1(n12327), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n12095) );
  OAI211_X1 U13670 ( .C1(n12320), .C2(n12097), .A(n12096), .B(n12095), .ZN(
        n12101) );
  OAI21_X1 U13671 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12099), .A(
        n12130), .ZN(n21507) );
  OR2_X1 U13672 ( .A1(n12315), .A2(n21507), .ZN(n12100) );
  NAND2_X1 U13673 ( .A1(n12101), .A2(n12100), .ZN(n15763) );
  AOI22_X1 U13674 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U13675 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U13676 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U13677 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12102) );
  NAND4_X1 U13678 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12111) );
  AOI22_X1 U13679 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U13680 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U13681 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U13682 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12106) );
  NAND4_X1 U13683 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  NOR2_X1 U13684 ( .A1(n12111), .A2(n12110), .ZN(n12114) );
  OAI21_X1 U13685 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15936), .A(n12315), 
        .ZN(n12112) );
  AOI21_X1 U13686 ( .B1(n12327), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12112), .ZN(
        n12113) );
  OAI21_X1 U13687 ( .B1(n12320), .B2(n12114), .A(n12113), .ZN(n12116) );
  XNOR2_X1 U13688 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12130), .ZN(
        n15937) );
  NAND2_X1 U13689 ( .A1(n12323), .A2(n15937), .ZN(n12115) );
  AOI22_X1 U13690 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U13691 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U13692 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U13693 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U13694 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12126) );
  AOI22_X1 U13695 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U13696 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U13697 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U13698 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U13699 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  NOR2_X1 U13700 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  OR2_X1 U13701 ( .A1(n12320), .A2(n12127), .ZN(n12134) );
  INV_X1 U13702 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14573) );
  OAI21_X1 U13703 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21829), .A(
        n11847), .ZN(n12128) );
  OAI21_X1 U13704 ( .B1(n12317), .B2(n14573), .A(n12128), .ZN(n12129) );
  INV_X1 U13705 ( .A(n12129), .ZN(n12133) );
  OAI21_X1 U13706 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12131), .A(
        n12179), .ZN(n21520) );
  NOR2_X1 U13707 ( .A1(n21520), .A2(n12315), .ZN(n12132) );
  AOI21_X1 U13708 ( .B1(n12134), .B2(n12133), .A(n12132), .ZN(n15752) );
  AOI22_X1 U13709 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U13710 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U13711 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U13712 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U13713 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12145) );
  AOI22_X1 U13714 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U13715 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U13716 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U13717 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12140) );
  NAND4_X1 U13718 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n12144) );
  NOR2_X1 U13719 ( .A1(n12145), .A2(n12144), .ZN(n12163) );
  AOI22_X1 U13720 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U13721 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U13722 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U13723 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U13724 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12156) );
  AOI22_X1 U13725 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13726 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11666), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U13727 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U13728 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12302), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U13729 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12155) );
  NOR2_X1 U13730 ( .A1(n12156), .A2(n12155), .ZN(n12164) );
  XNOR2_X1 U13731 ( .A(n12163), .B(n12164), .ZN(n12159) );
  INV_X1 U13732 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21545) );
  OAI21_X1 U13733 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21545), .A(n12315), 
        .ZN(n12157) );
  AOI21_X1 U13734 ( .B1(n12327), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12157), .ZN(
        n12158) );
  OAI21_X1 U13735 ( .B1(n12320), .B2(n12159), .A(n12158), .ZN(n12161) );
  XNOR2_X1 U13736 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12179), .ZN(
        n21531) );
  NAND2_X1 U13737 ( .A1(n21531), .A2(n12323), .ZN(n12160) );
  NOR2_X1 U13738 ( .A1(n12164), .A2(n12163), .ZN(n12198) );
  AOI22_X1 U13739 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U13740 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U13741 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U13742 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12165) );
  NAND4_X1 U13743 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12174) );
  AOI22_X1 U13744 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U13745 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U13746 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U13747 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12169) );
  NAND4_X1 U13748 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12173) );
  INV_X1 U13749 ( .A(n12197), .ZN(n12175) );
  XNOR2_X1 U13750 ( .A(n12198), .B(n12175), .ZN(n12178) );
  INV_X1 U13751 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15836) );
  NAND2_X1 U13752 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12176) );
  OAI211_X1 U13753 ( .C1(n12317), .C2(n15836), .A(n12315), .B(n12176), .ZN(
        n12177) );
  AOI21_X1 U13754 ( .B1(n12178), .B2(n12286), .A(n12177), .ZN(n12186) );
  INV_X1 U13755 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12183) );
  INV_X1 U13756 ( .A(n12181), .ZN(n12182) );
  NAND2_X1 U13757 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  NAND2_X1 U13758 ( .A1(n12222), .A2(n12184), .ZN(n15924) );
  NOR2_X1 U13759 ( .A1(n15924), .A2(n12315), .ZN(n12185) );
  AOI22_X1 U13760 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12271), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U13761 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11667), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U13762 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U13763 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11673), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U13764 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12196) );
  AOI22_X1 U13765 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U13766 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U13767 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U13768 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12191) );
  NAND4_X1 U13769 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12195) );
  NOR2_X1 U13770 ( .A1(n12196), .A2(n12195), .ZN(n12207) );
  NAND2_X1 U13771 ( .A1(n12198), .A2(n12197), .ZN(n12206) );
  XOR2_X1 U13772 ( .A(n12207), .B(n12206), .Z(n12199) );
  NAND2_X1 U13773 ( .A1(n12199), .A2(n12286), .ZN(n12202) );
  AOI21_X1 U13774 ( .B1(n15915), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12200) );
  AOI21_X1 U13775 ( .B1(n12327), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12200), .ZN(
        n12201) );
  NAND2_X1 U13776 ( .A1(n12202), .A2(n12201), .ZN(n12204) );
  XNOR2_X1 U13777 ( .A(n12222), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15917) );
  NAND2_X1 U13778 ( .A1(n15917), .A2(n12323), .ZN(n12203) );
  NAND2_X1 U13779 ( .A1(n12204), .A2(n12203), .ZN(n15673) );
  INV_X1 U13780 ( .A(n15673), .ZN(n12205) );
  NOR2_X1 U13781 ( .A1(n12207), .A2(n12206), .ZN(n12240) );
  AOI22_X1 U13782 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U13783 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U13784 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U13785 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12208) );
  NAND4_X1 U13786 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12217) );
  AOI22_X1 U13787 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U13788 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U13789 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U13790 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12212) );
  NAND4_X1 U13791 ( .A1(n12215), .A2(n12214), .A3(n12213), .A4(n12212), .ZN(
        n12216) );
  OR2_X1 U13792 ( .A1(n12217), .A2(n12216), .ZN(n12239) );
  INV_X1 U13793 ( .A(n12239), .ZN(n12218) );
  XNOR2_X1 U13794 ( .A(n12240), .B(n12218), .ZN(n12219) );
  NAND2_X1 U13795 ( .A1(n12219), .A2(n12286), .ZN(n12228) );
  INV_X1 U13796 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15825) );
  NAND2_X1 U13797 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12220) );
  OAI211_X1 U13798 ( .C1(n12317), .C2(n15825), .A(n12315), .B(n12220), .ZN(
        n12221) );
  INV_X1 U13799 ( .A(n12221), .ZN(n12227) );
  INV_X1 U13800 ( .A(n12223), .ZN(n12224) );
  INV_X1 U13801 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15662) );
  NAND2_X1 U13802 ( .A1(n12224), .A2(n15662), .ZN(n12225) );
  NAND2_X1 U13803 ( .A1(n12263), .A2(n12225), .ZN(n15906) );
  NOR2_X1 U13804 ( .A1(n15906), .A2(n12315), .ZN(n12226) );
  AOI21_X1 U13805 ( .B1(n12228), .B2(n12227), .A(n12226), .ZN(n15659) );
  AOI22_X1 U13806 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U13807 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U13808 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U13809 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U13810 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12238) );
  AOI22_X1 U13811 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U13812 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U13813 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U13814 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12233) );
  NAND4_X1 U13815 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12237) );
  NOR2_X1 U13816 ( .A1(n12238), .A2(n12237), .ZN(n12248) );
  NAND2_X1 U13817 ( .A1(n12240), .A2(n12239), .ZN(n12247) );
  XOR2_X1 U13818 ( .A(n12248), .B(n12247), .Z(n12241) );
  NAND2_X1 U13819 ( .A1(n12241), .A2(n12286), .ZN(n12246) );
  INV_X1 U13820 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15819) );
  NAND2_X1 U13821 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12242) );
  OAI211_X1 U13822 ( .C1(n12317), .C2(n15819), .A(n12315), .B(n12242), .ZN(
        n12243) );
  INV_X1 U13823 ( .A(n12243), .ZN(n12245) );
  XNOR2_X1 U13824 ( .A(n12263), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15897) );
  AND2_X1 U13825 ( .A1(n15897), .A2(n12323), .ZN(n12244) );
  AOI21_X1 U13826 ( .B1(n12246), .B2(n12245), .A(n12244), .ZN(n15646) );
  NOR2_X1 U13827 ( .A1(n12248), .A2(n12247), .ZN(n12283) );
  AOI22_X1 U13828 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U13829 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U13830 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U13831 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12249) );
  NAND4_X1 U13832 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12258) );
  AOI22_X1 U13833 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U13834 ( .A1(n11752), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U13835 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U13836 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12253) );
  NAND4_X1 U13837 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12257) );
  OR2_X1 U13838 ( .A1(n12258), .A2(n12257), .ZN(n12282) );
  INV_X1 U13839 ( .A(n12282), .ZN(n12259) );
  XNOR2_X1 U13840 ( .A(n12283), .B(n12259), .ZN(n12260) );
  NAND2_X1 U13841 ( .A1(n12260), .A2(n12286), .ZN(n12270) );
  INV_X1 U13842 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15812) );
  NAND2_X1 U13843 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12261) );
  OAI211_X1 U13844 ( .C1(n12317), .C2(n15812), .A(n12315), .B(n12261), .ZN(
        n12262) );
  INV_X1 U13845 ( .A(n12262), .ZN(n12269) );
  INV_X1 U13846 ( .A(n12263), .ZN(n12264) );
  INV_X1 U13847 ( .A(n12265), .ZN(n12266) );
  INV_X1 U13848 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15634) );
  NAND2_X1 U13849 ( .A1(n12266), .A2(n15634), .ZN(n12267) );
  NAND2_X1 U13850 ( .A1(n12322), .A2(n12267), .ZN(n15890) );
  NOR2_X1 U13851 ( .A1(n15890), .A2(n12315), .ZN(n12268) );
  AOI21_X1 U13852 ( .B1(n12270), .B2(n12269), .A(n12268), .ZN(n15633) );
  AOI22_X1 U13853 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U13854 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13855 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U13856 ( .A1(n11672), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12272) );
  NAND4_X1 U13857 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12281) );
  AOI22_X1 U13858 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U13859 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U13860 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12292), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U13861 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12276) );
  NAND4_X1 U13862 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12276), .ZN(
        n12280) );
  NOR2_X1 U13863 ( .A1(n12281), .A2(n12280), .ZN(n12312) );
  NAND2_X1 U13864 ( .A1(n12283), .A2(n12282), .ZN(n12311) );
  XOR2_X1 U13865 ( .A(n12312), .B(n12311), .Z(n12287) );
  INV_X1 U13866 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15805) );
  NAND2_X1 U13867 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12284) );
  OAI211_X1 U13868 ( .C1(n12317), .C2(n15805), .A(n12315), .B(n12284), .ZN(
        n12285) );
  AOI21_X1 U13869 ( .B1(n12287), .B2(n12286), .A(n12285), .ZN(n12288) );
  INV_X1 U13870 ( .A(n12288), .ZN(n12290) );
  XNOR2_X1 U13871 ( .A(n12322), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15879) );
  NAND2_X1 U13872 ( .A1(n15879), .A2(n12323), .ZN(n12289) );
  NAND2_X1 U13873 ( .A1(n12290), .A2(n12289), .ZN(n15620) );
  AOI22_X1 U13874 ( .A1(n12271), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U13875 ( .A1(n12292), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U13876 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U13877 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U13878 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12310) );
  AOI22_X1 U13879 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U13880 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U13881 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U13882 ( .A1(n12304), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11758), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U13883 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12309) );
  NOR2_X1 U13884 ( .A1(n12310), .A2(n12309), .ZN(n12314) );
  NOR2_X1 U13885 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  XOR2_X1 U13886 ( .A(n12314), .B(n12313), .Z(n12321) );
  INV_X1 U13887 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15799) );
  NAND2_X1 U13888 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12316) );
  OAI211_X1 U13889 ( .C1(n12317), .C2(n15799), .A(n12316), .B(n12315), .ZN(
        n12318) );
  INV_X1 U13890 ( .A(n12318), .ZN(n12319) );
  OAI21_X1 U13891 ( .B1(n12321), .B2(n12320), .A(n12319), .ZN(n12325) );
  INV_X1 U13892 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15881) );
  XNOR2_X1 U13893 ( .A(n13478), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15871) );
  NAND2_X1 U13894 ( .A1(n15871), .A2(n12323), .ZN(n12324) );
  NAND2_X1 U13895 ( .A1(n12325), .A2(n12324), .ZN(n15605) );
  AOI22_X1 U13896 ( .A1(n12327), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12326), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U13897 ( .A1(n21810), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12334) );
  XNOR2_X1 U13898 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U13899 ( .A1(n12342), .A2(n12340), .ZN(n12330) );
  NAND2_X1 U13900 ( .A1(n21823), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12329) );
  NAND2_X1 U13901 ( .A1(n12330), .A2(n12329), .ZN(n12351) );
  XNOR2_X1 U13902 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U13903 ( .A1(n12351), .A2(n12352), .ZN(n12332) );
  NAND2_X1 U13904 ( .A1(n21824), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12331) );
  XNOR2_X1 U13905 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12360) );
  INV_X1 U13906 ( .A(n12360), .ZN(n12333) );
  XNOR2_X1 U13907 ( .A(n12361), .B(n12333), .ZN(n12364) );
  OAI21_X1 U13908 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21810), .A(
        n12334), .ZN(n12336) );
  OAI21_X1 U13909 ( .B1(n12343), .B2(n14364), .A(n12392), .ZN(n12355) );
  AOI211_X1 U13910 ( .C1(n12335), .C2(n11645), .A(n12336), .B(n12355), .ZN(
        n12339) );
  INV_X1 U13911 ( .A(n12336), .ZN(n12337) );
  INV_X1 U13912 ( .A(n12375), .ZN(n12368) );
  AOI21_X1 U13913 ( .B1(n12379), .B2(n12337), .A(n12368), .ZN(n12338) );
  NOR2_X1 U13914 ( .A1(n12339), .A2(n12338), .ZN(n12346) );
  INV_X1 U13915 ( .A(n12340), .ZN(n12341) );
  XNOR2_X1 U13916 ( .A(n12342), .B(n12341), .ZN(n12383) );
  NOR3_X1 U13917 ( .A1(n12346), .A2(n13786), .A3(n12383), .ZN(n12350) );
  INV_X1 U13918 ( .A(n12383), .ZN(n12344) );
  AOI22_X1 U13919 ( .A1(n12345), .A2(n12344), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n12343), .ZN(n12349) );
  OAI21_X1 U13920 ( .B1(n14364), .B2(n12383), .A(n12346), .ZN(n12348) );
  NAND3_X1 U13921 ( .A1(n12379), .A2(n14364), .A3(n12383), .ZN(n12347) );
  OAI211_X1 U13922 ( .C1(n12350), .C2(n12349), .A(n12348), .B(n12347), .ZN(
        n12358) );
  XOR2_X1 U13923 ( .A(n12352), .B(n12351), .Z(n12384) );
  INV_X1 U13924 ( .A(n12355), .ZN(n12353) );
  NAND2_X1 U13925 ( .A1(n12379), .A2(n12384), .ZN(n12354) );
  OAI211_X1 U13926 ( .C1(n12384), .C2(n12366), .A(n12353), .B(n12354), .ZN(
        n12357) );
  INV_X1 U13927 ( .A(n12354), .ZN(n12356) );
  AOI22_X1 U13928 ( .A1(n12358), .A2(n12357), .B1(n12356), .B2(n12355), .ZN(
        n12359) );
  OAI21_X1 U13929 ( .B1(n12364), .B2(n12375), .A(n12359), .ZN(n12370) );
  NAND2_X1 U13930 ( .A1(n12361), .A2(n12360), .ZN(n12363) );
  NAND2_X1 U13931 ( .A1(n21825), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U13932 ( .A1(n12363), .A2(n12362), .ZN(n12372) );
  NOR2_X1 U13933 ( .A1(n12372), .A2(n12373), .ZN(n12367) );
  INV_X1 U13934 ( .A(n12364), .ZN(n12365) );
  OR2_X1 U13935 ( .A1(n12367), .A2(n12365), .ZN(n12386) );
  NAND2_X1 U13936 ( .A1(n12386), .A2(n12366), .ZN(n12369) );
  AOI222_X1 U13937 ( .A1(n12370), .A2(n12369), .B1(n12368), .B2(n12367), .C1(
        n11213), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12377) );
  INV_X1 U13938 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17062) );
  NOR2_X1 U13939 ( .A1(n12375), .A2(n12387), .ZN(n12376) );
  INV_X1 U13940 ( .A(n12387), .ZN(n12378) );
  AND2_X2 U13941 ( .A1(n11645), .A2(n14364), .ZN(n13785) );
  NAND3_X1 U13942 ( .A1(n15546), .A2(n14115), .A3(n13785), .ZN(n12389) );
  NAND2_X1 U13943 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  OR2_X1 U13944 ( .A1(n12386), .A2(n12385), .ZN(n12388) );
  NAND2_X1 U13945 ( .A1(n12388), .A2(n12387), .ZN(n13629) );
  NAND2_X1 U13946 ( .A1(n12389), .A2(n13654), .ZN(n12390) );
  NOR2_X1 U13947 ( .A1(n13874), .A2(n12392), .ZN(n14101) );
  NAND2_X1 U13948 ( .A1(n15546), .A2(n14101), .ZN(n13793) );
  INV_X1 U13949 ( .A(n14164), .ZN(n22131) );
  NOR2_X1 U13950 ( .A1(n21991), .A2(n22037), .ZN(n12391) );
  NAND4_X1 U13951 ( .A1(n13839), .A2(n22131), .A3(n12391), .A4(n11630), .ZN(
        n13873) );
  OR2_X1 U13952 ( .A1(n13873), .A2(n12392), .ZN(n12393) );
  AND2_X1 U13953 ( .A1(n15852), .A2(n22131), .ZN(n12396) );
  NOR4_X1 U13954 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12401) );
  NOR4_X1 U13955 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12400) );
  NOR4_X1 U13956 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12399) );
  NOR4_X1 U13957 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12398) );
  AND4_X1 U13958 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n12406) );
  NOR4_X1 U13959 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12404) );
  NOR4_X1 U13960 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12403) );
  NOR4_X1 U13961 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12402) );
  AND4_X1 U13962 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n19796), .ZN(
        n12405) );
  NAND2_X1 U13963 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  AOI22_X1 U13964 ( .A1(n21652), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n21649), .ZN(n12408) );
  INV_X1 U13965 ( .A(n12408), .ZN(n12412) );
  INV_X1 U13966 ( .A(DATAI_31_), .ZN(n12410) );
  NOR2_X1 U13967 ( .A1(n21657), .A2(n12410), .ZN(n12411) );
  NOR2_X1 U13968 ( .A1(n12412), .A2(n12411), .ZN(n12413) );
  NAND2_X1 U13969 ( .A1(n12414), .A2(n12413), .ZN(P1_U2873) );
  AOI22_X1 U13970 ( .A1(n10986), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12419) );
  AND2_X4 U13971 ( .A1(n12635), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12633) );
  AOI22_X1 U13972 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12418) );
  AND2_X4 U13973 ( .A1(n14293), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12628) );
  AOI22_X1 U13974 ( .A1(n12634), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U13975 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U13976 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U13977 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U13978 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U13979 ( .A1(n10965), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12420) );
  INV_X4 U13980 ( .A(n15470), .ZN(n12634) );
  AOI22_X1 U13981 ( .A1(n12634), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U13982 ( .A1(n12501), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U13983 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12425) );
  NAND3_X1 U13984 ( .A1(n12428), .A2(n12427), .A3(n11524), .ZN(n12436) );
  AOI22_X1 U13985 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U13986 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U13987 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12433) );
  INV_X1 U13988 ( .A(n12501), .ZN(n12627) );
  AOI22_X1 U13989 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12432) );
  NAND3_X1 U13990 ( .A1(n12434), .A2(n12433), .A3(n12432), .ZN(n12435) );
  NAND2_X2 U13991 ( .A1(n12436), .A2(n12435), .ZN(n14750) );
  AOI22_X1 U13992 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U13993 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U13994 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U13995 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U13996 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U13997 ( .A1(n15466), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U13998 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U13999 ( .A1(n12628), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U14000 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U14001 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U14002 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U14003 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12446) );
  NAND4_X1 U14004 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12451) );
  NAND2_X1 U14005 ( .A1(n12451), .A2(n12450), .ZN(n12458) );
  AOI22_X1 U14006 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U14007 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U14008 ( .A1(n12634), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U14009 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U14010 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12456) );
  NAND2_X1 U14011 ( .A1(n12456), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12457) );
  INV_X1 U14012 ( .A(n14750), .ZN(n13016) );
  AOI22_X1 U14013 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U14014 ( .A1(n10986), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U14015 ( .A1(n10965), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U14016 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12463) );
  NAND4_X1 U14017 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12472) );
  AOI22_X1 U14018 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U14019 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U14020 ( .A1(n12634), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U14021 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12467) );
  NAND4_X1 U14022 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12471) );
  AOI22_X1 U14023 ( .A1(n10965), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U14024 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U14025 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U14026 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12473) );
  NAND3_X1 U14027 ( .A1(n12476), .A2(n12475), .A3(n11519), .ZN(n12482) );
  AOI22_X1 U14028 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U14029 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U14030 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U14031 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12479) );
  NAND3_X1 U14032 ( .A1(n11035), .A2(n12480), .A3(n12479), .ZN(n12481) );
  NAND2_X2 U14033 ( .A1(n12482), .A2(n12481), .ZN(n18334) );
  INV_X2 U14034 ( .A(n18334), .ZN(n19594) );
  AOI22_X1 U14035 ( .A1(n10965), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U14036 ( .A1(n12501), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U14037 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U14038 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12502), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12483) );
  AND3_X1 U14039 ( .A1(n12484), .A2(n12450), .A3(n12483), .ZN(n12485) );
  NAND3_X1 U14040 ( .A1(n12487), .A2(n12486), .A3(n12485), .ZN(n12493) );
  AOI22_X1 U14041 ( .A1(n12634), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U14042 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U14043 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U14044 ( .A1(n10986), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12490) );
  NAND3_X1 U14045 ( .A1(n12491), .A2(n11520), .A3(n12490), .ZN(n12492) );
  NAND2_X1 U14046 ( .A1(n12494), .A2(n12519), .ZN(n12540) );
  NAND2_X1 U14047 ( .A1(n12495), .A2(n12540), .ZN(n12512) );
  NAND2_X1 U14048 ( .A1(n13975), .A2(n19437), .ZN(n12511) );
  AOI22_X1 U14049 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U14050 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U14051 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U14052 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12496) );
  NAND4_X1 U14053 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n12500) );
  NAND2_X1 U14054 ( .A1(n12500), .A2(n12450), .ZN(n12510) );
  AOI22_X1 U14055 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U14056 ( .A1(n12502), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12501), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U14057 ( .A1(n12634), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U14058 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12504) );
  NAND4_X1 U14059 ( .A1(n12507), .A2(n12506), .A3(n12505), .A4(n12504), .ZN(
        n12508) );
  NAND2_X1 U14060 ( .A1(n12508), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12509) );
  NAND2_X2 U14061 ( .A1(n12510), .A2(n12509), .ZN(n13001) );
  INV_X2 U14062 ( .A(n13001), .ZN(n13181) );
  NAND2_X1 U14063 ( .A1(n12521), .A2(n13181), .ZN(n12515) );
  NAND4_X1 U14064 ( .A1(n13001), .A2(n12519), .A3(n10981), .A4(n14750), .ZN(
        n12528) );
  INV_X1 U14065 ( .A(n12528), .ZN(n12513) );
  NAND3_X1 U14066 ( .A1(n12513), .A2(n12512), .A3(n12511), .ZN(n12514) );
  AND2_X1 U14067 ( .A1(n13975), .A2(n12516), .ZN(n12517) );
  NAND2_X1 U14068 ( .A1(n12560), .A2(n18334), .ZN(n12518) );
  NAND2_X1 U14069 ( .A1(n13192), .A2(n12518), .ZN(n12562) );
  INV_X1 U14070 ( .A(n12521), .ZN(n12522) );
  NAND2_X1 U14071 ( .A1(n12523), .A2(n12522), .ZN(n13041) );
  NAND3_X1 U14072 ( .A1(n13041), .A2(n13181), .A3(n18335), .ZN(n12524) );
  NOR2_X1 U14073 ( .A1(n12528), .A2(n19594), .ZN(n12529) );
  INV_X1 U14074 ( .A(n12537), .ZN(n12533) );
  OAI21_X1 U14075 ( .B1(n12537), .B2(n12536), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n12543) );
  MUX2_X1 U14076 ( .A(n12539), .B(n13974), .S(n19437), .Z(n12542) );
  INV_X1 U14077 ( .A(n12540), .ZN(n12541) );
  AOI22_X1 U14078 ( .A1(n12556), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12546) );
  INV_X1 U14079 ( .A(n12546), .ZN(n12550) );
  INV_X1 U14080 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12548) );
  INV_X1 U14081 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12555) );
  OAI21_X1 U14082 ( .B1(n12586), .B2(n12555), .A(n12554), .ZN(n12559) );
  INV_X1 U14083 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13775) );
  NAND2_X1 U14084 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12557) );
  NOR2_X1 U14085 ( .A1(n12559), .A2(n12558), .ZN(n12566) );
  NAND2_X1 U14086 ( .A1(n12561), .A2(n12560), .ZN(n13198) );
  INV_X1 U14087 ( .A(n12562), .ZN(n12563) );
  AOI21_X1 U14088 ( .B1(n13198), .B2(n12563), .A(n18340), .ZN(n12564) );
  INV_X1 U14089 ( .A(n12564), .ZN(n12565) );
  AND3_X1 U14090 ( .A1(n12567), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11287), 
        .ZN(n12568) );
  INV_X1 U14091 ( .A(n18637), .ZN(n12583) );
  NAND2_X1 U14092 ( .A1(n12583), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12569) );
  AND2_X1 U14093 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  AOI21_X1 U14094 ( .B1(n18340), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12572) );
  NAND2_X1 U14095 ( .A1(n12573), .A2(n12572), .ZN(n12578) );
  INV_X1 U14096 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12577) );
  NAND2_X1 U14097 ( .A1(n12574), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12576) );
  AND2_X2 U14098 ( .A1(n12580), .A2(n12579), .ZN(n12596) );
  NAND2_X1 U14099 ( .A1(n12582), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12585) );
  NAND2_X1 U14100 ( .A1(n12583), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U14101 ( .A1(n12585), .A2(n12584), .ZN(n12590) );
  INV_X1 U14102 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13263) );
  NAND2_X1 U14103 ( .A1(n12574), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12588) );
  AOI22_X1 U14104 ( .A1(n12556), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12587) );
  OAI211_X1 U14105 ( .C1(n12586), .C2(n13263), .A(n12588), .B(n12587), .ZN(
        n12589) );
  NAND2_X1 U14106 ( .A1(n12590), .A2(n12589), .ZN(n12591) );
  NAND2_X1 U14107 ( .A1(n18349), .A2(n12606), .ZN(n12618) );
  INV_X1 U14108 ( .A(n12618), .ZN(n12595) );
  INV_X1 U14109 ( .A(n12599), .ZN(n12601) );
  NAND2_X1 U14110 ( .A1(n12601), .A2(n12600), .ZN(n12620) );
  INV_X1 U14111 ( .A(n12620), .ZN(n12602) );
  AND2_X1 U14112 ( .A1(n14021), .A2(n12602), .ZN(n12603) );
  INV_X1 U14113 ( .A(n12605), .ZN(n12607) );
  NAND2_X1 U14114 ( .A1(n12607), .A2(n12606), .ZN(n12608) );
  INV_X1 U14115 ( .A(n12830), .ZN(n19203) );
  INV_X1 U14116 ( .A(n13945), .ZN(n12609) );
  OR2_X2 U14117 ( .A1(n14021), .A2(n12609), .ZN(n12621) );
  NAND2_X1 U14118 ( .A1(n16241), .A2(n18587), .ZN(n12610) );
  NOR2_X2 U14119 ( .A1(n12621), .A2(n12610), .ZN(n14741) );
  NAND2_X1 U14120 ( .A1(n13995), .A2(n18587), .ZN(n12611) );
  NOR2_X1 U14121 ( .A1(n18624), .A2(n13995), .ZN(n12612) );
  NAND2_X1 U14122 ( .A1(n12614), .A2(n12612), .ZN(n19173) );
  INV_X1 U14123 ( .A(n19173), .ZN(n12615) );
  AND2_X1 U14124 ( .A1(n18624), .A2(n16241), .ZN(n12613) );
  NAND2_X1 U14125 ( .A1(n12617), .A2(n18624), .ZN(n12711) );
  INV_X1 U14126 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12624) );
  NOR2_X2 U14127 ( .A1(n12619), .A2(n12618), .ZN(n19280) );
  NAND2_X1 U14128 ( .A1(n19280), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12623) );
  NOR2_X2 U14129 ( .A1(n12621), .A2(n12620), .ZN(n19208) );
  NAND2_X1 U14130 ( .A1(n19208), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12622) );
  OAI211_X1 U14131 ( .C1(n12711), .C2(n12624), .A(n12623), .B(n12622), .ZN(
        n12625) );
  INV_X1 U14132 ( .A(n12625), .ZN(n12626) );
  AND2_X2 U14133 ( .A1(n10986), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12684) );
  AND2_X2 U14134 ( .A1(n15466), .A2(n12450), .ZN(n12834) );
  AOI22_X1 U14135 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12632) );
  INV_X2 U14136 ( .A(n12627), .ZN(n15475) );
  AND2_X2 U14137 ( .A1(n15466), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12694) );
  AOI22_X1 U14138 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14139 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12630) );
  AND2_X2 U14140 ( .A1(n10989), .A2(n12450), .ZN(n15409) );
  AOI22_X1 U14141 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12629) );
  NAND4_X1 U14142 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n12642) );
  AND2_X2 U14143 ( .A1(n12633), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12725) );
  AND2_X2 U14144 ( .A1(n12633), .A2(n12450), .ZN(n15414) );
  AOI22_X1 U14145 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12640) );
  AND2_X2 U14146 ( .A1(n12634), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12699) );
  AND2_X2 U14147 ( .A1(n15462), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13274) );
  AOI22_X1 U14148 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12639) );
  AND2_X1 U14149 ( .A1(n12635), .A2(n15284), .ZN(n12672) );
  AOI22_X1 U14150 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12638) );
  AND2_X1 U14151 ( .A1(n12636), .A2(n15284), .ZN(n12661) );
  AOI22_X1 U14152 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12637) );
  NAND4_X1 U14153 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12641) );
  INV_X1 U14154 ( .A(n13260), .ZN(n12643) );
  NAND2_X1 U14155 ( .A1(n12643), .A2(n15436), .ZN(n12644) );
  AOI22_X1 U14156 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14741), .B1(
        n19236), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U14157 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19264), .B1(
        n19208), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U14158 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19280), .B1(
        n14881), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U14159 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19250), .B1(
        n19138), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12645) );
  INV_X1 U14160 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15312) );
  INV_X1 U14161 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12649) );
  OAI22_X1 U14162 ( .A1(n15312), .A2(n12711), .B1(n12830), .B2(n12649), .ZN(
        n12651) );
  INV_X1 U14163 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15314) );
  INV_X1 U14164 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14795) );
  OAI22_X1 U14165 ( .A1(n15314), .A2(n19173), .B1(n14774), .B2(n14795), .ZN(
        n12650) );
  NOR2_X1 U14166 ( .A1(n12651), .A2(n12650), .ZN(n12655) );
  NAND2_X1 U14167 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12654) );
  AOI21_X1 U14168 ( .B1(n19121), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n15436), .ZN(n12653) );
  AOI22_X1 U14169 ( .A1(n12834), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U14170 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U14171 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12656), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U14172 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12657) );
  NAND4_X1 U14173 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12667) );
  AOI22_X1 U14174 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12665) );
  INV_X1 U14175 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19708) );
  AOI22_X1 U14176 ( .A1(n13274), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U14177 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U14178 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U14179 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12666) );
  AND2_X1 U14180 ( .A1(n15436), .A2(n13233), .ZN(n13044) );
  AOI22_X1 U14181 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U14182 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12743), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U14183 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U14184 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12668) );
  NAND4_X1 U14185 ( .A1(n12671), .A2(n12670), .A3(n12669), .A4(n12668), .ZN(
        n12679) );
  AOI22_X1 U14186 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15414), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U14187 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U14188 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U14189 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12674) );
  NAND4_X1 U14190 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12678) );
  AOI22_X1 U14191 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U14192 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U14193 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U14194 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U14195 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12680) );
  NAND4_X1 U14196 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12689) );
  AOI22_X1 U14197 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U14198 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U14199 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12685) );
  NAND3_X1 U14200 ( .A1(n12687), .A2(n12686), .A3(n12685), .ZN(n12688) );
  AOI22_X1 U14201 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U14202 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U14203 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U14204 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12695) );
  NAND4_X1 U14205 ( .A1(n12698), .A2(n12697), .A3(n12696), .A4(n12695), .ZN(
        n12705) );
  AOI22_X1 U14206 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n15414), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U14207 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U14208 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U14209 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U14210 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12704) );
  INV_X1 U14211 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12706) );
  INV_X1 U14212 ( .A(n19121), .ZN(n19126) );
  INV_X1 U14213 ( .A(n19190), .ZN(n19187) );
  INV_X1 U14214 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15380) );
  OAI22_X1 U14215 ( .A1(n12706), .A2(n19126), .B1(n19187), .B2(n15380), .ZN(
        n12710) );
  INV_X1 U14216 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12708) );
  INV_X1 U14217 ( .A(n19160), .ZN(n19164) );
  INV_X1 U14218 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12707) );
  OAI22_X1 U14219 ( .A1(n12708), .A2(n19164), .B1(n14774), .B2(n12707), .ZN(
        n12709) );
  NOR2_X1 U14220 ( .A1(n12710), .A2(n12709), .ZN(n12715) );
  AOI22_X1 U14221 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14741), .B1(
        n14602), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U14222 ( .A1(n19203), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12713) );
  INV_X1 U14223 ( .A(n12711), .ZN(n19149) );
  NAND2_X1 U14224 ( .A1(n19149), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12712) );
  NAND4_X1 U14225 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12712), .ZN(
        n12724) );
  AOI22_X1 U14226 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19250), .B1(
        n14881), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U14227 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19280), .B1(
        n19208), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U14228 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19236), .B1(
        n19264), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12720) );
  INV_X1 U14229 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12717) );
  INV_X1 U14230 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12716) );
  OAI22_X1 U14231 ( .A1(n12717), .A2(n19173), .B1(n12820), .B2(n12716), .ZN(
        n12718) );
  INV_X1 U14232 ( .A(n12718), .ZN(n12719) );
  NAND4_X1 U14233 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12723) );
  AOI22_X1 U14234 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U14235 ( .A1(n12834), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U14236 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U14237 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U14238 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12736) );
  AOI22_X1 U14239 ( .A1(n15414), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U14240 ( .A1(n13274), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12656), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U14241 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U14242 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12673), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12731) );
  NAND4_X1 U14243 ( .A1(n12734), .A2(n12733), .A3(n12732), .A4(n12731), .ZN(
        n12735) );
  INV_X1 U14244 ( .A(n12781), .ZN(n12737) );
  NAND2_X1 U14245 ( .A1(n12737), .A2(n15436), .ZN(n12738) );
  NAND2_X1 U14246 ( .A1(n12740), .A2(n12741), .ZN(n12742) );
  AND2_X2 U14247 ( .A1(n12742), .A2(n13070), .ZN(n13056) );
  NAND2_X1 U14248 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12747) );
  NAND2_X1 U14249 ( .A1(n12834), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12746) );
  NAND2_X1 U14250 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12745) );
  NAND2_X1 U14251 ( .A1(n12694), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12744) );
  NAND2_X1 U14252 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12751) );
  NAND2_X1 U14253 ( .A1(n15414), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12750) );
  AOI22_X1 U14254 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U14255 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U14256 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U14257 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12755) );
  NAND2_X1 U14258 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12754) );
  INV_X1 U14259 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19296) );
  NAND2_X1 U14260 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12753) );
  NAND2_X1 U14261 ( .A1(n15409), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12752) );
  AND4_X2 U14262 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12935) );
  NAND2_X1 U14263 ( .A1(n13056), .A2(n12935), .ZN(n12789) );
  INV_X1 U14264 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12770) );
  NAND2_X1 U14265 ( .A1(n12985), .A2(n12795), .ZN(n12761) );
  NAND2_X1 U14266 ( .A1(n19272), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12760) );
  NAND2_X1 U14267 ( .A1(n12761), .A2(n12760), .ZN(n12765) );
  INV_X1 U14268 ( .A(n12765), .ZN(n12763) );
  MUX2_X1 U14269 ( .A(n19172), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12764) );
  INV_X1 U14270 ( .A(n12764), .ZN(n12762) );
  NAND2_X1 U14271 ( .A1(n12763), .A2(n12762), .ZN(n12766) );
  NAND2_X1 U14272 ( .A1(n12765), .A2(n12764), .ZN(n12773) );
  NAND2_X1 U14273 ( .A1(n12766), .A2(n12773), .ZN(n12988) );
  INV_X1 U14274 ( .A(n13027), .ZN(n12768) );
  NAND2_X1 U14275 ( .A1(n11287), .A2(n13248), .ZN(n12767) );
  NAND2_X1 U14276 ( .A1(n12768), .A2(n12767), .ZN(n12769) );
  NOR2_X1 U14277 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12771) );
  NAND2_X1 U14278 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19172), .ZN(
        n12772) );
  XNOR2_X1 U14279 ( .A(n12775), .B(n12776), .ZN(n13005) );
  MUX2_X1 U14280 ( .A(n13260), .B(n13005), .S(n12544), .Z(n12982) );
  INV_X1 U14281 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12774) );
  MUX2_X1 U14282 ( .A(n12982), .B(n12774), .S(n10975), .Z(n12790) );
  NAND3_X1 U14283 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12995), .A3(
        n18581), .ZN(n13008) );
  MUX2_X1 U14284 ( .A(n13229), .B(n13008), .S(n12544), .Z(n12983) );
  INV_X1 U14285 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12779) );
  MUX2_X1 U14286 ( .A(n12983), .B(n12779), .S(n10974), .Z(n12810) );
  INV_X1 U14287 ( .A(n12810), .ZN(n12780) );
  NAND2_X1 U14288 ( .A1(n13182), .A2(n12781), .ZN(n13222) );
  INV_X1 U14289 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U14290 ( .A1(n10975), .A2(n12782), .ZN(n12783) );
  NAND2_X1 U14291 ( .A1(n13222), .A2(n12783), .ZN(n12785) );
  NAND2_X1 U14292 ( .A1(n12784), .A2(n12785), .ZN(n12849) );
  INV_X1 U14293 ( .A(n12784), .ZN(n12787) );
  INV_X1 U14294 ( .A(n12785), .ZN(n12786) );
  NAND2_X1 U14295 ( .A1(n12787), .A2(n12786), .ZN(n12788) );
  NAND2_X1 U14296 ( .A1(n12849), .A2(n12788), .ZN(n18362) );
  NAND2_X1 U14297 ( .A1(n14533), .A2(n12935), .ZN(n12794) );
  INV_X1 U14298 ( .A(n12790), .ZN(n12792) );
  INV_X1 U14299 ( .A(n12791), .ZN(n12807) );
  NAND2_X1 U14300 ( .A1(n12792), .A2(n12807), .ZN(n12793) );
  NAND2_X1 U14301 ( .A1(n12809), .A2(n12793), .ZN(n14639) );
  NAND2_X1 U14302 ( .A1(n12794), .A2(n14639), .ZN(n14610) );
  INV_X1 U14303 ( .A(n12795), .ZN(n12984) );
  NAND2_X1 U14304 ( .A1(n12415), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12796) );
  AND2_X1 U14305 ( .A1(n12984), .A2(n12796), .ZN(n13006) );
  MUX2_X1 U14306 ( .A(n13006), .B(n13233), .S(n11287), .Z(n12797) );
  MUX2_X1 U14307 ( .A(n12797), .B(P2_EBX_REG_0__SCAN_IN), .S(n10975), .Z(
        n18351) );
  INV_X1 U14308 ( .A(n18351), .ZN(n12798) );
  INV_X1 U14309 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14627) );
  NOR2_X1 U14310 ( .A1(n12798), .A2(n14627), .ZN(n12800) );
  AND3_X1 U14311 ( .A1(n10975), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12799) );
  NOR2_X1 U14312 ( .A1(n12803), .A2(n12799), .ZN(n16233) );
  NOR2_X1 U14313 ( .A1(n12800), .A2(n16233), .ZN(n13852) );
  AND2_X1 U14314 ( .A1(n12800), .A2(n16233), .ZN(n13853) );
  NOR2_X1 U14315 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13853), .ZN(
        n12801) );
  NOR2_X1 U14316 ( .A1(n13852), .A2(n12801), .ZN(n15526) );
  INV_X1 U14317 ( .A(n12802), .ZN(n12805) );
  INV_X1 U14318 ( .A(n12803), .ZN(n12804) );
  NAND2_X1 U14319 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  NAND2_X1 U14320 ( .A1(n12807), .A2(n12806), .ZN(n14812) );
  XNOR2_X1 U14321 ( .A(n14812), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15524) );
  INV_X1 U14322 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18635) );
  NOR2_X1 U14323 ( .A1(n14812), .A2(n18635), .ZN(n12808) );
  AOI21_X1 U14324 ( .B1(n15526), .B2(n15524), .A(n12808), .ZN(n12811) );
  INV_X1 U14325 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14529) );
  XNOR2_X1 U14326 ( .A(n12810), .B(n12809), .ZN(n14764) );
  NOR2_X1 U14327 ( .A1(n14764), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12812) );
  AOI21_X1 U14328 ( .B1(n12811), .B2(n14529), .A(n12812), .ZN(n12817) );
  INV_X1 U14329 ( .A(n12811), .ZN(n14611) );
  INV_X1 U14330 ( .A(n12812), .ZN(n12813) );
  NAND3_X1 U14331 ( .A1(n14611), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n12813), .ZN(n12815) );
  NAND2_X1 U14332 ( .A1(n14764), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12814) );
  NAND2_X1 U14333 ( .A1(n12815), .A2(n12814), .ZN(n12816) );
  AOI21_X1 U14334 ( .B1(n14610), .B2(n12817), .A(n12816), .ZN(n14831) );
  INV_X1 U14335 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U14336 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19208), .B1(
        n19264), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U14337 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14741), .B1(
        n14602), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U14338 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19280), .B1(
        n19250), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12824) );
  INV_X1 U14339 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12821) );
  INV_X1 U14340 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12819) );
  OAI22_X1 U14341 ( .A1(n12821), .A2(n19173), .B1(n12820), .B2(n12819), .ZN(
        n12822) );
  INV_X1 U14342 ( .A(n12822), .ZN(n12823) );
  INV_X1 U14343 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U14344 ( .A1(n19236), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12828) );
  NAND2_X1 U14345 ( .A1(n14881), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12827) );
  OAI211_X1 U14346 ( .C1(n12830), .C2(n12829), .A(n12828), .B(n12827), .ZN(
        n12833) );
  INV_X1 U14347 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U14348 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19190), .B1(
        n19121), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U14349 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19160), .B1(
        n14778), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U14350 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U14351 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12743), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U14352 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U14353 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12836) );
  NAND4_X1 U14354 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        n12845) );
  AOI22_X1 U14355 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n15414), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U14356 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U14357 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U14358 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12840) );
  NAND4_X1 U14359 ( .A1(n12843), .A2(n12842), .A3(n12841), .A4(n12840), .ZN(
        n12844) );
  NAND2_X1 U14360 ( .A1(n12847), .A2(n15436), .ZN(n12846) );
  MUX2_X1 U14361 ( .A(n12847), .B(P2_EBX_REG_6__SCAN_IN), .S(n10975), .Z(
        n12850) );
  XNOR2_X1 U14362 ( .A(n12849), .B(n12850), .ZN(n18373) );
  INV_X1 U14363 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18597) );
  INV_X1 U14364 ( .A(n12850), .ZN(n12851) );
  INV_X1 U14365 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12852) );
  MUX2_X1 U14366 ( .A(n12969), .B(n12852), .S(n10974), .Z(n12853) );
  XNOR2_X1 U14367 ( .A(n12976), .B(n12853), .ZN(n18388) );
  NAND2_X1 U14368 ( .A1(n18388), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16634) );
  NAND2_X1 U14369 ( .A1(n10975), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12854) );
  INV_X1 U14370 ( .A(n12857), .ZN(n12864) );
  INV_X1 U14371 ( .A(n12854), .ZN(n12855) );
  NAND2_X1 U14372 ( .A1(n11076), .A2(n12855), .ZN(n12856) );
  NAND2_X1 U14373 ( .A1(n12864), .A2(n12856), .ZN(n14732) );
  NAND2_X1 U14374 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13076) );
  NOR2_X1 U14375 ( .A1(n14732), .A2(n13076), .ZN(n16609) );
  NAND2_X1 U14376 ( .A1(n10975), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12863) );
  NAND2_X1 U14377 ( .A1(n12857), .A2(n12863), .ZN(n12861) );
  INV_X1 U14378 ( .A(n12861), .ZN(n12859) );
  NAND2_X1 U14379 ( .A1(n12861), .A2(n12860), .ZN(n12862) );
  NAND2_X1 U14380 ( .A1(n12874), .A2(n12862), .ZN(n14808) );
  INV_X1 U14381 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16905) );
  OAI21_X1 U14382 ( .B1(n14808), .B2(n12935), .A(n16905), .ZN(n16612) );
  XNOR2_X1 U14383 ( .A(n12864), .B(n12863), .ZN(n18400) );
  NAND2_X1 U14384 ( .A1(n18400), .A2(n12969), .ZN(n12865) );
  INV_X1 U14385 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16888) );
  NAND2_X1 U14386 ( .A1(n12865), .A2(n16888), .ZN(n16622) );
  INV_X1 U14387 ( .A(n18388), .ZN(n12866) );
  INV_X1 U14388 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18595) );
  NAND2_X1 U14389 ( .A1(n12866), .A2(n18595), .ZN(n16635) );
  INV_X1 U14390 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18598) );
  OAI21_X1 U14391 ( .B1(n14732), .B2(n12935), .A(n18598), .ZN(n17287) );
  AND4_X1 U14392 ( .A1(n16612), .A2(n16622), .A3(n16635), .A4(n17287), .ZN(
        n12867) );
  INV_X1 U14393 ( .A(n14808), .ZN(n12869) );
  AND2_X1 U14394 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12868) );
  NAND2_X1 U14395 ( .A1(n12869), .A2(n12868), .ZN(n16611) );
  AND2_X1 U14396 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U14397 ( .A1(n18400), .A2(n12870), .ZN(n16621) );
  NAND2_X1 U14398 ( .A1(n10975), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12872) );
  INV_X1 U14399 ( .A(n12872), .ZN(n12873) );
  NAND2_X1 U14400 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  NAND2_X1 U14401 ( .A1(n12878), .A2(n12875), .ZN(n18409) );
  OR2_X1 U14402 ( .A1(n18409), .A2(n12935), .ZN(n12909) );
  INV_X1 U14403 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16891) );
  XNOR2_X1 U14404 ( .A(n12909), .B(n16891), .ZN(n16601) );
  NAND2_X1 U14405 ( .A1(n10974), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12877) );
  XNOR2_X1 U14406 ( .A(n12878), .B(n12877), .ZN(n14819) );
  AND2_X1 U14407 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12876) );
  NAND2_X1 U14408 ( .A1(n10974), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U14409 ( .A1(n10974), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12894) );
  OR2_X2 U14410 ( .A1(n12900), .A2(n12898), .ZN(n12907) );
  NOR2_X2 U14411 ( .A1(n12907), .A2(n12905), .ZN(n12902) );
  NAND2_X1 U14412 ( .A1(n10975), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12903) );
  NAND2_X1 U14413 ( .A1(n10975), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U14414 ( .A1(n12916), .A2(n11102), .ZN(n12879) );
  NAND2_X1 U14415 ( .A1(n12928), .A2(n12879), .ZN(n18510) );
  OR2_X1 U14416 ( .A1(n18510), .A2(n12935), .ZN(n12880) );
  INV_X1 U14417 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16494) );
  NAND2_X1 U14418 ( .A1(n12880), .A2(n16494), .ZN(n16489) );
  INV_X1 U14419 ( .A(n12881), .ZN(n12882) );
  XNOR2_X1 U14420 ( .A(n12883), .B(n12882), .ZN(n18452) );
  NAND2_X1 U14421 ( .A1(n18452), .A2(n12969), .ZN(n12884) );
  XNOR2_X1 U14422 ( .A(n12884), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16544) );
  INV_X1 U14423 ( .A(n12885), .ZN(n12887) );
  XNOR2_X1 U14424 ( .A(n12887), .B(n12886), .ZN(n14717) );
  NAND2_X1 U14425 ( .A1(n14717), .A2(n12969), .ZN(n12888) );
  INV_X1 U14426 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16854) );
  NAND2_X1 U14427 ( .A1(n12888), .A2(n16854), .ZN(n16557) );
  INV_X1 U14428 ( .A(n12889), .ZN(n12890) );
  XNOR2_X1 U14429 ( .A(n12891), .B(n12890), .ZN(n18423) );
  NAND2_X1 U14430 ( .A1(n18423), .A2(n12969), .ZN(n12892) );
  INV_X1 U14431 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16853) );
  NAND2_X1 U14432 ( .A1(n12892), .A2(n16853), .ZN(n16579) );
  AND2_X1 U14433 ( .A1(n16557), .A2(n16579), .ZN(n12897) );
  INV_X1 U14434 ( .A(n12893), .ZN(n12895) );
  XNOR2_X1 U14435 ( .A(n12895), .B(n12894), .ZN(n18440) );
  NAND2_X1 U14436 ( .A1(n18440), .A2(n12969), .ZN(n12896) );
  INV_X1 U14437 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16839) );
  NAND2_X1 U14438 ( .A1(n12896), .A2(n16839), .ZN(n16553) );
  AND2_X1 U14439 ( .A1(n12897), .A2(n16553), .ZN(n16528) );
  INV_X1 U14440 ( .A(n12898), .ZN(n12899) );
  XNOR2_X1 U14441 ( .A(n12900), .B(n12899), .ZN(n18464) );
  NAND2_X1 U14442 ( .A1(n18464), .A2(n12969), .ZN(n12901) );
  INV_X1 U14443 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16816) );
  NAND2_X1 U14444 ( .A1(n12901), .A2(n16816), .ZN(n16532) );
  INV_X1 U14445 ( .A(n12902), .ZN(n12904) );
  XNOR2_X1 U14446 ( .A(n12904), .B(n12903), .ZN(n18487) );
  NAND2_X1 U14447 ( .A1(n18487), .A2(n12969), .ZN(n12920) );
  INV_X1 U14448 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16783) );
  NAND2_X1 U14449 ( .A1(n12920), .A2(n16783), .ZN(n16507) );
  INV_X1 U14450 ( .A(n12905), .ZN(n12906) );
  XNOR2_X1 U14451 ( .A(n12907), .B(n12906), .ZN(n18476) );
  NAND2_X1 U14452 ( .A1(n18476), .A2(n12969), .ZN(n12908) );
  INV_X1 U14453 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16516) );
  NAND2_X1 U14454 ( .A1(n12908), .A2(n16516), .ZN(n16519) );
  AND2_X1 U14455 ( .A1(n16507), .A2(n16519), .ZN(n16482) );
  NAND2_X1 U14456 ( .A1(n12909), .A2(n16891), .ZN(n16476) );
  NAND2_X1 U14457 ( .A1(n16476), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12910) );
  NAND2_X1 U14458 ( .A1(n14819), .A2(n12969), .ZN(n16477) );
  NAND2_X1 U14459 ( .A1(n12910), .A2(n16477), .ZN(n12911) );
  AND4_X1 U14460 ( .A1(n16489), .A2(n16481), .A3(n16482), .A4(n12911), .ZN(
        n12912) );
  INV_X1 U14461 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16763) );
  NAND2_X1 U14462 ( .A1(n12918), .A2(n16763), .ZN(n12917) );
  INV_X1 U14463 ( .A(n12913), .ZN(n12914) );
  NAND2_X1 U14464 ( .A1(n11044), .A2(n12914), .ZN(n12915) );
  NAND2_X1 U14465 ( .A1(n12916), .A2(n12915), .ZN(n18499) );
  NOR2_X1 U14466 ( .A1(n18499), .A2(n12935), .ZN(n16486) );
  INV_X1 U14467 ( .A(n12918), .ZN(n12927) );
  NAND2_X1 U14468 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12919) );
  OR2_X1 U14469 ( .A1(n18510), .A2(n12919), .ZN(n16488) );
  OR2_X1 U14470 ( .A1(n12920), .A2(n16783), .ZN(n16508) );
  AND2_X1 U14471 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U14472 ( .A1(n18476), .A2(n12921), .ZN(n16518) );
  AND2_X1 U14473 ( .A1(n16508), .A2(n16518), .ZN(n16484) );
  AND2_X1 U14474 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12922) );
  NAND2_X1 U14475 ( .A1(n18464), .A2(n12922), .ZN(n16531) );
  INV_X1 U14476 ( .A(n18452), .ZN(n12923) );
  INV_X1 U14477 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16831) );
  OR3_X1 U14478 ( .A1(n12923), .A2(n12935), .A3(n16831), .ZN(n16530) );
  AND2_X1 U14479 ( .A1(n16531), .A2(n16530), .ZN(n16479) );
  AND2_X1 U14480 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12924) );
  NAND2_X1 U14481 ( .A1(n18440), .A2(n12924), .ZN(n16552) );
  AND2_X1 U14482 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12925) );
  NAND2_X1 U14483 ( .A1(n18423), .A2(n12925), .ZN(n16578) );
  INV_X1 U14484 ( .A(n14717), .ZN(n12926) );
  OR3_X1 U14485 ( .A1(n12926), .A2(n12935), .A3(n16854), .ZN(n16556) );
  AND3_X1 U14486 ( .A1(n16552), .A2(n16578), .A3(n16556), .ZN(n16478) );
  NAND2_X1 U14487 ( .A1(n10974), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12929) );
  XNOR2_X1 U14488 ( .A(n12928), .B(n12929), .ZN(n18530) );
  NAND2_X1 U14489 ( .A1(n18530), .A2(n12969), .ZN(n16467) );
  INV_X1 U14490 ( .A(n12928), .ZN(n12930) );
  NAND2_X1 U14491 ( .A1(n10974), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12932) );
  INV_X1 U14492 ( .A(n12931), .ZN(n12933) );
  NAND2_X1 U14493 ( .A1(n12933), .A2(n11249), .ZN(n12934) );
  NAND2_X1 U14494 ( .A1(n12938), .A2(n12934), .ZN(n16230) );
  OR2_X1 U14495 ( .A1(n16230), .A2(n12935), .ZN(n12936) );
  INV_X1 U14496 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16710) );
  NAND2_X1 U14497 ( .A1(n12936), .A2(n16710), .ZN(n16458) );
  NAND2_X1 U14498 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12937) );
  NOR2_X1 U14499 ( .A1(n16230), .A2(n12937), .ZN(n16459) );
  NAND2_X1 U14500 ( .A1(n10975), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12939) );
  XNOR2_X1 U14501 ( .A(n12938), .B(n12939), .ZN(n16212) );
  NAND2_X1 U14502 ( .A1(n16212), .A2(n12969), .ZN(n16443) );
  NAND2_X1 U14503 ( .A1(n10975), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U14504 ( .A1(n10974), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12946) );
  XNOR2_X1 U14505 ( .A(n12945), .B(n12946), .ZN(n16185) );
  NAND2_X1 U14506 ( .A1(n16185), .A2(n12969), .ZN(n12940) );
  INV_X1 U14507 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16674) );
  NAND2_X1 U14508 ( .A1(n12940), .A2(n16674), .ZN(n12942) );
  AND2_X1 U14509 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12941) );
  NAND2_X1 U14510 ( .A1(n16185), .A2(n12941), .ZN(n12961) );
  NAND2_X1 U14511 ( .A1(n12942), .A2(n12961), .ZN(n16419) );
  XNOR2_X1 U14512 ( .A(n11027), .B(n12943), .ZN(n18551) );
  NAND2_X1 U14513 ( .A1(n18551), .A2(n12969), .ZN(n12960) );
  INV_X1 U14514 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16675) );
  NOR2_X1 U14515 ( .A1(n16419), .A2(n16434), .ZN(n12944) );
  INV_X1 U14516 ( .A(n12945), .ZN(n12947) );
  NAND2_X1 U14517 ( .A1(n10975), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12949) );
  INV_X1 U14518 ( .A(n12948), .ZN(n12951) );
  INV_X1 U14519 ( .A(n12949), .ZN(n12950) );
  NAND2_X1 U14520 ( .A1(n12951), .A2(n12950), .ZN(n12952) );
  NAND2_X1 U14521 ( .A1(n12954), .A2(n12952), .ZN(n16184) );
  NOR2_X1 U14522 ( .A1(n16184), .A2(n12935), .ZN(n16396) );
  AND2_X1 U14523 ( .A1(n10974), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U14524 ( .A1(n12954), .A2(n12953), .ZN(n12955) );
  NAND2_X1 U14525 ( .A1(n12966), .A2(n12955), .ZN(n16169) );
  OAI21_X1 U14526 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16399), .ZN(n12956) );
  INV_X1 U14527 ( .A(n16399), .ZN(n12958) );
  INV_X1 U14528 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16653) );
  NAND2_X1 U14529 ( .A1(n12958), .A2(n16653), .ZN(n12959) );
  NAND2_X1 U14530 ( .A1(n12961), .A2(n16433), .ZN(n16395) );
  INV_X1 U14531 ( .A(n16395), .ZN(n12962) );
  NAND2_X1 U14532 ( .A1(n10975), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12964) );
  INV_X1 U14533 ( .A(n12966), .ZN(n12963) );
  XOR2_X1 U14534 ( .A(n12964), .B(n12963), .Z(n18573) );
  NAND2_X1 U14535 ( .A1(n18573), .A2(n12969), .ZN(n12971) );
  INV_X1 U14536 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15516) );
  NAND2_X1 U14537 ( .A1(n12971), .A2(n15516), .ZN(n15503) );
  NAND2_X1 U14538 ( .A1(n15504), .A2(n15503), .ZN(n13444) );
  INV_X1 U14539 ( .A(n12964), .ZN(n12965) );
  NAND2_X1 U14540 ( .A1(n10975), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12968) );
  XNOR2_X1 U14541 ( .A(n12973), .B(n12968), .ZN(n16142) );
  AOI21_X1 U14542 ( .B1(n16142), .B2(n12969), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13447) );
  AND2_X1 U14543 ( .A1(n12969), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12970) );
  NAND2_X1 U14544 ( .A1(n16142), .A2(n12970), .ZN(n13445) );
  INV_X1 U14545 ( .A(n12971), .ZN(n12972) );
  NAND2_X1 U14546 ( .A1(n12972), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15502) );
  INV_X1 U14547 ( .A(n12973), .ZN(n12975) );
  INV_X1 U14548 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U14549 ( .A1(n12975), .A2(n12974), .ZN(n12978) );
  INV_X1 U14550 ( .A(n12976), .ZN(n12977) );
  NOR2_X1 U14551 ( .A1(n16141), .A2(n12935), .ZN(n12979) );
  XOR2_X1 U14552 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12979), .Z(
        n12980) );
  XNOR2_X1 U14553 ( .A(n12981), .B(n12980), .ZN(n13432) );
  NAND2_X1 U14554 ( .A1(n12983), .A2(n12982), .ZN(n13029) );
  AND2_X1 U14555 ( .A1(n13008), .A2(n13005), .ZN(n12993) );
  AOI21_X1 U14556 ( .B1(n12998), .B2(n18335), .A(n13007), .ZN(n12991) );
  NAND2_X1 U14557 ( .A1(n13006), .A2(n12985), .ZN(n13025) );
  NAND2_X1 U14558 ( .A1(n11287), .A2(n13025), .ZN(n12987) );
  XNOR2_X1 U14559 ( .A(n12985), .B(n12984), .ZN(n13003) );
  OAI211_X1 U14560 ( .C1(n18335), .C2(n13006), .A(n18334), .B(n13003), .ZN(
        n12986) );
  OAI211_X1 U14561 ( .C1(n12989), .C2(n12988), .A(n12987), .B(n12986), .ZN(
        n12990) );
  OAI21_X1 U14562 ( .B1(n13027), .B2(n12991), .A(n12990), .ZN(n12992) );
  AOI22_X1 U14563 ( .A1(n13029), .A2(n12544), .B1(n12993), .B2(n12992), .ZN(
        n12996) );
  INV_X1 U14564 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17003) );
  NOR2_X1 U14565 ( .A1(n12996), .A2(n13030), .ZN(n12997) );
  MUX2_X1 U14566 ( .A(n12997), .B(n18581), .S(n18340), .Z(n13000) );
  INV_X1 U14567 ( .A(n14591), .ZN(n13969) );
  NAND2_X1 U14568 ( .A1(n13969), .A2(n18335), .ZN(n14275) );
  OAI211_X1 U14569 ( .C1(n19594), .C2(n13000), .A(n14275), .B(n13016), .ZN(
        n13039) );
  INV_X1 U14570 ( .A(n14275), .ZN(n13002) );
  NAND2_X1 U14571 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18655) );
  NOR2_X1 U14572 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n16996) );
  INV_X1 U14573 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21612) );
  INV_X2 U14574 ( .A(n17390), .ZN(n21598) );
  NOR2_X1 U14575 ( .A1(n21594), .A2(n21604), .ZN(n14335) );
  NAND3_X1 U14576 ( .A1(n13002), .A2(n14335), .A3(n13001), .ZN(n13038) );
  AND4_X1 U14577 ( .A1(n13008), .A2(n13007), .A3(n13005), .A4(n13003), .ZN(
        n13004) );
  OR2_X1 U14578 ( .A1(n13030), .A2(n13004), .ZN(n14338) );
  AND4_X1 U14579 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  OAI21_X1 U14580 ( .B1(n14338), .B2(n13009), .A(n16962), .ZN(n13011) );
  NAND2_X1 U14581 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15285) );
  OAI21_X1 U14582 ( .B1(n15285), .B2(n11243), .A(n18581), .ZN(n14330) );
  NOR2_X1 U14583 ( .A1(n16962), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n13010) );
  OAI21_X1 U14584 ( .B1(n12725), .B2(n14330), .A(n13010), .ZN(n17302) );
  NOR2_X1 U14585 ( .A1(n13041), .A2(n15436), .ZN(n13036) );
  MUX2_X1 U14586 ( .A(n14347), .B(n13001), .S(n15436), .Z(n13012) );
  NAND2_X1 U14587 ( .A1(n13012), .A2(n18655), .ZN(n13034) );
  INV_X1 U14588 ( .A(n14335), .ZN(n14345) );
  OR2_X1 U14589 ( .A1(n13013), .A2(n14345), .ZN(n13014) );
  OR2_X1 U14590 ( .A1(n14338), .A2(n13014), .ZN(n13024) );
  OAI21_X1 U14591 ( .B1(n13974), .B2(n14750), .A(n13181), .ZN(n13022) );
  NAND2_X1 U14592 ( .A1(n13017), .A2(n12519), .ZN(n13015) );
  AND2_X1 U14593 ( .A1(n19594), .A2(n15436), .ZN(n14346) );
  NAND2_X1 U14594 ( .A1(n13015), .A2(n14346), .ZN(n13187) );
  OR2_X1 U14595 ( .A1(n13017), .A2(n13016), .ZN(n13020) );
  NAND2_X1 U14596 ( .A1(n19594), .A2(n12519), .ZN(n13018) );
  OAI211_X1 U14597 ( .C1(n18335), .C2(n12540), .A(n13018), .B(n13181), .ZN(
        n13019) );
  NAND4_X1 U14598 ( .A1(n13187), .A2(n13197), .A3(n13020), .A4(n13019), .ZN(
        n13021) );
  AOI21_X1 U14599 ( .B1(n14332), .B2(n13022), .A(n13021), .ZN(n13023) );
  AND2_X1 U14600 ( .A1(n13024), .A2(n13023), .ZN(n14272) );
  INV_X1 U14601 ( .A(n13025), .ZN(n13026) );
  NOR2_X1 U14602 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  NOR2_X1 U14603 ( .A1(n13029), .A2(n13028), .ZN(n13031) );
  OR2_X1 U14604 ( .A1(n13031), .A2(n13030), .ZN(n14322) );
  INV_X1 U14605 ( .A(n14322), .ZN(n13033) );
  INV_X1 U14606 ( .A(n14346), .ZN(n13032) );
  NOR2_X1 U14607 ( .A1(n13041), .A2(n13032), .ZN(n14323) );
  NAND2_X1 U14608 ( .A1(n13033), .A2(n14323), .ZN(n13430) );
  OAI211_X1 U14609 ( .C1(n14338), .C2(n13034), .A(n14272), .B(n13430), .ZN(
        n13035) );
  AOI21_X1 U14610 ( .B1(n18645), .B2(n13036), .A(n13035), .ZN(n13037) );
  NAND3_X1 U14611 ( .A1(n13039), .A2(n13038), .A3(n13037), .ZN(n13040) );
  OR2_X1 U14612 ( .A1(n13041), .A2(n12544), .ZN(n14325) );
  OR2_X1 U14613 ( .A1(n13432), .A2(n18614), .ZN(n13428) );
  XOR2_X1 U14614 ( .A(n13248), .B(n13042), .Z(n15529) );
  INV_X1 U14615 ( .A(n13233), .ZN(n13043) );
  XOR2_X1 U14616 ( .A(n13243), .B(n13043), .Z(n13046) );
  INV_X1 U14617 ( .A(n13044), .ZN(n13748) );
  NAND2_X1 U14618 ( .A1(n13748), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13747) );
  NOR2_X1 U14619 ( .A1(n13046), .A2(n13747), .ZN(n13047) );
  INV_X1 U14620 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14628) );
  INV_X1 U14621 ( .A(n13747), .ZN(n13045) );
  XOR2_X1 U14622 ( .A(n13046), .B(n13045), .Z(n13851) );
  NOR2_X1 U14623 ( .A1(n14628), .A2(n13851), .ZN(n13850) );
  NOR2_X1 U14624 ( .A1(n13047), .A2(n13850), .ZN(n13048) );
  XOR2_X1 U14625 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13048), .Z(
        n15528) );
  NOR2_X1 U14626 ( .A1(n15529), .A2(n15528), .ZN(n15527) );
  NOR2_X1 U14627 ( .A1(n13048), .A2(n18635), .ZN(n13049) );
  XNOR2_X1 U14628 ( .A(n13050), .B(n14529), .ZN(n14532) );
  NAND2_X1 U14629 ( .A1(n13050), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13051) );
  OAI21_X1 U14630 ( .B1(n11007), .B2(n13229), .A(n12740), .ZN(n13053) );
  INV_X1 U14631 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14838) );
  INV_X1 U14632 ( .A(n13052), .ZN(n13054) );
  NAND2_X1 U14633 ( .A1(n13054), .A2(n13053), .ZN(n13055) );
  INV_X1 U14634 ( .A(n13057), .ZN(n13060) );
  OAI21_X1 U14635 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13056), .A(
        n13060), .ZN(n13061) );
  INV_X1 U14636 ( .A(n13071), .ZN(n13063) );
  MUX2_X1 U14637 ( .A(n13063), .B(n12818), .S(n13062), .Z(n13064) );
  OAI21_X1 U14638 ( .B1(n13057), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13064), .ZN(n13065) );
  NAND2_X1 U14639 ( .A1(n13066), .A2(n13067), .ZN(n13068) );
  NAND2_X1 U14640 ( .A1(n13068), .A2(n13057), .ZN(n13069) );
  NAND2_X1 U14641 ( .A1(n16945), .A2(n13069), .ZN(n16639) );
  INV_X1 U14642 ( .A(n13070), .ZN(n13072) );
  XNOR2_X1 U14643 ( .A(n13077), .B(n12935), .ZN(n13073) );
  XNOR2_X1 U14644 ( .A(n13073), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16638) );
  NAND2_X1 U14645 ( .A1(n16639), .A2(n16638), .ZN(n16640) );
  INV_X1 U14646 ( .A(n13073), .ZN(n13074) );
  NAND2_X1 U14647 ( .A1(n13074), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13075) );
  OAI21_X1 U14648 ( .B1(n13077), .B2(n12935), .A(n18598), .ZN(n13078) );
  NAND3_X1 U14649 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16847) );
  INV_X1 U14650 ( .A(n16847), .ZN(n16845) );
  NAND4_X1 U14651 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(n16845), .ZN(n16752) );
  NAND2_X1 U14652 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16760) );
  NOR2_X1 U14653 ( .A1(n16752), .A2(n16760), .ZN(n13080) );
  NOR3_X1 U14654 ( .A1(n16831), .A2(n16839), .A3(n16816), .ZN(n16754) );
  NAND2_X1 U14655 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16754), .ZN(
        n16751) );
  INV_X1 U14656 ( .A(n16751), .ZN(n16777) );
  AND2_X1 U14657 ( .A1(n13080), .A2(n16777), .ZN(n13208) );
  INV_X1 U14658 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16733) );
  NOR2_X4 U14659 ( .A1(n16492), .A2(n16733), .ZN(n16470) );
  AND2_X1 U14660 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16660) );
  INV_X1 U14661 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16666) );
  NAND2_X1 U14662 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13452) );
  NAND2_X1 U14663 ( .A1(n15507), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13081) );
  XNOR2_X1 U14664 ( .A(n13081), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13441) );
  INV_X1 U14665 ( .A(n14323), .ZN(n13082) );
  INV_X1 U14666 ( .A(n13084), .ZN(n13085) );
  AOI22_X1 U14667 ( .A1(n10978), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13088) );
  NAND2_X1 U14668 ( .A1(n13171), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n13087) );
  OAI211_X1 U14669 ( .C1(n13174), .C2(n14838), .A(n13088), .B(n13087), .ZN(
        n14035) );
  INV_X2 U14670 ( .A(n13174), .ZN(n13138) );
  INV_X1 U14671 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U14672 ( .A1(n10978), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13089) );
  OAI21_X1 U14673 ( .B1(n13169), .B2(n13225), .A(n13089), .ZN(n13090) );
  AOI21_X1 U14674 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13138), .A(
        n13090), .ZN(n14040) );
  AOI22_X1 U14675 ( .A1(n13161), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13092) );
  NAND2_X1 U14676 ( .A1(n13171), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n13091) );
  OAI211_X1 U14677 ( .C1(n13174), .C2(n18597), .A(n13092), .B(n13091), .ZN(
        n14158) );
  INV_X1 U14678 ( .A(n14156), .ZN(n14130) );
  NAND2_X1 U14679 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13098) );
  INV_X1 U14680 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n13095) );
  NAND2_X1 U14681 ( .A1(n13161), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13094) );
  NAND2_X1 U14682 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13093) );
  OAI211_X1 U14683 ( .C1(n13169), .C2(n13095), .A(n13094), .B(n13093), .ZN(
        n13096) );
  INV_X1 U14684 ( .A(n13096), .ZN(n13097) );
  NAND2_X1 U14685 ( .A1(n13098), .A2(n13097), .ZN(n14131) );
  NAND2_X1 U14686 ( .A1(n14130), .A2(n14131), .ZN(n14224) );
  INV_X1 U14687 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n18601) );
  NAND2_X1 U14688 ( .A1(n13161), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13101) );
  NAND2_X1 U14689 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13100) );
  OAI211_X1 U14690 ( .C1(n13169), .C2(n18601), .A(n13101), .B(n13100), .ZN(
        n13102) );
  AOI21_X1 U14691 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n13102), .ZN(n14223) );
  INV_X1 U14692 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n18402) );
  NAND2_X1 U14693 ( .A1(n13161), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13104) );
  NAND2_X1 U14694 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13103) );
  OAI211_X1 U14695 ( .C1(n13169), .C2(n18402), .A(n13104), .B(n13103), .ZN(
        n13105) );
  AOI21_X1 U14696 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n13105), .ZN(n14264) );
  INV_X1 U14697 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n16615) );
  NAND2_X1 U14698 ( .A1(n13161), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U14699 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13106) );
  OAI211_X1 U14700 ( .C1(n13169), .C2(n16615), .A(n13107), .B(n13106), .ZN(
        n13108) );
  AOI21_X1 U14701 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n13108), .ZN(n14415) );
  NOR2_X2 U14702 ( .A1(n14416), .A2(n14415), .ZN(n14459) );
  INV_X1 U14703 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16597) );
  NAND2_X1 U14704 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13110) );
  AOI22_X1 U14705 ( .A1(n13161), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n13109) );
  OAI211_X1 U14706 ( .C1(n13169), .C2(n16597), .A(n13110), .B(n13109), .ZN(
        n14458) );
  INV_X1 U14707 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n16590) );
  NAND2_X1 U14708 ( .A1(n13161), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U14709 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13111) );
  OAI211_X1 U14710 ( .C1(n13169), .C2(n16590), .A(n13112), .B(n13111), .ZN(
        n13113) );
  AOI21_X1 U14711 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n13113), .ZN(n14507) );
  INV_X1 U14712 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U14713 ( .A1(n13161), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U14714 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13114) );
  OAI211_X1 U14715 ( .C1(n13169), .C2(n13351), .A(n13115), .B(n13114), .ZN(
        n13116) );
  AOI21_X1 U14716 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n13116), .ZN(n14545) );
  INV_X1 U14717 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U14718 ( .A1(n13161), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13118) );
  NAND2_X1 U14719 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13117) );
  OAI211_X1 U14720 ( .C1(n13169), .C2(n16570), .A(n13118), .B(n13117), .ZN(
        n13119) );
  AOI21_X1 U14721 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n13119), .ZN(n14648) );
  INV_X1 U14722 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n18442) );
  NAND2_X1 U14723 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13121) );
  AOI22_X1 U14724 ( .A1(n10978), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n13120) );
  OAI211_X1 U14725 ( .C1(n13169), .C2(n18442), .A(n13121), .B(n13120), .ZN(
        n14687) );
  INV_X1 U14726 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U14727 ( .A1(n13161), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U14728 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13122) );
  OAI211_X1 U14729 ( .C1(n13169), .C2(n13124), .A(n13123), .B(n13122), .ZN(
        n13125) );
  AOI21_X1 U14730 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n13125), .ZN(n14865) );
  INV_X1 U14731 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n16535) );
  NAND2_X1 U14732 ( .A1(n13161), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U14733 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13126) );
  OAI211_X1 U14734 ( .C1(n13169), .C2(n16535), .A(n13127), .B(n13126), .ZN(
        n13128) );
  AOI21_X1 U14735 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n13128), .ZN(n14930) );
  INV_X1 U14736 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n16522) );
  NAND2_X1 U14737 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13130) );
  AOI22_X1 U14738 ( .A1(n13161), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n13129) );
  OAI211_X1 U14739 ( .C1(n13169), .C2(n16522), .A(n13130), .B(n13129), .ZN(
        n14970) );
  INV_X1 U14740 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18490) );
  NAND2_X1 U14741 ( .A1(n13161), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13132) );
  NAND2_X1 U14742 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13131) );
  OAI211_X1 U14743 ( .C1(n13169), .C2(n18490), .A(n13132), .B(n13131), .ZN(
        n13133) );
  AOI21_X1 U14744 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n13133), .ZN(n15016) );
  INV_X1 U14745 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n13136) );
  NAND2_X1 U14746 ( .A1(n13161), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13135) );
  NAND2_X1 U14747 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13134) );
  OAI211_X1 U14748 ( .C1(n13169), .C2(n13136), .A(n13135), .B(n13134), .ZN(
        n13137) );
  AOI21_X1 U14749 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n13137), .ZN(n16304) );
  INV_X1 U14750 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n18513) );
  NAND2_X1 U14751 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13140) );
  AOI22_X1 U14752 ( .A1(n13161), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n13139) );
  OAI211_X1 U14753 ( .C1(n13169), .C2(n18513), .A(n13140), .B(n13139), .ZN(
        n16297) );
  AND2_X2 U14754 ( .A1(n16303), .A2(n16297), .ZN(n16299) );
  INV_X1 U14755 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n13143) );
  NAND2_X1 U14756 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13142) );
  AOI22_X1 U14757 ( .A1(n13161), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n13141) );
  OAI211_X1 U14758 ( .C1(n13169), .C2(n13143), .A(n13142), .B(n13141), .ZN(
        n16289) );
  INV_X1 U14759 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17380) );
  NAND2_X1 U14760 ( .A1(n10978), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13145) );
  NAND2_X1 U14761 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13144) );
  OAI211_X1 U14762 ( .C1(n13169), .C2(n17380), .A(n13145), .B(n13144), .ZN(
        n13146) );
  AOI21_X1 U14763 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n13146), .ZN(n16220) );
  INV_X1 U14764 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U14765 ( .A1(n10978), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13148) );
  NAND2_X1 U14766 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13147) );
  OAI211_X1 U14767 ( .C1(n13169), .C2(n13149), .A(n13148), .B(n13147), .ZN(
        n13150) );
  AOI21_X1 U14768 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n13150), .ZN(n16201) );
  INV_X1 U14769 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n18547) );
  NAND2_X1 U14770 ( .A1(n10978), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U14771 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13151) );
  OAI211_X1 U14772 ( .C1(n13169), .C2(n18547), .A(n13152), .B(n13151), .ZN(
        n13153) );
  AOI21_X1 U14773 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n13153), .ZN(n16275) );
  INV_X1 U14774 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n13156) );
  NAND2_X1 U14775 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13155) );
  AOI22_X1 U14776 ( .A1(n10978), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n13154) );
  OAI211_X1 U14777 ( .C1(n13169), .C2(n13156), .A(n13155), .B(n13154), .ZN(
        n16186) );
  NAND2_X1 U14778 ( .A1(n16273), .A2(n16186), .ZN(n16188) );
  INV_X1 U14779 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U14780 ( .A1(n13161), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13158) );
  NAND2_X1 U14781 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13157) );
  OAI211_X1 U14782 ( .C1(n13169), .C2(n17384), .A(n13158), .B(n13157), .ZN(
        n13159) );
  AOI21_X1 U14783 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13159), .ZN(n16171) );
  INV_X1 U14784 ( .A(n13160), .ZN(n16170) );
  INV_X1 U14785 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17385) );
  NAND2_X1 U14786 ( .A1(n10978), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13163) );
  NAND2_X1 U14787 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13162) );
  OAI211_X1 U14788 ( .C1(n13169), .C2(n17385), .A(n13163), .B(n13162), .ZN(
        n13164) );
  AOI21_X1 U14789 ( .B1(n13138), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n13164), .ZN(n16156) );
  INV_X1 U14790 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n18563) );
  NAND2_X1 U14791 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13166) );
  AOI22_X1 U14792 ( .A1(n10978), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n13165) );
  OAI211_X1 U14793 ( .C1(n13169), .C2(n18563), .A(n13166), .B(n13165), .ZN(
        n15514) );
  NAND2_X1 U14794 ( .A1(n16155), .A2(n15514), .ZN(n15513) );
  INV_X1 U14795 ( .A(n15513), .ZN(n13170) );
  INV_X1 U14796 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17386) );
  NAND2_X1 U14797 ( .A1(n13138), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13168) );
  AOI22_X1 U14798 ( .A1(n13161), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13167) );
  OAI211_X1 U14799 ( .C1(n13169), .C2(n17386), .A(n13168), .B(n13167), .ZN(
        n13450) );
  INV_X1 U14800 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U14801 ( .A1(n10978), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13173) );
  NAND2_X1 U14802 ( .A1(n13171), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13172) );
  OAI211_X1 U14803 ( .C1(n13174), .C2(n14626), .A(n13173), .B(n13172), .ZN(
        n13175) );
  INV_X1 U14804 ( .A(n13175), .ZN(n13176) );
  AOI21_X1 U14805 ( .B1(n13178), .B2(n15436), .A(n14280), .ZN(n13179) );
  NAND3_X1 U14806 ( .A1(n13182), .A2(n15436), .A3(n13181), .ZN(n13183) );
  INV_X1 U14807 ( .A(n14327), .ZN(n13184) );
  INV_X1 U14808 ( .A(n18615), .ZN(n13185) );
  NAND2_X1 U14809 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U14810 ( .A1(n18635), .A2(n14526), .ZN(n18617) );
  INV_X1 U14811 ( .A(n18617), .ZN(n14528) );
  NOR2_X1 U14812 ( .A1(n14838), .A2(n12818), .ZN(n16947) );
  NAND3_X1 U14813 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n16947), .ZN(n16931) );
  OR3_X1 U14814 ( .A1(n18598), .A2(n18595), .A3(n16931), .ZN(n13200) );
  NOR2_X1 U14815 ( .A1(n14528), .A2(n13200), .ZN(n13206) );
  NAND2_X1 U14816 ( .A1(n13185), .A2(n13206), .ZN(n13202) );
  NAND2_X1 U14817 ( .A1(n13186), .A2(n18335), .ZN(n14289) );
  NAND2_X1 U14818 ( .A1(n14289), .A2(n13187), .ZN(n13195) );
  NAND2_X1 U14819 ( .A1(n13197), .A2(n14750), .ZN(n13189) );
  INV_X1 U14820 ( .A(n13188), .ZN(n13615) );
  AOI22_X1 U14821 ( .A1(n13189), .A2(n13615), .B1(n19594), .B2(n13001), .ZN(
        n13193) );
  NAND2_X1 U14822 ( .A1(n13191), .A2(n13190), .ZN(n13970) );
  NAND3_X1 U14823 ( .A1(n13193), .A2(n13192), .A3(n13970), .ZN(n13194) );
  AOI21_X1 U14824 ( .B1(n19437), .B2(n13195), .A(n13194), .ZN(n13196) );
  OAI21_X1 U14825 ( .B1(n13198), .B2(n13197), .A(n13196), .ZN(n14315) );
  NOR2_X1 U14826 ( .A1(n14315), .A2(n14279), .ZN(n13199) );
  INV_X1 U14827 ( .A(n14526), .ZN(n18619) );
  NAND2_X1 U14828 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18619), .ZN(
        n18616) );
  NOR2_X1 U14829 ( .A1(n13200), .A2(n18616), .ZN(n16804) );
  NAND2_X1 U14830 ( .A1(n16807), .A2(n16804), .ZN(n13201) );
  NAND2_X1 U14831 ( .A1(n13202), .A2(n13201), .ZN(n16890) );
  INV_X1 U14832 ( .A(n16752), .ZN(n16803) );
  NAND2_X1 U14833 ( .A1(n16890), .A2(n16803), .ZN(n16813) );
  NAND2_X1 U14834 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16777), .ZN(
        n13203) );
  NOR2_X1 U14835 ( .A1(n16813), .A2(n13203), .ZN(n16738) );
  AND2_X1 U14836 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U14837 ( .A1(n16738), .A2(n13204), .ZN(n16715) );
  AND2_X1 U14838 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U14839 ( .A1(n16698), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13205) );
  OR2_X1 U14840 ( .A1(n16691), .A2(n16660), .ZN(n13211) );
  INV_X1 U14841 ( .A(n13205), .ZN(n13210) );
  NAND2_X1 U14842 ( .A1(n13423), .A2(n18600), .ZN(n13996) );
  OAI21_X1 U14843 ( .B1(n18615), .B2(n13206), .A(n13996), .ZN(n16750) );
  NOR2_X1 U14844 ( .A1(n16755), .A2(n16804), .ZN(n13207) );
  OR2_X1 U14845 ( .A1(n16750), .A2(n13207), .ZN(n16924) );
  INV_X1 U14846 ( .A(n16924), .ZN(n13209) );
  NAND2_X1 U14847 ( .A1(n13209), .A2(n13208), .ZN(n16742) );
  NAND2_X1 U14848 ( .A1(n18593), .A2(n13996), .ZN(n16887) );
  OAI21_X1 U14849 ( .B1(n16494), .B2(n16742), .A(n16887), .ZN(n16729) );
  OAI21_X1 U14850 ( .B1(n18593), .B2(n13210), .A(n16729), .ZN(n16689) );
  INV_X1 U14851 ( .A(n16689), .ZN(n16702) );
  NAND2_X1 U14852 ( .A1(n13211), .A2(n16702), .ZN(n16680) );
  NOR2_X1 U14853 ( .A1(n18593), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13212) );
  NOR2_X1 U14854 ( .A1(n16680), .A2(n13212), .ZN(n16654) );
  INV_X1 U14855 ( .A(n18593), .ZN(n16930) );
  INV_X1 U14856 ( .A(n13452), .ZN(n13213) );
  NAND2_X1 U14857 ( .A1(n13213), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13216) );
  NAND2_X1 U14858 ( .A1(n16930), .A2(n13216), .ZN(n13214) );
  NAND2_X1 U14859 ( .A1(n16654), .A2(n13214), .ZN(n13453) );
  INV_X1 U14860 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n13416) );
  NOR2_X1 U14861 ( .A1(n18488), .A2(n13416), .ZN(n13438) );
  INV_X1 U14862 ( .A(n16691), .ZN(n13215) );
  NAND3_X1 U14863 ( .A1(n13215), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16660), .ZN(n15515) );
  NOR3_X1 U14864 ( .A1(n15515), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13216), .ZN(n13217) );
  AOI211_X1 U14865 ( .C1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13453), .A(
        n13438), .B(n13217), .ZN(n13425) );
  INV_X1 U14866 ( .A(n13228), .ZN(n13223) );
  NOR2_X1 U14867 ( .A1(n12519), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13218) );
  NAND2_X1 U14868 ( .A1(n13273), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n13221) );
  NAND2_X1 U14869 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13220) );
  OAI211_X1 U14870 ( .C1(n13223), .C2(n13222), .A(n13221), .B(n13220), .ZN(
        n13227) );
  NOR2_X1 U14871 ( .A1(n13417), .A2(n13225), .ZN(n13226) );
  OR2_X1 U14872 ( .A1(n13227), .A2(n13226), .ZN(n14835) );
  INV_X2 U14873 ( .A(n13391), .ZN(n13379) );
  AOI22_X1 U14874 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U14875 ( .A1(n13375), .A2(n13229), .ZN(n13231) );
  INV_X1 U14876 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n14618) );
  OR2_X1 U14877 ( .A1(n13417), .A2(n14618), .ZN(n13230) );
  NAND2_X1 U14878 ( .A1(n13375), .A2(n13233), .ZN(n13235) );
  MUX2_X1 U14879 ( .A(n12519), .B(n19274), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13234) );
  NAND2_X1 U14880 ( .A1(n13219), .A2(n13974), .ZN(n13249) );
  NAND3_X1 U14881 ( .A1(n13235), .A2(n13234), .A3(n13249), .ZN(n13968) );
  INV_X1 U14882 ( .A(n12519), .ZN(n13976) );
  NAND2_X1 U14883 ( .A1(n13976), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n13236) );
  OAI211_X1 U14884 ( .C1(n15436), .C2(n14627), .A(n13236), .B(n19262), .ZN(
        n13237) );
  INV_X1 U14885 ( .A(n13237), .ZN(n13238) );
  AOI22_X1 U14886 ( .A1(n13219), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13218), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13240) );
  OR2_X1 U14887 ( .A1(n13417), .A2(n12548), .ZN(n13239) );
  NAND2_X1 U14888 ( .A1(n13240), .A2(n13239), .ZN(n13246) );
  INV_X1 U14889 ( .A(n13246), .ZN(n13241) );
  NOR2_X1 U14890 ( .A1(n13974), .A2(n13976), .ZN(n13242) );
  MUX2_X1 U14891 ( .A(n13242), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n13245) );
  AND2_X1 U14892 ( .A1(n13375), .A2(n13243), .ZN(n13244) );
  NOR2_X1 U14893 ( .A1(n13245), .A2(n13244), .ZN(n13982) );
  NAND2_X1 U14894 ( .A1(n13981), .A2(n13982), .ZN(n13986) );
  NAND2_X1 U14895 ( .A1(n13375), .A2(n13248), .ZN(n13250) );
  OAI211_X1 U14896 ( .C1(n19262), .C2(n19172), .A(n13250), .B(n13249), .ZN(
        n13251) );
  AND3_X1 U14897 ( .A1(n13986), .A2(n11514), .A3(n13251), .ZN(n13252) );
  AOI22_X1 U14898 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13254) );
  OR2_X1 U14899 ( .A1(n13417), .A2(n12577), .ZN(n13253) );
  NAND2_X1 U14900 ( .A1(n13254), .A2(n13253), .ZN(n14472) );
  NOR2_X1 U14901 ( .A1(n14473), .A2(n14472), .ZN(n13255) );
  NAND2_X1 U14902 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13259) );
  AND2_X1 U14903 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13257) );
  AOI21_X1 U14904 ( .B1(n13273), .B2(P2_EAX_REG_3__SCAN_IN), .A(n13257), .ZN(
        n13258) );
  AND2_X1 U14905 ( .A1(n13259), .A2(n13258), .ZN(n13262) );
  NAND2_X1 U14906 ( .A1(n13375), .A2(n13260), .ZN(n13261) );
  OAI211_X1 U14907 ( .C1(n13417), .C2(n13263), .A(n13262), .B(n13261), .ZN(
        n14468) );
  NAND2_X1 U14908 ( .A1(n14469), .A2(n14468), .ZN(n14470) );
  NAND2_X1 U14909 ( .A1(n14835), .A2(n14834), .ZN(n13266) );
  NAND2_X1 U14910 ( .A1(n13375), .A2(n13264), .ZN(n13265) );
  INV_X1 U14911 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n18372) );
  NAND2_X1 U14912 ( .A1(n13273), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U14913 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13267) );
  OAI211_X1 U14914 ( .C1(n13417), .C2(n18372), .A(n13268), .B(n13267), .ZN(
        n14079) );
  NAND2_X1 U14915 ( .A1(n14078), .A2(n14079), .ZN(n13270) );
  NAND2_X1 U14916 ( .A1(n13375), .A2(n12969), .ZN(n13269) );
  NAND2_X1 U14917 ( .A1(n13270), .A2(n13269), .ZN(n14081) );
  AOI22_X1 U14918 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13272) );
  OR2_X1 U14919 ( .A1(n13417), .A2(n13095), .ZN(n13271) );
  NAND2_X1 U14920 ( .A1(n13272), .A2(n13271), .ZN(n14080) );
  NAND2_X1 U14921 ( .A1(n14081), .A2(n14080), .ZN(n14083) );
  AOI22_X1 U14922 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U14923 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U14924 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U14925 ( .A1(n13274), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13276) );
  AOI22_X1 U14926 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13275) );
  NAND4_X1 U14927 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13284) );
  AOI22_X1 U14928 ( .A1(n12834), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U14929 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12656), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U14930 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U14931 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12673), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13279) );
  NAND4_X1 U14932 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  NAND2_X1 U14933 ( .A1(n13375), .A2(n14229), .ZN(n13286) );
  OR2_X1 U14934 ( .A1(n13417), .A2(n18601), .ZN(n13285) );
  AOI22_X1 U14935 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U14936 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12684), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13291) );
  AOI22_X1 U14937 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13290) );
  AOI22_X1 U14938 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U14939 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13288) );
  NAND4_X1 U14940 ( .A1(n13291), .A2(n13290), .A3(n13289), .A4(n13288), .ZN(
        n13297) );
  AOI22_X1 U14941 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15414), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U14942 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n13274), .B1(
        n12699), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U14943 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U14944 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13292) );
  NAND4_X1 U14945 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        n13296) );
  NAND2_X1 U14946 ( .A1(n13375), .A2(n14261), .ZN(n13298) );
  OAI211_X1 U14947 ( .C1(n13417), .C2(n18402), .A(n13299), .B(n13298), .ZN(
        n14076) );
  AOI22_X1 U14948 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U14949 ( .A1(n15414), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U14950 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U14951 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U14952 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13300) );
  NAND4_X1 U14953 ( .A1(n13303), .A2(n13302), .A3(n13301), .A4(n13300), .ZN(
        n13309) );
  AOI22_X1 U14954 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U14955 ( .A1(n13274), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12656), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U14956 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U14957 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13304) );
  NAND4_X1 U14958 ( .A1(n13307), .A2(n13306), .A3(n13305), .A4(n13304), .ZN(
        n13308) );
  NAND2_X1 U14959 ( .A1(n13375), .A2(n14422), .ZN(n13311) );
  NAND2_X1 U14960 ( .A1(n13410), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U14961 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U14962 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U14963 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U14964 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U14965 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13313) );
  NAND4_X1 U14966 ( .A1(n13316), .A2(n13315), .A3(n13314), .A4(n13313), .ZN(
        n13322) );
  AOI22_X1 U14967 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13320) );
  AOI22_X1 U14968 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U14969 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U14970 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13317) );
  NAND4_X1 U14971 ( .A1(n13320), .A2(n13319), .A3(n13318), .A4(n13317), .ZN(
        n13321) );
  NAND2_X1 U14972 ( .A1(n13375), .A2(n14462), .ZN(n13324) );
  NAND2_X1 U14973 ( .A1(n13410), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U14974 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n15414), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U14975 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U14976 ( .A1(n13274), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13327) );
  AOI22_X1 U14977 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13326) );
  NAND4_X1 U14978 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n13335) );
  AOI22_X1 U14979 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12684), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13333) );
  AOI22_X1 U14980 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12656), .B1(
        n12699), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U14981 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12661), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13331) );
  AOI22_X1 U14982 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12672), .B1(
        n12673), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13330) );
  NAND4_X1 U14983 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        n13334) );
  INV_X1 U14984 ( .A(n13375), .ZN(n13338) );
  AOI22_X1 U14985 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13337) );
  NAND2_X1 U14986 ( .A1(n13410), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n13336) );
  OAI211_X1 U14987 ( .C1(n14509), .C2(n13338), .A(n13337), .B(n13336), .ZN(
        n14179) );
  AND2_X2 U14988 ( .A1(n16893), .A2(n14179), .ZN(n14220) );
  AOI22_X1 U14989 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U14990 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U14991 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U14992 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U14993 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13339) );
  NAND4_X1 U14994 ( .A1(n13342), .A2(n13341), .A3(n13340), .A4(n13339), .ZN(
        n13348) );
  AOI22_X1 U14995 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U14996 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U14997 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U14998 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13343) );
  NAND4_X1 U14999 ( .A1(n13346), .A2(n13345), .A3(n13344), .A4(n13343), .ZN(
        n13347) );
  NAND2_X1 U15000 ( .A1(n13375), .A2(n14548), .ZN(n13349) );
  OAI211_X1 U15001 ( .C1(n13417), .C2(n13351), .A(n13350), .B(n13349), .ZN(
        n14219) );
  AOI22_X1 U15002 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U15003 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12834), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13355) );
  AOI22_X1 U15004 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13354) );
  AOI22_X1 U15005 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n15409), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U15006 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13352) );
  NAND4_X1 U15007 ( .A1(n13355), .A2(n13354), .A3(n13353), .A4(n13352), .ZN(
        n13361) );
  AOI22_X1 U15008 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n15414), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U15009 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13358) );
  AOI22_X1 U15010 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12661), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13357) );
  AOI22_X1 U15011 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12672), .B1(
        n12673), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13356) );
  NAND4_X1 U15012 ( .A1(n13359), .A2(n13358), .A3(n13357), .A4(n13356), .ZN(
        n13360) );
  NAND2_X1 U15013 ( .A1(n13375), .A2(n14656), .ZN(n13363) );
  NAND2_X1 U15014 ( .A1(n13410), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U15015 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U15016 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U15017 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12743), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U15018 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12835), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U15019 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13365) );
  NAND4_X1 U15020 ( .A1(n13368), .A2(n13367), .A3(n13366), .A4(n13365), .ZN(
        n13374) );
  AOI22_X1 U15021 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12725), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U15022 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U15023 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U15024 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13369) );
  NAND4_X1 U15025 ( .A1(n13372), .A2(n13371), .A3(n13370), .A4(n13369), .ZN(
        n13373) );
  NAND2_X1 U15026 ( .A1(n13375), .A2(n14686), .ZN(n13377) );
  NAND2_X1 U15027 ( .A1(n13410), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U15028 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U15029 ( .A1(n13410), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n13380) );
  NAND2_X1 U15030 ( .A1(n13381), .A2(n13380), .ZN(n16822) );
  NOR2_X1 U15031 ( .A1(n13417), .A2(n16535), .ZN(n13383) );
  INV_X1 U15032 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13933) );
  OAI22_X1 U15033 ( .A1(n13391), .A2(n16816), .B1(n13390), .B2(n13933), .ZN(
        n13382) );
  OR2_X1 U15034 ( .A1(n13383), .A2(n13382), .ZN(n16381) );
  NAND2_X1 U15035 ( .A1(n16380), .A2(n16381), .ZN(n16791) );
  AOI22_X1 U15036 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13385) );
  NAND2_X1 U15037 ( .A1(n13410), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n13384) );
  OR2_X2 U15038 ( .A1(n16791), .A2(n16790), .ZN(n16793) );
  AOI22_X1 U15039 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U15040 ( .A1(n13410), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13386) );
  NOR2_X4 U15041 ( .A1(n16793), .A2(n16370), .ZN(n16766) );
  AOI22_X1 U15042 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U15043 ( .A1(n13410), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U15044 ( .A1(n13389), .A2(n13388), .ZN(n16765) );
  NOR2_X1 U15045 ( .A1(n13417), .A2(n18513), .ZN(n13393) );
  INV_X1 U15046 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16363) );
  OAI22_X1 U15047 ( .A1(n13391), .A2(n16494), .B1(n13390), .B2(n16363), .ZN(
        n13392) );
  OR2_X1 U15048 ( .A1(n13393), .A2(n13392), .ZN(n16361) );
  AOI22_X1 U15049 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U15050 ( .A1(n13410), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13394) );
  AND2_X1 U15051 ( .A1(n13395), .A2(n13394), .ZN(n16726) );
  AOI22_X1 U15052 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13397) );
  NAND2_X1 U15053 ( .A1(n13410), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n13396) );
  AND2_X1 U15054 ( .A1(n13397), .A2(n13396), .ZN(n16223) );
  AOI22_X1 U15055 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13399) );
  NAND2_X1 U15056 ( .A1(n13410), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15057 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n13218), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13401) );
  NAND2_X1 U15058 ( .A1(n13410), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n13400) );
  NAND2_X1 U15059 ( .A1(n13401), .A2(n13400), .ZN(n16332) );
  NAND2_X1 U15060 ( .A1(n16333), .A2(n16332), .ZN(n16335) );
  AOI22_X1 U15061 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n13218), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n13403) );
  NAND2_X1 U15062 ( .A1(n13410), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13402) );
  AND2_X1 U15063 ( .A1(n13403), .A2(n13402), .ZN(n16189) );
  AOI22_X1 U15064 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U15065 ( .A1(n13410), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U15066 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13407) );
  NAND2_X1 U15067 ( .A1(n13410), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n13406) );
  NAND2_X1 U15068 ( .A1(n13407), .A2(n13406), .ZN(n16161) );
  AOI22_X1 U15069 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U15070 ( .A1(n13410), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U15071 ( .A1(n13409), .A2(n13408), .ZN(n15509) );
  AOI22_X1 U15072 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n13273), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U15073 ( .A1(n13410), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U15074 ( .A1(n13412), .A2(n13411), .ZN(n13451) );
  INV_X1 U15075 ( .A(n13451), .ZN(n13413) );
  NAND2_X1 U15076 ( .A1(n13379), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13415) );
  NAND2_X1 U15077 ( .A1(n13218), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n13414) );
  OAI211_X1 U15078 ( .C1(n13417), .C2(n13416), .A(n13415), .B(n13414), .ZN(
        n13418) );
  INV_X1 U15079 ( .A(n14337), .ZN(n14321) );
  INV_X1 U15080 ( .A(n13180), .ZN(n13421) );
  AND2_X1 U15081 ( .A1(n13421), .A2(n13420), .ZN(n14320) );
  AOI21_X1 U15082 ( .B1(n14321), .B2(n18335), .A(n14320), .ZN(n13422) );
  NAND2_X1 U15083 ( .A1(n19110), .A2(n18628), .ZN(n13424) );
  OAI211_X1 U15084 ( .C1(n16104), .C2(n18607), .A(n13425), .B(n13424), .ZN(
        n13426) );
  AOI21_X1 U15085 ( .B1(n13441), .B2(n18623), .A(n13426), .ZN(n13427) );
  NAND2_X1 U15086 ( .A1(n13428), .A2(n13427), .ZN(P2_U3015) );
  INV_X1 U15087 ( .A(n14325), .ZN(n13429) );
  NAND2_X1 U15088 ( .A1(n18645), .A2(n13429), .ZN(n13431) );
  NAND2_X1 U15089 ( .A1(n13431), .A2(n13430), .ZN(n14333) );
  OR2_X1 U15090 ( .A1(n13432), .A2(n17295), .ZN(n13443) );
  NAND2_X1 U15091 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17303) );
  NAND2_X1 U15092 ( .A1(n19262), .A2(n17303), .ZN(n18344) );
  OR2_X1 U15093 ( .A1(n18344), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13433) );
  AND2_X1 U15094 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17000) );
  INV_X1 U15095 ( .A(n14022), .ZN(n14349) );
  NAND2_X1 U15096 ( .A1(n21569), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U15097 ( .A1(n14349), .A2(n13434), .ZN(n13751) );
  INV_X1 U15098 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16641) );
  INV_X1 U15099 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U15100 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14629) );
  NOR2_X2 U15101 ( .A1(n17269), .A2(n14629), .ZN(n14702) );
  NAND2_X1 U15102 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n14702), .ZN(
        n14701) );
  NOR2_X2 U15103 ( .A1(n16641), .A2(n14703), .ZN(n14706) );
  NOR2_X2 U15104 ( .A1(n16116), .A2(n16511), .ZN(n16118) );
  INV_X1 U15105 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16121) );
  NOR2_X2 U15106 ( .A1(n16124), .A2(n16457), .ZN(n16125) );
  INV_X1 U15107 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16128) );
  NOR2_X2 U15108 ( .A1(n16132), .A2(n18565), .ZN(n16105) );
  NAND2_X1 U15109 ( .A1(n16105), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13436) );
  NOR2_X1 U15110 ( .A1(n17301), .A2(n14625), .ZN(n13437) );
  AOI211_X1 U15111 ( .C1(n17286), .C2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13438), .B(n13437), .ZN(n13439) );
  OAI21_X1 U15112 ( .B1(n16104), .B2(n17296), .A(n13439), .ZN(n13440) );
  AOI21_X1 U15113 ( .B1(n13441), .B2(n17270), .A(n13440), .ZN(n13442) );
  NAND2_X1 U15114 ( .A1(n13443), .A2(n13442), .ZN(P2_U2983) );
  NAND2_X1 U15115 ( .A1(n13444), .A2(n15502), .ZN(n13449) );
  INV_X1 U15116 ( .A(n13445), .ZN(n13446) );
  NOR2_X1 U15117 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  XNOR2_X1 U15118 ( .A(n13449), .B(n13448), .ZN(n13467) );
  XNOR2_X1 U15119 ( .A(n15513), .B(n13450), .ZN(n16152) );
  XOR2_X1 U15120 ( .A(n13451), .B(n15511), .Z(n16149) );
  NOR2_X1 U15121 ( .A1(n15515), .A2(n13452), .ZN(n13454) );
  OAI21_X1 U15122 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13454), .A(
        n13453), .ZN(n13455) );
  NAND2_X1 U15123 ( .A1(n18427), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13461) );
  OAI211_X1 U15124 ( .C1(n16149), .C2(n18603), .A(n13455), .B(n13461), .ZN(
        n13456) );
  XNOR2_X1 U15125 ( .A(n15507), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13459) );
  OAI211_X1 U15126 ( .C1(n13467), .C2(n18614), .A(n11515), .B(n11513), .ZN(
        P2_U3016) );
  NOR2_X1 U15127 ( .A1(n13459), .A2(n17294), .ZN(n13466) );
  XNOR2_X1 U15128 ( .A(n16105), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16144) );
  NAND2_X1 U15129 ( .A1(n17286), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13460) );
  OAI211_X1 U15130 ( .C1(n17301), .C2(n16144), .A(n13461), .B(n13460), .ZN(
        n13462) );
  INV_X1 U15131 ( .A(n13462), .ZN(n13463) );
  INV_X1 U15132 ( .A(n13467), .ZN(n13468) );
  NAND2_X1 U15133 ( .A1(n13470), .A2(n13469), .ZN(P2_U2984) );
  NAND3_X1 U15134 ( .A1(n11213), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17057) );
  INV_X1 U15135 ( .A(n17057), .ZN(n13471) );
  NAND2_X1 U15136 ( .A1(n13472), .A2(n22037), .ZN(n13473) );
  NAND2_X1 U15137 ( .A1(n11078), .A2(n13473), .ZN(n13803) );
  NOR2_X1 U15138 ( .A1(n13803), .A2(n11648), .ZN(n13475) );
  NAND2_X1 U15139 ( .A1(n16089), .A2(n21667), .ZN(n13474) );
  NAND2_X1 U15140 ( .A1(n13475), .A2(n13474), .ZN(n13789) );
  INV_X1 U15141 ( .A(n21852), .ZN(n21850) );
  NAND2_X1 U15142 ( .A1(n21850), .A2(n13480), .ZN(n21228) );
  NAND2_X1 U15143 ( .A1(n21228), .A2(n11213), .ZN(n13476) );
  NAND2_X1 U15144 ( .A1(n11213), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17049) );
  NAND2_X1 U15145 ( .A1(n21829), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U15146 ( .A1(n17049), .A2(n13477), .ZN(n14009) );
  INV_X1 U15147 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15873) );
  XNOR2_X1 U15148 ( .A(n13479), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14379) );
  INV_X1 U15149 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n19839) );
  NOR2_X1 U15150 ( .A1(n21401), .A2(n19839), .ZN(n15990) );
  AOI21_X1 U15151 ( .B1(n19943), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15990), .ZN(n13481) );
  OAI21_X1 U15152 ( .B1(n19952), .B2(n14379), .A(n13481), .ZN(n13482) );
  AOI21_X1 U15153 ( .B1(n15549), .B2(n19948), .A(n13482), .ZN(n13594) );
  AND2_X1 U15154 ( .A1(n21667), .A2(n21946), .ZN(n13501) );
  AOI21_X1 U15155 ( .B1(n13486), .B2(n14114), .A(n13501), .ZN(n13483) );
  XNOR2_X1 U15156 ( .A(n13486), .B(n13497), .ZN(n13487) );
  NAND2_X1 U15157 ( .A1(n13487), .A2(n14114), .ZN(n13489) );
  AND3_X1 U15158 ( .A1(n13489), .A2(n13488), .A3(n22037), .ZN(n13490) );
  NAND2_X1 U15159 ( .A1(n13491), .A2(n13490), .ZN(n13492) );
  NAND2_X1 U15160 ( .A1(n13940), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13495) );
  INV_X1 U15161 ( .A(n13492), .ZN(n13493) );
  OR2_X1 U15162 ( .A1(n14008), .A2(n13493), .ZN(n13494) );
  NAND2_X1 U15163 ( .A1(n13495), .A2(n13494), .ZN(n13505) );
  INV_X1 U15164 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14209) );
  XNOR2_X1 U15165 ( .A(n13505), .B(n14209), .ZN(n14044) );
  NAND2_X1 U15166 ( .A1(n21752), .A2(n13786), .ZN(n13504) );
  INV_X1 U15167 ( .A(n13496), .ZN(n13500) );
  NAND2_X1 U15168 ( .A1(n13498), .A2(n13497), .ZN(n13499) );
  NAND2_X1 U15169 ( .A1(n13499), .A2(n13500), .ZN(n13516) );
  OAI21_X1 U15170 ( .B1(n13500), .B2(n13499), .A(n13516), .ZN(n13502) );
  AOI21_X1 U15171 ( .B1(n13502), .B2(n14114), .A(n13501), .ZN(n13503) );
  NAND2_X1 U15172 ( .A1(n13504), .A2(n13503), .ZN(n14043) );
  NAND2_X1 U15173 ( .A1(n14044), .A2(n14043), .ZN(n13507) );
  NAND2_X1 U15174 ( .A1(n13505), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13506) );
  NAND2_X1 U15175 ( .A1(n13507), .A2(n13506), .ZN(n13511) );
  INV_X1 U15176 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14211) );
  XNOR2_X1 U15177 ( .A(n13511), .B(n14211), .ZN(n14203) );
  INV_X1 U15178 ( .A(n14114), .ZN(n21232) );
  XNOR2_X1 U15179 ( .A(n13516), .B(n13515), .ZN(n13509) );
  OAI22_X1 U15180 ( .A1(n13508), .A2(n13510), .B1(n21232), .B2(n13509), .ZN(
        n14202) );
  NAND2_X1 U15181 ( .A1(n14203), .A2(n14202), .ZN(n13513) );
  NAND2_X1 U15182 ( .A1(n13511), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13512) );
  NAND2_X1 U15183 ( .A1(n13513), .A2(n13512), .ZN(n14245) );
  NAND2_X1 U15184 ( .A1(n13514), .A2(n13786), .ZN(n13519) );
  NAND2_X1 U15185 ( .A1(n13516), .A2(n13515), .ZN(n13525) );
  XNOR2_X1 U15186 ( .A(n13525), .B(n13523), .ZN(n13517) );
  NAND2_X1 U15187 ( .A1(n13517), .A2(n14114), .ZN(n13518) );
  NAND2_X1 U15188 ( .A1(n13519), .A2(n13518), .ZN(n13520) );
  INV_X1 U15189 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14187) );
  XNOR2_X1 U15190 ( .A(n13520), .B(n14187), .ZN(n14244) );
  NAND2_X1 U15191 ( .A1(n13520), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13521) );
  NAND2_X1 U15192 ( .A1(n13522), .A2(n13786), .ZN(n13528) );
  INV_X1 U15193 ( .A(n13523), .ZN(n13524) );
  OR2_X1 U15194 ( .A1(n13525), .A2(n13524), .ZN(n13534) );
  XNOR2_X1 U15195 ( .A(n13534), .B(n13532), .ZN(n13526) );
  NAND2_X1 U15196 ( .A1(n13526), .A2(n14114), .ZN(n13527) );
  NAND2_X1 U15197 ( .A1(n13528), .A2(n13527), .ZN(n13529) );
  XNOR2_X1 U15198 ( .A(n13529), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19871) );
  INV_X1 U15199 ( .A(n13532), .ZN(n13533) );
  NOR2_X1 U15200 ( .A1(n13534), .A2(n13533), .ZN(n13536) );
  NAND2_X1 U15201 ( .A1(n13536), .A2(n13535), .ZN(n13553) );
  OAI211_X1 U15202 ( .C1(n13536), .C2(n13535), .A(n13553), .B(n14114), .ZN(
        n13537) );
  XNOR2_X1 U15203 ( .A(n13540), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14583) );
  NAND2_X1 U15204 ( .A1(n13540), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13541) );
  NAND2_X1 U15205 ( .A1(n13542), .A2(n13786), .ZN(n13545) );
  XNOR2_X1 U15206 ( .A(n13553), .B(n13551), .ZN(n13543) );
  NAND2_X1 U15207 ( .A1(n13543), .A2(n14114), .ZN(n13544) );
  NAND2_X1 U15208 ( .A1(n13545), .A2(n13544), .ZN(n13547) );
  INV_X1 U15209 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13546) );
  XNOR2_X1 U15210 ( .A(n13547), .B(n13546), .ZN(n19879) );
  NAND2_X2 U15211 ( .A1(n13550), .A2(n13549), .ZN(n13560) );
  NAND2_X1 U15212 ( .A1(n14114), .A2(n13551), .ZN(n13552) );
  OR2_X1 U15213 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  NAND2_X1 U15214 ( .A1(n19883), .A2(n13554), .ZN(n13557) );
  XNOR2_X1 U15215 ( .A(n13557), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14872) );
  INV_X1 U15216 ( .A(n14872), .ZN(n13555) );
  INV_X1 U15217 ( .A(n13557), .ZN(n13558) );
  INV_X1 U15218 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14484) );
  NAND2_X1 U15219 ( .A1(n13558), .A2(n14484), .ZN(n13559) );
  INV_X1 U15220 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14913) );
  XNOR2_X1 U15221 ( .A(n19945), .B(n14913), .ZN(n14900) );
  NAND2_X1 U15222 ( .A1(n19894), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13562) );
  INV_X1 U15223 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13569) );
  INV_X1 U15224 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13572) );
  INV_X1 U15225 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15552) );
  NAND3_X1 U15226 ( .A1(n13569), .A2(n13572), .A3(n15552), .ZN(n13563) );
  NAND2_X1 U15227 ( .A1(n19894), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19910) );
  INV_X1 U15228 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21254) );
  NAND2_X1 U15229 ( .A1(n19883), .A2(n21254), .ZN(n13564) );
  NAND2_X1 U15230 ( .A1(n19910), .A2(n13564), .ZN(n15967) );
  INV_X1 U15231 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21255) );
  NOR2_X1 U15232 ( .A1(n15967), .A2(n15966), .ZN(n19908) );
  NAND3_X1 U15233 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U15234 ( .A1(n19883), .A2(n13565), .ZN(n13566) );
  NAND2_X1 U15235 ( .A1(n19908), .A2(n13566), .ZN(n19918) );
  NAND2_X1 U15236 ( .A1(n19894), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13567) );
  NAND2_X1 U15237 ( .A1(n19910), .A2(n13567), .ZN(n13574) );
  NOR2_X1 U15238 ( .A1(n19883), .A2(n13569), .ZN(n19921) );
  NOR2_X1 U15239 ( .A1(n13574), .A2(n19921), .ZN(n15953) );
  NAND2_X1 U15240 ( .A1(n19918), .A2(n15953), .ZN(n13571) );
  NAND2_X1 U15241 ( .A1(n19894), .A2(n15552), .ZN(n15955) );
  NAND2_X1 U15242 ( .A1(n19883), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13568) );
  NAND2_X1 U15243 ( .A1(n15955), .A2(n13568), .ZN(n19932) );
  NAND2_X1 U15244 ( .A1(n19883), .A2(n13569), .ZN(n19930) );
  AND2_X1 U15245 ( .A1(n19932), .A2(n19930), .ZN(n13570) );
  NAND2_X1 U15246 ( .A1(n13571), .A2(n13570), .ZN(n15952) );
  NOR2_X1 U15247 ( .A1(n15952), .A2(n13572), .ZN(n13575) );
  NOR2_X1 U15248 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15963) );
  AND2_X1 U15249 ( .A1(n15963), .A2(n21255), .ZN(n13573) );
  NOR2_X1 U15250 ( .A1(n19883), .A2(n13573), .ZN(n15951) );
  NAND3_X1 U15251 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21378) );
  NAND2_X1 U15252 ( .A1(n13576), .A2(n19945), .ZN(n19944) );
  NOR2_X1 U15253 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13577) );
  INV_X1 U15254 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19936) );
  INV_X1 U15255 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15558) );
  NAND3_X1 U15256 ( .A1(n13577), .A2(n19936), .A3(n15558), .ZN(n13578) );
  AND3_X1 U15257 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15987) );
  NAND2_X1 U15258 ( .A1(n13580), .A2(n16043), .ZN(n13582) );
  AND2_X1 U15259 ( .A1(n15911), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13581) );
  NAND2_X1 U15260 ( .A1(n13582), .A2(n13581), .ZN(n13584) );
  INV_X1 U15261 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21404) );
  INV_X1 U15262 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16052) );
  INV_X1 U15263 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16066) );
  AND3_X1 U15264 ( .A1(n21404), .A2(n16052), .A3(n16066), .ZN(n15885) );
  NAND2_X1 U15265 ( .A1(n13583), .A2(n15941), .ZN(n15903) );
  INV_X1 U15266 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15887) );
  INV_X1 U15267 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16038) );
  NAND2_X1 U15268 ( .A1(n15887), .A2(n16038), .ZN(n16026) );
  NAND2_X1 U15269 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16025) );
  INV_X1 U15270 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16010) );
  AND2_X1 U15271 ( .A1(n19883), .A2(n16010), .ZN(n13585) );
  XNOR2_X1 U15272 ( .A(n19945), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13591) );
  INV_X1 U15273 ( .A(n13591), .ZN(n13587) );
  INV_X1 U15274 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16002) );
  AOI21_X1 U15275 ( .B1(n16002), .B2(n16010), .A(n19945), .ZN(n13589) );
  INV_X1 U15276 ( .A(n13589), .ZN(n13586) );
  NAND2_X1 U15277 ( .A1(n19883), .A2(n16002), .ZN(n13590) );
  INV_X1 U15278 ( .A(n13590), .ZN(n13588) );
  INV_X1 U15279 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15988) );
  OAI21_X1 U15280 ( .B1(n13589), .B2(n13588), .A(n15988), .ZN(n13592) );
  NAND2_X1 U15281 ( .A1(n13594), .A2(n13593), .ZN(P1_U2968) );
  NOR2_X1 U15282 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n13596) );
  NOR4_X1 U15283 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13595) );
  NAND4_X1 U15284 ( .A1(n13596), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n13595), .ZN(n13608) );
  NOR3_X1 U15285 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22244), .ZN(n13598) );
  NOR4_X1 U15286 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13597) );
  NAND4_X1 U15287 ( .A1(n21663), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n13598), .A4(
        n13597), .ZN(U214) );
  NOR4_X1 U15288 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13602) );
  NOR4_X1 U15289 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13601) );
  NOR4_X1 U15290 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13600) );
  NOR4_X1 U15291 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13599) );
  NAND4_X1 U15292 ( .A1(n13602), .A2(n13601), .A3(n13600), .A4(n13599), .ZN(
        n13607) );
  NOR4_X1 U15293 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13605) );
  NOR4_X1 U15294 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13604) );
  NOR4_X1 U15295 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13603) );
  NAND4_X1 U15296 ( .A1(n13605), .A2(n13604), .A3(n13603), .A4(n17375), .ZN(
        n13606) );
  OAI21_X4 U15297 ( .B1(n13607), .B2(n13606), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13649) );
  INV_X2 U15298 ( .A(U214), .ZN(n19993) );
  INV_X1 U15299 ( .A(n18345), .ZN(n18661) );
  INV_X1 U15300 ( .A(n13612), .ZN(n13610) );
  INV_X1 U15301 ( .A(n14332), .ZN(n13609) );
  NAND2_X1 U15302 ( .A1(n13610), .A2(n13609), .ZN(n16244) );
  NOR2_X1 U15303 ( .A1(n19276), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13613) );
  AOI211_X1 U15304 ( .C1(P2_MEMORYFETCH_REG_SCAN_IN), .C2(n16244), .A(n13613), 
        .B(n14635), .ZN(n13611) );
  INV_X1 U15305 ( .A(n13611), .ZN(P2_U2814) );
  INV_X1 U15306 ( .A(n16244), .ZN(n18358) );
  NOR4_X1 U15307 ( .A1(n18358), .A2(n14635), .A3(P2_READREQUEST_REG_SCAN_IN), 
        .A4(n13613), .ZN(n13614) );
  AOI21_X1 U15308 ( .B1(n18341), .B2(n13615), .A(n13614), .ZN(P2_U3612) );
  INV_X1 U15309 ( .A(n14635), .ZN(n13616) );
  INV_X1 U15310 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13618) );
  NAND3_X1 U15311 ( .A1(n14635), .A2(n18335), .A3(n18655), .ZN(n13754) );
  AOI22_X1 U15312 ( .A1(n15486), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13649), .ZN(n16365) );
  NOR2_X1 U15313 ( .A1(n13754), .A2(n16365), .ZN(n13722) );
  AOI21_X1 U15314 ( .B1(n13743), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13722), .ZN(
        n13617) );
  OAI21_X1 U15315 ( .B1(n13631), .B2(n13618), .A(n13617), .ZN(P2_U2957) );
  INV_X1 U15316 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13620) );
  AOI22_X1 U15317 ( .A1(n15486), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13649), .ZN(n19436) );
  NOR2_X1 U15318 ( .A1(n13754), .A2(n19436), .ZN(n13706) );
  AOI21_X1 U15319 ( .B1(n13743), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13706), .ZN(
        n13619) );
  OAI21_X1 U15320 ( .B1(n13631), .B2(n13620), .A(n13619), .ZN(P2_U2955) );
  INV_X1 U15321 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13622) );
  INV_X1 U15322 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n19967) );
  INV_X1 U15323 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20534) );
  AOI22_X1 U15324 ( .A1(n15486), .A2(n19967), .B1(n20534), .B2(n13649), .ZN(
        n19297) );
  INV_X1 U15325 ( .A(n19297), .ZN(n14754) );
  NOR2_X1 U15326 ( .A1(n13754), .A2(n14754), .ZN(n13725) );
  AOI21_X1 U15327 ( .B1(n13743), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13725), .ZN(
        n13621) );
  OAI21_X1 U15328 ( .B1(n13631), .B2(n13622), .A(n13621), .ZN(P2_U2958) );
  INV_X1 U15329 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13624) );
  INV_X1 U15330 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n19964) );
  INV_X1 U15331 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20543) );
  AOI22_X1 U15332 ( .A1(n15486), .A2(n19964), .B1(n20543), .B2(n13649), .ZN(
        n19393) );
  INV_X1 U15333 ( .A(n19393), .ZN(n14748) );
  NOR2_X1 U15334 ( .A1(n13754), .A2(n14748), .ZN(n13703) );
  AOI21_X1 U15335 ( .B1(n13743), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13703), .ZN(
        n13623) );
  OAI21_X1 U15336 ( .B1(n13631), .B2(n13624), .A(n13623), .ZN(P2_U2956) );
  INV_X1 U15337 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U15338 ( .A1(n15486), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13649), .ZN(n16352) );
  NOR2_X1 U15339 ( .A1(n13754), .A2(n16352), .ZN(n13731) );
  AOI21_X1 U15340 ( .B1(n13743), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13731), .ZN(
        n13625) );
  OAI21_X1 U15341 ( .B1(n13631), .B2(n13626), .A(n13625), .ZN(P2_U2959) );
  NAND2_X1 U15342 ( .A1(n21852), .A2(n21549), .ZN(n19955) );
  INV_X1 U15343 ( .A(n19955), .ZN(n14356) );
  INV_X1 U15344 ( .A(n13629), .ZN(n15540) );
  AND2_X1 U15345 ( .A1(n15538), .A2(n15540), .ZN(n15544) );
  INV_X1 U15346 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22245) );
  AOI21_X1 U15347 ( .B1(n15544), .B2(n14250), .A(n22245), .ZN(n13630) );
  OR3_X1 U15348 ( .A1(n13664), .A2(n14356), .A3(n13630), .ZN(P1_U2801) );
  INV_X1 U15349 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14144) );
  INV_X1 U15350 ( .A(n13631), .ZN(n13698) );
  NAND2_X1 U15351 ( .A1(n13698), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13634) );
  INV_X1 U15352 ( .A(n13754), .ZN(n13652) );
  INV_X1 U15353 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n19974) );
  OR2_X1 U15354 ( .A1(n13649), .A2(n19974), .ZN(n13633) );
  NAND2_X1 U15355 ( .A1(n13649), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13632) );
  NAND2_X1 U15356 ( .A1(n13633), .A2(n13632), .ZN(n19113) );
  NAND2_X1 U15357 ( .A1(n13652), .A2(n19113), .ZN(n13640) );
  OAI211_X1 U15358 ( .C1(n14633), .C2(n14144), .A(n13634), .B(n13640), .ZN(
        P2_U2963) );
  INV_X1 U15359 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14151) );
  NAND2_X1 U15360 ( .A1(n13698), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13637) );
  INV_X1 U15361 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n19972) );
  OR2_X1 U15362 ( .A1(n13649), .A2(n19972), .ZN(n13636) );
  NAND2_X1 U15363 ( .A1(n13649), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13635) );
  NAND2_X1 U15364 ( .A1(n13636), .A2(n13635), .ZN(n19116) );
  NAND2_X1 U15365 ( .A1(n13652), .A2(n19116), .ZN(n13638) );
  OAI211_X1 U15366 ( .C1(n14151), .C2(n14633), .A(n13637), .B(n13638), .ZN(
        P2_U2962) );
  INV_X1 U15367 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17360) );
  NAND2_X1 U15368 ( .A1(n13698), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13639) );
  OAI211_X1 U15369 ( .C1(n17360), .C2(n14633), .A(n13639), .B(n13638), .ZN(
        P2_U2977) );
  INV_X1 U15370 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17362) );
  NAND2_X1 U15371 ( .A1(n13698), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13641) );
  OAI211_X1 U15372 ( .C1(n17362), .C2(n14633), .A(n13641), .B(n13640), .ZN(
        P2_U2978) );
  INV_X1 U15373 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U15374 ( .A1(n13698), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13644) );
  INV_X1 U15375 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n19976) );
  OR2_X1 U15376 ( .A1(n13649), .A2(n19976), .ZN(n13643) );
  NAND2_X1 U15377 ( .A1(n13649), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13642) );
  NAND2_X1 U15378 ( .A1(n13643), .A2(n13642), .ZN(n16316) );
  NAND2_X1 U15379 ( .A1(n13652), .A2(n16316), .ZN(n13738) );
  OAI211_X1 U15380 ( .C1(n14633), .C2(n14139), .A(n13644), .B(n13738), .ZN(
        P2_U2964) );
  INV_X1 U15381 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14147) );
  NAND2_X1 U15382 ( .A1(n13698), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U15383 ( .A1(n15486), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13649), .ZN(n14222) );
  INV_X1 U15384 ( .A(n14222), .ZN(n16310) );
  NAND2_X1 U15385 ( .A1(n13652), .A2(n16310), .ZN(n13745) );
  OAI211_X1 U15386 ( .C1(n14633), .C2(n14147), .A(n13645), .B(n13745), .ZN(
        P2_U2965) );
  INV_X1 U15387 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U15388 ( .A1(n13698), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13648) );
  INV_X1 U15389 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n19979) );
  OR2_X1 U15390 ( .A1(n13649), .A2(n19979), .ZN(n13647) );
  NAND2_X1 U15391 ( .A1(n13649), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U15392 ( .A1(n13647), .A2(n13646), .ZN(n15490) );
  NAND2_X1 U15393 ( .A1(n13652), .A2(n15490), .ZN(n13741) );
  OAI211_X1 U15394 ( .C1(n14633), .C2(n14155), .A(n13648), .B(n13741), .ZN(
        P2_U2966) );
  INV_X1 U15395 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14137) );
  NAND2_X1 U15396 ( .A1(n13698), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13653) );
  INV_X1 U15397 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13661) );
  OR2_X1 U15398 ( .A1(n13649), .A2(n13661), .ZN(n13651) );
  NAND2_X1 U15399 ( .A1(n13649), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13650) );
  NAND2_X1 U15400 ( .A1(n13651), .A2(n13650), .ZN(n16336) );
  NAND2_X1 U15401 ( .A1(n13652), .A2(n16336), .ZN(n13735) );
  OAI211_X1 U15402 ( .C1(n14633), .C2(n14137), .A(n13653), .B(n13735), .ZN(
        P2_U2961) );
  NAND2_X1 U15403 ( .A1(n15546), .A2(n17021), .ZN(n13655) );
  NAND2_X1 U15404 ( .A1(n13655), .A2(n13654), .ZN(n13780) );
  NAND2_X1 U15405 ( .A1(n13780), .A2(n14250), .ZN(n13656) );
  INV_X1 U15406 ( .A(n21227), .ZN(n13658) );
  OAI21_X1 U15407 ( .B1(n14356), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13658), 
        .ZN(n13657) );
  OAI21_X1 U15408 ( .B1(n13659), .B2(n13658), .A(n13657), .ZN(P1_U3487) );
  INV_X1 U15409 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U15410 ( .A1(n14364), .A2(n21229), .ZN(n14088) );
  OR2_X1 U15411 ( .A1(n21662), .A2(n13661), .ZN(n13663) );
  NAND2_X1 U15412 ( .A1(n21662), .A2(DATAI_9_), .ZN(n13662) );
  NAND2_X1 U15413 ( .A1(n13663), .A2(n13662), .ZN(n14559) );
  NAND2_X1 U15414 ( .A1(n13934), .A2(n14559), .ZN(n13671) );
  OAI21_X4 U15415 ( .B1(n14114), .B2(n21229), .A(n13664), .ZN(n13922) );
  NAND2_X1 U15416 ( .A1(n13922), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13665) );
  OAI211_X1 U15417 ( .C1(n14565), .C2(n13884), .A(n13671), .B(n13665), .ZN(
        P1_U2946) );
  INV_X1 U15418 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13666) );
  OR2_X1 U15419 ( .A1(n21662), .A2(n13666), .ZN(n13668) );
  NAND2_X1 U15420 ( .A1(n21662), .A2(DATAI_8_), .ZN(n13667) );
  NAND2_X1 U15421 ( .A1(n13668), .A2(n13667), .ZN(n14501) );
  NAND2_X1 U15422 ( .A1(n13934), .A2(n14501), .ZN(n13870) );
  NAND2_X1 U15423 ( .A1(n13922), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13669) );
  OAI211_X1 U15424 ( .C1(n15836), .C2(n13884), .A(n13870), .B(n13669), .ZN(
        P1_U2945) );
  INV_X1 U15425 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19783) );
  NAND2_X1 U15426 ( .A1(n13922), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13670) );
  OAI211_X1 U15427 ( .C1(n19783), .C2(n13884), .A(n13671), .B(n13670), .ZN(
        P1_U2961) );
  OR2_X1 U15428 ( .A1(n21662), .A2(n19976), .ZN(n13673) );
  NAND2_X1 U15429 ( .A1(n21662), .A2(DATAI_12_), .ZN(n13672) );
  NAND2_X1 U15430 ( .A1(n13673), .A2(n13672), .ZN(n15025) );
  NAND2_X1 U15431 ( .A1(n13934), .A2(n15025), .ZN(n13909) );
  NAND2_X1 U15432 ( .A1(n13922), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n13674) );
  OAI211_X1 U15433 ( .C1(n15026), .C2(n13884), .A(n13909), .B(n13674), .ZN(
        P1_U2964) );
  INV_X1 U15434 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14576) );
  INV_X1 U15435 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13675) );
  OR2_X1 U15436 ( .A1(n21662), .A2(n13675), .ZN(n13677) );
  NAND2_X1 U15437 ( .A1(n21662), .A2(DATAI_5_), .ZN(n13676) );
  AND2_X1 U15438 ( .A1(n13677), .A2(n13676), .ZN(n22035) );
  INV_X1 U15439 ( .A(n22035), .ZN(n13678) );
  NAND2_X1 U15440 ( .A1(n13934), .A2(n13678), .ZN(n13861) );
  NAND2_X1 U15441 ( .A1(n13922), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13679) );
  OAI211_X1 U15442 ( .C1(n14576), .C2(n13884), .A(n13861), .B(n13679), .ZN(
        P1_U2942) );
  INV_X1 U15443 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13680) );
  OR2_X1 U15444 ( .A1(n21662), .A2(n13680), .ZN(n13682) );
  NAND2_X1 U15445 ( .A1(n21662), .A2(DATAI_13_), .ZN(n13681) );
  NAND2_X1 U15446 ( .A1(n13682), .A2(n13681), .ZN(n15000) );
  NAND2_X1 U15447 ( .A1(n13934), .A2(n15000), .ZN(n13911) );
  NAND2_X1 U15448 ( .A1(n13922), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13683) );
  OAI211_X1 U15449 ( .C1(n15001), .C2(n13884), .A(n13911), .B(n13683), .ZN(
        P1_U2965) );
  INV_X1 U15450 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19788) );
  OR2_X1 U15451 ( .A1(n21662), .A2(n19974), .ZN(n13685) );
  NAND2_X1 U15452 ( .A1(n21662), .A2(DATAI_11_), .ZN(n13684) );
  NAND2_X1 U15453 ( .A1(n13685), .A2(n13684), .ZN(n14968) );
  NAND2_X1 U15454 ( .A1(n13934), .A2(n14968), .ZN(n13921) );
  NAND2_X1 U15455 ( .A1(n13922), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13686) );
  OAI211_X1 U15456 ( .C1(n19788), .C2(n13884), .A(n13921), .B(n13686), .ZN(
        P1_U2963) );
  INV_X1 U15457 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14562) );
  INV_X1 U15458 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13687) );
  OR2_X1 U15459 ( .A1(n21662), .A2(n13687), .ZN(n13689) );
  NAND2_X1 U15460 ( .A1(n21662), .A2(DATAI_7_), .ZN(n13688) );
  AND2_X1 U15461 ( .A1(n13689), .A2(n13688), .ZN(n22128) );
  INV_X1 U15462 ( .A(n22128), .ZN(n13690) );
  NAND2_X1 U15463 ( .A1(n13934), .A2(n13690), .ZN(n13905) );
  NAND2_X1 U15464 ( .A1(n13922), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13691) );
  OAI211_X1 U15465 ( .C1(n14562), .C2(n13884), .A(n13905), .B(n13691), .ZN(
        P1_U2944) );
  INV_X1 U15466 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19786) );
  OR2_X1 U15467 ( .A1(n21662), .A2(n19972), .ZN(n13693) );
  NAND2_X1 U15468 ( .A1(n21662), .A2(DATAI_10_), .ZN(n13692) );
  NAND2_X1 U15469 ( .A1(n13693), .A2(n13692), .ZN(n14694) );
  NAND2_X1 U15470 ( .A1(n13934), .A2(n14694), .ZN(n13924) );
  NAND2_X1 U15471 ( .A1(n13922), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13694) );
  OAI211_X1 U15472 ( .C1(n19786), .C2(n13884), .A(n13924), .B(n13694), .ZN(
        P1_U2962) );
  INV_X1 U15473 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19792) );
  OR2_X1 U15474 ( .A1(n21662), .A2(n19979), .ZN(n13696) );
  NAND2_X1 U15475 ( .A1(n21662), .A2(DATAI_14_), .ZN(n13695) );
  NAND2_X1 U15476 ( .A1(n13696), .A2(n13695), .ZN(n15002) );
  NAND2_X1 U15477 ( .A1(n13934), .A2(n15002), .ZN(n13913) );
  NAND2_X1 U15478 ( .A1(n13922), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13697) );
  OAI211_X1 U15479 ( .C1(n19792), .C2(n13884), .A(n13913), .B(n13697), .ZN(
        P1_U2966) );
  INV_X1 U15480 ( .A(n13698), .ZN(n13756) );
  INV_X1 U15481 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13700) );
  OAI22_X1 U15482 ( .A1(n13649), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15486), .ZN(n19592) );
  NOR2_X1 U15483 ( .A1(n13754), .A2(n19592), .ZN(n13728) );
  AOI21_X1 U15484 ( .B1(n13743), .B2(P2_EAX_REG_0__SCAN_IN), .A(n13728), .ZN(
        n13699) );
  OAI21_X1 U15485 ( .B1(n13756), .B2(n13700), .A(n13699), .ZN(P2_U2967) );
  INV_X1 U15486 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13702) );
  OAI22_X1 U15487 ( .A1(n13649), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15486), .ZN(n19497) );
  NOR2_X1 U15488 ( .A1(n13754), .A2(n19497), .ZN(n13713) );
  AOI21_X1 U15489 ( .B1(n13743), .B2(P2_EAX_REG_2__SCAN_IN), .A(n13713), .ZN(
        n13701) );
  OAI21_X1 U15490 ( .B1(n13756), .B2(n13702), .A(n13701), .ZN(P2_U2969) );
  INV_X1 U15491 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13705) );
  AOI21_X1 U15492 ( .B1(n13743), .B2(P2_EAX_REG_4__SCAN_IN), .A(n13703), .ZN(
        n13704) );
  OAI21_X1 U15493 ( .B1(n13756), .B2(n13705), .A(n13704), .ZN(P2_U2971) );
  INV_X1 U15494 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13708) );
  AOI21_X1 U15495 ( .B1(n13743), .B2(P2_EAX_REG_3__SCAN_IN), .A(n13706), .ZN(
        n13707) );
  OAI21_X1 U15496 ( .B1(n13756), .B2(n13708), .A(n13707), .ZN(P2_U2970) );
  INV_X1 U15497 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13710) );
  AOI22_X1 U15498 ( .A1(n15486), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13649), .ZN(n14744) );
  NOR2_X1 U15499 ( .A1(n13754), .A2(n14744), .ZN(n13716) );
  AOI21_X1 U15500 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n13743), .A(n13716), .ZN(
        n13709) );
  OAI21_X1 U15501 ( .B1(n13756), .B2(n13710), .A(n13709), .ZN(P2_U2968) );
  INV_X1 U15502 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U15503 ( .A1(n15486), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13649), .ZN(n16347) );
  NOR2_X1 U15504 ( .A1(n13754), .A2(n16347), .ZN(n13719) );
  AOI21_X1 U15505 ( .B1(P2_EAX_REG_8__SCAN_IN), .B2(n13743), .A(n13719), .ZN(
        n13711) );
  OAI21_X1 U15506 ( .B1(n13756), .B2(n13712), .A(n13711), .ZN(P2_U2975) );
  INV_X1 U15507 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13715) );
  AOI21_X1 U15508 ( .B1(n13743), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13713), .ZN(
        n13714) );
  OAI21_X1 U15509 ( .B1(n13756), .B2(n13715), .A(n13714), .ZN(P2_U2954) );
  INV_X1 U15510 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13718) );
  AOI21_X1 U15511 ( .B1(n13743), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13716), .ZN(
        n13717) );
  OAI21_X1 U15512 ( .B1(n13756), .B2(n13718), .A(n13717), .ZN(P2_U2953) );
  INV_X1 U15513 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n13721) );
  AOI21_X1 U15514 ( .B1(n13743), .B2(P2_EAX_REG_24__SCAN_IN), .A(n13719), .ZN(
        n13720) );
  OAI21_X1 U15515 ( .B1(n13756), .B2(n13721), .A(n13720), .ZN(P2_U2960) );
  INV_X1 U15516 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13724) );
  AOI21_X1 U15517 ( .B1(n13743), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13722), .ZN(
        n13723) );
  OAI21_X1 U15518 ( .B1(n13756), .B2(n13724), .A(n13723), .ZN(P2_U2972) );
  INV_X1 U15519 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13727) );
  AOI21_X1 U15520 ( .B1(n13743), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13725), .ZN(
        n13726) );
  OAI21_X1 U15521 ( .B1(n13756), .B2(n13727), .A(n13726), .ZN(P2_U2973) );
  INV_X1 U15522 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13730) );
  AOI21_X1 U15523 ( .B1(n13743), .B2(P2_EAX_REG_16__SCAN_IN), .A(n13728), .ZN(
        n13729) );
  OAI21_X1 U15524 ( .B1(n13756), .B2(n13730), .A(n13729), .ZN(P2_U2952) );
  INV_X1 U15525 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13733) );
  AOI21_X1 U15526 ( .B1(n13743), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13731), .ZN(
        n13732) );
  OAI21_X1 U15527 ( .B1(n13756), .B2(n13733), .A(n13732), .ZN(P2_U2974) );
  INV_X1 U15528 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U15529 ( .A1(n13743), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n13734) );
  OAI211_X1 U15530 ( .C1(n13756), .C2(n13736), .A(n13735), .B(n13734), .ZN(
        P2_U2976) );
  INV_X1 U15531 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n13739) );
  NAND2_X1 U15532 ( .A1(n13743), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n13737) );
  OAI211_X1 U15533 ( .C1(n13756), .C2(n13739), .A(n13738), .B(n13737), .ZN(
        P2_U2979) );
  INV_X1 U15534 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n13742) );
  NAND2_X1 U15535 ( .A1(n13743), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n13740) );
  OAI211_X1 U15536 ( .C1(n13756), .C2(n13742), .A(n13741), .B(n13740), .ZN(
        P2_U2981) );
  INV_X1 U15537 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13746) );
  NAND2_X1 U15538 ( .A1(n13743), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13744) );
  OAI211_X1 U15539 ( .C1(n13756), .C2(n13746), .A(n13745), .B(n13744), .ZN(
        P2_U2980) );
  XNOR2_X1 U15540 ( .A(n18351), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18584) );
  INV_X1 U15541 ( .A(n18584), .ZN(n13750) );
  NOR2_X1 U15542 ( .A1(n18600), .A2(n12555), .ZN(n18589) );
  OAI21_X1 U15543 ( .B1(n13748), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13747), .ZN(n18586) );
  NOR2_X1 U15544 ( .A1(n17294), .A2(n18586), .ZN(n13749) );
  AOI211_X1 U15545 ( .C1(n17274), .C2(n13750), .A(n18589), .B(n13749), .ZN(
        n13753) );
  OAI21_X1 U15546 ( .B1(n17286), .B2(n13751), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13752) );
  OAI211_X1 U15547 ( .C1(n17296), .C2(n18587), .A(n13753), .B(n13752), .ZN(
        P2_U3014) );
  INV_X1 U15548 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13755) );
  AOI22_X1 U15549 ( .A1(n15486), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13649), .ZN(n14467) );
  INV_X1 U15550 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17372) );
  OAI222_X1 U15551 ( .A1(n13756), .A2(n13755), .B1(n13754), .B2(n14467), .C1(
        n14633), .C2(n17372), .ZN(P2_U2982) );
  NAND2_X1 U15552 ( .A1(n12532), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13757) );
  NOR2_X1 U15553 ( .A1(n19276), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13758) );
  AOI21_X1 U15554 ( .B1(n14019), .B2(n16959), .A(n13758), .ZN(n13759) );
  INV_X1 U15555 ( .A(n13761), .ZN(n13762) );
  INV_X1 U15556 ( .A(n19243), .ZN(n14299) );
  OAI21_X1 U15557 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n14299), .ZN(n19146) );
  NAND2_X1 U15558 ( .A1(n14019), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13763) );
  OAI21_X1 U15559 ( .B1(n19146), .B2(n19276), .A(n13763), .ZN(n13764) );
  NAND2_X1 U15560 ( .A1(n14591), .A2(n14320), .ZN(n14271) );
  INV_X1 U15561 ( .A(n14279), .ZN(n13768) );
  NAND2_X1 U15562 ( .A1(n14271), .A2(n13768), .ZN(n13769) );
  INV_X1 U15563 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13770) );
  MUX2_X1 U15564 ( .A(n13770), .B(n13995), .S(n16284), .Z(n13771) );
  OAI21_X1 U15565 ( .B1(n17320), .B2(n16302), .A(n13771), .ZN(P2_U2886) );
  AND2_X1 U15566 ( .A1(n19262), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13773) );
  OAI211_X1 U15567 ( .C1(n15436), .C2(n19708), .A(n15487), .B(n13773), .ZN(
        n13774) );
  MUX2_X1 U15568 ( .A(n13775), .B(n18587), .S(n16284), .Z(n13776) );
  OAI21_X1 U15569 ( .B1(n17305), .B2(n16302), .A(n13776), .ZN(P2_U2887) );
  INV_X1 U15570 ( .A(n21587), .ZN(n13778) );
  NAND2_X1 U15571 ( .A1(n13778), .A2(n21229), .ZN(n17050) );
  NAND2_X1 U15572 ( .A1(n13779), .A2(n17050), .ZN(n13784) );
  INV_X1 U15573 ( .A(n13780), .ZN(n13782) );
  NAND2_X1 U15574 ( .A1(n15546), .A2(n14115), .ZN(n13781) );
  NAND2_X1 U15575 ( .A1(n13782), .A2(n13781), .ZN(n13783) );
  NAND2_X1 U15576 ( .A1(n13784), .A2(n13783), .ZN(n13797) );
  NOR2_X1 U15577 ( .A1(n13874), .A2(n13878), .ZN(n15535) );
  INV_X1 U15578 ( .A(n15535), .ZN(n13794) );
  AOI21_X1 U15579 ( .B1(n13786), .B2(n11656), .A(n21667), .ZN(n13787) );
  AND2_X1 U15580 ( .A1(n13788), .A2(n13787), .ZN(n13811) );
  NOR2_X1 U15581 ( .A1(n13789), .A2(n13811), .ZN(n13790) );
  OR2_X1 U15582 ( .A1(n15538), .A2(n13790), .ZN(n14096) );
  OAI21_X1 U15583 ( .B1(n13805), .B2(n14093), .A(n14096), .ZN(n13791) );
  INV_X1 U15584 ( .A(n13791), .ZN(n13792) );
  OAI211_X1 U15585 ( .C1(n15546), .C2(n13794), .A(n13793), .B(n13792), .ZN(
        n13795) );
  INV_X1 U15586 ( .A(n13795), .ZN(n13796) );
  NAND2_X1 U15587 ( .A1(n17044), .A2(n14250), .ZN(n13801) );
  INV_X1 U15588 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21547) );
  NAND2_X1 U15589 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16083), .ZN(n21552) );
  NOR2_X1 U15590 ( .A1(n21547), .A2(n21552), .ZN(n13799) );
  INV_X1 U15591 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21805) );
  NOR2_X1 U15592 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21805), .ZN(n13798) );
  NOR2_X1 U15593 ( .A1(n13799), .A2(n13798), .ZN(n13800) );
  NAND2_X1 U15594 ( .A1(n13801), .A2(n13800), .ZN(n16984) );
  NAND2_X1 U15595 ( .A1(n13803), .A2(n10968), .ZN(n13810) );
  INV_X1 U15596 ( .A(n14093), .ZN(n21902) );
  OAI21_X1 U15597 ( .B1(n21902), .B2(n11630), .A(n14164), .ZN(n13804) );
  OAI21_X1 U15598 ( .B1(n13804), .B2(n13839), .A(n14364), .ZN(n13809) );
  NAND2_X1 U15599 ( .A1(n11648), .A2(n11645), .ZN(n13808) );
  INV_X1 U15600 ( .A(n13805), .ZN(n14371) );
  NAND2_X1 U15601 ( .A1(n13806), .A2(n14371), .ZN(n13807) );
  NAND4_X1 U15602 ( .A1(n13810), .A2(n13809), .A3(n13808), .A4(n13807), .ZN(
        n13812) );
  NOR2_X1 U15603 ( .A1(n13812), .A2(n13811), .ZN(n13814) );
  AND2_X1 U15604 ( .A1(n13814), .A2(n13813), .ZN(n14107) );
  NAND2_X1 U15605 ( .A1(n13815), .A2(n14108), .ZN(n13816) );
  NOR2_X1 U15606 ( .A1(n14115), .A2(n13816), .ZN(n13817) );
  AND3_X1 U15607 ( .A1(n12382), .A2(n14107), .A3(n13817), .ZN(n16090) );
  NOR2_X1 U15608 ( .A1(n13818), .A2(n13833), .ZN(n13821) );
  NOR2_X1 U15609 ( .A1(n14371), .A2(n14114), .ZN(n15547) );
  INV_X1 U15610 ( .A(n15547), .ZN(n13819) );
  NOR2_X1 U15611 ( .A1(n13874), .A2(n13819), .ZN(n13832) );
  XNOR2_X1 U15612 ( .A(n16097), .B(n13830), .ZN(n13824) );
  INV_X1 U15613 ( .A(n13824), .ZN(n13820) );
  AOI22_X1 U15614 ( .A1(n17021), .A2(n13821), .B1(n13832), .B2(n13820), .ZN(
        n13823) );
  NAND3_X1 U15615 ( .A1(n16090), .A2(n13839), .A3(n13824), .ZN(n13822) );
  OAI211_X1 U15616 ( .C1(n13802), .C2(n16090), .A(n13823), .B(n13822), .ZN(
        n17018) );
  INV_X1 U15617 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14119) );
  NOR2_X1 U15618 ( .A1(n21549), .A2(n14119), .ZN(n16100) );
  INV_X1 U15619 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14208) );
  OAI22_X1 U15620 ( .A1(n14208), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n15988), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16095) );
  INV_X1 U15621 ( .A(n16096), .ZN(n21555) );
  AOI222_X1 U15622 ( .A1(n17018), .A2(n16094), .B1(n16100), .B2(n16095), .C1(
        n21555), .C2(n13824), .ZN(n13826) );
  NAND2_X1 U15623 ( .A1(n16982), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13825) );
  OAI21_X1 U15624 ( .B1(n16982), .B2(n13826), .A(n13825), .ZN(P1_U3472) );
  INV_X1 U15625 ( .A(n16090), .ZN(n13828) );
  NAND2_X1 U15626 ( .A1(n21753), .A2(n13828), .ZN(n13845) );
  INV_X1 U15627 ( .A(n13833), .ZN(n13829) );
  NAND2_X1 U15628 ( .A1(n17021), .A2(n13829), .ZN(n13835) );
  INV_X1 U15629 ( .A(n16097), .ZN(n13841) );
  NAND2_X1 U15630 ( .A1(n13841), .A2(n13830), .ZN(n13831) );
  AOI22_X1 U15631 ( .A1(n17021), .A2(n13833), .B1(n13832), .B2(n13831), .ZN(
        n13834) );
  MUX2_X1 U15632 ( .A(n13835), .B(n13834), .S(n11427), .Z(n13844) );
  NAND2_X1 U15633 ( .A1(n16097), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13836) );
  NAND2_X1 U15634 ( .A1(n13836), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13837) );
  NAND2_X1 U15635 ( .A1(n13838), .A2(n13837), .ZN(n13846) );
  NAND3_X1 U15636 ( .A1(n16090), .A2(n13839), .A3(n13846), .ZN(n13843) );
  NAND2_X1 U15637 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  NAND4_X1 U15638 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n17019) );
  AOI22_X1 U15639 ( .A1(n17019), .A2(n16094), .B1(n21555), .B2(n13846), .ZN(
        n13848) );
  NAND2_X1 U15640 ( .A1(n16982), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13847) );
  OAI21_X1 U15641 ( .B1(n16982), .B2(n13848), .A(n13847), .ZN(P1_U3469) );
  INV_X1 U15642 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13849) );
  MUX2_X1 U15643 ( .A(n17286), .B(n17260), .S(n13849), .Z(n13858) );
  AOI21_X1 U15644 ( .B1(n14628), .B2(n13851), .A(n13850), .ZN(n13997) );
  INV_X1 U15645 ( .A(n13997), .ZN(n13856) );
  NOR2_X1 U15646 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  XOR2_X1 U15647 ( .A(n13854), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13992) );
  NAND2_X1 U15648 ( .A1(n13992), .A2(n17274), .ZN(n13855) );
  NAND2_X1 U15649 ( .A1(n18427), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13998) );
  OAI211_X1 U15650 ( .C1(n17294), .C2(n13856), .A(n13855), .B(n13998), .ZN(
        n13857) );
  AOI211_X1 U15651 ( .C1(n17273), .C2(n16241), .A(n13858), .B(n13857), .ZN(
        n13859) );
  INV_X1 U15652 ( .A(n13859), .ZN(P2_U3013) );
  INV_X1 U15653 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19776) );
  NAND2_X1 U15654 ( .A1(n13922), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n13860) );
  OAI211_X1 U15655 ( .C1(n19776), .C2(n13884), .A(n13861), .B(n13860), .ZN(
        P1_U2957) );
  INV_X1 U15656 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13862) );
  OR2_X1 U15657 ( .A1(n21662), .A2(n13862), .ZN(n13864) );
  NAND2_X1 U15658 ( .A1(n21662), .A2(DATAI_2_), .ZN(n13863) );
  INV_X1 U15659 ( .A(n21900), .ZN(n21641) );
  NAND2_X1 U15660 ( .A1(n13934), .A2(n21641), .ZN(n13898) );
  NAND2_X1 U15661 ( .A1(n13922), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13865) );
  OAI211_X1 U15662 ( .C1(n12062), .C2(n13884), .A(n13898), .B(n13865), .ZN(
        P1_U2939) );
  INV_X1 U15663 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19774) );
  OR2_X1 U15664 ( .A1(n21662), .A2(n19964), .ZN(n13867) );
  NAND2_X1 U15665 ( .A1(n21662), .A2(DATAI_4_), .ZN(n13866) );
  AND2_X1 U15666 ( .A1(n13867), .A2(n13866), .ZN(n21989) );
  INV_X1 U15667 ( .A(n21989), .ZN(n21645) );
  NAND2_X1 U15668 ( .A1(n13934), .A2(n21645), .ZN(n13891) );
  NAND2_X1 U15669 ( .A1(n13922), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n13868) );
  OAI211_X1 U15670 ( .C1(n19774), .C2(n13884), .A(n13891), .B(n13868), .ZN(
        P1_U2956) );
  NAND2_X1 U15671 ( .A1(n13922), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13869) );
  OAI211_X1 U15672 ( .C1(n14502), .C2(n13884), .A(n13870), .B(n13869), .ZN(
        P1_U2960) );
  XNOR2_X1 U15673 ( .A(n13872), .B(n13871), .ZN(n14397) );
  OAI21_X1 U15674 ( .B1(n15546), .B2(n13874), .A(n13873), .ZN(n13876) );
  AND2_X2 U15675 ( .A1(n15588), .A2(n13785), .ZN(n15591) );
  INV_X1 U15676 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U15677 ( .A1(n15591), .A2(n13879), .ZN(n13881) );
  INV_X1 U15678 ( .A(n21946), .ZN(n13877) );
  NAND2_X1 U15679 ( .A1(n13877), .A2(n11645), .ZN(n14056) );
  NAND2_X1 U15680 ( .A1(n14056), .A2(n14208), .ZN(n13880) );
  NAND2_X1 U15681 ( .A1(n14056), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13882) );
  OAI21_X1 U15682 ( .B1(n10968), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13882), .ZN(
        n14072) );
  XNOR2_X1 U15683 ( .A(n14053), .B(n14072), .ZN(n14055) );
  XNOR2_X1 U15684 ( .A(n14055), .B(n13785), .ZN(n14394) );
  AOI22_X1 U15685 ( .A1(n19865), .A2(n14394), .B1(n15794), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13883) );
  OAI21_X1 U15686 ( .B1(n14397), .B2(n15796), .A(n13883), .ZN(P1_U2871) );
  OR2_X1 U15687 ( .A1(n21662), .A2(n19967), .ZN(n13886) );
  NAND2_X1 U15688 ( .A1(n21662), .A2(DATAI_6_), .ZN(n13885) );
  AND2_X1 U15689 ( .A1(n13886), .A2(n13885), .ZN(n22083) );
  INV_X1 U15690 ( .A(n22083), .ZN(n21650) );
  NAND2_X1 U15691 ( .A1(n13934), .A2(n21650), .ZN(n13889) );
  NAND2_X1 U15692 ( .A1(n13922), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n13887) );
  OAI211_X1 U15693 ( .C1(n13884), .C2(n19778), .A(n13889), .B(n13887), .ZN(
        P1_U2958) );
  NAND2_X1 U15694 ( .A1(n13922), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13888) );
  OAI211_X1 U15695 ( .C1(n13884), .C2(n14573), .A(n13889), .B(n13888), .ZN(
        P1_U2943) );
  INV_X1 U15696 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14579) );
  NAND2_X1 U15697 ( .A1(n13922), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13890) );
  OAI211_X1 U15698 ( .C1(n13884), .C2(n14579), .A(n13891), .B(n13890), .ZN(
        P1_U2941) );
  INV_X1 U15699 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13892) );
  OR2_X1 U15700 ( .A1(n21662), .A2(n13892), .ZN(n13894) );
  NAND2_X1 U15701 ( .A1(n21662), .A2(DATAI_1_), .ZN(n13893) );
  AND2_X1 U15702 ( .A1(n13894), .A2(n13893), .ZN(n21857) );
  INV_X1 U15703 ( .A(n21857), .ZN(n13895) );
  NAND2_X1 U15704 ( .A1(n13934), .A2(n13895), .ZN(n13919) );
  NAND2_X1 U15705 ( .A1(n13922), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n13896) );
  OAI211_X1 U15706 ( .C1(n11838), .C2(n13884), .A(n13919), .B(n13896), .ZN(
        P1_U2953) );
  INV_X1 U15707 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19771) );
  NAND2_X1 U15708 ( .A1(n13922), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n13897) );
  OAI211_X1 U15709 ( .C1(n19771), .C2(n13884), .A(n13898), .B(n13897), .ZN(
        P1_U2954) );
  INV_X1 U15710 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13899) );
  OR2_X1 U15711 ( .A1(n21662), .A2(n13899), .ZN(n13901) );
  NAND2_X1 U15712 ( .A1(n21662), .A2(DATAI_3_), .ZN(n13900) );
  AND2_X1 U15713 ( .A1(n13901), .A2(n13900), .ZN(n21944) );
  INV_X1 U15714 ( .A(n21944), .ZN(n13902) );
  NAND2_X1 U15715 ( .A1(n13934), .A2(n13902), .ZN(n13907) );
  NAND2_X1 U15716 ( .A1(n13922), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n13903) );
  OAI211_X1 U15717 ( .C1(n11864), .C2(n13884), .A(n13907), .B(n13903), .ZN(
        P1_U2955) );
  NAND2_X1 U15718 ( .A1(n13922), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n13904) );
  OAI211_X1 U15719 ( .C1(n11828), .C2(n13884), .A(n13905), .B(n13904), .ZN(
        P1_U2959) );
  INV_X1 U15720 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14567) );
  NAND2_X1 U15721 ( .A1(n13922), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13906) );
  OAI211_X1 U15722 ( .C1(n14567), .C2(n13884), .A(n13907), .B(n13906), .ZN(
        P1_U2940) );
  NAND2_X1 U15723 ( .A1(n13922), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13908) );
  OAI211_X1 U15724 ( .C1(n15812), .C2(n13884), .A(n13909), .B(n13908), .ZN(
        P1_U2949) );
  NAND2_X1 U15725 ( .A1(n13922), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13910) );
  OAI211_X1 U15726 ( .C1(n15805), .C2(n13884), .A(n13911), .B(n13910), .ZN(
        P1_U2950) );
  NAND2_X1 U15727 ( .A1(n13922), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U15728 ( .C1(n15799), .C2(n13884), .A(n13913), .B(n13912), .ZN(
        P1_U2951) );
  INV_X1 U15729 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13914) );
  OR2_X1 U15730 ( .A1(n21662), .A2(n13914), .ZN(n13916) );
  NAND2_X1 U15731 ( .A1(n21662), .A2(DATAI_0_), .ZN(n13915) );
  AND2_X1 U15732 ( .A1(n13916), .A2(n13915), .ZN(n21661) );
  INV_X1 U15733 ( .A(n21661), .ZN(n21637) );
  NAND2_X1 U15734 ( .A1(n13934), .A2(n21637), .ZN(n13926) );
  NAND2_X1 U15735 ( .A1(n13922), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U15736 ( .C1(n12026), .C2(n13884), .A(n13926), .B(n13917), .ZN(
        P1_U2937) );
  INV_X1 U15737 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U15738 ( .A1(n13922), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13918) );
  OAI211_X1 U15739 ( .C1(n14253), .C2(n13884), .A(n13919), .B(n13918), .ZN(
        P1_U2938) );
  NAND2_X1 U15740 ( .A1(n13922), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13920) );
  OAI211_X1 U15741 ( .C1(n15819), .C2(n13884), .A(n13921), .B(n13920), .ZN(
        P1_U2948) );
  NAND2_X1 U15742 ( .A1(n13922), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13923) );
  OAI211_X1 U15743 ( .C1(n15825), .C2(n13884), .A(n13924), .B(n13923), .ZN(
        P1_U2947) );
  NAND2_X1 U15744 ( .A1(n13922), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n13925) );
  OAI211_X1 U15745 ( .C1(n11848), .C2(n13884), .A(n13926), .B(n13925), .ZN(
        P1_U2952) );
  INV_X1 U15746 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13931) );
  OR2_X1 U15747 ( .A1(n14332), .A2(n18661), .ZN(n13927) );
  OAI21_X1 U15748 ( .B1(n14275), .B2(n13927), .A(n14633), .ZN(n13929) );
  INV_X1 U15749 ( .A(n21604), .ZN(n13928) );
  NOR2_X4 U15750 ( .A1(n17337), .A2(n17369), .ZN(n17357) );
  AOI22_X1 U15751 ( .A1(n17358), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13930) );
  OAI21_X1 U15752 ( .B1(n13931), .B2(n14154), .A(n13930), .ZN(P2_U2933) );
  AOI22_X1 U15753 ( .A1(n17358), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13932) );
  OAI21_X1 U15754 ( .B1(n13933), .B2(n14154), .A(n13932), .ZN(P2_U2934) );
  INV_X1 U15755 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19795) );
  INV_X1 U15756 ( .A(n13934), .ZN(n13939) );
  INV_X1 U15757 ( .A(DATAI_15_), .ZN(n13935) );
  NOR2_X1 U15758 ( .A1(n21663), .A2(n13935), .ZN(n13936) );
  AOI21_X1 U15759 ( .B1(n21663), .B2(BUF1_REG_15__SCAN_IN), .A(n13936), .ZN(
        n15862) );
  INV_X1 U15760 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13937) );
  OAI222_X1 U15761 ( .A1(n13884), .A2(n19795), .B1(n13939), .B2(n15862), .C1(
        n13938), .C2(n13937), .ZN(P1_U2967) );
  XNOR2_X1 U15762 ( .A(n13940), .B(n14208), .ZN(n14177) );
  NAND2_X1 U15763 ( .A1(n14177), .A2(n19949), .ZN(n13944) );
  INV_X1 U15764 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13941) );
  OAI22_X1 U15765 ( .A1(n19901), .A2(n14390), .B1(n21401), .B2(n13941), .ZN(
        n13942) );
  AOI21_X1 U15766 ( .B1(n19927), .B2(n14390), .A(n13942), .ZN(n13943) );
  OAI211_X1 U15767 ( .C1(n19915), .C2(n14397), .A(n13944), .B(n13943), .ZN(
        P1_U2998) );
  NAND2_X1 U15768 ( .A1(n13945), .A2(n14022), .ZN(n13949) );
  NAND2_X1 U15769 ( .A1(n19243), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14880) );
  NAND2_X1 U15770 ( .A1(n14299), .A2(n19172), .ZN(n13946) );
  NAND2_X1 U15771 ( .A1(n14880), .A2(n13946), .ZN(n19145) );
  NOR2_X1 U15772 ( .A1(n19145), .A2(n19276), .ZN(n13947) );
  AOI21_X1 U15773 ( .B1(n14019), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13947), .ZN(n13948) );
  NAND2_X1 U15774 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  NAND2_X1 U15775 ( .A1(n13955), .A2(n13954), .ZN(n14017) );
  MUX2_X1 U15776 ( .A(n12609), .B(n12770), .S(n14161), .Z(n13957) );
  OAI21_X1 U15777 ( .B1(n17309), .B2(n16302), .A(n13957), .ZN(P2_U2885) );
  OR2_X1 U15778 ( .A1(n21687), .A2(n21829), .ZN(n21786) );
  NOR2_X1 U15779 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21556) );
  INV_X1 U15780 ( .A(n13958), .ZN(n13959) );
  OAI21_X1 U15781 ( .B1(n13959), .B2(n16098), .A(n14443), .ZN(n13960) );
  NAND2_X1 U15782 ( .A1(n13960), .A2(n21547), .ZN(n16084) );
  NAND2_X1 U15783 ( .A1(n16084), .A2(n21547), .ZN(n13962) );
  INV_X1 U15784 ( .A(n21552), .ZN(n13961) );
  NAND2_X1 U15785 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  NAND2_X1 U15786 ( .A1(n22129), .A2(n13963), .ZN(n17061) );
  NAND2_X1 U15787 ( .A1(n17061), .A2(n21852), .ZN(n14070) );
  AOI211_X1 U15788 ( .C1(n21829), .C2(n21687), .A(n21701), .B(n14070), .ZN(
        n13966) );
  NAND2_X1 U15789 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21805), .ZN(n16085) );
  NAND2_X1 U15790 ( .A1(n17061), .A2(n16085), .ZN(n14071) );
  OAI22_X1 U15791 ( .A1(n14071), .A2(n13964), .B1(n21823), .B2(n17061), .ZN(
        n13965) );
  OR2_X1 U15792 ( .A1(n13966), .A2(n13965), .ZN(P1_U3477) );
  XNOR2_X1 U15793 ( .A(n13968), .B(n13967), .ZN(n18583) );
  XNOR2_X1 U15794 ( .A(n17305), .B(n18583), .ZN(n13980) );
  NAND2_X1 U15795 ( .A1(n13969), .A2(n14327), .ZN(n14273) );
  NAND2_X1 U15796 ( .A1(n14273), .A2(n13970), .ZN(n13971) );
  AND2_X1 U15797 ( .A1(n13188), .A2(n18655), .ZN(n14336) );
  NAND2_X1 U15798 ( .A1(n18341), .A2(n14336), .ZN(n13972) );
  AND2_X1 U15799 ( .A1(n19496), .A2(n12519), .ZN(n15489) );
  INV_X1 U15800 ( .A(n14684), .ZN(n19489) );
  INV_X1 U15801 ( .A(n19592), .ZN(n19580) );
  NAND2_X1 U15802 ( .A1(n19489), .A2(n19580), .ZN(n13979) );
  NAND2_X1 U15803 ( .A1(n19496), .A2(n13976), .ZN(n16373) );
  INV_X1 U15804 ( .A(n18583), .ZN(n13977) );
  AOI22_X1 U15805 ( .A1(n19585), .A2(n13977), .B1(n19579), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13978) );
  OAI211_X1 U15806 ( .C1(n13980), .C2(n19342), .A(n13979), .B(n13978), .ZN(
        P2_U2919) );
  NOR2_X1 U15807 ( .A1(n17305), .A2(n18583), .ZN(n13988) );
  INV_X1 U15808 ( .A(n13981), .ZN(n13984) );
  INV_X1 U15809 ( .A(n13982), .ZN(n13983) );
  NAND2_X1 U15810 ( .A1(n13984), .A2(n13983), .ZN(n13985) );
  NAND2_X1 U15811 ( .A1(n13986), .A2(n13985), .ZN(n16236) );
  XOR2_X1 U15812 ( .A(n16236), .B(n17320), .Z(n13987) );
  NOR2_X1 U15813 ( .A1(n13987), .A2(n13988), .ZN(n14474) );
  AOI21_X1 U15814 ( .B1(n13988), .B2(n13987), .A(n14474), .ZN(n13991) );
  AOI22_X1 U15815 ( .A1(n19585), .A2(n16236), .B1(n19579), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13990) );
  INV_X1 U15816 ( .A(n14744), .ZN(n16383) );
  NAND2_X1 U15817 ( .A1(n19489), .A2(n16383), .ZN(n13989) );
  OAI211_X1 U15818 ( .C1(n13991), .C2(n19342), .A(n13990), .B(n13989), .ZN(
        P2_U2918) );
  OAI211_X1 U15819 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16930), .B(n14526), .ZN(n13994) );
  NAND2_X1 U15820 ( .A1(n18627), .A2(n13992), .ZN(n13993) );
  OAI211_X1 U15821 ( .C1(n13995), .C2(n18607), .A(n13994), .B(n13993), .ZN(
        n14001) );
  INV_X1 U15822 ( .A(n16236), .ZN(n17313) );
  INV_X1 U15823 ( .A(n13996), .ZN(n18590) );
  AOI22_X1 U15824 ( .A1(n18623), .A2(n13997), .B1(n18590), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13999) );
  OAI211_X1 U15825 ( .C1(n17313), .C2(n18603), .A(n13999), .B(n13998), .ZN(
        n14000) );
  OR2_X1 U15826 ( .A1(n14001), .A2(n14000), .ZN(P2_U3045) );
  XNOR2_X1 U15827 ( .A(n21701), .B(n21752), .ZN(n14002) );
  OAI222_X1 U15828 ( .A1(n14071), .A2(n13802), .B1(n14070), .B2(n14002), .C1(
        n21824), .C2(n17061), .ZN(P1_U3476) );
  OAI21_X1 U15829 ( .B1(n14005), .B2(n14004), .A(n14003), .ZN(n14518) );
  OR2_X1 U15830 ( .A1(n14006), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14007) );
  AND2_X1 U15831 ( .A1(n14008), .A2(n14007), .ZN(n21410) );
  OAI21_X1 U15832 ( .B1(n19943), .B2(n14009), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14010) );
  INV_X1 U15833 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14525) );
  OR2_X1 U15834 ( .A1(n21401), .A2(n14525), .ZN(n21417) );
  NAND2_X1 U15835 ( .A1(n14010), .A2(n21417), .ZN(n14011) );
  AOI21_X1 U15836 ( .B1(n19949), .B2(n21410), .A(n14011), .ZN(n14012) );
  OAI21_X1 U15837 ( .B1(n19915), .B2(n14518), .A(n14012), .ZN(P1_U2999) );
  INV_X1 U15838 ( .A(n14013), .ZN(n14014) );
  NAND2_X1 U15839 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  NAND2_X1 U15840 ( .A1(n14880), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14018) );
  NOR2_X1 U15841 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19172), .ZN(
        n19225) );
  NAND2_X1 U15842 ( .A1(n19243), .A2(n19225), .ZN(n19209) );
  AOI21_X1 U15843 ( .B1(n14018), .B2(n19209), .A(n19276), .ZN(n19144) );
  AOI21_X1 U15844 ( .B1(n14019), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19144), .ZN(n14025) );
  INV_X1 U15845 ( .A(n14025), .ZN(n14020) );
  INV_X1 U15846 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19480) );
  NAND2_X1 U15847 ( .A1(n14020), .A2(n14023), .ZN(n14028) );
  INV_X1 U15848 ( .A(n14023), .ZN(n14024) );
  AND2_X1 U15849 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  NAND2_X1 U15850 ( .A1(n12532), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14027) );
  AND2_X1 U15851 ( .A1(n14028), .A2(n14027), .ZN(n14029) );
  INV_X1 U15852 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14895) );
  OR2_X1 U15853 ( .A1(n14033), .A2(n14032), .ZN(n14034) );
  NAND2_X1 U15854 ( .A1(n14129), .A2(n14034), .ZN(n19343) );
  OAI21_X1 U15855 ( .B1(n14036), .B2(n14035), .A(n14039), .ZN(n14763) );
  NOR2_X1 U15856 ( .A1(n14763), .A2(n14161), .ZN(n14037) );
  AOI21_X1 U15857 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n14161), .A(n14037), .ZN(
        n14038) );
  OAI21_X1 U15858 ( .B1(n19343), .B2(n16302), .A(n14038), .ZN(P2_U2883) );
  XOR2_X1 U15859 ( .A(n14129), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14042)
         );
  AOI21_X1 U15860 ( .B1(n14040), .B2(n14039), .A(n14157), .ZN(n18368) );
  INV_X1 U15861 ( .A(n18368), .ZN(n14845) );
  MUX2_X1 U15862 ( .A(n12782), .B(n14845), .S(n16284), .Z(n14041) );
  OAI21_X1 U15863 ( .B1(n14042), .B2(n16302), .A(n14041), .ZN(P2_U2882) );
  XNOR2_X1 U15864 ( .A(n14044), .B(n14043), .ZN(n14125) );
  INV_X1 U15865 ( .A(n14045), .ZN(n14046) );
  AOI21_X1 U15866 ( .B1(n14048), .B2(n14047), .A(n14046), .ZN(n14052) );
  INV_X2 U15867 ( .A(n21401), .ZN(n21390) );
  AOI22_X1 U15868 ( .A1(n19943), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21390), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14049) );
  OAI21_X1 U15869 ( .B1(n19952), .B2(n14404), .A(n14049), .ZN(n14050) );
  AOI21_X1 U15870 ( .B1(n14052), .B2(n19948), .A(n14050), .ZN(n14051) );
  OAI21_X1 U15871 ( .B1(n14125), .B2(n21546), .A(n14051), .ZN(P1_U2997) );
  INV_X1 U15872 ( .A(n14052), .ZN(n14409) );
  INV_X1 U15873 ( .A(n14053), .ZN(n14054) );
  AOI21_X1 U15874 ( .B1(n14055), .B2(n13785), .A(n14054), .ZN(n14062) );
  INV_X1 U15875 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U15876 ( .A1(n15591), .A2(n14399), .ZN(n14060) );
  NAND2_X1 U15877 ( .A1(n14056), .A2(n14209), .ZN(n14058) );
  NAND2_X1 U15878 ( .A1(n13785), .A2(n14399), .ZN(n14057) );
  NAND3_X1 U15879 ( .A1(n14058), .A2(n15607), .A3(n14057), .ZN(n14059) );
  NAND2_X1 U15880 ( .A1(n14060), .A2(n14059), .ZN(n14061) );
  NOR2_X1 U15881 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  OR2_X1 U15882 ( .A1(n14214), .A2(n14063), .ZN(n14398) );
  INV_X1 U15883 ( .A(n14398), .ZN(n14064) );
  AOI22_X1 U15884 ( .A1(n19865), .A2(n14064), .B1(n15794), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14065) );
  OAI21_X1 U15885 ( .B1(n14409), .B2(n15783), .A(n14065), .ZN(P1_U2870) );
  INV_X1 U15886 ( .A(n21753), .ZN(n14385) );
  INV_X1 U15887 ( .A(n13508), .ZN(n14068) );
  NAND2_X1 U15888 ( .A1(n21822), .A2(n21701), .ZN(n21846) );
  NAND2_X1 U15889 ( .A1(n21742), .A2(n21701), .ZN(n21746) );
  INV_X1 U15890 ( .A(n21746), .ZN(n14067) );
  AOI21_X1 U15891 ( .B1(n14068), .B2(n21846), .A(n14067), .ZN(n14069) );
  OAI222_X1 U15892 ( .A1(n17061), .A2(n21825), .B1(n14071), .B2(n14385), .C1(
        n14070), .C2(n14069), .ZN(P1_U3475) );
  INV_X1 U15893 ( .A(n14072), .ZN(n14073) );
  AOI21_X1 U15894 ( .B1(n15580), .B2(n14119), .A(n14073), .ZN(n21408) );
  INV_X1 U15895 ( .A(n21408), .ZN(n14075) );
  INV_X1 U15896 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14074) );
  OAI222_X1 U15897 ( .A1(n14075), .A2(n15785), .B1(n14074), .B2(n19870), .C1(
        n14518), .C2(n15783), .ZN(P1_U2872) );
  OAI21_X1 U15898 ( .B1(n14076), .B2(n14085), .A(n14801), .ZN(n18403) );
  INV_X1 U15899 ( .A(n16336), .ZN(n14077) );
  INV_X1 U15900 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17356) );
  OAI222_X1 U15901 ( .A1(n18403), .A2(n19348), .B1(n14684), .B2(n14077), .C1(
        n19496), .C2(n17356), .ZN(P2_U2910) );
  XNOR2_X1 U15902 ( .A(n14078), .B(n14079), .ZN(n18384) );
  INV_X1 U15903 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17350) );
  OAI222_X1 U15904 ( .A1(n14684), .A2(n14754), .B1(n18384), .B2(n19348), .C1(
        n19496), .C2(n17350), .ZN(P2_U2913) );
  OR2_X1 U15905 ( .A1(n14081), .A2(n14080), .ZN(n14082) );
  AND2_X1 U15906 ( .A1(n14082), .A2(n14083), .ZN(n16934) );
  INV_X1 U15907 ( .A(n16934), .ZN(n18390) );
  INV_X1 U15908 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17352) );
  OAI222_X1 U15909 ( .A1(n14684), .A2(n16352), .B1(n18390), .B2(n19348), .C1(
        n19496), .C2(n17352), .ZN(P2_U2912) );
  NAND2_X1 U15910 ( .A1(n14084), .A2(n14083), .ZN(n14087) );
  INV_X1 U15911 ( .A(n14085), .ZN(n14086) );
  NAND2_X1 U15912 ( .A1(n14087), .A2(n14086), .ZN(n18602) );
  INV_X1 U15913 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17354) );
  OAI222_X1 U15914 ( .A1(n14684), .A2(n16347), .B1(n18602), .B2(n19348), .C1(
        n19496), .C2(n17354), .ZN(P2_U2911) );
  NAND2_X1 U15915 ( .A1(n14088), .A2(n17050), .ZN(n14363) );
  NAND2_X1 U15916 ( .A1(n14115), .A2(n14363), .ZN(n14090) );
  NAND3_X1 U15917 ( .A1(n14090), .A2(n11645), .A3(n14089), .ZN(n14091) );
  NAND2_X1 U15918 ( .A1(n15546), .A2(n14091), .ZN(n14095) );
  INV_X1 U15919 ( .A(n21229), .ZN(n21586) );
  AOI21_X1 U15920 ( .B1(n14364), .B2(n21587), .A(n21586), .ZN(n14092) );
  NAND2_X1 U15921 ( .A1(n15540), .A2(n14092), .ZN(n14094) );
  MUX2_X1 U15922 ( .A(n14095), .B(n14094), .S(n14093), .Z(n14100) );
  OR2_X1 U15923 ( .A1(n16089), .A2(n21859), .ZN(n14097) );
  OAI21_X1 U15924 ( .B1(n15546), .B2(n14097), .A(n14096), .ZN(n14098) );
  INV_X1 U15925 ( .A(n14098), .ZN(n14099) );
  NOR2_X1 U15926 ( .A1(n14102), .A2(n14101), .ZN(n15537) );
  OAI21_X1 U15927 ( .B1(n15538), .B2(n15545), .A(n15547), .ZN(n14104) );
  NAND2_X1 U15928 ( .A1(n14113), .A2(n21991), .ZN(n14103) );
  NAND3_X1 U15929 ( .A1(n15537), .A2(n14104), .A3(n14103), .ZN(n14105) );
  OAI211_X1 U15930 ( .C1(n14108), .C2(n11645), .A(n14107), .B(n14106), .ZN(
        n14109) );
  NAND2_X1 U15931 ( .A1(n14118), .A2(n14109), .ZN(n21238) );
  NOR2_X1 U15932 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21238), .ZN(
        n14110) );
  NOR2_X1 U15933 ( .A1(n21390), .A2(n14118), .ZN(n21242) );
  INV_X1 U15934 ( .A(n21327), .ZN(n21414) );
  NAND2_X1 U15935 ( .A1(n14118), .A2(n17021), .ZN(n21239) );
  NAND2_X1 U15936 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14111) );
  OAI22_X1 U15937 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21328), .B1(
        n14111), .B2(n21367), .ZN(n14122) );
  NAND2_X1 U15938 ( .A1(n14113), .A2(n14112), .ZN(n14116) );
  NAND2_X1 U15939 ( .A1(n14115), .A2(n14114), .ZN(n17051) );
  NAND2_X1 U15940 ( .A1(n14116), .A2(n17051), .ZN(n14117) );
  NAND2_X1 U15941 ( .A1(n21390), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n14120) );
  OAI21_X1 U15942 ( .B1(n14119), .B2(n14208), .A(n14209), .ZN(n21276) );
  OR2_X1 U15943 ( .A1(n21367), .A2(n21276), .ZN(n14210) );
  OAI211_X1 U15944 ( .C1(n21389), .C2(n14398), .A(n14120), .B(n14210), .ZN(
        n14121) );
  AOI221_X1 U15945 ( .B1(n21414), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n14122), .C2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n14121), .ZN(
        n14124) );
  NAND3_X1 U15946 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21310), .A3(
        n14209), .ZN(n14123) );
  OAI211_X1 U15947 ( .C1(n21335), .C2(n14125), .A(n14124), .B(n14123), .ZN(
        P1_U3029) );
  INV_X1 U15948 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U15949 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17357), .B1(n17369), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14126) );
  OAI21_X1 U15950 ( .B1(n14127), .B2(n14154), .A(n14126), .ZN(P2_U2935) );
  INV_X1 U15951 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19340) );
  XNOR2_X1 U15952 ( .A(n14226), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14134) );
  OR2_X1 U15953 ( .A1(n14131), .A2(n14130), .ZN(n14132) );
  NAND2_X1 U15954 ( .A1(n14224), .A2(n14132), .ZN(n18391) );
  MUX2_X1 U15955 ( .A(n12852), .B(n18391), .S(n16284), .Z(n14133) );
  OAI21_X1 U15956 ( .B1(n14134), .B2(n16302), .A(n14133), .ZN(P2_U2880) );
  INV_X1 U15957 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U15958 ( .A1(n17369), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14135) );
  OAI21_X1 U15959 ( .B1(n16342), .B2(n14154), .A(n14135), .ZN(P2_U2927) );
  AOI22_X1 U15960 ( .A1(n17369), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14136) );
  OAI21_X1 U15961 ( .B1(n14137), .B2(n14154), .A(n14136), .ZN(P2_U2926) );
  AOI22_X1 U15962 ( .A1(n17369), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14138) );
  OAI21_X1 U15963 ( .B1(n14139), .B2(n14154), .A(n14138), .ZN(P2_U2923) );
  INV_X1 U15964 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U15965 ( .A1(n17369), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14140) );
  OAI21_X1 U15966 ( .B1(n14141), .B2(n14154), .A(n14140), .ZN(P2_U2929) );
  AOI22_X1 U15967 ( .A1(n17369), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14142) );
  OAI21_X1 U15968 ( .B1(n16363), .B2(n14154), .A(n14142), .ZN(P2_U2930) );
  AOI22_X1 U15969 ( .A1(n17369), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14143) );
  OAI21_X1 U15970 ( .B1(n14144), .B2(n14154), .A(n14143), .ZN(P2_U2924) );
  INV_X1 U15971 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16354) );
  AOI22_X1 U15972 ( .A1(n17369), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14145) );
  OAI21_X1 U15973 ( .B1(n16354), .B2(n14154), .A(n14145), .ZN(P2_U2928) );
  AOI22_X1 U15974 ( .A1(n17369), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14146) );
  OAI21_X1 U15975 ( .B1(n14147), .B2(n14154), .A(n14146), .ZN(P2_U2922) );
  INV_X1 U15976 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U15977 ( .A1(n17369), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14148) );
  OAI21_X1 U15978 ( .B1(n14149), .B2(n14154), .A(n14148), .ZN(P2_U2931) );
  AOI22_X1 U15979 ( .A1(n17369), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14150) );
  OAI21_X1 U15980 ( .B1(n14151), .B2(n14154), .A(n14150), .ZN(P2_U2925) );
  INV_X1 U15981 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16372) );
  AOI22_X1 U15982 ( .A1(n17358), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14152) );
  OAI21_X1 U15983 ( .B1(n16372), .B2(n14154), .A(n14152), .ZN(P2_U2932) );
  AOI22_X1 U15984 ( .A1(n17358), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14153) );
  OAI21_X1 U15985 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(P2_U2921) );
  OAI21_X1 U15986 ( .B1(n14158), .B2(n14157), .A(n14156), .ZN(n17280) );
  NOR2_X1 U15987 ( .A1(n14129), .A2(n15371), .ZN(n14160) );
  INV_X1 U15988 ( .A(n14226), .ZN(n14159) );
  OAI211_X1 U15989 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14160), .A(
        n14159), .B(n16307), .ZN(n14163) );
  NAND2_X1 U15990 ( .A1(n14161), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14162) );
  OAI211_X1 U15991 ( .C1(n17280), .C2(n14161), .A(n14163), .B(n14162), .ZN(
        P2_U2881) );
  NAND2_X1 U15992 ( .A1(n14165), .A2(n14164), .ZN(n14166) );
  INV_X1 U15993 ( .A(n14166), .ZN(n14167) );
  OAI222_X1 U15994 ( .A1(n15866), .A2(n14397), .B1(n15852), .B2(n11838), .C1(
        n15863), .C2(n21857), .ZN(P1_U2903) );
  OAI222_X1 U15995 ( .A1(n15866), .A2(n14409), .B1(n15864), .B2(n19771), .C1(
        n15863), .C2(n21900), .ZN(P1_U2902) );
  OAI222_X1 U15996 ( .A1(n15866), .A2(n14518), .B1(n15852), .B2(n11848), .C1(
        n15863), .C2(n21661), .ZN(P1_U2904) );
  OAI21_X1 U15997 ( .B1(n14170), .B2(n14169), .A(n14168), .ZN(n14389) );
  OAI222_X1 U15998 ( .A1(n15866), .A2(n14389), .B1(n15864), .B2(n11864), .C1(
        n15863), .C2(n21944), .ZN(P1_U2901) );
  NOR2_X1 U15999 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21367), .ZN(
        n21412) );
  OAI21_X1 U16000 ( .B1(n21412), .B2(n21414), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14173) );
  NOR2_X1 U16001 ( .A1(n21401), .A2(n13941), .ZN(n14171) );
  AOI21_X1 U16002 ( .B1(n21409), .B2(n14394), .A(n14171), .ZN(n14172) );
  NAND2_X1 U16003 ( .A1(n14173), .A2(n14172), .ZN(n14176) );
  NAND2_X1 U16004 ( .A1(n21328), .A2(n21367), .ZN(n21337) );
  INV_X1 U16005 ( .A(n21337), .ZN(n21385) );
  NOR3_X1 U16006 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14174), .A3(
        n21385), .ZN(n14175) );
  AOI211_X1 U16007 ( .C1(n21411), .C2(n14177), .A(n14176), .B(n14175), .ZN(
        n14178) );
  INV_X1 U16008 ( .A(n14178), .ZN(P1_U3030) );
  INV_X1 U16009 ( .A(n16316), .ZN(n14181) );
  NOR2_X1 U16010 ( .A1(n16893), .A2(n14179), .ZN(n14180) );
  OR2_X1 U16011 ( .A1(n14220), .A2(n14180), .ZN(n16880) );
  INV_X1 U16012 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17364) );
  OAI222_X1 U16013 ( .A1(n14684), .A2(n14181), .B1(n16880), .B2(n19348), .C1(
        n19496), .C2(n17364), .ZN(P2_U2907) );
  AOI21_X1 U16014 ( .B1(n14183), .B2(n14168), .A(n14182), .ZN(n14248) );
  INV_X1 U16015 ( .A(n14248), .ZN(n14457) );
  INV_X1 U16016 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14449) );
  INV_X1 U16017 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n19869) );
  NAND2_X1 U16018 ( .A1(n14193), .A2(n19869), .ZN(n14186) );
  NAND2_X1 U16019 ( .A1(n13785), .A2(n19869), .ZN(n14184) );
  OAI211_X1 U16020 ( .C1(n10968), .C2(n14211), .A(n14184), .B(n14056), .ZN(
        n14185) );
  AND2_X1 U16021 ( .A1(n14186), .A2(n14185), .ZN(n14213) );
  OAI21_X1 U16022 ( .B1(n10968), .B2(n14187), .A(n14056), .ZN(n14188) );
  OAI21_X1 U16023 ( .B1(n13878), .B2(P1_EBX_REG_4__SCAN_IN), .A(n14188), .ZN(
        n14190) );
  NAND2_X1 U16024 ( .A1(n15591), .A2(n14449), .ZN(n14189) );
  XNOR2_X1 U16025 ( .A(n14212), .B(n14198), .ZN(n14450) );
  OAI222_X1 U16026 ( .A1(n15783), .A2(n14457), .B1(n19870), .B2(n14449), .C1(
        n15785), .C2(n14450), .ZN(P1_U2868) );
  OAI222_X1 U16027 ( .A1(n15866), .A2(n14457), .B1(n15852), .B2(n19774), .C1(
        n15863), .C2(n21989), .ZN(P1_U2900) );
  OAI21_X1 U16028 ( .B1(n14182), .B2(n14192), .A(n14191), .ZN(n19874) );
  INV_X1 U16029 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21265) );
  INV_X1 U16030 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14194) );
  NAND2_X1 U16031 ( .A1(n13785), .A2(n14194), .ZN(n14195) );
  OAI211_X1 U16032 ( .C1(n10968), .C2(n21265), .A(n14195), .B(n14056), .ZN(
        n14196) );
  OAI21_X1 U16033 ( .B1(n15590), .B2(P1_EBX_REG_5__SCAN_IN), .A(n14196), .ZN(
        n14197) );
  OAI21_X1 U16034 ( .B1(n14212), .B2(n14198), .A(n14197), .ZN(n14199) );
  NAND2_X1 U16035 ( .A1(n14199), .A2(n14241), .ZN(n21272) );
  INV_X1 U16036 ( .A(n21272), .ZN(n14200) );
  AOI22_X1 U16037 ( .A1(n19865), .A2(n14200), .B1(n15794), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14201) );
  OAI21_X1 U16038 ( .B1(n19874), .B2(n15796), .A(n14201), .ZN(P1_U2867) );
  XNOR2_X1 U16039 ( .A(n14203), .B(n14202), .ZN(n14218) );
  INV_X1 U16040 ( .A(n14389), .ZN(n19867) );
  INV_X1 U16041 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14204) );
  NOR2_X1 U16042 ( .A1(n21401), .A2(n14204), .ZN(n14215) );
  AOI21_X1 U16043 ( .B1(n19943), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14215), .ZN(n14205) );
  OAI21_X1 U16044 ( .B1(n19952), .B2(n14381), .A(n14205), .ZN(n14206) );
  AOI21_X1 U16045 ( .B1(n19867), .B2(n19948), .A(n14206), .ZN(n14207) );
  OAI21_X1 U16046 ( .B1(n14218), .B2(n21546), .A(n14207), .ZN(P1_U2996) );
  NOR2_X1 U16047 ( .A1(n14209), .A2(n14208), .ZN(n21277) );
  OAI211_X1 U16048 ( .C1(n21277), .C2(n21328), .A(n21327), .B(n14210), .ZN(
        n16074) );
  AOI22_X1 U16049 ( .A1(n21277), .A2(n21310), .B1(n21325), .B2(n21276), .ZN(
        n21287) );
  INV_X1 U16050 ( .A(n21287), .ZN(n21282) );
  AOI22_X1 U16051 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16074), .B1(
        n21282), .B2(n14211), .ZN(n14217) );
  OAI21_X1 U16052 ( .B1(n14214), .B2(n14213), .A(n14212), .ZN(n14370) );
  INV_X1 U16053 ( .A(n14370), .ZN(n19864) );
  AOI21_X1 U16054 ( .B1(n21409), .B2(n19864), .A(n14215), .ZN(n14216) );
  OAI211_X1 U16055 ( .C1(n14218), .C2(n21335), .A(n14217), .B(n14216), .ZN(
        P1_U3028) );
  OR2_X1 U16056 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  NAND2_X1 U16057 ( .A1(n14411), .A2(n14221), .ZN(n18436) );
  INV_X1 U16058 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17366) );
  OAI222_X1 U16059 ( .A1(n14684), .A2(n14222), .B1(n18436), .B2(n19348), .C1(
        n19496), .C2(n17366), .ZN(P2_U2906) );
  OAI222_X1 U16060 ( .A1(n15866), .A2(n19874), .B1(n15852), .B2(n19776), .C1(
        n15863), .C2(n22035), .ZN(P1_U2899) );
  NAND2_X1 U16061 ( .A1(n14224), .A2(n14223), .ZN(n14225) );
  NAND2_X1 U16062 ( .A1(n14263), .A2(n14225), .ZN(n18606) );
  INV_X1 U16063 ( .A(n14260), .ZN(n14228) );
  OAI211_X1 U16064 ( .C1(n11098), .C2(n14229), .A(n14228), .B(n16307), .ZN(
        n14231) );
  NAND2_X1 U16065 ( .A1(n14161), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14230) );
  OAI211_X1 U16066 ( .C1(n18606), .C2(n14161), .A(n14231), .B(n14230), .ZN(
        P2_U2879) );
  INV_X1 U16067 ( .A(n14232), .ZN(n14433) );
  NAND2_X1 U16068 ( .A1(n14191), .A2(n14233), .ZN(n14234) );
  NAND2_X1 U16069 ( .A1(n14433), .A2(n14234), .ZN(n21423) );
  INV_X1 U16070 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21421) );
  NAND2_X1 U16071 ( .A1(n15591), .A2(n21421), .ZN(n14239) );
  INV_X1 U16072 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14235) );
  NAND2_X1 U16073 ( .A1(n14056), .A2(n14235), .ZN(n14237) );
  NAND2_X1 U16074 ( .A1(n13785), .A2(n21421), .ZN(n14236) );
  NAND3_X1 U16075 ( .A1(n14237), .A2(n15607), .A3(n14236), .ZN(n14238) );
  AND2_X1 U16076 ( .A1(n14239), .A2(n14238), .ZN(n14240) );
  AND2_X1 U16077 ( .A1(n14241), .A2(n14240), .ZN(n14242) );
  OR2_X1 U16078 ( .A1(n14242), .A2(n14438), .ZN(n21420) );
  INV_X1 U16079 ( .A(n21420), .ZN(n16072) );
  AOI22_X1 U16080 ( .A1(n19865), .A2(n16072), .B1(n15794), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n14243) );
  OAI21_X1 U16081 ( .B1(n21423), .B2(n15783), .A(n14243), .ZN(P1_U2866) );
  XNOR2_X1 U16082 ( .A(n14245), .B(n14244), .ZN(n14259) );
  INV_X1 U16083 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n19801) );
  NOR2_X1 U16084 ( .A1(n21401), .A2(n19801), .ZN(n14256) );
  AOI21_X1 U16085 ( .B1(n19943), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14256), .ZN(n14246) );
  OAI21_X1 U16086 ( .B1(n19952), .B2(n14451), .A(n14246), .ZN(n14247) );
  AOI21_X1 U16087 ( .B1(n14248), .B2(n19948), .A(n14247), .ZN(n14249) );
  OAI21_X1 U16088 ( .B1(n14259), .B2(n21546), .A(n14249), .ZN(P1_U2995) );
  NAND3_X1 U16089 ( .A1(n15546), .A2(n14250), .A3(n17021), .ZN(n14251) );
  INV_X1 U16090 ( .A(n16083), .ZN(n17059) );
  NOR2_X1 U16091 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17059), .ZN(n19780) );
  NOR2_X4 U16092 ( .A1(n19767), .A2(n21230), .ZN(n19784) );
  AOI22_X1 U16093 ( .A1(n19780), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14252) );
  OAI21_X1 U16094 ( .B1(n14253), .B2(n14578), .A(n14252), .ZN(P1_U2919) );
  AOI22_X1 U16095 ( .A1(n21230), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14254) );
  OAI21_X1 U16096 ( .B1(n12062), .B2(n14578), .A(n14254), .ZN(P1_U2918) );
  NAND2_X1 U16097 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21263) );
  OAI211_X1 U16098 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21282), .B(n21263), .ZN(n14258) );
  NOR2_X1 U16099 ( .A1(n21389), .A2(n14450), .ZN(n14255) );
  AOI211_X1 U16100 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n16074), .A(
        n14256), .B(n14255), .ZN(n14257) );
  OAI211_X1 U16101 ( .C1(n14259), .C2(n21335), .A(n14258), .B(n14257), .ZN(
        P1_U3027) );
  INV_X1 U16102 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n14267) );
  OAI211_X1 U16103 ( .C1(n14260), .C2(n14261), .A(n14418), .B(n16307), .ZN(
        n14266) );
  INV_X1 U16104 ( .A(n14416), .ZN(n14262) );
  AOI21_X1 U16105 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(n16920) );
  NAND2_X1 U16106 ( .A1(n16920), .A2(n16284), .ZN(n14265) );
  OAI211_X1 U16107 ( .C1(n16284), .C2(n14267), .A(n14266), .B(n14265), .ZN(
        P2_U2878) );
  INV_X1 U16108 ( .A(n14336), .ZN(n14268) );
  OR2_X1 U16109 ( .A1(n14337), .A2(n14268), .ZN(n14269) );
  OR2_X1 U16110 ( .A1(n14269), .A2(n14338), .ZN(n14270) );
  AND4_X1 U16111 ( .A1(n14273), .A2(n14272), .A3(n14271), .A4(n14270), .ZN(
        n14277) );
  OR2_X1 U16112 ( .A1(n14332), .A2(n14345), .ZN(n14274) );
  OR2_X1 U16113 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  INV_X1 U16114 ( .A(n16957), .ZN(n14317) );
  NAND2_X1 U16115 ( .A1(n18624), .A2(n14315), .ZN(n14287) );
  NOR2_X1 U16116 ( .A1(n14327), .A2(n14320), .ZN(n14311) );
  NOR2_X1 U16117 ( .A1(n14293), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14310) );
  NOR2_X1 U16118 ( .A1(n14310), .A2(n10989), .ZN(n14284) );
  OR2_X1 U16119 ( .A1(n14280), .A2(n14279), .ZN(n14304) );
  NAND2_X1 U16120 ( .A1(n14304), .A2(n14284), .ZN(n14283) );
  NAND2_X1 U16121 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14308) );
  NAND2_X1 U16122 ( .A1(n13178), .A2(n14308), .ZN(n14306) );
  NOR2_X1 U16123 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14281) );
  OR2_X1 U16124 ( .A1(n14306), .A2(n14281), .ZN(n14282) );
  OAI211_X1 U16125 ( .C1(n14311), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        n14285) );
  INV_X1 U16126 ( .A(n14285), .ZN(n14286) );
  NAND2_X1 U16127 ( .A1(n14287), .A2(n14286), .ZN(n14288) );
  OAI22_X1 U16128 ( .A1(n14317), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n14288), .B2(n16957), .ZN(n14342) );
  INV_X1 U16129 ( .A(n14342), .ZN(n14303) );
  INV_X1 U16130 ( .A(n14288), .ZN(n16970) );
  NAND2_X1 U16131 ( .A1(n18349), .A2(n14315), .ZN(n14291) );
  INV_X1 U16132 ( .A(n13178), .ZN(n14309) );
  AND2_X1 U16133 ( .A1(n14289), .A2(n13180), .ZN(n14294) );
  MUX2_X1 U16134 ( .A(n14309), .B(n14294), .S(n12415), .Z(n14290) );
  NAND2_X1 U16135 ( .A1(n14291), .A2(n14290), .ZN(n16956) );
  INV_X1 U16136 ( .A(n16956), .ZN(n14292) );
  AOI21_X1 U16137 ( .B1(n14292), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14300) );
  NAND2_X1 U16138 ( .A1(n16241), .A2(n14315), .ZN(n14298) );
  NOR2_X1 U16139 ( .A1(n12636), .A2(n14293), .ZN(n14296) );
  INV_X1 U16140 ( .A(n14294), .ZN(n14295) );
  AOI22_X1 U16141 ( .A1(n14296), .A2(n14295), .B1(n13178), .B2(n11243), .ZN(
        n14297) );
  NAND2_X1 U16142 ( .A1(n14298), .A2(n14297), .ZN(n16965) );
  OAI22_X1 U16143 ( .A1(n14300), .A2(n16965), .B1(n14299), .B2(n16956), .ZN(
        n14301) );
  AOI211_X1 U16144 ( .C1(n16970), .C2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16957), .B(n14301), .ZN(n14302) );
  AOI21_X1 U16145 ( .B1(n19172), .B2(n14303), .A(n14302), .ZN(n14319) );
  NAND2_X1 U16146 ( .A1(n14304), .A2(n14278), .ZN(n14307) );
  INV_X1 U16147 ( .A(n14310), .ZN(n14305) );
  NAND3_X1 U16148 ( .A1(n14307), .A2(n14306), .A3(n14305), .ZN(n14313) );
  OAI22_X1 U16149 ( .A1(n14311), .A2(n14310), .B1(n14309), .B2(n14308), .ZN(
        n14312) );
  MUX2_X1 U16150 ( .A(n14313), .B(n14312), .S(n12450), .Z(n14314) );
  AOI211_X1 U16151 ( .C1(n14021), .C2(n14315), .A(n15409), .B(n14314), .ZN(
        n16974) );
  NAND2_X1 U16152 ( .A1(n16974), .A2(n14317), .ZN(n14316) );
  OAI21_X1 U16153 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14317), .A(
        n14316), .ZN(n14341) );
  OR2_X1 U16154 ( .A1(n14341), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14318) );
  AOI221_X1 U16155 ( .B1(n14319), .B2(n14318), .C1(n14341), .C2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14344) );
  INV_X1 U16156 ( .A(n14320), .ZN(n14329) );
  AOI22_X1 U16157 ( .A1(n14323), .A2(n14322), .B1(n14338), .B2(n14321), .ZN(
        n14324) );
  OAI21_X1 U16158 ( .B1(n18645), .B2(n14325), .A(n14324), .ZN(n14326) );
  AOI21_X1 U16159 ( .B1(n14591), .B2(n14327), .A(n14326), .ZN(n14328) );
  OAI21_X1 U16160 ( .B1(n14591), .B2(n14329), .A(n14328), .ZN(n18663) );
  INV_X1 U16161 ( .A(n14330), .ZN(n14331) );
  OR3_X1 U16162 ( .A1(n14332), .A2(n14331), .A3(n18335), .ZN(n18578) );
  INV_X1 U16163 ( .A(n18578), .ZN(n14334) );
  NOR3_X1 U16164 ( .A1(n18663), .A2(n14334), .A3(n14333), .ZN(n14340) );
  NOR4_X1 U16165 ( .A1(n14338), .A2(n14337), .A3(n14336), .A4(n14335), .ZN(
        n18662) );
  OAI21_X1 U16166 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18662), .ZN(n14339) );
  OAI211_X1 U16167 ( .C1(n14342), .C2(n14341), .A(n14340), .B(n14339), .ZN(
        n14343) );
  AOI211_X1 U16168 ( .C1(n16957), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n14344), .B(n14343), .ZN(n18660) );
  NAND3_X1 U16169 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18660), .A3(n16962), 
        .ZN(n14350) );
  NOR2_X1 U16170 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14345), .ZN(n14632) );
  AND2_X1 U16171 ( .A1(n14346), .A2(n14632), .ZN(n14631) );
  AND2_X1 U16172 ( .A1(n14347), .A2(n14631), .ZN(n14348) );
  AOI21_X1 U16173 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n18652) );
  OAI21_X1 U16174 ( .B1(n18652), .B2(n18340), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14351) );
  NOR2_X1 U16175 ( .A1(n18340), .A2(n17303), .ZN(n17001) );
  INV_X1 U16176 ( .A(n17001), .ZN(n18647) );
  NAND2_X1 U16177 ( .A1(n14351), .A2(n18647), .ZN(P2_U3593) );
  INV_X1 U16178 ( .A(n19162), .ZN(n19245) );
  MUX2_X1 U16179 ( .A(n14021), .B(P2_EBX_REG_3__SCAN_IN), .S(n14161), .Z(
        n14354) );
  AOI21_X1 U16180 ( .B1(n19245), .B2(n16307), .A(n14354), .ZN(n14355) );
  INV_X1 U16181 ( .A(n14355), .ZN(P2_U2884) );
  OAI222_X1 U16182 ( .A1(n15866), .A2(n21423), .B1(n15863), .B2(n22083), .C1(
        n19778), .C2(n15852), .ZN(P1_U2898) );
  NOR2_X1 U16183 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21549), .ZN(n14357) );
  AOI211_X1 U16184 ( .C1(n14357), .C2(n11847), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n14356), .ZN(n14358) );
  AOI21_X1 U16185 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21556), .A(n11213), 
        .ZN(n17055) );
  NOR2_X1 U16186 ( .A1(n14358), .A2(n17055), .ZN(n14359) );
  NOR2_X1 U16187 ( .A1(n14379), .A2(n21549), .ZN(n14360) );
  INV_X1 U16188 ( .A(n14362), .ZN(n14372) );
  NAND2_X1 U16189 ( .A1(n14364), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14368) );
  INV_X1 U16190 ( .A(n14368), .ZN(n14365) );
  NOR2_X1 U16191 ( .A1(n14373), .A2(n14365), .ZN(n14366) );
  AND2_X1 U16192 ( .A1(n21229), .A2(n21829), .ZN(n14367) );
  NOR2_X1 U16193 ( .A1(n14368), .A2(n14367), .ZN(n14369) );
  OAI22_X1 U16194 ( .A1(n19869), .A2(n21505), .B1(n21535), .B2(n14370), .ZN(
        n14387) );
  NAND2_X1 U16195 ( .A1(n14372), .A2(n14371), .ZN(n14445) );
  AND2_X2 U16196 ( .A1(n14663), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21517) );
  NAND2_X4 U16197 ( .A1(n14374), .A2(n14373), .ZN(n21453) );
  INV_X1 U16198 ( .A(n21453), .ZN(n21509) );
  NAND3_X1 U16199 ( .A1(n21509), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14377) );
  OAI221_X1 U16200 ( .B1(n21453), .B2(P1_REIP_REG_2__SCAN_IN), .C1(n21453), 
        .C2(P1_REIP_REG_1__SCAN_IN), .A(n14663), .ZN(n14375) );
  NAND2_X1 U16201 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n14375), .ZN(n14376) );
  OAI21_X1 U16202 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n14377), .A(n14376), .ZN(
        n14378) );
  AOI21_X1 U16203 ( .B1(n21517), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14378), .ZN(n14384) );
  AND2_X1 U16204 ( .A1(n14379), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14380) );
  INV_X1 U16205 ( .A(n14381), .ZN(n14382) );
  NAND2_X1 U16206 ( .A1(n21530), .A2(n14382), .ZN(n14383) );
  OAI211_X1 U16207 ( .C1(n14445), .C2(n14385), .A(n14384), .B(n14383), .ZN(
        n14386) );
  NOR2_X1 U16208 ( .A1(n14387), .A2(n14386), .ZN(n14388) );
  OAI21_X1 U16209 ( .B1(n14519), .B2(n14389), .A(n14388), .ZN(P1_U2837) );
  NOR2_X1 U16210 ( .A1(n21453), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U16211 ( .A1(n21530), .A2(n14390), .B1(n15550), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U16212 ( .A1(n21517), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14391) );
  OAI211_X1 U16213 ( .C1(n14445), .C2(n13964), .A(n14392), .B(n14391), .ZN(
        n14393) );
  NOR2_X1 U16214 ( .A1(n14406), .A2(n14393), .ZN(n14396) );
  AOI22_X1 U16215 ( .A1(n21490), .A2(n14394), .B1(n21529), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n14395) );
  OAI211_X1 U16216 ( .C1(n14519), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        P1_U2839) );
  INV_X1 U16217 ( .A(n14445), .ZN(n14522) );
  NOR2_X1 U16218 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n21453), .ZN(n14401) );
  OAI22_X1 U16219 ( .A1(n14399), .A2(n21505), .B1(n21535), .B2(n14398), .ZN(
        n14400) );
  AOI21_X1 U16220 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n14401), .A(n14400), .ZN(
        n14403) );
  NAND2_X1 U16221 ( .A1(n21517), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14402) );
  OAI211_X1 U16222 ( .C1(n21519), .C2(n14404), .A(n14403), .B(n14402), .ZN(
        n14405) );
  AOI21_X1 U16223 ( .B1(n11214), .B2(n14522), .A(n14405), .ZN(n14408) );
  OAI21_X1 U16224 ( .B1(n14406), .B2(n15550), .A(P1_REIP_REG_2__SCAN_IN), .ZN(
        n14407) );
  OAI211_X1 U16225 ( .C1(n14409), .C2(n14519), .A(n14408), .B(n14407), .ZN(
        P1_U2838) );
  INV_X1 U16226 ( .A(n15490), .ZN(n14414) );
  NAND2_X1 U16227 ( .A1(n14411), .A2(n14410), .ZN(n14412) );
  AND2_X1 U16228 ( .A1(n14465), .A2(n14412), .ZN(n16849) );
  INV_X1 U16229 ( .A(n16849), .ZN(n14413) );
  INV_X1 U16230 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17368) );
  OAI222_X1 U16231 ( .A1(n14684), .A2(n14414), .B1(n14413), .B2(n19348), .C1(
        n19496), .C2(n17368), .ZN(P2_U2905) );
  AND2_X1 U16232 ( .A1(n14416), .A2(n14415), .ZN(n14417) );
  OR2_X1 U16233 ( .A1(n14417), .A2(n14459), .ZN(n16911) );
  INV_X1 U16234 ( .A(n14418), .ZN(n14423) );
  INV_X1 U16235 ( .A(n14461), .ZN(n14421) );
  OAI211_X1 U16236 ( .C1(n14423), .C2(n14422), .A(n14421), .B(n16307), .ZN(
        n14425) );
  NAND2_X1 U16237 ( .A1(n14161), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14424) );
  OAI211_X1 U16238 ( .C1(n16911), .C2(n14161), .A(n14425), .B(n14424), .ZN(
        P2_U2877) );
  NAND3_X1 U16239 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n14447) );
  NOR2_X1 U16240 ( .A1(n14447), .A2(n19801), .ZN(n21424) );
  OAI21_X1 U16241 ( .B1(n21424), .B2(n21453), .A(n14663), .ZN(n14454) );
  NAND2_X1 U16242 ( .A1(n21509), .A2(n21424), .ZN(n14426) );
  OAI22_X1 U16243 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n14426), .B1(n21535), 
        .B2(n21272), .ZN(n14429) );
  AOI22_X1 U16244 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n21517), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(n21529), .ZN(n14427) );
  INV_X1 U16245 ( .A(n21495), .ZN(n15728) );
  OAI211_X1 U16246 ( .C1(n21519), .C2(n19873), .A(n14427), .B(n15728), .ZN(
        n14428) );
  AOI211_X1 U16247 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n14454), .A(n14429), .B(
        n14428), .ZN(n14430) );
  OAI21_X1 U16248 ( .B1(n14519), .B2(n19874), .A(n14430), .ZN(P1_U2835) );
  NAND2_X1 U16249 ( .A1(n14433), .A2(n14432), .ZN(n14434) );
  AND2_X1 U16250 ( .A1(n14431), .A2(n14434), .ZN(n21440) );
  INV_X1 U16251 ( .A(n21440), .ZN(n14441) );
  INV_X1 U16252 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14440) );
  NAND2_X1 U16253 ( .A1(n15580), .A2(n13546), .ZN(n14436) );
  MUX2_X1 U16254 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n14435) );
  AND2_X1 U16255 ( .A1(n14436), .A2(n14435), .ZN(n14437) );
  NOR2_X1 U16256 ( .A1(n14438), .A2(n14437), .ZN(n14439) );
  OR2_X1 U16257 ( .A1(n14490), .A2(n14439), .ZN(n21273) );
  OAI222_X1 U16258 ( .A1(n14441), .A2(n15783), .B1(n14440), .B2(n19870), .C1(
        n15785), .C2(n21273), .ZN(P1_U2865) );
  OAI222_X1 U16259 ( .A1(n15866), .A2(n14441), .B1(n15852), .B2(n11828), .C1(
        n15863), .C2(n22128), .ZN(P1_U2897) );
  OR2_X1 U16260 ( .A1(n21453), .A2(n21424), .ZN(n14446) );
  INV_X1 U16261 ( .A(n21715), .ZN(n21797) );
  OR2_X1 U16262 ( .A1(n14442), .A2(n21797), .ZN(n14444) );
  XNOR2_X1 U16263 ( .A(n14444), .B(n14443), .ZN(n17039) );
  OAI22_X1 U16264 ( .A1(n14447), .A2(n14446), .B1(n17039), .B2(n14445), .ZN(
        n14448) );
  AOI211_X1 U16265 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21495), .B(n14448), .ZN(n14456) );
  NOR2_X1 U16266 ( .A1(n14449), .A2(n21505), .ZN(n14453) );
  OAI22_X1 U16267 ( .A1(n14451), .A2(n21519), .B1(n21535), .B2(n14450), .ZN(
        n14452) );
  AOI211_X1 U16268 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n14454), .A(n14453), .B(
        n14452), .ZN(n14455) );
  OAI211_X1 U16269 ( .C1(n14519), .C2(n14457), .A(n14456), .B(n14455), .ZN(
        P1_U2836) );
  OR2_X1 U16270 ( .A1(n14459), .A2(n14458), .ZN(n14460) );
  NAND2_X1 U16271 ( .A1(n14506), .A2(n14460), .ZN(n18414) );
  NAND2_X1 U16272 ( .A1(n14461), .A2(n14462), .ZN(n14510) );
  OAI211_X1 U16273 ( .C1(n14461), .C2(n14462), .A(n14508), .B(n16307), .ZN(
        n14464) );
  NAND2_X1 U16274 ( .A1(n14161), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14463) );
  OAI211_X1 U16275 ( .C1(n18414), .C2(n14161), .A(n14464), .B(n14463), .ZN(
        P2_U2876) );
  AOI21_X1 U16276 ( .B1(n14466), .B2(n14465), .A(n11062), .ZN(n16834) );
  INV_X1 U16277 ( .A(n16834), .ZN(n18443) );
  OAI222_X1 U16278 ( .A1(n18443), .A2(n19348), .B1(n14684), .B2(n14467), .C1(
        n19496), .C2(n17372), .ZN(P2_U2904) );
  OR2_X1 U16279 ( .A1(n14469), .A2(n14468), .ZN(n14471) );
  NAND2_X1 U16280 ( .A1(n14471), .A2(n14470), .ZN(n14679) );
  XNOR2_X1 U16281 ( .A(n19162), .B(n14679), .ZN(n14478) );
  XNOR2_X1 U16282 ( .A(n14473), .B(n14472), .ZN(n19487) );
  AOI21_X1 U16283 ( .B1(n17313), .B2(n17320), .A(n14474), .ZN(n14475) );
  XOR2_X1 U16284 ( .A(n19487), .B(n14475), .Z(n19492) );
  NAND2_X1 U16285 ( .A1(n19492), .A2(n19491), .ZN(n19490) );
  NAND2_X1 U16286 ( .A1(n14475), .A2(n19487), .ZN(n14476) );
  NAND2_X1 U16287 ( .A1(n19490), .A2(n14476), .ZN(n14477) );
  NOR2_X1 U16288 ( .A1(n14477), .A2(n14478), .ZN(n14678) );
  AOI21_X1 U16289 ( .B1(n14478), .B2(n14477), .A(n14678), .ZN(n14481) );
  INV_X1 U16290 ( .A(n19436), .ZN(n16375) );
  AOI22_X1 U16291 ( .A1(n19489), .A2(n16375), .B1(n19579), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n14480) );
  INV_X1 U16292 ( .A(n14679), .ZN(n17318) );
  NAND2_X1 U16293 ( .A1(n17318), .A2(n19585), .ZN(n14479) );
  OAI211_X1 U16294 ( .C1(n14481), .C2(n19342), .A(n14480), .B(n14479), .ZN(
        P2_U2916) );
  AOI21_X1 U16295 ( .B1(n14483), .B2(n14431), .A(n14482), .ZN(n14876) );
  INV_X1 U16296 ( .A(n14876), .ZN(n14503) );
  INV_X1 U16297 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14497) );
  NAND2_X1 U16298 ( .A1(n15591), .A2(n14497), .ZN(n14488) );
  NAND2_X1 U16299 ( .A1(n14056), .A2(n14484), .ZN(n14486) );
  NAND2_X1 U16300 ( .A1(n13785), .A2(n14497), .ZN(n14485) );
  NAND3_X1 U16301 ( .A1(n14486), .A2(n15607), .A3(n14485), .ZN(n14487) );
  NAND2_X1 U16302 ( .A1(n14488), .A2(n14487), .ZN(n14489) );
  NAND2_X1 U16303 ( .A1(n14490), .A2(n14489), .ZN(n14542) );
  OR2_X1 U16304 ( .A1(n14490), .A2(n14489), .ZN(n14491) );
  NAND2_X1 U16305 ( .A1(n14542), .A2(n14491), .ZN(n21295) );
  INV_X1 U16306 ( .A(n21295), .ZN(n14492) );
  AOI22_X1 U16307 ( .A1(n19865), .A2(n14492), .B1(n15794), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14493) );
  OAI21_X1 U16308 ( .B1(n14503), .B2(n15796), .A(n14493), .ZN(P1_U2864) );
  NAND4_X1 U16309 ( .A1(n21424), .A2(P1_REIP_REG_7__SCAN_IN), .A3(
        P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14495) );
  INV_X1 U16310 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n19806) );
  NOR2_X1 U16311 ( .A1(n14495), .A2(n19806), .ZN(n14662) );
  OAI21_X1 U16312 ( .B1(n14662), .B2(n21453), .A(n14663), .ZN(n14555) );
  OR2_X1 U16313 ( .A1(n21453), .A2(n14662), .ZN(n14494) );
  OAI22_X1 U16314 ( .A1(n21535), .A2(n21295), .B1(n14495), .B2(n14494), .ZN(
        n14499) );
  AOI22_X1 U16315 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n21517), .B1(
        n14875), .B2(n21530), .ZN(n14496) );
  OAI211_X1 U16316 ( .C1(n21505), .C2(n14497), .A(n14496), .B(n15728), .ZN(
        n14498) );
  AOI211_X1 U16317 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n14555), .A(n14499), .B(
        n14498), .ZN(n14500) );
  OAI21_X1 U16318 ( .B1(n14503), .B2(n21537), .A(n14500), .ZN(P1_U2832) );
  INV_X1 U16319 ( .A(n14501), .ZN(n15837) );
  OAI222_X1 U16320 ( .A1(n14503), .A2(n15866), .B1(n14502), .B2(n15852), .C1(
        n15863), .C2(n15837), .ZN(P1_U2896) );
  INV_X1 U16321 ( .A(n14504), .ZN(n14505) );
  AOI21_X1 U16322 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n16877) );
  INV_X1 U16323 ( .A(n16877), .ZN(n14516) );
  INV_X1 U16324 ( .A(n14508), .ZN(n14513) );
  INV_X1 U16325 ( .A(n14547), .ZN(n14511) );
  OAI211_X1 U16326 ( .C1(n14513), .C2(n14512), .A(n14511), .B(n16307), .ZN(
        n14515) );
  NAND2_X1 U16327 ( .A1(n14161), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14514) );
  OAI211_X1 U16328 ( .C1(n14516), .C2(n14161), .A(n14515), .B(n14514), .ZN(
        P2_U2875) );
  NAND2_X2 U16329 ( .A1(n21453), .A2(n14663), .ZN(n21485) );
  AOI21_X1 U16330 ( .B1(n21544), .B2(n21519), .A(n14517), .ZN(n14521) );
  NOR2_X1 U16331 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  AOI211_X1 U16332 ( .C1(n14522), .C2(n16086), .A(n14521), .B(n14520), .ZN(
        n14524) );
  AOI22_X1 U16333 ( .A1(n21408), .A2(n21490), .B1(n21529), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n14523) );
  OAI211_X1 U16334 ( .C1(n15720), .C2(n14525), .A(n14524), .B(n14523), .ZN(
        P1_U2840) );
  XNOR2_X1 U16335 ( .A(n14610), .B(n14529), .ZN(n14612) );
  XNOR2_X1 U16336 ( .A(n14612), .B(n14611), .ZN(n17263) );
  NAND2_X1 U16337 ( .A1(n17318), .A2(n18628), .ZN(n14531) );
  AOI21_X1 U16338 ( .B1(n16807), .B2(n14526), .A(n18590), .ZN(n18636) );
  NOR2_X1 U16339 ( .A1(n16755), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18620) );
  INV_X1 U16340 ( .A(n18620), .ZN(n14527) );
  OAI211_X1 U16341 ( .C1(n18617), .C2(n18615), .A(n18636), .B(n14527), .ZN(
        n16929) );
  AOI211_X1 U16342 ( .C1(n18615), .C2(n18616), .A(n14528), .B(n18593), .ZN(
        n16937) );
  AOI22_X1 U16343 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16929), .B1(
        n16937), .B2(n14529), .ZN(n14530) );
  OAI211_X1 U16344 ( .C1(n13263), .C2(n18600), .A(n14531), .B(n14530), .ZN(
        n14536) );
  NOR2_X1 U16345 ( .A1(n14533), .A2(n14532), .ZN(n17262) );
  INV_X1 U16346 ( .A(n14534), .ZN(n17261) );
  NOR3_X1 U16347 ( .A1(n17262), .A2(n17261), .A3(n18608), .ZN(n14535) );
  AOI211_X1 U16348 ( .C1(n18625), .C2(n14021), .A(n14536), .B(n14535), .ZN(
        n14537) );
  OAI21_X1 U16349 ( .B1(n18614), .B2(n17263), .A(n14537), .ZN(P2_U3043) );
  OR2_X1 U16350 ( .A1(n14482), .A2(n14539), .ZN(n14540) );
  AND2_X1 U16351 ( .A1(n14538), .A2(n14540), .ZN(n14908) );
  MUX2_X1 U16352 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n14541) );
  NAND2_X1 U16353 ( .A1(n11517), .A2(n14541), .ZN(n14543) );
  INV_X1 U16354 ( .A(n14948), .ZN(n14965) );
  AOI21_X1 U16355 ( .B1(n14543), .B2(n14542), .A(n14965), .ZN(n14915) );
  AOI22_X1 U16356 ( .A1(n19865), .A2(n14915), .B1(n15794), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14544) );
  OAI21_X1 U16357 ( .B1(n14560), .B2(n15783), .A(n14544), .ZN(P1_U2863) );
  NAND2_X1 U16358 ( .A1(n14504), .A2(n14545), .ZN(n14546) );
  NAND2_X1 U16359 ( .A1(n14649), .A2(n14546), .ZN(n18431) );
  NAND2_X1 U16360 ( .A1(n14547), .A2(n14548), .ZN(n14654) );
  OAI211_X1 U16361 ( .C1(n14547), .C2(n14548), .A(n14652), .B(n16307), .ZN(
        n14550) );
  NAND2_X1 U16362 ( .A1(n14161), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14549) );
  OAI211_X1 U16363 ( .C1(n18431), .C2(n14161), .A(n14550), .B(n14549), .ZN(
        P2_U2874) );
  NOR2_X1 U16364 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21453), .ZN(n14554) );
  AOI22_X1 U16365 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n21529), .B1(n21490), .B2(
        n14915), .ZN(n14551) );
  OAI211_X1 U16366 ( .C1(n21544), .C2(n14552), .A(n14551), .B(n15728), .ZN(
        n14553) );
  AOI21_X1 U16367 ( .B1(n14554), .B2(n14662), .A(n14553), .ZN(n14557) );
  AOI22_X1 U16368 ( .A1(n14555), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n21530), 
        .B2(n14904), .ZN(n14556) );
  OAI211_X1 U16369 ( .C1(n14560), .C2(n21537), .A(n14557), .B(n14556), .ZN(
        P1_U2831) );
  AOI22_X1 U16370 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n19784), .B1(n19780), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14558) );
  OAI21_X1 U16371 ( .B1(n12026), .B2(n14578), .A(n14558), .ZN(P1_U2920) );
  INV_X1 U16372 ( .A(n14559), .ZN(n15831) );
  OAI222_X1 U16373 ( .A1(n14560), .A2(n15866), .B1(n19783), .B2(n15864), .C1(
        n15863), .C2(n15831), .ZN(P1_U2895) );
  AOI22_X1 U16374 ( .A1(n19780), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14561) );
  OAI21_X1 U16375 ( .B1(n14562), .B2(n14578), .A(n14561), .ZN(P1_U2913) );
  AOI22_X1 U16376 ( .A1(n21230), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14563) );
  OAI21_X1 U16377 ( .B1(n15825), .B2(n14578), .A(n14563), .ZN(P1_U2910) );
  AOI22_X1 U16378 ( .A1(n21230), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14564) );
  OAI21_X1 U16379 ( .B1(n14565), .B2(n14578), .A(n14564), .ZN(P1_U2911) );
  AOI22_X1 U16380 ( .A1(n21230), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14566) );
  OAI21_X1 U16381 ( .B1(n14567), .B2(n14578), .A(n14566), .ZN(P1_U2917) );
  AOI22_X1 U16382 ( .A1(n21230), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14568) );
  OAI21_X1 U16383 ( .B1(n15805), .B2(n14578), .A(n14568), .ZN(P1_U2907) );
  AOI22_X1 U16384 ( .A1(n21230), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14569) );
  OAI21_X1 U16385 ( .B1(n15812), .B2(n14578), .A(n14569), .ZN(P1_U2908) );
  AOI22_X1 U16386 ( .A1(n21230), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14570) );
  OAI21_X1 U16387 ( .B1(n15799), .B2(n14578), .A(n14570), .ZN(P1_U2906) );
  AOI22_X1 U16388 ( .A1(n21230), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14571) );
  OAI21_X1 U16389 ( .B1(n15819), .B2(n14578), .A(n14571), .ZN(P1_U2909) );
  AOI22_X1 U16390 ( .A1(n21230), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14572) );
  OAI21_X1 U16391 ( .B1(n14573), .B2(n14578), .A(n14572), .ZN(P1_U2914) );
  AOI22_X1 U16392 ( .A1(n21230), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14574) );
  OAI21_X1 U16393 ( .B1(n15836), .B2(n14578), .A(n14574), .ZN(P1_U2912) );
  AOI22_X1 U16394 ( .A1(n21230), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14575) );
  OAI21_X1 U16395 ( .B1(n14576), .B2(n14578), .A(n14575), .ZN(P1_U2915) );
  AOI22_X1 U16396 ( .A1(n21230), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14577) );
  OAI21_X1 U16397 ( .B1(n14579), .B2(n14578), .A(n14577), .ZN(P1_U2916) );
  INV_X1 U16398 ( .A(n14580), .ZN(n14581) );
  AOI21_X1 U16399 ( .B1(n14583), .B2(n14582), .A(n14581), .ZN(n16070) );
  INV_X1 U16400 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21426) );
  NOR2_X1 U16401 ( .A1(n21401), .A2(n21426), .ZN(n16071) );
  AOI21_X1 U16402 ( .B1(n19943), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16071), .ZN(n14586) );
  INV_X1 U16403 ( .A(n21432), .ZN(n14584) );
  NAND2_X1 U16404 ( .A1(n19927), .A2(n14584), .ZN(n14585) );
  OAI211_X1 U16405 ( .C1(n21423), .C2(n19915), .A(n14586), .B(n14585), .ZN(
        n14587) );
  AOI21_X1 U16406 ( .B1(n16070), .B2(n19949), .A(n14587), .ZN(n14588) );
  INV_X1 U16407 ( .A(n14588), .ZN(P1_U2993) );
  NAND2_X1 U16408 ( .A1(n17320), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19278) );
  OR2_X1 U16409 ( .A1(n17321), .A2(n19278), .ZN(n14590) );
  AND2_X1 U16410 ( .A1(n19225), .A2(n19272), .ZN(n14601) );
  INV_X1 U16411 ( .A(n14601), .ZN(n14589) );
  NAND2_X1 U16412 ( .A1(n14590), .A2(n14589), .ZN(n14599) );
  AOI21_X1 U16413 ( .B1(n16962), .B2(n19263), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18656) );
  AND2_X1 U16414 ( .A1(n17303), .A2(n18656), .ZN(n14592) );
  NAND2_X1 U16415 ( .A1(n14592), .A2(n19262), .ZN(n19284) );
  INV_X1 U16416 ( .A(n19284), .ZN(n19133) );
  NAND2_X1 U16417 ( .A1(n14602), .A2(n19133), .ZN(n14597) );
  INV_X1 U16418 ( .A(n14592), .ZN(n14593) );
  NAND3_X1 U16419 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19225), .A3(
        n19272), .ZN(n14606) );
  NAND2_X1 U16420 ( .A1(n19276), .A2(n14606), .ZN(n14595) );
  NAND2_X1 U16421 ( .A1(n19281), .A2(n14595), .ZN(n14596) );
  NAND2_X1 U16422 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  NAND2_X1 U16423 ( .A1(n14599), .A2(n14598), .ZN(n19666) );
  INV_X1 U16424 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15373) );
  NAND2_X1 U16425 ( .A1(n14601), .A2(n19282), .ZN(n14604) );
  INV_X1 U16426 ( .A(n14606), .ZN(n19664) );
  OAI21_X1 U16427 ( .B1(n14602), .B2(n19664), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14603) );
  NAND2_X1 U16428 ( .A1(n14604), .A2(n14603), .ZN(n19665) );
  INV_X1 U16429 ( .A(n19256), .ZN(n14605) );
  INV_X1 U16430 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20559) );
  INV_X1 U16431 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n22039) );
  OAI22_X1 U16432 ( .A1(n20559), .A2(n14782), .B1(n22039), .B2(n14783), .ZN(
        n19384) );
  INV_X1 U16433 ( .A(n19388), .ZN(n19380) );
  OAI22_X1 U16434 ( .A1(n19669), .A2(n19392), .B1(n19380), .B2(n14606), .ZN(
        n14608) );
  NOR2_X1 U16435 ( .A1(n19387), .A2(n19564), .ZN(n14607) );
  AOI211_X1 U16436 ( .C1(n14600), .C2(n19665), .A(n14608), .B(n14607), .ZN(
        n14609) );
  OAI21_X1 U16437 ( .B1(n19524), .B2(n15373), .A(n14609), .ZN(P2_U3093) );
  AOI22_X1 U16438 ( .A1(n14612), .A2(n14611), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14610), .ZN(n14614) );
  XNOR2_X1 U16439 ( .A(n14764), .B(n14838), .ZN(n14613) );
  XNOR2_X1 U16440 ( .A(n14614), .B(n14613), .ZN(n17275) );
  INV_X1 U16441 ( .A(n17275), .ZN(n14624) );
  XNOR2_X1 U16442 ( .A(n14615), .B(n14838), .ZN(n17271) );
  INV_X1 U16443 ( .A(n16929), .ZN(n14616) );
  OAI21_X1 U16444 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18593), .A(
        n14616), .ZN(n14841) );
  NAND2_X1 U16445 ( .A1(n14841), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14621) );
  AOI21_X1 U16446 ( .B1(n14617), .B2(n14470), .A(n14834), .ZN(n14767) );
  NAND2_X1 U16447 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16937), .ZN(
        n16948) );
  OAI22_X1 U16448 ( .A1(n18488), .A2(n14618), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16948), .ZN(n14619) );
  AOI21_X1 U16449 ( .B1(n18628), .B2(n14767), .A(n14619), .ZN(n14620) );
  OAI211_X1 U16450 ( .C1(n14763), .C2(n18607), .A(n14621), .B(n14620), .ZN(
        n14622) );
  AOI21_X1 U16451 ( .B1(n17271), .B2(n18623), .A(n14622), .ZN(n14623) );
  OAI21_X1 U16452 ( .B1(n14624), .B2(n18614), .A(n14623), .ZN(P2_U3042) );
  AOI21_X1 U16453 ( .B1(n17269), .B2(n14629), .A(n14702), .ZN(n17259) );
  INV_X1 U16454 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U16455 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14627), .B1(n18356), 
        .B2(n18340), .ZN(n18348) );
  AOI22_X1 U16456 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14628), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18340), .ZN(n16232) );
  NOR2_X1 U16457 ( .A1(n18348), .A2(n16232), .ZN(n16231) );
  OAI21_X1 U16458 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n14629), .ZN(n15532) );
  NAND2_X1 U16459 ( .A1(n16231), .A2(n15532), .ZN(n14700) );
  NAND2_X1 U16460 ( .A1(n10997), .A2(n14700), .ZN(n14630) );
  XNOR2_X1 U16461 ( .A(n17259), .B(n14630), .ZN(n14646) );
  NAND4_X1 U16462 ( .A1(n18340), .A2(n19263), .A3(n21569), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n18643) );
  NAND2_X1 U16463 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19263), .ZN(n18646) );
  NOR3_X1 U16464 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19262), .A3(n18646), 
        .ZN(n18649) );
  NOR4_X4 U16465 ( .A1(n18427), .A2(n18341), .A3(n18558), .A4(n18649), .ZN(
        n18528) );
  OAI22_X1 U16466 ( .A1(n17269), .A2(n18564), .B1(n13263), .B2(n18562), .ZN(
        n14645) );
  OR2_X1 U16467 ( .A1(n14633), .A2(n14632), .ZN(n16134) );
  INV_X1 U16468 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16247) );
  NAND2_X1 U16469 ( .A1(n21569), .A2(n18655), .ZN(n14637) );
  AND2_X1 U16470 ( .A1(n16247), .A2(n14637), .ZN(n14634) );
  NAND2_X1 U16471 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  NAND2_X2 U16472 ( .A1(n16134), .A2(n14636), .ZN(n18568) );
  NAND2_X1 U16473 ( .A1(n18341), .A2(n11287), .ZN(n14641) );
  INV_X1 U16474 ( .A(n14637), .ZN(n14638) );
  INV_X1 U16475 ( .A(n14639), .ZN(n14640) );
  AOI22_X1 U16476 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(n18568), .B1(n18572), .B2(
        n14640), .ZN(n14643) );
  NAND2_X1 U16477 ( .A1(n14021), .A2(n18570), .ZN(n14642) );
  OAI211_X1 U16478 ( .C1(n14679), .C2(n18576), .A(n14643), .B(n14642), .ZN(
        n14644) );
  AOI211_X1 U16479 ( .C1(n14646), .C2(n18558), .A(n14645), .B(n14644), .ZN(
        n14647) );
  OAI21_X1 U16480 ( .B1(n19162), .B2(n16244), .A(n14647), .ZN(P2_U2852) );
  INV_X1 U16481 ( .A(n14688), .ZN(n14651) );
  NAND2_X1 U16482 ( .A1(n14649), .A2(n14648), .ZN(n14650) );
  NAND2_X1 U16483 ( .A1(n14651), .A2(n14650), .ZN(n16851) );
  INV_X1 U16484 ( .A(n14652), .ZN(n14657) );
  INV_X1 U16485 ( .A(n14685), .ZN(n14655) );
  OAI211_X1 U16486 ( .C1(n14657), .C2(n14656), .A(n14655), .B(n16307), .ZN(
        n14659) );
  NAND2_X1 U16487 ( .A1(n14161), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14658) );
  OAI211_X1 U16488 ( .C1(n16851), .C2(n14161), .A(n14659), .B(n14658), .ZN(
        P2_U2873) );
  AOI21_X1 U16489 ( .B1(n14661), .B2(n14538), .A(n14660), .ZN(n19891) );
  INV_X1 U16490 ( .A(n19891), .ZN(n14695) );
  NAND2_X1 U16491 ( .A1(n14662), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14664) );
  INV_X1 U16492 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21297) );
  NOR2_X1 U16493 ( .A1(n14664), .A2(n21297), .ZN(n21444) );
  OAI21_X1 U16494 ( .B1(n21444), .B2(n21453), .A(n14663), .ZN(n21458) );
  OAI21_X1 U16495 ( .B1(n14664), .B2(n21453), .A(n21297), .ZN(n14674) );
  INV_X1 U16496 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U16497 ( .A1(n15591), .A2(n14670), .ZN(n14668) );
  INV_X1 U16498 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19885) );
  NAND2_X1 U16499 ( .A1(n14056), .A2(n19885), .ZN(n14666) );
  NAND2_X1 U16500 ( .A1(n13785), .A2(n14670), .ZN(n14665) );
  NAND3_X1 U16501 ( .A1(n14666), .A2(n15607), .A3(n14665), .ZN(n14667) );
  NAND2_X1 U16502 ( .A1(n14668), .A2(n14667), .ZN(n14964) );
  INV_X1 U16503 ( .A(n14964), .ZN(n14669) );
  XNOR2_X1 U16504 ( .A(n14948), .B(n14669), .ZN(n21296) );
  OAI22_X1 U16505 ( .A1(n14670), .A2(n21505), .B1(n21535), .B2(n21296), .ZN(
        n14671) );
  AOI211_X1 U16506 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n14671), .B(n21495), .ZN(n14672) );
  OAI21_X1 U16507 ( .B1(n19889), .B2(n21519), .A(n14672), .ZN(n14673) );
  AOI21_X1 U16508 ( .B1(n21458), .B2(n14674), .A(n14673), .ZN(n14675) );
  OAI21_X1 U16509 ( .B1(n14695), .B2(n21537), .A(n14675), .ZN(P1_U2830) );
  INV_X1 U16510 ( .A(n21296), .ZN(n14676) );
  AOI22_X1 U16511 ( .A1(n19865), .A2(n14676), .B1(n15794), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14677) );
  OAI21_X1 U16512 ( .B1(n14695), .B2(n15796), .A(n14677), .ZN(P1_U2862) );
  AOI21_X1 U16513 ( .B1(n19162), .B2(n14679), .A(n14678), .ZN(n14680) );
  NOR2_X1 U16514 ( .A1(n14680), .A2(n14767), .ZN(n19344) );
  XOR2_X1 U16515 ( .A(n19343), .B(n19344), .Z(n14681) );
  NAND2_X1 U16516 ( .A1(n14681), .A2(n19586), .ZN(n14683) );
  AOI22_X1 U16517 ( .A1(n19585), .A2(n14767), .B1(n19579), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14682) );
  OAI211_X1 U16518 ( .C1(n14748), .C2(n14684), .A(n14683), .B(n14682), .ZN(
        P2_U2915) );
  INV_X1 U16519 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14693) );
  OAI211_X1 U16520 ( .C1(n14685), .C2(n14686), .A(n14862), .B(n16307), .ZN(
        n14692) );
  OR2_X1 U16521 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  NAND2_X1 U16522 ( .A1(n14864), .A2(n14689), .ZN(n18444) );
  INV_X1 U16523 ( .A(n18444), .ZN(n14690) );
  NAND2_X1 U16524 ( .A1(n14690), .A2(n16284), .ZN(n14691) );
  OAI211_X1 U16525 ( .C1(n16284), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        P2_U2872) );
  INV_X1 U16526 ( .A(n14694), .ZN(n15826) );
  OAI222_X1 U16527 ( .A1(n14695), .A2(n15866), .B1(n19786), .B2(n15864), .C1(
        n15863), .C2(n15826), .ZN(P1_U2894) );
  INV_X1 U16528 ( .A(n14714), .ZN(n14696) );
  AOI21_X1 U16529 ( .B1(n18425), .B2(n14712), .A(n14696), .ZN(n18429) );
  NOR2_X1 U16530 ( .A1(n14709), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14697) );
  OR2_X1 U16531 ( .A1(n14710), .A2(n14697), .ZN(n18422) );
  INV_X1 U16532 ( .A(n18422), .ZN(n16604) );
  AND2_X1 U16533 ( .A1(n14705), .A2(n14698), .ZN(n14699) );
  NOR2_X1 U16534 ( .A1(n14707), .A2(n14699), .ZN(n18397) );
  AOI21_X1 U16535 ( .B1(n16641), .B2(n14703), .A(n14706), .ZN(n18386) );
  AOI21_X1 U16536 ( .B1(n14846), .B2(n14701), .A(n14704), .ZN(n18367) );
  NOR2_X1 U16537 ( .A1(n17259), .A2(n14700), .ZN(n14759) );
  OAI21_X1 U16538 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14702), .A(
        n14701), .ZN(n17278) );
  NAND2_X1 U16539 ( .A1(n14759), .A2(n17278), .ZN(n18365) );
  NOR2_X1 U16540 ( .A1(n18367), .A2(n18365), .ZN(n18377) );
  OAI21_X1 U16541 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n14704), .A(
        n14703), .ZN(n18378) );
  NAND2_X1 U16542 ( .A1(n18377), .A2(n18378), .ZN(n18385) );
  NOR2_X1 U16543 ( .A1(n18386), .A2(n18385), .ZN(n14725) );
  OAI21_X1 U16544 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n14706), .A(
        n14705), .ZN(n17300) );
  NAND2_X1 U16545 ( .A1(n14725), .A2(n17300), .ZN(n18396) );
  NOR2_X1 U16546 ( .A1(n18397), .A2(n18396), .ZN(n14797) );
  NOR2_X1 U16547 ( .A1(n14707), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14708) );
  OR2_X1 U16548 ( .A1(n14709), .A2(n14708), .ZN(n16618) );
  NAND2_X1 U16549 ( .A1(n14797), .A2(n16618), .ZN(n18417) );
  NOR2_X1 U16550 ( .A1(n16604), .A2(n18417), .ZN(n14825) );
  OR2_X1 U16551 ( .A1(n14710), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14711) );
  NAND2_X1 U16552 ( .A1(n14712), .A2(n14711), .ZN(n16592) );
  NAND2_X1 U16553 ( .A1(n14825), .A2(n16592), .ZN(n18428) );
  NOR2_X1 U16554 ( .A1(n18429), .A2(n18428), .ZN(n16112) );
  NOR2_X1 U16555 ( .A1(n18535), .A2(n16112), .ZN(n14716) );
  AND2_X1 U16556 ( .A1(n14714), .A2(n14713), .ZN(n14715) );
  OR2_X1 U16557 ( .A1(n14715), .A2(n16110), .ZN(n16571) );
  XNOR2_X1 U16558 ( .A(n14716), .B(n16571), .ZN(n14723) );
  AOI22_X1 U16559 ( .A1(n14717), .A2(n18572), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n18568), .ZN(n14718) );
  OAI211_X1 U16560 ( .C1(n16570), .C2(n18562), .A(n14718), .B(n18488), .ZN(
        n14719) );
  AOI21_X1 U16561 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18529), .A(
        n14719), .ZN(n14721) );
  NAND2_X1 U16562 ( .A1(n18531), .A2(n16849), .ZN(n14720) );
  OAI211_X1 U16563 ( .C1(n18511), .C2(n16851), .A(n14721), .B(n14720), .ZN(
        n14722) );
  AOI21_X1 U16564 ( .B1(n14723), .B2(n18558), .A(n14722), .ZN(n14724) );
  INV_X1 U16565 ( .A(n14724), .ZN(P2_U2841) );
  NOR2_X1 U16566 ( .A1(n18535), .A2(n14725), .ZN(n14726) );
  XNOR2_X1 U16567 ( .A(n14726), .B(n17300), .ZN(n14734) );
  NOR2_X1 U16568 ( .A1(n18511), .A2(n18606), .ZN(n14729) );
  AOI22_X1 U16569 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18528), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18529), .ZN(n14727) );
  OAI211_X1 U16570 ( .C1(n18576), .C2(n18602), .A(n14727), .B(n18600), .ZN(
        n14728) );
  NOR2_X1 U16571 ( .A1(n14729), .A2(n14728), .ZN(n14731) );
  NAND2_X1 U16572 ( .A1(n18568), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14730) );
  OAI211_X1 U16573 ( .C1(n18509), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14733) );
  AOI21_X1 U16574 ( .B1(n14734), .B2(n18558), .A(n14733), .ZN(n14735) );
  INV_X1 U16575 ( .A(n14735), .ZN(P2_U2847) );
  INV_X1 U16576 ( .A(n17320), .ZN(n14736) );
  NAND2_X1 U16577 ( .A1(n14736), .A2(n17305), .ZN(n19119) );
  NOR2_X2 U16578 ( .A1(n17321), .A2(n19119), .ZN(n19658) );
  OAI21_X1 U16579 ( .B1(n19658), .B2(n19659), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14740) );
  INV_X1 U16580 ( .A(n19146), .ZN(n19259) );
  NAND2_X1 U16581 ( .A1(n19259), .A2(n19225), .ZN(n14739) );
  NAND2_X1 U16582 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19225), .ZN(
        n19211) );
  NOR2_X1 U16583 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19211), .ZN(
        n19656) );
  AOI21_X1 U16584 ( .B1(n19656), .B2(n19281), .A(n19231), .ZN(n14738) );
  NAND2_X1 U16585 ( .A1(n14741), .A2(n19133), .ZN(n14737) );
  INV_X1 U16586 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14747) );
  INV_X1 U16587 ( .A(n19572), .ZN(n19575) );
  AOI22_X1 U16588 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n19598), .B1(
        BUF1_REG_17__SCAN_IN), .B2(n19597), .ZN(n19578) );
  AOI22_X1 U16589 ( .A1(n19659), .A2(n19575), .B1(n19658), .B2(n19569), .ZN(
        n14746) );
  OAI21_X1 U16590 ( .B1(n14741), .B2(n19656), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14743) );
  NAND3_X1 U16591 ( .A1(n19259), .A2(n19282), .A3(n19225), .ZN(n14742) );
  NAND2_X1 U16592 ( .A1(n14743), .A2(n14742), .ZN(n19657) );
  NOR2_X2 U16593 ( .A1(n14744), .A2(n19591), .ZN(n19574) );
  NOR2_X2 U16594 ( .A1(n15436), .A2(n14781), .ZN(n19573) );
  AOI22_X1 U16595 ( .A1(n19657), .A2(n19574), .B1(n19656), .B2(n19573), .ZN(
        n14745) );
  OAI211_X1 U16596 ( .C1(n19663), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        P2_U3097) );
  INV_X1 U16597 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U16598 ( .A1(n19659), .A2(n19432), .B1(n19658), .B2(n19427), .ZN(
        n14752) );
  NOR2_X2 U16599 ( .A1(n14750), .A2(n14781), .ZN(n19431) );
  AOI22_X1 U16600 ( .A1(n19657), .A2(n14749), .B1(n19656), .B2(n19431), .ZN(
        n14751) );
  OAI211_X1 U16601 ( .C1(n19663), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        P2_U3100) );
  INV_X1 U16602 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14758) );
  AOI22_X1 U16603 ( .A1(n19659), .A2(n19336), .B1(n19658), .B2(n19337), .ZN(
        n14757) );
  NOR2_X2 U16604 ( .A1(n15487), .A2(n14781), .ZN(n19335) );
  AOI22_X1 U16605 ( .A1(n19657), .A2(n14755), .B1(n19656), .B2(n19335), .ZN(
        n14756) );
  OAI211_X1 U16606 ( .C1(n19663), .C2(n14758), .A(n14757), .B(n14756), .ZN(
        P2_U3102) );
  INV_X1 U16607 ( .A(n17278), .ZN(n14762) );
  NOR2_X1 U16608 ( .A1(n18535), .A2(n14759), .ZN(n14761) );
  AOI21_X1 U16609 ( .B1(n14762), .B2(n14761), .A(n18643), .ZN(n14760) );
  OAI21_X1 U16610 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14772) );
  INV_X1 U16611 ( .A(n14763), .ZN(n17272) );
  INV_X1 U16612 ( .A(n14764), .ZN(n14769) );
  AOI22_X1 U16613 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18568), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18529), .ZN(n14765) );
  OAI211_X1 U16614 ( .C1(n14618), .C2(n18562), .A(n18600), .B(n14765), .ZN(
        n14766) );
  AOI21_X1 U16615 ( .B1(n18531), .B2(n14767), .A(n14766), .ZN(n14768) );
  OAI21_X1 U16616 ( .B1(n14769), .B2(n18509), .A(n14768), .ZN(n14770) );
  AOI21_X1 U16617 ( .B1(n17272), .B2(n18570), .A(n14770), .ZN(n14771) );
  OAI211_X1 U16618 ( .C1(n19343), .C2(n16244), .A(n14772), .B(n14771), .ZN(
        P2_U2851) );
  NOR2_X1 U16619 ( .A1(n19124), .A2(n19278), .ZN(n14777) );
  NAND3_X1 U16620 ( .A1(n19272), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19148) );
  INV_X1 U16621 ( .A(n19148), .ZN(n14776) );
  NOR2_X1 U16622 ( .A1(n19274), .A2(n19148), .ZN(n19609) );
  AOI21_X1 U16623 ( .B1(n19609), .B2(n19281), .A(n19231), .ZN(n14773) );
  OAI21_X1 U16624 ( .B1(n14774), .B2(n19284), .A(n14773), .ZN(n14775) );
  INV_X1 U16625 ( .A(n19611), .ZN(n14796) );
  INV_X1 U16626 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14787) );
  OAI21_X1 U16627 ( .B1(n14778), .B2(n19609), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14779) );
  OAI21_X1 U16628 ( .B1(n19148), .B2(n19276), .A(n14779), .ZN(n19610) );
  NAND2_X1 U16629 ( .A1(n12519), .A2(n19593), .ZN(n19226) );
  INV_X1 U16630 ( .A(n19609), .ZN(n19135) );
  NOR2_X2 U16631 ( .A1(n19124), .A2(n19182), .ZN(n19617) );
  INV_X1 U16632 ( .A(n19614), .ZN(n19500) );
  INV_X1 U16633 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n22135) );
  INV_X1 U16634 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n20636) );
  OAI22_X1 U16635 ( .A1(n22135), .A2(n14783), .B1(n20636), .B2(n14782), .ZN(
        n19292) );
  AOI22_X1 U16636 ( .A1(n19617), .A2(n19293), .B1(n19500), .B2(n19292), .ZN(
        n14784) );
  OAI21_X1 U16637 ( .B1(n19226), .B2(n19135), .A(n14784), .ZN(n14785) );
  AOI21_X1 U16638 ( .B1(n19610), .B2(n14780), .A(n14785), .ZN(n14786) );
  OAI21_X1 U16639 ( .B1(n14796), .B2(n14787), .A(n14786), .ZN(P2_U3159) );
  INV_X1 U16640 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14791) );
  INV_X1 U16641 ( .A(n19335), .ZN(n19316) );
  AOI22_X1 U16642 ( .A1(n19617), .A2(n19336), .B1(n19500), .B2(n19337), .ZN(
        n14788) );
  OAI21_X1 U16643 ( .B1(n19316), .B2(n19135), .A(n14788), .ZN(n14789) );
  AOI21_X1 U16644 ( .B1(n19610), .B2(n14755), .A(n14789), .ZN(n14790) );
  OAI21_X1 U16645 ( .B1(n14796), .B2(n14791), .A(n14790), .ZN(P2_U3158) );
  INV_X1 U16646 ( .A(n19573), .ZN(n19556) );
  AOI22_X1 U16647 ( .A1(n19617), .A2(n19575), .B1(n19500), .B2(n19569), .ZN(
        n14792) );
  OAI21_X1 U16648 ( .B1(n19556), .B2(n19135), .A(n14792), .ZN(n14793) );
  AOI21_X1 U16649 ( .B1(n19610), .B2(n19574), .A(n14793), .ZN(n14794) );
  OAI21_X1 U16650 ( .B1(n14796), .B2(n14795), .A(n14794), .ZN(P2_U3153) );
  NOR2_X1 U16651 ( .A1(n18535), .A2(n14797), .ZN(n14798) );
  XNOR2_X1 U16652 ( .A(n14798), .B(n16618), .ZN(n14799) );
  NAND2_X1 U16653 ( .A1(n14799), .A2(n18558), .ZN(n14807) );
  NAND2_X1 U16654 ( .A1(n14801), .A2(n14800), .ZN(n14802) );
  AND2_X1 U16655 ( .A1(n11070), .A2(n14802), .ZN(n16908) );
  INV_X1 U16656 ( .A(n16908), .ZN(n19118) );
  AOI22_X1 U16657 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n18528), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18529), .ZN(n14803) );
  OAI211_X1 U16658 ( .C1(n18576), .C2(n19118), .A(n14803), .B(n18600), .ZN(
        n14805) );
  NOR2_X1 U16659 ( .A1(n16911), .A2(n18511), .ZN(n14804) );
  AOI211_X1 U16660 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n18568), .A(n14805), .B(
        n14804), .ZN(n14806) );
  OAI211_X1 U16661 ( .C1(n18509), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        P2_U2845) );
  NOR2_X1 U16662 ( .A1(n18535), .A2(n16231), .ZN(n14809) );
  XNOR2_X1 U16663 ( .A(n14809), .B(n15532), .ZN(n14810) );
  NAND2_X1 U16664 ( .A1(n14810), .A2(n18558), .ZN(n14818) );
  AOI22_X1 U16665 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18529), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n18528), .ZN(n14811) );
  INV_X1 U16666 ( .A(n14811), .ZN(n14816) );
  INV_X1 U16667 ( .A(n18568), .ZN(n18516) );
  OAI22_X1 U16668 ( .A1(n18516), .A2(n12770), .B1(n14812), .B2(n18509), .ZN(
        n14813) );
  AOI21_X1 U16669 ( .B1(n18531), .B2(n19487), .A(n14813), .ZN(n14814) );
  OAI21_X1 U16670 ( .B1(n12609), .B2(n18511), .A(n14814), .ZN(n14815) );
  NOR2_X1 U16671 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  OAI211_X1 U16672 ( .C1(n16244), .C2(n17309), .A(n14818), .B(n14817), .ZN(
        P2_U2853) );
  NOR3_X1 U16673 ( .A1(n18535), .A2(n14825), .A3(n18643), .ZN(n18418) );
  INV_X1 U16674 ( .A(n14819), .ZN(n14824) );
  NOR2_X1 U16675 ( .A1(n18576), .A2(n16880), .ZN(n14822) );
  AOI22_X1 U16676 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18529), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18568), .ZN(n14820) );
  OAI211_X1 U16677 ( .C1(n16590), .C2(n18562), .A(n18600), .B(n14820), .ZN(
        n14821) );
  AOI211_X1 U16678 ( .C1(n16877), .C2(n18570), .A(n14822), .B(n14821), .ZN(
        n14823) );
  OAI21_X1 U16679 ( .B1(n14824), .B2(n18509), .A(n14823), .ZN(n14828) );
  NOR2_X1 U16680 ( .A1(n18535), .A2(n14825), .ZN(n14826) );
  NOR3_X1 U16681 ( .A1(n14826), .A2(n18643), .A3(n16592), .ZN(n14827) );
  AOI211_X1 U16682 ( .C1(n18418), .C2(n16592), .A(n14828), .B(n14827), .ZN(
        n14829) );
  INV_X1 U16683 ( .A(n14829), .ZN(P2_U2843) );
  XNOR2_X1 U16684 ( .A(n14830), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14832) );
  XNOR2_X1 U16685 ( .A(n14832), .B(n14831), .ZN(n14851) );
  NAND2_X1 U16686 ( .A1(n14833), .A2(n12818), .ZN(n14844) );
  NAND3_X1 U16687 ( .A1(n13066), .A2(n18623), .A3(n14844), .ZN(n14843) );
  XNOR2_X1 U16688 ( .A(n14835), .B(n14834), .ZN(n19347) );
  INV_X1 U16689 ( .A(n19347), .ZN(n14836) );
  AOI22_X1 U16690 ( .A1(n18628), .A2(n14836), .B1(n18427), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n14837) );
  OAI21_X1 U16691 ( .B1(n18607), .B2(n14845), .A(n14837), .ZN(n14840) );
  AOI211_X1 U16692 ( .C1(n14838), .C2(n12818), .A(n16947), .B(n16948), .ZN(
        n14839) );
  AOI211_X1 U16693 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n14841), .A(
        n14840), .B(n14839), .ZN(n14842) );
  OAI211_X1 U16694 ( .C1(n14851), .C2(n18614), .A(n14843), .B(n14842), .ZN(
        P2_U3041) );
  NAND3_X1 U16695 ( .A1(n13066), .A2(n17270), .A3(n14844), .ZN(n14850) );
  NOR2_X1 U16696 ( .A1(n17296), .A2(n14845), .ZN(n14848) );
  OAI22_X1 U16697 ( .A1(n14846), .A2(n17268), .B1(n13225), .B2(n18488), .ZN(
        n14847) );
  AOI211_X1 U16698 ( .C1(n17260), .C2(n18367), .A(n14848), .B(n14847), .ZN(
        n14849) );
  OAI211_X1 U16699 ( .C1(n17295), .C2(n14851), .A(n14850), .B(n14849), .ZN(
        P2_U3009) );
  INV_X1 U16700 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U16701 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U16702 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U16703 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14853) );
  AOI22_X1 U16704 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14852) );
  NAND4_X1 U16705 ( .A1(n14855), .A2(n14854), .A3(n14853), .A4(n14852), .ZN(
        n14861) );
  AOI22_X1 U16706 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14859) );
  AOI22_X1 U16707 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14858) );
  AOI22_X1 U16708 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14857) );
  AOI22_X1 U16709 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14856) );
  NAND4_X1 U16710 ( .A1(n14859), .A2(n14858), .A3(n14857), .A4(n14856), .ZN(
        n14860) );
  NOR2_X1 U16711 ( .A1(n14861), .A2(n14860), .ZN(n14863) );
  AOI21_X1 U16712 ( .B1(n14863), .B2(n14862), .A(n11061), .ZN(n19587) );
  NAND2_X1 U16713 ( .A1(n19587), .A2(n16307), .ZN(n14867) );
  XOR2_X1 U16714 ( .A(n14865), .B(n14864), .Z(n18457) );
  NAND2_X1 U16715 ( .A1(n18457), .A2(n16284), .ZN(n14866) );
  OAI211_X1 U16716 ( .C1(n16284), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        P2_U2871) );
  INV_X1 U16717 ( .A(n14869), .ZN(n14870) );
  AOI21_X1 U16718 ( .B1(n14872), .B2(n14871), .A(n14870), .ZN(n21285) );
  OAI22_X1 U16719 ( .A1(n19901), .A2(n14873), .B1(n21401), .B2(n19806), .ZN(
        n14874) );
  AOI21_X1 U16720 ( .B1(n14875), .B2(n19927), .A(n14874), .ZN(n14878) );
  NAND2_X1 U16721 ( .A1(n14876), .A2(n19948), .ZN(n14877) );
  OAI211_X1 U16722 ( .C1(n21285), .C2(n21546), .A(n14878), .B(n14877), .ZN(
        P1_U2991) );
  INV_X1 U16723 ( .A(n19257), .ZN(n19279) );
  OAI21_X1 U16724 ( .B1(n19701), .B2(n19705), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14879) );
  NAND2_X1 U16725 ( .A1(n14879), .A2(n19282), .ZN(n14888) );
  NOR2_X1 U16726 ( .A1(n14880), .A2(n19154), .ZN(n19595) );
  INV_X1 U16727 ( .A(n14881), .ZN(n14882) );
  NOR2_X1 U16728 ( .A1(n14882), .A2(n19284), .ZN(n14883) );
  OAI22_X1 U16729 ( .A1(n14888), .A2(n19595), .B1(n19231), .B2(n14883), .ZN(
        n14884) );
  NOR2_X1 U16730 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19224) );
  NOR2_X1 U16731 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19273) );
  NAND2_X1 U16732 ( .A1(n19224), .A2(n19273), .ZN(n14885) );
  INV_X1 U16733 ( .A(n14885), .ZN(n19699) );
  NOR2_X1 U16734 ( .A1(n19595), .A2(n19699), .ZN(n14887) );
  OAI21_X1 U16735 ( .B1(n14881), .B2(n19699), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14886) );
  INV_X1 U16736 ( .A(n19701), .ZN(n14897) );
  AOI22_X1 U16737 ( .A1(n19705), .A2(n19389), .B1(n19699), .B2(n19388), .ZN(
        n14889) );
  OAI21_X1 U16738 ( .B1(n14897), .B2(n19392), .A(n14889), .ZN(n14890) );
  AOI21_X1 U16739 ( .B1(n19703), .B2(n14600), .A(n14890), .ZN(n14891) );
  OAI21_X1 U16740 ( .B1(n19709), .B2(n15371), .A(n14891), .ZN(P2_U3053) );
  AOI22_X1 U16741 ( .A1(n19705), .A2(n19432), .B1(n19431), .B2(n19699), .ZN(
        n14892) );
  OAI21_X1 U16742 ( .B1(n14897), .B2(n19435), .A(n14892), .ZN(n14893) );
  AOI21_X1 U16743 ( .B1(n19703), .B2(n14749), .A(n14893), .ZN(n14894) );
  OAI21_X1 U16744 ( .B1(n19709), .B2(n14895), .A(n14894), .ZN(P2_U3052) );
  INV_X1 U16745 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U16746 ( .A1(n19705), .A2(n19575), .B1(n19573), .B2(n19699), .ZN(
        n14896) );
  OAI21_X1 U16747 ( .B1(n14897), .B2(n19578), .A(n14896), .ZN(n14898) );
  AOI21_X1 U16748 ( .B1(n19703), .B2(n19574), .A(n14898), .ZN(n14899) );
  OAI21_X1 U16749 ( .B1(n19709), .B2(n15304), .A(n14899), .ZN(P2_U3049) );
  NAND2_X1 U16750 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  NAND2_X1 U16751 ( .A1(n19884), .A2(n14902), .ZN(n14918) );
  INV_X1 U16752 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14903) );
  NOR2_X1 U16753 ( .A1(n21401), .A2(n14903), .ZN(n14914) );
  AOI21_X1 U16754 ( .B1(n19943), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n14914), .ZN(n14906) );
  NAND2_X1 U16755 ( .A1(n19927), .A2(n14904), .ZN(n14905) );
  NAND2_X1 U16756 ( .A1(n14906), .A2(n14905), .ZN(n14907) );
  AOI21_X1 U16757 ( .B1(n14908), .B2(n19948), .A(n14907), .ZN(n14909) );
  OAI21_X1 U16758 ( .B1(n14918), .B2(n21546), .A(n14909), .ZN(P1_U2990) );
  INV_X1 U16759 ( .A(n21263), .ZN(n16073) );
  NAND2_X1 U16760 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16073), .ZN(
        n16076) );
  NOR2_X1 U16761 ( .A1(n14235), .A2(n16076), .ZN(n21283) );
  NAND2_X1 U16762 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21283), .ZN(
        n21286) );
  NOR2_X1 U16763 ( .A1(n14484), .A2(n21286), .ZN(n14912) );
  NAND2_X1 U16764 ( .A1(n14912), .A2(n21276), .ZN(n15979) );
  NAND3_X1 U16765 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14912), .ZN(n15976) );
  INV_X1 U16766 ( .A(n21328), .ZN(n14910) );
  AOI22_X1 U16767 ( .A1(n21325), .A2(n15979), .B1(n15976), .B2(n14910), .ZN(
        n14911) );
  NAND2_X1 U16768 ( .A1(n21327), .A2(n14911), .ZN(n21299) );
  AND2_X1 U16769 ( .A1(n21282), .A2(n14912), .ZN(n21301) );
  AOI22_X1 U16770 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21299), .B1(
        n21301), .B2(n14913), .ZN(n14917) );
  AOI21_X1 U16771 ( .B1(n21409), .B2(n14915), .A(n14914), .ZN(n14916) );
  OAI211_X1 U16772 ( .C1(n14918), .C2(n21335), .A(n14917), .B(n14916), .ZN(
        P1_U3022) );
  AOI22_X1 U16773 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U16774 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U16775 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14920) );
  AOI22_X1 U16776 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14919) );
  NAND4_X1 U16777 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        n14928) );
  AOI22_X1 U16778 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12725), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14926) );
  AOI22_X1 U16779 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n13274), .B1(
        n12699), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U16780 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U16781 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14923) );
  NAND4_X1 U16782 ( .A1(n14926), .A2(n14925), .A3(n14924), .A4(n14923), .ZN(
        n14927) );
  OR2_X1 U16783 ( .A1(n14928), .A2(n14927), .ZN(n14929) );
  OAI21_X1 U16784 ( .B1(n11061), .B2(n14929), .A(n14983), .ZN(n16379) );
  AND2_X1 U16785 ( .A1(n11081), .A2(n14930), .ZN(n14931) );
  OR2_X1 U16786 ( .A1(n14931), .A2(n14971), .ZN(n18467) );
  NOR2_X1 U16787 ( .A1(n18467), .A2(n14161), .ZN(n14932) );
  AOI21_X1 U16788 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n14161), .A(n14932), .ZN(
        n14933) );
  OAI21_X1 U16789 ( .B1(n16379), .B2(n16302), .A(n14933), .ZN(P2_U2870) );
  INV_X1 U16790 ( .A(n14660), .ZN(n14935) );
  NAND2_X1 U16791 ( .A1(n14935), .A2(n11450), .ZN(n14936) );
  NAND2_X1 U16792 ( .A1(n14937), .A2(n14936), .ZN(n14961) );
  OAI21_X1 U16793 ( .B1(n14961), .B2(n14962), .A(n14937), .ZN(n15020) );
  AND2_X1 U16794 ( .A1(n15020), .A2(n15021), .ZN(n15022) );
  INV_X1 U16795 ( .A(n14938), .ZN(n14939) );
  INV_X1 U16796 ( .A(n14941), .ZN(n15972) );
  INV_X1 U16797 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U16798 ( .A1(n21444), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n21454) );
  INV_X1 U16799 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21305) );
  NOR2_X1 U16800 ( .A1(n21454), .A2(n21305), .ZN(n14942) );
  NAND2_X1 U16801 ( .A1(n14942), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15708) );
  OAI211_X1 U16802 ( .C1(n14942), .C2(P1_REIP_REG_13__SCAN_IN), .A(n21509), 
        .B(n15708), .ZN(n14943) );
  OAI21_X1 U16803 ( .B1(n21505), .B2(n14944), .A(n14943), .ZN(n14959) );
  INV_X1 U16804 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21309) );
  NAND2_X1 U16805 ( .A1(n15580), .A2(n21309), .ZN(n14946) );
  MUX2_X1 U16806 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14945) );
  AND2_X1 U16807 ( .A1(n14946), .A2(n14945), .ZN(n14963) );
  NAND2_X1 U16808 ( .A1(n14963), .A2(n14964), .ZN(n14947) );
  MUX2_X1 U16809 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14949) );
  NAND2_X1 U16810 ( .A1(n11521), .A2(n14949), .ZN(n14953) );
  OAI21_X1 U16811 ( .B1(n10968), .B2(n21255), .A(n14056), .ZN(n14950) );
  OAI21_X1 U16812 ( .B1(n13878), .B2(P1_EBX_REG_12__SCAN_IN), .A(n14950), .ZN(
        n14952) );
  INV_X1 U16813 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U16814 ( .A1(n15591), .A2(n15030), .ZN(n14951) );
  INV_X1 U16815 ( .A(n15027), .ZN(n14955) );
  INV_X1 U16816 ( .A(n14953), .ZN(n14954) );
  AOI21_X1 U16817 ( .B1(n15028), .B2(n14955), .A(n14954), .ZN(n14956) );
  OR2_X1 U16818 ( .A1(n14995), .A2(n14956), .ZN(n14999) );
  INV_X1 U16819 ( .A(n14999), .ZN(n21247) );
  AOI22_X1 U16820 ( .A1(n15550), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n21490), 
        .B2(n21247), .ZN(n14957) );
  OAI211_X1 U16821 ( .C1(n21544), .C2(n15970), .A(n14957), .B(n15728), .ZN(
        n14958) );
  AOI211_X1 U16822 ( .C1(n21530), .C2(n15972), .A(n14959), .B(n14958), .ZN(
        n14960) );
  OAI21_X1 U16823 ( .B1(n15975), .B2(n21537), .A(n14960), .ZN(P1_U2827) );
  XOR2_X1 U16824 ( .A(n14962), .B(n14961), .Z(n21448) );
  INV_X1 U16825 ( .A(n21448), .ZN(n14969) );
  INV_X1 U16826 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14967) );
  AOI21_X1 U16827 ( .B1(n14965), .B2(n14964), .A(n14963), .ZN(n14966) );
  OR2_X1 U16828 ( .A1(n14966), .A2(n15028), .ZN(n21445) );
  OAI222_X1 U16829 ( .A1(n14969), .A2(n15783), .B1(n14967), .B2(n19870), .C1(
        n15785), .C2(n21445), .ZN(P1_U2861) );
  INV_X1 U16830 ( .A(n14968), .ZN(n15820) );
  OAI222_X1 U16831 ( .A1(n14969), .A2(n15866), .B1(n19788), .B2(n15852), .C1(
        n15863), .C2(n15820), .ZN(P1_U2893) );
  OR2_X1 U16832 ( .A1(n14971), .A2(n14970), .ZN(n14972) );
  NAND2_X1 U16833 ( .A1(n11074), .A2(n14972), .ZN(n18479) );
  AOI22_X1 U16834 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14976) );
  AOI22_X1 U16835 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16836 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U16837 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14973) );
  NAND4_X1 U16838 ( .A1(n14976), .A2(n14975), .A3(n14974), .A4(n14973), .ZN(
        n14982) );
  AOI22_X1 U16839 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14980) );
  AOI22_X1 U16840 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14979) );
  AOI22_X1 U16841 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16842 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14977) );
  NAND4_X1 U16843 ( .A1(n14980), .A2(n14979), .A3(n14978), .A4(n14977), .ZN(
        n14981) );
  NOR2_X1 U16844 ( .A1(n14982), .A2(n14981), .ZN(n14984) );
  AOI21_X1 U16845 ( .B1(n14984), .B2(n14983), .A(n15014), .ZN(n19483) );
  NAND2_X1 U16846 ( .A1(n19483), .A2(n16307), .ZN(n14986) );
  NAND2_X1 U16847 ( .A1(n14161), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14985) );
  OAI211_X1 U16848 ( .C1(n18479), .C2(n14161), .A(n14986), .B(n14985), .ZN(
        P2_U2869) );
  OR2_X1 U16849 ( .A1(n14938), .A2(n14988), .ZN(n14989) );
  AND2_X1 U16850 ( .A1(n14987), .A2(n14989), .ZN(n21468) );
  INV_X1 U16851 ( .A(n21468), .ZN(n15003) );
  INV_X1 U16852 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21465) );
  NAND2_X1 U16853 ( .A1(n15591), .A2(n21465), .ZN(n14993) );
  INV_X1 U16854 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21261) );
  NAND2_X1 U16855 ( .A1(n14056), .A2(n21261), .ZN(n14991) );
  NAND2_X1 U16856 ( .A1(n13785), .A2(n21465), .ZN(n14990) );
  NAND3_X1 U16857 ( .A1(n14991), .A2(n15607), .A3(n14990), .ZN(n14992) );
  NAND2_X1 U16858 ( .A1(n14993), .A2(n14992), .ZN(n14994) );
  OR2_X1 U16859 ( .A1(n14995), .A2(n14994), .ZN(n14996) );
  NAND2_X1 U16860 ( .A1(n11012), .A2(n14996), .ZN(n21464) );
  INV_X1 U16861 ( .A(n21464), .ZN(n14997) );
  AOI22_X1 U16862 ( .A1(n19865), .A2(n14997), .B1(n15794), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14998) );
  OAI21_X1 U16863 ( .B1(n15003), .B2(n15783), .A(n14998), .ZN(P1_U2858) );
  OAI222_X1 U16864 ( .A1(n15975), .A2(n15783), .B1(n14944), .B2(n19870), .C1(
        n15785), .C2(n14999), .ZN(P1_U2859) );
  INV_X1 U16865 ( .A(n15000), .ZN(n15806) );
  OAI222_X1 U16866 ( .A1(n15866), .A2(n15975), .B1(n15863), .B2(n15806), .C1(
        n15001), .C2(n15852), .ZN(P1_U2891) );
  INV_X1 U16867 ( .A(n15002), .ZN(n15800) );
  OAI222_X1 U16868 ( .A1(n15003), .A2(n15866), .B1(n19792), .B2(n15864), .C1(
        n15863), .C2(n15800), .ZN(P1_U2890) );
  AOI22_X1 U16869 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U16870 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16871 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U16872 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15004) );
  NAND4_X1 U16873 ( .A1(n15007), .A2(n15006), .A3(n15005), .A4(n15004), .ZN(
        n15013) );
  AOI22_X1 U16874 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15011) );
  AOI22_X1 U16875 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15010) );
  AOI22_X1 U16876 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U16877 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15008) );
  NAND4_X1 U16878 ( .A1(n15011), .A2(n15010), .A3(n15009), .A4(n15008), .ZN(
        n15012) );
  NAND2_X2 U16879 ( .A1(n15014), .A2(n15015), .ZN(n16305) );
  OAI21_X1 U16880 ( .B1(n15014), .B2(n15015), .A(n16305), .ZN(n16378) );
  NAND2_X1 U16881 ( .A1(n14161), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U16882 ( .A1(n11074), .A2(n15016), .ZN(n15017) );
  NAND2_X1 U16883 ( .A1(n11018), .A2(n15017), .ZN(n18493) );
  INV_X1 U16884 ( .A(n18493), .ZN(n16781) );
  NAND2_X1 U16885 ( .A1(n16781), .A2(n16284), .ZN(n15018) );
  OAI211_X1 U16886 ( .C1(n16378), .C2(n16302), .A(n15019), .B(n15018), .ZN(
        P2_U2868) );
  INV_X1 U16887 ( .A(n15020), .ZN(n15024) );
  INV_X1 U16888 ( .A(n15021), .ZN(n15023) );
  AOI21_X1 U16889 ( .B1(n15024), .B2(n15023), .A(n15022), .ZN(n21456) );
  INV_X1 U16890 ( .A(n21456), .ZN(n15031) );
  INV_X1 U16891 ( .A(n15025), .ZN(n15813) );
  OAI222_X1 U16892 ( .A1(n15031), .A2(n15866), .B1(n15026), .B2(n15864), .C1(
        n15863), .C2(n15813), .ZN(P1_U2892) );
  XNOR2_X1 U16893 ( .A(n15028), .B(n15027), .ZN(n21452) );
  INV_X1 U16894 ( .A(n21452), .ZN(n15029) );
  OAI222_X1 U16895 ( .A1(n15031), .A2(n15783), .B1(n15030), .B2(n19870), .C1(
        n15785), .C2(n15029), .ZN(P1_U2860) );
  INV_X1 U16896 ( .A(n15788), .ZN(n15032) );
  AOI21_X1 U16897 ( .B1(n15033), .B2(n14987), .A(n15032), .ZN(n21480) );
  INV_X1 U16898 ( .A(n21480), .ZN(n15865) );
  MUX2_X1 U16899 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n15034) );
  NAND2_X1 U16900 ( .A1(n11518), .A2(n15034), .ZN(n15035) );
  AOI21_X1 U16901 ( .B1(n15035), .B2(n11012), .A(n11401), .ZN(n21479) );
  AOI22_X1 U16902 ( .A1(n21479), .A2(n19865), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15794), .ZN(n15036) );
  OAI21_X1 U16903 ( .B1(n15865), .B2(n15783), .A(n15036), .ZN(P1_U2857) );
  NOR2_X2 U16904 ( .A1(n20727), .A2(n15038), .ZN(n15054) );
  AOI22_X1 U16905 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15037) );
  OAI21_X1 U16906 ( .B1(n11019), .B2(n17712), .A(n15037), .ZN(n15047) );
  AOI22_X1 U16907 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15045) );
  AOI22_X1 U16908 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15044) );
  AOI22_X1 U16909 ( .A1(n10970), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U16910 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15042) );
  NAND4_X1 U16911 ( .A1(n15045), .A2(n15044), .A3(n15043), .A4(n15042), .ZN(
        n15046) );
  AOI22_X1 U16912 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15063) );
  AOI22_X1 U16913 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15062) );
  INV_X1 U16914 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15053) );
  AOI22_X1 U16915 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15052) );
  OAI21_X1 U16916 ( .B1(n11019), .B2(n15053), .A(n15052), .ZN(n15060) );
  AOI22_X1 U16917 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15058) );
  BUF_X4 U16918 ( .A(n15054), .Z(n17764) );
  AOI22_X1 U16919 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U16920 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U16921 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15055) );
  NAND4_X1 U16922 ( .A1(n15058), .A2(n15057), .A3(n15056), .A4(n15055), .ZN(
        n15059) );
  INV_X2 U16923 ( .A(n11021), .ZN(n17736) );
  AOI22_X1 U16924 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15064) );
  OAI21_X1 U16925 ( .B1(n11019), .B2(n17414), .A(n15064), .ZN(n15072) );
  AOI22_X1 U16926 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U16927 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U16928 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15068) );
  AOI22_X1 U16929 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15067) );
  NAND4_X1 U16930 ( .A1(n15070), .A2(n15069), .A3(n15068), .A4(n15067), .ZN(
        n15071) );
  AOI22_X1 U16931 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U16932 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U16933 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15078) );
  OAI21_X1 U16934 ( .B1(n11019), .B2(n17725), .A(n15078), .ZN(n15085) );
  AOI22_X1 U16935 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U16936 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15082) );
  AOI22_X1 U16937 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15081) );
  AOI22_X1 U16938 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15080) );
  NAND4_X1 U16939 ( .A1(n15083), .A2(n15082), .A3(n15081), .A4(n15080), .ZN(
        n15084) );
  AOI211_X1 U16940 ( .C1(n17764), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15085), .B(n15084), .ZN(n15086) );
  NAND3_X1 U16941 ( .A1(n15088), .A2(n15087), .A3(n15086), .ZN(n15128) );
  AOI22_X1 U16942 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15098) );
  AOI22_X1 U16943 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U16944 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15090) );
  OAI21_X1 U16945 ( .B1(n11019), .B2(n17739), .A(n15090), .ZN(n15096) );
  AOI22_X1 U16946 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U16947 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U16948 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U16949 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U16950 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15107) );
  AOI22_X1 U16951 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15106) );
  AOI22_X1 U16952 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15099) );
  OAI21_X1 U16953 ( .B1(n11019), .B2(n17420), .A(n15099), .ZN(n15105) );
  AOI22_X1 U16954 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U16955 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U16956 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U16957 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15100) );
  NAND4_X1 U16958 ( .A1(n15103), .A2(n15102), .A3(n15101), .A4(n15100), .ZN(
        n15104) );
  AOI22_X1 U16959 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15079), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15111) );
  AOI22_X1 U16960 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U16961 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U16962 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15108) );
  NAND4_X1 U16963 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15117) );
  AOI22_X1 U16964 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16965 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U16966 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U16967 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15112) );
  NAND4_X1 U16968 ( .A1(n15115), .A2(n15114), .A3(n15113), .A4(n15112), .ZN(
        n15116) );
  AOI22_X1 U16969 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15066), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15127) );
  AOI22_X1 U16970 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15126) );
  INV_X1 U16971 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U16972 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15118) );
  OAI21_X1 U16973 ( .B1(n11019), .B2(n17396), .A(n15118), .ZN(n15124) );
  AOI22_X1 U16974 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15122) );
  AOI22_X1 U16975 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U16976 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U16977 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15119) );
  NAND4_X1 U16978 ( .A1(n15122), .A2(n15121), .A3(n15120), .A4(n15119), .ZN(
        n15123) );
  AOI211_X1 U16979 ( .C1(n15079), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n15124), .B(n15123), .ZN(n15125) );
  NAND3_X1 U16980 ( .A1(n15127), .A2(n15126), .A3(n15125), .ZN(n15245) );
  INV_X1 U16981 ( .A(n15245), .ZN(n18883) );
  NAND2_X1 U16982 ( .A1(n20746), .A2(n18883), .ZN(n20690) );
  NOR2_X1 U16983 ( .A1(n15260), .A2(n20690), .ZN(n15244) );
  AND3_X1 U16984 ( .A1(n20671), .A2(n20748), .A3(n15244), .ZN(n15142) );
  NAND2_X1 U16985 ( .A1(n20557), .A2(n20746), .ZN(n20737) );
  NAND2_X1 U16986 ( .A1(n15128), .A2(n20736), .ZN(n20691) );
  AOI21_X1 U16987 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20680), .A(
        n15256), .ZN(n17786) );
  INV_X1 U16988 ( .A(n17786), .ZN(n15141) );
  OAI22_X1 U16989 ( .A1(n20712), .A2(n21169), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15255) );
  AOI22_X1 U16990 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n21174), .B2(n21165), .ZN(
        n15138) );
  AND2_X1 U16991 ( .A1(n15256), .A2(n15255), .ZN(n15129) );
  OR2_X1 U16992 ( .A1(n15138), .A2(n15139), .ZN(n15130) );
  OAI21_X1 U16993 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21165), .A(
        n15130), .ZN(n15131) );
  OAI22_X1 U16994 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21176), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15131), .ZN(n15133) );
  NOR2_X1 U16995 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21176), .ZN(
        n15132) );
  NAND2_X1 U16996 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15131), .ZN(
        n15134) );
  AOI22_X1 U16997 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15133), .B1(
        n15132), .B2(n15134), .ZN(n15136) );
  NAND2_X1 U16998 ( .A1(n15255), .A2(n15136), .ZN(n15140) );
  AOI21_X1 U16999 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15134), .A(
        n15133), .ZN(n15135) );
  OAI21_X1 U17000 ( .B1(n15139), .B2(n15138), .A(n15136), .ZN(n15137) );
  AOI21_X1 U17001 ( .B1(n15139), .B2(n15138), .A(n15137), .ZN(n17787) );
  INV_X1 U17002 ( .A(n17787), .ZN(n15258) );
  OAI221_X1 U17003 ( .B1(n15142), .B2(n17785), .C1(n15142), .C2(n17788), .A(
        n21221), .ZN(n20494) );
  NOR3_X1 U17004 ( .A1(n20063), .A2(n20055), .A3(n20494), .ZN(n17655) );
  INV_X1 U17005 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20304) );
  INV_X1 U17006 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20125) );
  NAND2_X1 U17007 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n17433) );
  NAND4_X1 U17008 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_13__SCAN_IN), .ZN(n15144)
         );
  AND4_X1 U17009 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n17393) );
  AND2_X1 U17010 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17393), .ZN(n17392) );
  AND3_X1 U17011 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .ZN(n17412) );
  NAND4_X1 U17012 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(n17392), .A4(n17412), .ZN(n15143) );
  NOR4_X1 U17013 ( .A1(n20125), .A2(n17433), .A3(n15144), .A4(n15143), .ZN(
        n17651) );
  NAND2_X1 U17014 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17651), .ZN(n17649) );
  NOR2_X1 U17015 ( .A1(n20304), .A2(n17649), .ZN(n17610) );
  AND2_X1 U17016 ( .A1(n17655), .A2(n17610), .ZN(n17623) );
  NAND3_X1 U17017 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17623), .ZN(n17535) );
  NAND4_X1 U17018 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .A4(P3_EBX_REG_25__SCAN_IN), .ZN(n15146)
         );
  NAND4_X1 U17019 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n15145)
         );
  NOR3_X1 U17020 ( .A1(n17535), .A2(n15146), .A3(n15145), .ZN(n17552) );
  NAND3_X1 U17021 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(P3_EBX_REG_29__SCAN_IN), 
        .A3(n17552), .ZN(n17534) );
  INV_X1 U17022 ( .A(n17534), .ZN(n17533) );
  AOI21_X1 U17023 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17552), .A(
        P3_EBX_REG_30__SCAN_IN), .ZN(n15147) );
  NOR2_X1 U17024 ( .A1(n17533), .A2(n15147), .ZN(n15241) );
  AOI22_X1 U17025 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U17026 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U17027 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15149) );
  AOI22_X1 U17028 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15148) );
  NAND4_X1 U17029 ( .A1(n15151), .A2(n15150), .A3(n15149), .A4(n15148), .ZN(
        n15157) );
  AOI22_X1 U17030 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U17031 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U17032 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U17033 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15152) );
  NAND4_X1 U17034 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15156) );
  NOR2_X1 U17035 ( .A1(n15157), .A2(n15156), .ZN(n17555) );
  AOI22_X1 U17036 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U17037 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15160) );
  AOI22_X1 U17038 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U17039 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15158) );
  NAND4_X1 U17040 ( .A1(n15161), .A2(n15160), .A3(n15159), .A4(n15158), .ZN(
        n15167) );
  AOI22_X1 U17041 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U17042 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U17043 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U17044 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15162) );
  NAND4_X1 U17045 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15166) );
  NOR2_X1 U17046 ( .A1(n15167), .A2(n15166), .ZN(n17549) );
  AOI22_X1 U17047 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15171) );
  AOI22_X1 U17048 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15170) );
  AOI22_X1 U17049 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U17050 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15168) );
  NAND4_X1 U17051 ( .A1(n15171), .A2(n15170), .A3(n15169), .A4(n15168), .ZN(
        n15177) );
  AOI22_X1 U17052 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U17053 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U17054 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U17055 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15172) );
  NAND4_X1 U17056 ( .A1(n15175), .A2(n15174), .A3(n15173), .A4(n15172), .ZN(
        n15176) );
  NOR2_X1 U17057 ( .A1(n15177), .A2(n15176), .ZN(n17570) );
  AOI22_X1 U17058 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U17059 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15180) );
  AOI22_X1 U17060 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15179) );
  AOI22_X1 U17061 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15178) );
  NAND4_X1 U17062 ( .A1(n15181), .A2(n15180), .A3(n15179), .A4(n15178), .ZN(
        n15187) );
  AOI22_X1 U17063 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15185) );
  AOI22_X1 U17064 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15184) );
  AOI22_X1 U17065 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U17066 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15182) );
  NAND4_X1 U17067 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15186) );
  NOR2_X1 U17068 ( .A1(n15187), .A2(n15186), .ZN(n17580) );
  AOI22_X1 U17069 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U17070 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U17071 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10993), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U17072 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15188) );
  NAND4_X1 U17073 ( .A1(n15191), .A2(n15190), .A3(n15189), .A4(n15188), .ZN(
        n15197) );
  AOI22_X1 U17074 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U17075 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U17076 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U17077 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15192) );
  NAND4_X1 U17078 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        n15196) );
  NOR2_X1 U17079 ( .A1(n15197), .A2(n15196), .ZN(n17581) );
  NOR2_X1 U17080 ( .A1(n17580), .A2(n17581), .ZN(n17579) );
  AOI22_X1 U17081 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10993), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17741), .ZN(n15207) );
  AOI22_X1 U17082 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17722), .ZN(n15206) );
  AOI22_X1 U17083 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10969), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15198) );
  OAI21_X1 U17084 ( .B1(n11021), .B2(n17712), .A(n15198), .ZN(n15204) );
  AOI22_X1 U17085 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15202) );
  AOI22_X1 U17086 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15201) );
  AOI22_X1 U17087 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17737), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U17088 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10971), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17687), .ZN(n15199) );
  NAND4_X1 U17089 ( .A1(n15202), .A2(n15201), .A3(n15200), .A4(n15199), .ZN(
        n15203) );
  AOI211_X1 U17090 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n10976), .A(
        n15204), .B(n15203), .ZN(n15205) );
  NAND3_X1 U17091 ( .A1(n15207), .A2(n15206), .A3(n15205), .ZN(n17575) );
  NAND2_X1 U17092 ( .A1(n17579), .A2(n17575), .ZN(n17574) );
  NOR2_X1 U17093 ( .A1(n17570), .A2(n17574), .ZN(n17569) );
  AOI22_X1 U17094 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15218) );
  AOI22_X1 U17095 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15217) );
  AOI22_X1 U17096 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15209) );
  OAI21_X1 U17097 ( .B1(n11021), .B2(n17396), .A(n15209), .ZN(n15215) );
  AOI22_X1 U17098 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15213) );
  AOI22_X1 U17099 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15212) );
  AOI22_X1 U17100 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15211) );
  AOI22_X1 U17101 ( .A1(n15066), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15210) );
  NAND4_X1 U17102 ( .A1(n15213), .A2(n15212), .A3(n15211), .A4(n15210), .ZN(
        n15214) );
  AOI211_X1 U17103 ( .C1(n17759), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15215), .B(n15214), .ZN(n15216) );
  NAND3_X1 U17104 ( .A1(n15218), .A2(n15217), .A3(n15216), .ZN(n17566) );
  NAND2_X1 U17105 ( .A1(n17569), .A2(n17566), .ZN(n17565) );
  NOR2_X1 U17106 ( .A1(n17549), .A2(n17565), .ZN(n17561) );
  AOI22_X1 U17107 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U17108 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U17109 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15219) );
  OAI21_X1 U17110 ( .B1(n11021), .B2(n17420), .A(n15219), .ZN(n15225) );
  AOI22_X1 U17111 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15223) );
  AOI22_X1 U17112 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15222) );
  AOI22_X1 U17113 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15221) );
  AOI22_X1 U17114 ( .A1(n10969), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15220) );
  NAND4_X1 U17115 ( .A1(n15223), .A2(n15222), .A3(n15221), .A4(n15220), .ZN(
        n15224) );
  AOI211_X1 U17116 ( .C1(n17759), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15225), .B(n15224), .ZN(n15226) );
  NAND3_X1 U17117 ( .A1(n15228), .A2(n15227), .A3(n15226), .ZN(n17560) );
  NAND2_X1 U17118 ( .A1(n17561), .A2(n17560), .ZN(n17559) );
  NOR2_X1 U17119 ( .A1(n17555), .A2(n17559), .ZN(n17554) );
  AOI22_X1 U17120 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15232) );
  AOI22_X1 U17121 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15231) );
  AOI22_X1 U17122 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U17123 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15229) );
  NAND4_X1 U17124 ( .A1(n15232), .A2(n15231), .A3(n15230), .A4(n15229), .ZN(
        n15238) );
  AOI22_X1 U17125 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15236) );
  AOI22_X1 U17126 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U17127 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U17128 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15233) );
  NAND4_X1 U17129 ( .A1(n15236), .A2(n15235), .A3(n15234), .A4(n15233), .ZN(
        n15237) );
  NOR2_X1 U17130 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  XOR2_X1 U17131 ( .A(n17554), .B(n15239), .Z(n20608) );
  INV_X1 U17132 ( .A(n20608), .ZN(n15240) );
  NOR2_X2 U17133 ( .A1(n17657), .A2(n20671), .ZN(n17658) );
  MUX2_X1 U17134 ( .A(n15241), .B(n15240), .S(n17658), .Z(P3_U2673) );
  NAND2_X1 U17135 ( .A1(n20557), .A2(n20558), .ZN(n20734) );
  NAND4_X1 U17136 ( .A1(n18883), .A2(n20748), .A3(n15246), .A4(n15249), .ZN(
        n20719) );
  NAND2_X1 U17137 ( .A1(n20738), .A2(n20055), .ZN(n15247) );
  NOR2_X1 U17138 ( .A1(n20719), .A2(n20746), .ZN(n15262) );
  AOI21_X1 U17139 ( .B1(n20055), .B2(n20746), .A(n20678), .ZN(n15269) );
  NAND2_X1 U17140 ( .A1(n20746), .A2(n20748), .ZN(n15268) );
  OAI211_X1 U17141 ( .C1(n20558), .C2(n15268), .A(n15245), .B(n20737), .ZN(
        n15242) );
  NAND2_X1 U17142 ( .A1(n20063), .A2(n15243), .ZN(n21196) );
  NAND3_X1 U17143 ( .A1(n20063), .A2(n15246), .A3(n15244), .ZN(n17784) );
  NAND2_X1 U17144 ( .A1(n20592), .A2(n20506), .ZN(n20499) );
  NAND3_X1 U17145 ( .A1(n20063), .A2(n20495), .A3(n20499), .ZN(n15267) );
  OAI21_X1 U17146 ( .B1(n15246), .B2(n15245), .A(n15267), .ZN(n15252) );
  NOR2_X1 U17147 ( .A1(n20671), .A2(n15249), .ZN(n15250) );
  NAND2_X1 U17148 ( .A1(n15247), .A2(n20746), .ZN(n15265) );
  INV_X1 U17149 ( .A(n15265), .ZN(n15248) );
  OAI22_X1 U17150 ( .A1(n20748), .A2(n15250), .B1(n15249), .B2(n15248), .ZN(
        n15251) );
  NOR3_X1 U17151 ( .A1(n15253), .A2(n15252), .A3(n15251), .ZN(n17783) );
  INV_X1 U17152 ( .A(n17783), .ZN(n20717) );
  INV_X1 U17153 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20100) );
  OAI21_X1 U17154 ( .B1(n15254), .B2(n20712), .A(n20100), .ZN(n16977) );
  NAND2_X1 U17155 ( .A1(n20681), .A2(n16977), .ZN(n21161) );
  NOR2_X1 U17156 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20728) );
  INV_X1 U17157 ( .A(n20728), .ZN(n20703) );
  NOR2_X1 U17158 ( .A1(n21161), .A2(n20703), .ZN(n15272) );
  INV_X1 U17159 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21625) );
  OR2_X2 U17160 ( .A1(n21625), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18326) );
  INV_X1 U17161 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21622) );
  NOR2_X1 U17162 ( .A1(n21622), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n21615) );
  INV_X1 U17163 ( .A(n21615), .ZN(n21619) );
  NAND2_X1 U17164 ( .A1(n20739), .A2(n16992), .ZN(n16990) );
  NAND2_X1 U17165 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21198) );
  INV_X1 U17166 ( .A(n21198), .ZN(n21628) );
  XNOR2_X1 U17167 ( .A(n15256), .B(n15255), .ZN(n15259) );
  AOI211_X1 U17168 ( .C1(n20497), .C2(n16990), .A(n21628), .B(n20741), .ZN(
        n15270) );
  INV_X1 U17169 ( .A(n17782), .ZN(n15261) );
  OAI211_X1 U17170 ( .C1(n20678), .C2(n20748), .A(n15261), .B(n15260), .ZN(
        n15264) );
  INV_X1 U17171 ( .A(n15262), .ZN(n15263) );
  OAI21_X1 U17172 ( .B1(n15265), .B2(n15264), .A(n15263), .ZN(n15266) );
  OAI211_X1 U17173 ( .C1(n15269), .C2(n15268), .A(n15267), .B(n15266), .ZN(
        n20743) );
  NOR2_X1 U17174 ( .A1(n21208), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18692) );
  INV_X1 U17175 ( .A(n18692), .ZN(n15271) );
  INV_X1 U17176 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20685) );
  INV_X1 U17177 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21075) );
  NAND2_X1 U17178 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17662), .ZN(n21206) );
  INV_X1 U17179 ( .A(n21206), .ZN(n16988) );
  NAND2_X1 U17180 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n16988), .ZN(n16978) );
  INV_X1 U17181 ( .A(n20730), .ZN(n20733) );
  MUX2_X1 U17182 ( .A(n15272), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20733), .Z(P3_U3284) );
  AOI22_X1 U17183 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12684), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15276) );
  AOI22_X1 U17184 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12743), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15275) );
  AOI22_X1 U17185 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n12835), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U17186 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15273) );
  NAND4_X1 U17187 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15282) );
  AOI22_X1 U17188 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U17189 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15279) );
  AOI22_X1 U17190 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U17191 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15277) );
  NAND4_X1 U17192 ( .A1(n15280), .A2(n15279), .A3(n15278), .A4(n15277), .ZN(
        n15281) );
  OR2_X1 U17193 ( .A1(n15282), .A2(n15281), .ZN(n15422) );
  AOI22_X1 U17194 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15293) );
  AOI22_X1 U17195 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U17196 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15291) );
  INV_X1 U17197 ( .A(n15466), .ZN(n15450) );
  INV_X1 U17198 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15288) );
  NAND2_X1 U17199 ( .A1(n10983), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n15287) );
  INV_X1 U17200 ( .A(n15284), .ZN(n15286) );
  NAND2_X1 U17201 ( .A1(n15286), .A2(n15285), .ZN(n15474) );
  OAI211_X1 U17202 ( .C1(n15450), .C2(n15288), .A(n15287), .B(n15474), .ZN(
        n15289) );
  INV_X1 U17203 ( .A(n15289), .ZN(n15290) );
  NAND4_X1 U17204 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15302) );
  AOI22_X1 U17205 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U17206 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U17207 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15298) );
  INV_X1 U17208 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15295) );
  INV_X1 U17209 ( .A(n15474), .ZN(n15465) );
  NAND2_X1 U17210 ( .A1(n12503), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n15294) );
  OAI211_X1 U17211 ( .C1(n15450), .C2(n15295), .A(n15465), .B(n15294), .ZN(
        n15296) );
  INV_X1 U17212 ( .A(n15296), .ZN(n15297) );
  NAND4_X1 U17213 ( .A1(n15300), .A2(n15299), .A3(n15298), .A4(n15297), .ZN(
        n15301) );
  NAND2_X1 U17214 ( .A1(n15302), .A2(n15301), .ZN(n15423) );
  INV_X1 U17215 ( .A(n15423), .ZN(n15303) );
  NAND2_X1 U17216 ( .A1(n15422), .A2(n15303), .ZN(n15424) );
  AOI22_X1 U17217 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15475), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15311) );
  AOI22_X1 U17218 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15310) );
  AOI22_X1 U17219 ( .A1(n10983), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15309) );
  INV_X1 U17220 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15306) );
  OR2_X1 U17221 ( .A1(n12431), .A2(n15304), .ZN(n15305) );
  OAI211_X1 U17222 ( .C1(n15450), .C2(n15306), .A(n15305), .B(n15474), .ZN(
        n15307) );
  INV_X1 U17223 ( .A(n15307), .ZN(n15308) );
  NAND4_X1 U17224 ( .A1(n15311), .A2(n15310), .A3(n15309), .A4(n15308), .ZN(
        n15321) );
  AOI22_X1 U17225 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15475), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U17226 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15318) );
  AOI22_X1 U17227 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15317) );
  OR2_X1 U17228 ( .A1(n15470), .A2(n15312), .ZN(n15313) );
  OAI211_X1 U17229 ( .C1(n15450), .C2(n15314), .A(n15313), .B(n15465), .ZN(
        n15315) );
  INV_X1 U17230 ( .A(n15315), .ZN(n15316) );
  NAND4_X1 U17231 ( .A1(n15319), .A2(n15318), .A3(n15317), .A4(n15316), .ZN(
        n15320) );
  NAND2_X1 U17232 ( .A1(n15321), .A2(n15320), .ZN(n15427) );
  NOR2_X1 U17233 ( .A1(n15424), .A2(n15427), .ZN(n15428) );
  AOI22_X1 U17234 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15328) );
  AOI22_X1 U17235 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15327) );
  AOI22_X1 U17236 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15326) );
  INV_X1 U17237 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15323) );
  NAND2_X1 U17238 ( .A1(n10983), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n15322) );
  OAI211_X1 U17239 ( .C1(n15450), .C2(n15323), .A(n15474), .B(n15322), .ZN(
        n15324) );
  INV_X1 U17240 ( .A(n15324), .ZN(n15325) );
  NAND4_X1 U17241 ( .A1(n15328), .A2(n15327), .A3(n15326), .A4(n15325), .ZN(
        n15337) );
  AOI22_X1 U17242 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15335) );
  AOI22_X1 U17243 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15334) );
  AOI22_X1 U17244 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15333) );
  INV_X1 U17245 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15330) );
  NAND2_X1 U17246 ( .A1(n12503), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n15329) );
  OAI211_X1 U17247 ( .C1(n15450), .C2(n15330), .A(n15465), .B(n15329), .ZN(
        n15331) );
  INV_X1 U17248 ( .A(n15331), .ZN(n15332) );
  NAND4_X1 U17249 ( .A1(n15335), .A2(n15334), .A3(n15333), .A4(n15332), .ZN(
        n15336) );
  AND2_X1 U17250 ( .A1(n15337), .A2(n15336), .ZN(n15430) );
  NAND2_X1 U17251 ( .A1(n15428), .A2(n15430), .ZN(n15433) );
  AOI22_X1 U17252 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15344) );
  AOI22_X1 U17253 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15343) );
  AOI22_X1 U17254 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15342) );
  INV_X1 U17255 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15339) );
  NAND2_X1 U17256 ( .A1(n12503), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n15338) );
  OAI211_X1 U17257 ( .C1(n15450), .C2(n15339), .A(n15474), .B(n15338), .ZN(
        n15340) );
  INV_X1 U17258 ( .A(n15340), .ZN(n15341) );
  NAND4_X1 U17259 ( .A1(n15344), .A2(n15343), .A3(n15342), .A4(n15341), .ZN(
        n15353) );
  AOI22_X1 U17260 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U17261 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15350) );
  AOI22_X1 U17262 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15349) );
  INV_X1 U17263 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15346) );
  NAND2_X1 U17264 ( .A1(n10983), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n15345) );
  OAI211_X1 U17265 ( .C1(n15450), .C2(n15346), .A(n15465), .B(n15345), .ZN(
        n15347) );
  INV_X1 U17266 ( .A(n15347), .ZN(n15348) );
  NAND4_X1 U17267 ( .A1(n15351), .A2(n15350), .A3(n15349), .A4(n15348), .ZN(
        n15352) );
  AND2_X1 U17268 ( .A1(n15353), .A2(n15352), .ZN(n15435) );
  INV_X1 U17269 ( .A(n15435), .ZN(n15354) );
  OR2_X1 U17270 ( .A1(n15433), .A2(n15354), .ZN(n15438) );
  AOI22_X1 U17271 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U17272 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15360) );
  AOI22_X1 U17273 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15359) );
  INV_X1 U17274 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15356) );
  NAND2_X1 U17275 ( .A1(n12503), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n15355) );
  OAI211_X1 U17276 ( .C1(n15450), .C2(n15356), .A(n15355), .B(n15474), .ZN(
        n15357) );
  INV_X1 U17277 ( .A(n15357), .ZN(n15358) );
  NAND4_X1 U17278 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15370) );
  AOI22_X1 U17279 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U17280 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15367) );
  AOI22_X1 U17281 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15366) );
  INV_X1 U17282 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U17283 ( .A1(n10982), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n15362) );
  OAI211_X1 U17284 ( .C1(n15450), .C2(n15363), .A(n15465), .B(n15362), .ZN(
        n15364) );
  INV_X1 U17285 ( .A(n15364), .ZN(n15365) );
  NAND4_X1 U17286 ( .A1(n15368), .A2(n15367), .A3(n15366), .A4(n15365), .ZN(
        n15369) );
  NAND2_X1 U17287 ( .A1(n15370), .A2(n15369), .ZN(n15442) );
  AOI22_X1 U17288 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15378) );
  AOI22_X1 U17289 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15377) );
  AOI22_X1 U17290 ( .A1(n12503), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15376) );
  OR2_X1 U17291 ( .A1(n12431), .A2(n15371), .ZN(n15372) );
  OAI211_X1 U17292 ( .C1(n12627), .C2(n15373), .A(n15372), .B(n15474), .ZN(
        n15374) );
  INV_X1 U17293 ( .A(n15374), .ZN(n15375) );
  NAND4_X1 U17294 ( .A1(n15378), .A2(n15377), .A3(n15376), .A4(n15375), .ZN(
        n15387) );
  AOI22_X1 U17295 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15475), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U17296 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U17297 ( .A1(n15466), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15383) );
  NAND2_X1 U17298 ( .A1(n10983), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n15379) );
  OAI211_X1 U17299 ( .C1(n10991), .C2(n15380), .A(n15465), .B(n15379), .ZN(
        n15381) );
  INV_X1 U17300 ( .A(n15381), .ZN(n15382) );
  NAND4_X1 U17301 ( .A1(n15385), .A2(n15384), .A3(n15383), .A4(n15382), .ZN(
        n15386) );
  AND2_X1 U17302 ( .A1(n15387), .A2(n15386), .ZN(n16256) );
  NAND2_X1 U17303 ( .A1(n18335), .A2(n16256), .ZN(n15388) );
  NOR2_X1 U17304 ( .A1(n16255), .A2(n15388), .ZN(n16251) );
  AOI22_X1 U17305 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15392) );
  AOI22_X1 U17306 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U17307 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U17308 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15389) );
  NAND4_X1 U17309 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        n15398) );
  AOI22_X1 U17310 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12725), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U17311 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15395) );
  AOI22_X1 U17312 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U17313 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15393) );
  NAND4_X1 U17314 ( .A1(n15396), .A2(n15395), .A3(n15394), .A4(n15393), .ZN(
        n15397) );
  NOR2_X1 U17315 ( .A1(n15398), .A2(n15397), .ZN(n16306) );
  AOI22_X1 U17316 ( .A1(n12684), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U17317 ( .A1(n12743), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12694), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15401) );
  AOI22_X1 U17318 ( .A1(n12835), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U17319 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15399) );
  NAND4_X1 U17320 ( .A1(n15402), .A2(n15401), .A3(n15400), .A4(n15399), .ZN(
        n15408) );
  AOI22_X1 U17321 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15406) );
  AOI22_X1 U17322 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15405) );
  AOI22_X1 U17323 ( .A1(n12672), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U17324 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15403) );
  NAND4_X1 U17325 ( .A1(n15406), .A2(n15405), .A3(n15404), .A4(n15403), .ZN(
        n15407) );
  OR2_X1 U17326 ( .A1(n15408), .A2(n15407), .ZN(n16296) );
  AOI22_X1 U17327 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12834), .B1(
        n12684), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U17328 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12694), .B1(
        n12743), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U17329 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12726), .B1(
        n12835), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15411) );
  AOI22_X1 U17330 ( .A1(n12656), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15409), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15410) );
  NAND4_X1 U17331 ( .A1(n15413), .A2(n15412), .A3(n15411), .A4(n15410), .ZN(
        n15421) );
  AOI22_X1 U17332 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12725), .B1(
        n15414), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U17333 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12699), .B1(
        n13274), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U17334 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12672), .B1(
        n15415), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U17335 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12673), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15416) );
  NAND4_X1 U17336 ( .A1(n15419), .A2(n15418), .A3(n15417), .A4(n15416), .ZN(
        n15420) );
  XOR2_X1 U17337 ( .A(n15423), .B(n15422), .Z(n16283) );
  INV_X1 U17338 ( .A(n15424), .ZN(n15425) );
  NAND2_X1 U17339 ( .A1(n15439), .A2(n15425), .ZN(n15426) );
  AOI22_X1 U17340 ( .A1(n15427), .A2(n15426), .B1(n15428), .B2(n18335), .ZN(
        n16279) );
  OAI211_X1 U17341 ( .C1(n15428), .C2(n15430), .A(n15439), .B(n15433), .ZN(
        n15432) );
  INV_X1 U17342 ( .A(n15430), .ZN(n15431) );
  NOR2_X1 U17343 ( .A1(n18335), .A2(n15431), .ZN(n16271) );
  NAND2_X1 U17344 ( .A1(n16272), .A2(n16271), .ZN(n16270) );
  NAND2_X1 U17345 ( .A1(n16270), .A2(n11526), .ZN(n15437) );
  XNOR2_X1 U17346 ( .A(n15433), .B(n15435), .ZN(n15434) );
  NAND2_X1 U17347 ( .A1(n15436), .A2(n15435), .ZN(n16266) );
  INV_X1 U17348 ( .A(n15438), .ZN(n15441) );
  INV_X1 U17349 ( .A(n15442), .ZN(n15440) );
  OAI211_X1 U17350 ( .C1(n15441), .C2(n15440), .A(n15439), .B(n16255), .ZN(
        n15443) );
  NOR2_X1 U17351 ( .A1(n18335), .A2(n15442), .ZN(n16262) );
  AOI22_X1 U17352 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15445) );
  AOI22_X1 U17353 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U17354 ( .A1(n15445), .A2(n15444), .ZN(n15459) );
  AOI22_X1 U17355 ( .A1(n15462), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15447) );
  AOI21_X1 U17356 ( .B1(n15475), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n15474), .ZN(n15446) );
  OAI211_X1 U17357 ( .C1(n15470), .C2(n15448), .A(n15447), .B(n15446), .ZN(
        n15458) );
  INV_X1 U17358 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15449) );
  OAI21_X1 U17359 ( .B1(n15450), .B2(n15449), .A(n15474), .ZN(n15453) );
  INV_X1 U17360 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15451) );
  OAI22_X1 U17361 ( .A1(n12431), .A2(n19340), .B1(n14278), .B2(n15451), .ZN(
        n15452) );
  AOI211_X1 U17362 ( .C1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .C2(n10965), .A(
        n15453), .B(n15452), .ZN(n15456) );
  AOI22_X1 U17363 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15471), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U17364 ( .A1(n15475), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15454) );
  NAND3_X1 U17365 ( .A1(n15456), .A2(n15455), .A3(n15454), .ZN(n15457) );
  OAI21_X1 U17366 ( .B1(n15459), .B2(n15458), .A(n15457), .ZN(n15460) );
  NOR2_X1 U17367 ( .A1(n15461), .A2(n15460), .ZN(n16250) );
  AOI21_X1 U17368 ( .B1(n16251), .B2(n16248), .A(n16250), .ZN(n15484) );
  INV_X1 U17369 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U17370 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15462), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15464) );
  NAND2_X1 U17371 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n15463) );
  OAI211_X1 U17372 ( .C1(n19222), .C2(n12627), .A(n15464), .B(n15463), .ZN(
        n15482) );
  INV_X1 U17373 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15469) );
  AOI21_X1 U17374 ( .B1(n15466), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15465), .ZN(n15468) );
  AOI22_X1 U17375 ( .A1(n10983), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15467) );
  OAI211_X1 U17376 ( .C1(n15470), .C2(n15469), .A(n15468), .B(n15467), .ZN(
        n15481) );
  AOI22_X1 U17377 ( .A1(n15283), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15466), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15473) );
  AOI22_X1 U17378 ( .A1(n15471), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15472) );
  NAND2_X1 U17379 ( .A1(n15473), .A2(n15472), .ZN(n15480) );
  INV_X1 U17380 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U17381 ( .A1(n12503), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12628), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15477) );
  AOI21_X1 U17382 ( .B1(n15475), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n15474), .ZN(n15476) );
  OAI211_X1 U17383 ( .C1(n12431), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15479) );
  OAI22_X1 U17384 ( .A1(n15482), .A2(n15481), .B1(n15480), .B2(n15479), .ZN(
        n15483) );
  XNOR2_X1 U17385 ( .A(n15484), .B(n15483), .ZN(n15497) );
  NOR2_X1 U17386 ( .A1(n15487), .A2(n13649), .ZN(n15485) );
  AOI22_X1 U17387 ( .A1(n19583), .A2(BUF1_REG_30__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n15492) );
  NOR2_X1 U17388 ( .A1(n15487), .A2(n15486), .ZN(n15488) );
  AOI22_X1 U17389 ( .A1(n19582), .A2(BUF2_REG_30__SCAN_IN), .B1(n19581), .B2(
        n15490), .ZN(n15491) );
  OAI211_X1 U17390 ( .C1(n16149), .C2(n16373), .A(n15492), .B(n15491), .ZN(
        n15493) );
  INV_X1 U17391 ( .A(n15493), .ZN(n15494) );
  OAI21_X1 U17392 ( .B1(n15497), .B2(n19342), .A(n15494), .ZN(P2_U2889) );
  NAND2_X1 U17393 ( .A1(n16152), .A2(n16284), .ZN(n15496) );
  NAND2_X1 U17394 ( .A1(n14161), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15495) );
  OAI211_X1 U17395 ( .C1(n15497), .C2(n16302), .A(n15496), .B(n15495), .ZN(
        P2_U2857) );
  AOI21_X1 U17396 ( .B1(n17021), .B2(n16094), .A(n16982), .ZN(n15501) );
  OR2_X1 U17397 ( .A1(n21699), .A2(n16090), .ZN(n17024) );
  OAI21_X1 U17398 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16089), .A(
        n17024), .ZN(n15499) );
  OAI22_X1 U17399 ( .A1(n21549), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16096), .ZN(n15498) );
  AOI21_X1 U17400 ( .B1(n15499), .B2(n16094), .A(n15498), .ZN(n15500) );
  OAI22_X1 U17401 ( .A1(n15501), .A2(n11541), .B1(n16982), .B2(n15500), .ZN(
        P1_U3474) );
  NAND2_X1 U17402 ( .A1(n15503), .A2(n15502), .ZN(n15505) );
  XOR2_X1 U17403 ( .A(n15505), .B(n15504), .Z(n16394) );
  INV_X1 U17404 ( .A(n16414), .ZN(n15506) );
  AOI21_X1 U17405 ( .B1(n15506), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15508) );
  NOR2_X1 U17406 ( .A1(n15508), .A2(n15507), .ZN(n16392) );
  OR2_X1 U17407 ( .A1(n16164), .A2(n15509), .ZN(n15510) );
  NAND2_X1 U17408 ( .A1(n18427), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16388) );
  OAI21_X1 U17409 ( .B1(n18577), .B2(n18603), .A(n16388), .ZN(n15512) );
  INV_X1 U17410 ( .A(n15512), .ZN(n15521) );
  NOR2_X1 U17411 ( .A1(n16654), .A2(n15516), .ZN(n15519) );
  INV_X1 U17412 ( .A(n15515), .ZN(n16650) );
  XNOR2_X1 U17413 ( .A(n15516), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15517) );
  AND2_X1 U17414 ( .A1(n16650), .A2(n15517), .ZN(n15518) );
  AOI21_X1 U17415 ( .B1(n16392), .B2(n18623), .A(n15522), .ZN(n15523) );
  OAI21_X1 U17416 ( .B1(n16394), .B2(n18614), .A(n15523), .ZN(P2_U3017) );
  INV_X1 U17417 ( .A(n15524), .ZN(n15525) );
  XNOR2_X1 U17418 ( .A(n15526), .B(n15525), .ZN(n18626) );
  NOR2_X1 U17419 ( .A1(n18600), .A2(n12577), .ZN(n18621) );
  AOI21_X1 U17420 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n18621), .ZN(n15531) );
  AOI21_X1 U17421 ( .B1(n15529), .B2(n15528), .A(n15527), .ZN(n18622) );
  NAND2_X1 U17422 ( .A1(n18622), .A2(n17270), .ZN(n15530) );
  OAI211_X1 U17423 ( .C1(n17301), .C2(n15532), .A(n15531), .B(n15530), .ZN(
        n15533) );
  AOI21_X1 U17424 ( .B1(n17274), .B2(n18626), .A(n15533), .ZN(n15534) );
  OAI21_X1 U17425 ( .B1(n12609), .B2(n17296), .A(n15534), .ZN(P2_U3012) );
  NAND2_X1 U17426 ( .A1(n15546), .A2(n15535), .ZN(n15536) );
  OAI21_X1 U17427 ( .B1(n15546), .B2(n15537), .A(n15536), .ZN(n15543) );
  INV_X1 U17428 ( .A(n15545), .ZN(n15541) );
  INV_X1 U17429 ( .A(n15538), .ZN(n15539) );
  OAI22_X1 U17430 ( .A1(n15546), .A2(n15541), .B1(n15540), .B2(n15539), .ZN(
        n15542) );
  OR2_X1 U17431 ( .A1(n15543), .A2(n15542), .ZN(n17036) );
  NAND2_X1 U17432 ( .A1(n15547), .A2(n21229), .ZN(n15548) );
  NAND2_X1 U17433 ( .A1(n15548), .A2(n17050), .ZN(n21231) );
  NOR2_X1 U17434 ( .A1(n19953), .A2(n21231), .ZN(n17034) );
  NOR2_X1 U17435 ( .A1(n17034), .A2(n21561), .ZN(n21548) );
  MUX2_X1 U17436 ( .A(P1_MORE_REG_SCAN_IN), .B(n17036), .S(n21548), .Z(
        P1_U3484) );
  INV_X1 U17437 ( .A(n15549), .ZN(n15603) );
  NAND3_X1 U17438 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .ZN(n15709) );
  NAND2_X1 U17439 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15710) );
  INV_X1 U17440 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n19817) );
  NOR4_X1 U17441 ( .A1(n15708), .A2(n15709), .A3(n15710), .A4(n19817), .ZN(
        n21508) );
  NAND2_X1 U17442 ( .A1(n21508), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15700) );
  OAI21_X1 U17443 ( .B1(n15550), .B2(n15700), .A(n21485), .ZN(n21510) );
  OAI21_X1 U17444 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21453), .A(n21510), 
        .ZN(n21522) );
  NOR2_X1 U17445 ( .A1(n21453), .A2(n21522), .ZN(n21524) );
  NAND2_X1 U17446 ( .A1(n21524), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n21533) );
  INV_X1 U17447 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21534) );
  NAND2_X1 U17448 ( .A1(n15690), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U17449 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15551) );
  INV_X1 U17450 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n17139) );
  NAND2_X1 U17451 ( .A1(n15614), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15601) );
  AND2_X1 U17452 ( .A1(n15601), .A2(n21485), .ZN(n15613) );
  OAI22_X1 U17453 ( .A1(n15596), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n13878), .ZN(n15599) );
  OAI22_X1 U17454 ( .A1(n15596), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n13878), .ZN(n15608) );
  INV_X1 U17455 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21486) );
  NAND2_X1 U17456 ( .A1(n15591), .A2(n21486), .ZN(n15556) );
  NAND2_X1 U17457 ( .A1(n14056), .A2(n15552), .ZN(n15554) );
  NAND2_X1 U17458 ( .A1(n13785), .A2(n21486), .ZN(n15553) );
  NAND3_X1 U17459 ( .A1(n15554), .A2(n15607), .A3(n15553), .ZN(n15555) );
  AND2_X1 U17460 ( .A1(n15556), .A2(n15555), .ZN(n15790) );
  MUX2_X1 U17461 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n15557) );
  NAND2_X1 U17462 ( .A1(n11522), .A2(n15557), .ZN(n15726) );
  INV_X1 U17463 ( .A(n15591), .ZN(n15586) );
  OAI21_X1 U17464 ( .B1(n10968), .B2(n15558), .A(n14056), .ZN(n15560) );
  INV_X1 U17465 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15781) );
  NAND2_X1 U17466 ( .A1(n13785), .A2(n15781), .ZN(n15559) );
  NAND2_X1 U17467 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  OAI21_X1 U17468 ( .B1(n15586), .B2(P1_EBX_REG_18__SCAN_IN), .A(n15561), .ZN(
        n15779) );
  NAND2_X1 U17469 ( .A1(n15780), .A2(n15779), .ZN(n15778) );
  INV_X1 U17470 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21361) );
  INV_X1 U17471 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15712) );
  NAND2_X1 U17472 ( .A1(n13785), .A2(n15712), .ZN(n15562) );
  OAI211_X1 U17473 ( .C1(n10968), .C2(n21361), .A(n15562), .B(n14056), .ZN(
        n15563) );
  OAI21_X1 U17474 ( .B1(n15590), .B2(P1_EBX_REG_19__SCAN_IN), .A(n15563), .ZN(
        n15714) );
  INV_X1 U17475 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21506) );
  NAND2_X1 U17476 ( .A1(n15591), .A2(n21506), .ZN(n15567) );
  NAND2_X1 U17477 ( .A1(n14056), .A2(n19936), .ZN(n15565) );
  NAND2_X1 U17478 ( .A1(n13785), .A2(n21506), .ZN(n15564) );
  NAND3_X1 U17479 ( .A1(n15565), .A2(n15607), .A3(n15564), .ZN(n15566) );
  INV_X1 U17480 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15568) );
  NAND2_X1 U17481 ( .A1(n15580), .A2(n15568), .ZN(n15570) );
  MUX2_X1 U17482 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n15569) );
  AND2_X1 U17483 ( .A1(n15570), .A2(n15569), .ZN(n15698) );
  INV_X1 U17484 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15759) );
  NAND2_X1 U17485 ( .A1(n15591), .A2(n15759), .ZN(n15574) );
  INV_X1 U17486 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U17487 ( .A1(n14056), .A2(n15977), .ZN(n15572) );
  NAND2_X1 U17488 ( .A1(n13785), .A2(n15759), .ZN(n15571) );
  NAND3_X1 U17489 ( .A1(n15572), .A2(n15607), .A3(n15571), .ZN(n15573) );
  NAND2_X1 U17490 ( .A1(n15574), .A2(n15573), .ZN(n15756) );
  MUX2_X1 U17491 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n15576) );
  NAND2_X1 U17492 ( .A1(n15580), .A2(n21404), .ZN(n15575) );
  NAND2_X1 U17493 ( .A1(n15576), .A2(n15575), .ZN(n15749) );
  OAI21_X1 U17494 ( .B1(n10968), .B2(n16066), .A(n14056), .ZN(n15577) );
  OAI21_X1 U17495 ( .B1(n13878), .B2(P1_EBX_REG_24__SCAN_IN), .A(n15577), .ZN(
        n15579) );
  INV_X1 U17496 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15746) );
  NAND2_X1 U17497 ( .A1(n15591), .A2(n15746), .ZN(n15578) );
  MUX2_X1 U17498 ( .A(n15590), .B(n15607), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n15582) );
  NAND2_X1 U17499 ( .A1(n15580), .A2(n16052), .ZN(n15581) );
  AND2_X1 U17500 ( .A1(n15582), .A2(n15581), .ZN(n15674) );
  INV_X1 U17501 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16042) );
  NAND2_X1 U17502 ( .A1(n14056), .A2(n16042), .ZN(n15584) );
  INV_X1 U17503 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15741) );
  NAND2_X1 U17504 ( .A1(n13785), .A2(n15741), .ZN(n15583) );
  NAND3_X1 U17505 ( .A1(n15584), .A2(n15607), .A3(n15583), .ZN(n15585) );
  OAI21_X1 U17506 ( .B1(n15586), .B2(P1_EBX_REG_26__SCAN_IN), .A(n15585), .ZN(
        n15664) );
  INV_X1 U17507 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15740) );
  NAND2_X1 U17508 ( .A1(n13785), .A2(n15740), .ZN(n15587) );
  OAI211_X1 U17509 ( .C1(n10968), .C2(n16038), .A(n15587), .B(n14056), .ZN(
        n15589) );
  OAI21_X1 U17510 ( .B1(n15590), .B2(P1_EBX_REG_27__SCAN_IN), .A(n15589), .ZN(
        n15648) );
  INV_X1 U17511 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U17512 ( .A1(n15591), .A2(n15739), .ZN(n15595) );
  NAND2_X1 U17513 ( .A1(n14056), .A2(n15887), .ZN(n15593) );
  NAND2_X1 U17514 ( .A1(n13785), .A2(n15739), .ZN(n15592) );
  NAND3_X1 U17515 ( .A1(n15593), .A2(n15607), .A3(n15592), .ZN(n15594) );
  AND2_X1 U17516 ( .A1(n15595), .A2(n15594), .ZN(n15635) );
  INV_X1 U17517 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15737) );
  NAND2_X1 U17518 ( .A1(n13785), .A2(n15737), .ZN(n15597) );
  OAI21_X1 U17519 ( .B1(n15596), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15597), .ZN(n15606) );
  MUX2_X1 U17520 ( .A(n15597), .B(n15606), .S(n15607), .Z(n15622) );
  MUX2_X1 U17521 ( .A(n15607), .B(n15608), .S(n15621), .Z(n15598) );
  AOI22_X1 U17522 ( .A1(n21529), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21517), .ZN(n15600) );
  OAI21_X1 U17523 ( .B1(n15603), .B2(n21537), .A(n15602), .ZN(P1_U2809) );
  INV_X1 U17524 ( .A(n15875), .ZN(n15736) );
  OAI22_X1 U17525 ( .A1(n15621), .A2(n15607), .B1(n15637), .B2(n15606), .ZN(
        n15609) );
  XNOR2_X1 U17526 ( .A(n15609), .B(n15608), .ZN(n16004) );
  NAND2_X1 U17527 ( .A1(n21529), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n15611) );
  AOI22_X1 U17528 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21517), .B1(
        n21530), .B2(n15871), .ZN(n15610) );
  NAND2_X1 U17529 ( .A1(n15611), .A2(n15610), .ZN(n15612) );
  AOI21_X1 U17530 ( .B1(n16004), .B2(n21490), .A(n15612), .ZN(n15616) );
  OAI21_X1 U17531 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n15614), .A(n15613), 
        .ZN(n15615) );
  OAI211_X1 U17532 ( .C1(n15736), .C2(n21537), .A(n15616), .B(n15615), .ZN(
        P1_U2810) );
  INV_X1 U17533 ( .A(n15618), .ZN(n15619) );
  INV_X1 U17534 ( .A(n15883), .ZN(n15738) );
  INV_X1 U17535 ( .A(n15629), .ZN(n15640) );
  AND2_X1 U17536 ( .A1(n21485), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15628) );
  INV_X1 U17537 ( .A(n15621), .ZN(n15624) );
  NAND2_X1 U17538 ( .A1(n15637), .A2(n15622), .ZN(n15623) );
  NAND2_X1 U17539 ( .A1(n15624), .A2(n15623), .ZN(n16008) );
  AOI22_X1 U17540 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n21517), .B1(
        n21530), .B2(n15879), .ZN(n15626) );
  NAND2_X1 U17541 ( .A1(n21529), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n15625) );
  OAI211_X1 U17542 ( .C1(n16008), .C2(n21535), .A(n15626), .B(n15625), .ZN(
        n15627) );
  AOI21_X1 U17543 ( .B1(n15640), .B2(n15628), .A(n15627), .ZN(n15631) );
  INV_X1 U17544 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n19835) );
  NAND2_X1 U17545 ( .A1(n15629), .A2(n19835), .ZN(n15630) );
  OAI211_X1 U17546 ( .C1(n15738), .C2(n21537), .A(n15631), .B(n15630), .ZN(
        P1_U2811) );
  OAI21_X1 U17547 ( .B1(n15632), .B2(n15633), .A(n15617), .ZN(n15894) );
  OAI22_X1 U17548 ( .A1(n15634), .A2(n21544), .B1(n21519), .B2(n15890), .ZN(
        n15639) );
  NAND2_X1 U17549 ( .A1(n15650), .A2(n15635), .ZN(n15636) );
  NAND2_X1 U17550 ( .A1(n15637), .A2(n15636), .ZN(n16018) );
  NOR2_X1 U17551 ( .A1(n16018), .A2(n21535), .ZN(n15638) );
  AOI211_X1 U17552 ( .C1(n21529), .C2(P1_EBX_REG_28__SCAN_IN), .A(n15639), .B(
        n15638), .ZN(n15643) );
  INV_X1 U17553 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15889) );
  NOR2_X1 U17554 ( .A1(n15720), .A2(n15889), .ZN(n15641) );
  OAI21_X1 U17555 ( .B1(n15647), .B2(n15641), .A(n15640), .ZN(n15642) );
  OAI211_X1 U17556 ( .C1(n15894), .C2(n21537), .A(n15643), .B(n15642), .ZN(
        P1_U2812) );
  INV_X1 U17557 ( .A(n15632), .ZN(n15645) );
  INV_X1 U17558 ( .A(n15647), .ZN(n15655) );
  OAI21_X1 U17559 ( .B1(n15720), .B2(n17139), .A(n15657), .ZN(n15654) );
  NAND2_X1 U17560 ( .A1(n15663), .A2(n15648), .ZN(n15649) );
  NAND2_X1 U17561 ( .A1(n15650), .A2(n15649), .ZN(n16035) );
  AOI22_X1 U17562 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n21517), .B1(
        n21530), .B2(n15897), .ZN(n15652) );
  NAND2_X1 U17563 ( .A1(n21529), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n15651) );
  OAI211_X1 U17564 ( .C1(n16035), .C2(n21535), .A(n15652), .B(n15651), .ZN(
        n15653) );
  AOI21_X1 U17565 ( .B1(n15655), .B2(n15654), .A(n15653), .ZN(n15656) );
  OAI21_X1 U17566 ( .B1(n15901), .B2(n21537), .A(n15656), .ZN(P1_U2813) );
  INV_X1 U17567 ( .A(n15657), .ZN(n15670) );
  INV_X1 U17568 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n17152) );
  INV_X1 U17569 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n17157) );
  NOR2_X1 U17570 ( .A1(n17152), .A2(n17157), .ZN(n15658) );
  AOI22_X1 U17571 ( .A1(n15690), .A2(n15658), .B1(P1_REIP_REG_26__SCAN_IN), 
        .B2(n21485), .ZN(n15669) );
  INV_X1 U17572 ( .A(n15659), .ZN(n15661) );
  INV_X1 U17573 ( .A(n15672), .ZN(n15660) );
  NAND2_X1 U17574 ( .A1(n15908), .A2(n21525), .ZN(n15668) );
  OAI22_X1 U17575 ( .A1(n15662), .A2(n21544), .B1(n21519), .B2(n15906), .ZN(
        n15666) );
  OAI21_X1 U17576 ( .B1(n15676), .B2(n15664), .A(n15663), .ZN(n16045) );
  NOR2_X1 U17577 ( .A1(n16045), .A2(n21535), .ZN(n15665) );
  AOI211_X1 U17578 ( .C1(n21529), .C2(P1_EBX_REG_26__SCAN_IN), .A(n15666), .B(
        n15665), .ZN(n15667) );
  OAI211_X1 U17579 ( .C1(n15670), .C2(n15669), .A(n15668), .B(n15667), .ZN(
        P1_U2814) );
  AOI21_X1 U17580 ( .B1(n15673), .B2(n15684), .A(n15672), .ZN(n15914) );
  INV_X1 U17581 ( .A(n15914), .ZN(n15744) );
  OR2_X1 U17582 ( .A1(n15690), .A2(n15720), .ZN(n21532) );
  OAI21_X1 U17583 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n21453), .A(n21532), 
        .ZN(n15682) );
  NOR2_X1 U17584 ( .A1(n15688), .A2(n15674), .ZN(n15675) );
  OR2_X1 U17585 ( .A1(n15676), .A2(n15675), .ZN(n16054) );
  AOI22_X1 U17586 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n21517), .B1(
        n21530), .B2(n15917), .ZN(n15678) );
  NAND2_X1 U17587 ( .A1(n21529), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n15677) );
  OAI211_X1 U17588 ( .C1(n16054), .C2(n21535), .A(n15678), .B(n15677), .ZN(
        n15681) );
  NOR2_X1 U17589 ( .A1(n15679), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15680) );
  AOI211_X1 U17590 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n15682), .A(n15681), 
        .B(n15680), .ZN(n15683) );
  OAI21_X1 U17591 ( .B1(n15744), .B2(n21537), .A(n15683), .ZN(P1_U2815) );
  AOI21_X1 U17592 ( .B1(n15685), .B2(n15748), .A(n15671), .ZN(n15926) );
  NAND2_X1 U17593 ( .A1(n15926), .A2(n21525), .ZN(n15695) );
  AND2_X1 U17594 ( .A1(n11023), .A2(n15686), .ZN(n15687) );
  NOR2_X1 U17595 ( .A1(n15688), .A2(n15687), .ZN(n16065) );
  AOI22_X1 U17596 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n21517), .B1(
        P1_EBX_REG_24__SCAN_IN), .B2(n21529), .ZN(n15689) );
  OAI21_X1 U17597 ( .B1(n15924), .B2(n21519), .A(n15689), .ZN(n15693) );
  INV_X1 U17598 ( .A(n15690), .ZN(n15691) );
  NOR2_X1 U17599 ( .A1(n15691), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15692) );
  AOI211_X1 U17600 ( .C1(n21490), .C2(n16065), .A(n15693), .B(n15692), .ZN(
        n15694) );
  OAI211_X1 U17601 ( .C1(n21532), .C2(n17157), .A(n15695), .B(n15694), .ZN(
        P1_U2816) );
  INV_X1 U17602 ( .A(n15753), .ZN(n15696) );
  OAI21_X1 U17603 ( .B1(n15697), .B2(n15765), .A(n15696), .ZN(n15939) );
  INV_X1 U17604 ( .A(n21510), .ZN(n15706) );
  NOR2_X1 U17605 ( .A1(n15769), .A2(n15698), .ZN(n15699) );
  OR2_X1 U17606 ( .A1(n15757), .A2(n15699), .ZN(n21394) );
  NOR3_X1 U17607 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n21453), .A3(n15700), 
        .ZN(n15703) );
  AOI22_X1 U17608 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n21517), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(n21529), .ZN(n15701) );
  INV_X1 U17609 ( .A(n15701), .ZN(n15702) );
  AOI211_X1 U17610 ( .C1(n21530), .C2(n15937), .A(n15703), .B(n15702), .ZN(
        n15704) );
  OAI21_X1 U17611 ( .B1(n21394), .B2(n21535), .A(n15704), .ZN(n15705) );
  AOI21_X1 U17612 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15706), .A(n15705), 
        .ZN(n15707) );
  OAI21_X1 U17613 ( .B1(n15939), .B2(n21537), .A(n15707), .ZN(P1_U2819) );
  OAI21_X1 U17614 ( .B1(n12084), .B2(n11094), .A(n15764), .ZN(n15949) );
  NOR2_X1 U17615 ( .A1(n15709), .A2(n21473), .ZN(n21494) );
  NAND2_X1 U17616 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n21494), .ZN(n21498) );
  OAI21_X1 U17617 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(P1_REIP_REG_19__SCAN_IN), 
        .A(n15710), .ZN(n15711) );
  OAI22_X1 U17618 ( .A1(n15712), .A2(n21505), .B1(n21498), .B2(n15711), .ZN(
        n15719) );
  OAI21_X1 U17619 ( .B1(n21544), .B2(n15944), .A(n15728), .ZN(n15718) );
  INV_X1 U17620 ( .A(n15768), .ZN(n15713) );
  AOI21_X1 U17621 ( .B1(n15714), .B2(n15778), .A(n15713), .ZN(n21375) );
  INV_X1 U17622 ( .A(n21375), .ZN(n15716) );
  INV_X1 U17623 ( .A(n15946), .ZN(n15715) );
  OAI22_X1 U17624 ( .A1(n15716), .A2(n21535), .B1(n15715), .B2(n21519), .ZN(
        n15717) );
  NOR3_X1 U17625 ( .A1(n15719), .A2(n15718), .A3(n15717), .ZN(n15723) );
  INV_X1 U17626 ( .A(n21498), .ZN(n15721) );
  NOR2_X1 U17627 ( .A1(n15721), .A2(n15720), .ZN(n21501) );
  NAND2_X1 U17628 ( .A1(n21501), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15722) );
  OAI211_X1 U17629 ( .C1(n15949), .C2(n21537), .A(n15723), .B(n15722), .ZN(
        P1_U2821) );
  INV_X1 U17630 ( .A(n15775), .ZN(n15724) );
  OAI21_X1 U17631 ( .B1(n11060), .B2(n15725), .A(n15724), .ZN(n15962) );
  OAI21_X1 U17632 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21494), .A(n21501), 
        .ZN(n15732) );
  AND2_X1 U17633 ( .A1(n15793), .A2(n15726), .ZN(n15727) );
  OR2_X1 U17634 ( .A1(n15727), .A2(n15780), .ZN(n15786) );
  INV_X1 U17635 ( .A(n15786), .ZN(n21345) );
  AOI22_X1 U17636 ( .A1(n15959), .A2(n21530), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n21529), .ZN(n15729) );
  OAI211_X1 U17637 ( .C1(n21544), .C2(n15957), .A(n15729), .B(n15728), .ZN(
        n15730) );
  AOI21_X1 U17638 ( .B1(n21490), .B2(n21345), .A(n15730), .ZN(n15731) );
  OAI211_X1 U17639 ( .C1(n15962), .C2(n21537), .A(n15732), .B(n15731), .ZN(
        P1_U2823) );
  INV_X1 U17640 ( .A(n15993), .ZN(n15734) );
  INV_X1 U17641 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15733) );
  OAI22_X1 U17642 ( .A1(n15734), .A2(n15785), .B1(n19870), .B2(n15733), .ZN(
        P1_U2841) );
  AOI22_X1 U17643 ( .A1(n16004), .A2(n19865), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15794), .ZN(n15735) );
  OAI21_X1 U17644 ( .B1(n15736), .B2(n15796), .A(n15735), .ZN(P1_U2842) );
  OAI222_X1 U17645 ( .A1(n15796), .A2(n15738), .B1(n15737), .B2(n19870), .C1(
        n16008), .C2(n15785), .ZN(P1_U2843) );
  OAI222_X1 U17646 ( .A1(n15796), .A2(n15894), .B1(n15739), .B2(n19870), .C1(
        n16018), .C2(n15785), .ZN(P1_U2844) );
  OAI222_X1 U17647 ( .A1(n15796), .A2(n15901), .B1(n15740), .B2(n19870), .C1(
        n16035), .C2(n15785), .ZN(P1_U2845) );
  INV_X1 U17648 ( .A(n15908), .ZN(n15742) );
  OAI222_X1 U17649 ( .A1(n15796), .A2(n15742), .B1(n15741), .B2(n19870), .C1(
        n16045), .C2(n15785), .ZN(P1_U2846) );
  INV_X1 U17650 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15743) );
  OAI222_X1 U17651 ( .A1(n15796), .A2(n15744), .B1(n15743), .B2(n19870), .C1(
        n16054), .C2(n15785), .ZN(P1_U2847) );
  INV_X1 U17652 ( .A(n15926), .ZN(n15747) );
  INV_X1 U17653 ( .A(n16065), .ZN(n15745) );
  OAI222_X1 U17654 ( .A1(n15796), .A2(n15747), .B1(n15746), .B2(n19870), .C1(
        n15745), .C2(n15785), .ZN(P1_U2848) );
  OAI21_X1 U17655 ( .B1(n12162), .B2(n11095), .A(n15748), .ZN(n21538) );
  INV_X1 U17656 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15751) );
  NAND2_X1 U17657 ( .A1(n11071), .A2(n15749), .ZN(n15750) );
  AND2_X1 U17658 ( .A1(n11023), .A2(n15750), .ZN(n21399) );
  INV_X1 U17659 ( .A(n21399), .ZN(n21536) );
  OAI222_X1 U17660 ( .A1(n15783), .A2(n21538), .B1(n15751), .B2(n19870), .C1(
        n21536), .C2(n15785), .ZN(P1_U2849) );
  OR2_X1 U17661 ( .A1(n15753), .A2(n15752), .ZN(n15754) );
  AND2_X1 U17662 ( .A1(n15755), .A2(n15754), .ZN(n21654) );
  OR2_X1 U17663 ( .A1(n15757), .A2(n15756), .ZN(n15758) );
  NAND2_X1 U17664 ( .A1(n11071), .A2(n15758), .ZN(n21528) );
  OAI22_X1 U17665 ( .A1(n21528), .A2(n15785), .B1(n15759), .B2(n19870), .ZN(
        n15760) );
  AOI21_X1 U17666 ( .B1(n21654), .B2(n19866), .A(n15760), .ZN(n15761) );
  INV_X1 U17667 ( .A(n15761), .ZN(P1_U2850) );
  INV_X1 U17668 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15762) );
  OAI222_X1 U17669 ( .A1(n15939), .A2(n15783), .B1(n15762), .B2(n19870), .C1(
        n15785), .C2(n21394), .ZN(P1_U2851) );
  AND2_X1 U17670 ( .A1(n15764), .A2(n15763), .ZN(n15766) );
  OR2_X1 U17671 ( .A1(n15766), .A2(n15765), .ZN(n21512) );
  AND2_X1 U17672 ( .A1(n15768), .A2(n15767), .ZN(n15770) );
  OR2_X1 U17673 ( .A1(n15770), .A2(n15769), .ZN(n21516) );
  OAI22_X1 U17674 ( .A1(n21516), .A2(n15785), .B1(n21506), .B2(n19870), .ZN(
        n15771) );
  AOI21_X1 U17675 ( .B1(n21646), .B2(n19866), .A(n15771), .ZN(n15772) );
  INV_X1 U17676 ( .A(n15772), .ZN(P1_U2852) );
  AOI22_X1 U17677 ( .A1(n21375), .A2(n19865), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15794), .ZN(n15773) );
  OAI21_X1 U17678 ( .B1(n15949), .B2(n15796), .A(n15773), .ZN(P1_U2853) );
  OR2_X1 U17679 ( .A1(n15775), .A2(n15774), .ZN(n15776) );
  AND2_X1 U17680 ( .A1(n15777), .A2(n15776), .ZN(n21642) );
  INV_X1 U17681 ( .A(n21642), .ZN(n15782) );
  OAI21_X1 U17682 ( .B1(n15780), .B2(n15779), .A(n15778), .ZN(n21504) );
  OAI222_X1 U17683 ( .A1(n15782), .A2(n15783), .B1(n15781), .B2(n19870), .C1(
        n15785), .C2(n21504), .ZN(P1_U2854) );
  INV_X1 U17684 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15784) );
  OAI222_X1 U17685 ( .A1(n15786), .A2(n15785), .B1(n15784), .B2(n19870), .C1(
        n15962), .C2(n15783), .ZN(P1_U2855) );
  AND2_X1 U17686 ( .A1(n15788), .A2(n15787), .ZN(n15789) );
  NOR2_X1 U17687 ( .A1(n11060), .A2(n15789), .ZN(n21638) );
  INV_X1 U17688 ( .A(n21638), .ZN(n15797) );
  NAND2_X1 U17689 ( .A1(n15791), .A2(n15790), .ZN(n15792) );
  NAND2_X1 U17690 ( .A1(n15793), .A2(n15792), .ZN(n21357) );
  INV_X1 U17691 ( .A(n21357), .ZN(n21489) );
  AOI22_X1 U17692 ( .A1(n21489), .A2(n19865), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n15794), .ZN(n15795) );
  OAI21_X1 U17693 ( .B1(n15797), .B2(n15796), .A(n15795), .ZN(P1_U2856) );
  INV_X1 U17694 ( .A(DATAI_30_), .ZN(n15804) );
  NAND2_X1 U17695 ( .A1(n15875), .A2(n21653), .ZN(n15803) );
  OAI22_X1 U17696 ( .A1(n21636), .A2(n15800), .B1(n15852), .B2(n15799), .ZN(
        n15801) );
  AOI21_X1 U17697 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n21652), .A(n15801), .ZN(
        n15802) );
  OAI211_X1 U17698 ( .C1(n21657), .C2(n15804), .A(n15803), .B(n15802), .ZN(
        P1_U2874) );
  INV_X1 U17699 ( .A(DATAI_29_), .ZN(n15810) );
  NAND2_X1 U17700 ( .A1(n15883), .A2(n21653), .ZN(n15809) );
  OAI22_X1 U17701 ( .A1(n21636), .A2(n15806), .B1(n15852), .B2(n15805), .ZN(
        n15807) );
  AOI21_X1 U17702 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n21652), .A(n15807), .ZN(
        n15808) );
  OAI211_X1 U17703 ( .C1(n21657), .C2(n15810), .A(n15809), .B(n15808), .ZN(
        P1_U2875) );
  INV_X1 U17704 ( .A(DATAI_28_), .ZN(n15817) );
  INV_X1 U17705 ( .A(n15894), .ZN(n15811) );
  NAND2_X1 U17706 ( .A1(n15811), .A2(n21653), .ZN(n15816) );
  OAI22_X1 U17707 ( .A1(n21636), .A2(n15813), .B1(n15852), .B2(n15812), .ZN(
        n15814) );
  AOI21_X1 U17708 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n21652), .A(n15814), .ZN(
        n15815) );
  OAI211_X1 U17709 ( .C1(n21657), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        P1_U2876) );
  INV_X1 U17710 ( .A(DATAI_27_), .ZN(n15824) );
  INV_X1 U17711 ( .A(n15901), .ZN(n15818) );
  NAND2_X1 U17712 ( .A1(n15818), .A2(n21653), .ZN(n15823) );
  OAI22_X1 U17713 ( .A1(n21636), .A2(n15820), .B1(n15852), .B2(n15819), .ZN(
        n15821) );
  AOI21_X1 U17714 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n21652), .A(n15821), .ZN(
        n15822) );
  OAI211_X1 U17715 ( .C1(n21657), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        P1_U2877) );
  INV_X1 U17716 ( .A(DATAI_26_), .ZN(n15830) );
  NAND2_X1 U17717 ( .A1(n15908), .A2(n21653), .ZN(n15829) );
  OAI22_X1 U17718 ( .A1(n21636), .A2(n15826), .B1(n15852), .B2(n15825), .ZN(
        n15827) );
  AOI21_X1 U17719 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n21652), .A(n15827), .ZN(
        n15828) );
  OAI211_X1 U17720 ( .C1(n21657), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        P1_U2878) );
  INV_X1 U17721 ( .A(DATAI_25_), .ZN(n15835) );
  NAND2_X1 U17722 ( .A1(n15914), .A2(n21653), .ZN(n15834) );
  OAI22_X1 U17723 ( .A1(n21636), .A2(n15831), .B1(n15864), .B2(n14565), .ZN(
        n15832) );
  AOI21_X1 U17724 ( .B1(n21652), .B2(BUF1_REG_25__SCAN_IN), .A(n15832), .ZN(
        n15833) );
  OAI211_X1 U17725 ( .C1(n21657), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        P1_U2879) );
  INV_X1 U17726 ( .A(DATAI_24_), .ZN(n21665) );
  NAND2_X1 U17727 ( .A1(n15926), .A2(n21653), .ZN(n15840) );
  OAI22_X1 U17728 ( .A1(n21636), .A2(n15837), .B1(n15864), .B2(n15836), .ZN(
        n15838) );
  AOI21_X1 U17729 ( .B1(n21652), .B2(BUF1_REG_24__SCAN_IN), .A(n15838), .ZN(
        n15839) );
  OAI211_X1 U17730 ( .C1(n21657), .C2(n21665), .A(n15840), .B(n15839), .ZN(
        P1_U2880) );
  INV_X1 U17731 ( .A(DATAI_23_), .ZN(n15845) );
  INV_X1 U17732 ( .A(n21538), .ZN(n15841) );
  NAND2_X1 U17733 ( .A1(n15841), .A2(n21653), .ZN(n15844) );
  OAI22_X1 U17734 ( .A1(n21636), .A2(n22128), .B1(n15864), .B2(n14562), .ZN(
        n15842) );
  AOI21_X1 U17735 ( .B1(n21652), .B2(BUF1_REG_23__SCAN_IN), .A(n15842), .ZN(
        n15843) );
  OAI211_X1 U17736 ( .C1(n21657), .C2(n15845), .A(n15844), .B(n15843), .ZN(
        P1_U2881) );
  INV_X1 U17737 ( .A(DATAI_21_), .ZN(n15850) );
  INV_X1 U17738 ( .A(n15939), .ZN(n15846) );
  NAND2_X1 U17739 ( .A1(n15846), .A2(n21653), .ZN(n15849) );
  OAI22_X1 U17740 ( .A1(n21636), .A2(n22035), .B1(n15864), .B2(n14576), .ZN(
        n15847) );
  AOI21_X1 U17741 ( .B1(n21652), .B2(BUF1_REG_21__SCAN_IN), .A(n15847), .ZN(
        n15848) );
  OAI211_X1 U17742 ( .C1(n21657), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        P1_U2883) );
  INV_X1 U17743 ( .A(DATAI_19_), .ZN(n15856) );
  INV_X1 U17744 ( .A(n15949), .ZN(n15851) );
  NAND2_X1 U17745 ( .A1(n15851), .A2(n21653), .ZN(n15855) );
  OAI22_X1 U17746 ( .A1(n21636), .A2(n21944), .B1(n15852), .B2(n14567), .ZN(
        n15853) );
  AOI21_X1 U17747 ( .B1(n21652), .B2(BUF1_REG_19__SCAN_IN), .A(n15853), .ZN(
        n15854) );
  OAI211_X1 U17748 ( .C1(n21657), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        P1_U2885) );
  INV_X1 U17749 ( .A(DATAI_17_), .ZN(n15861) );
  INV_X1 U17750 ( .A(n15962), .ZN(n15857) );
  NAND2_X1 U17751 ( .A1(n15857), .A2(n21653), .ZN(n15860) );
  OAI22_X1 U17752 ( .A1(n21636), .A2(n21857), .B1(n15864), .B2(n14253), .ZN(
        n15858) );
  AOI21_X1 U17753 ( .B1(n21652), .B2(BUF1_REG_17__SCAN_IN), .A(n15858), .ZN(
        n15859) );
  OAI211_X1 U17754 ( .C1(n21657), .C2(n15861), .A(n15860), .B(n15859), .ZN(
        P1_U2887) );
  OAI222_X1 U17755 ( .A1(n15866), .A2(n15865), .B1(n15864), .B2(n19795), .C1(
        n15863), .C2(n15862), .ZN(P1_U2889) );
  NAND2_X1 U17756 ( .A1(n15867), .A2(n16010), .ZN(n15869) );
  XNOR2_X1 U17757 ( .A(n19945), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15878) );
  NAND3_X1 U17758 ( .A1(n15869), .A2(n15878), .A3(n15868), .ZN(n15870) );
  XNOR2_X1 U17759 ( .A(n15870), .B(n16002), .ZN(n16007) );
  NAND2_X1 U17760 ( .A1(n19927), .A2(n15871), .ZN(n15872) );
  NAND2_X1 U17761 ( .A1(n21390), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15999) );
  OAI211_X1 U17762 ( .C1(n15873), .C2(n19901), .A(n15872), .B(n15999), .ZN(
        n15874) );
  AOI21_X1 U17763 ( .B1(n15875), .B2(n19948), .A(n15874), .ZN(n15876) );
  OAI21_X1 U17764 ( .B1(n16007), .B2(n21546), .A(n15876), .ZN(P1_U2969) );
  NAND2_X1 U17765 ( .A1(n19927), .A2(n15879), .ZN(n15880) );
  NAND2_X1 U17766 ( .A1(n21390), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16009) );
  OAI211_X1 U17767 ( .C1(n19901), .C2(n15881), .A(n15880), .B(n16009), .ZN(
        n15882) );
  AOI21_X1 U17768 ( .B1(n15883), .B2(n19948), .A(n15882), .ZN(n15884) );
  OAI21_X1 U17769 ( .B1(n21546), .B2(n16016), .A(n15884), .ZN(P1_U2970) );
  INV_X1 U17770 ( .A(n15987), .ZN(n16043) );
  MUX2_X1 U17771 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n16042), .S(
        n19883), .Z(n15886) );
  XNOR2_X1 U17772 ( .A(n15888), .B(n15887), .ZN(n16017) );
  NAND2_X1 U17773 ( .A1(n16017), .A2(n19949), .ZN(n15893) );
  NOR2_X1 U17774 ( .A1(n21401), .A2(n15889), .ZN(n16019) );
  NOR2_X1 U17775 ( .A1(n19952), .A2(n15890), .ZN(n15891) );
  AOI211_X1 U17776 ( .C1(n19943), .C2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16019), .B(n15891), .ZN(n15892) );
  OAI211_X1 U17777 ( .C1(n19915), .C2(n15894), .A(n15893), .B(n15892), .ZN(
        P1_U2971) );
  NOR2_X1 U17778 ( .A1(n21401), .A2(n17139), .ZN(n16033) );
  INV_X1 U17779 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15895) );
  NOR2_X1 U17780 ( .A1(n19901), .A2(n15895), .ZN(n15896) );
  AOI211_X1 U17781 ( .C1(n19927), .C2(n15897), .A(n16033), .B(n15896), .ZN(
        n15900) );
  XNOR2_X1 U17782 ( .A(n19945), .B(n16038), .ZN(n15898) );
  NAND2_X1 U17783 ( .A1(n16030), .A2(n19949), .ZN(n15899) );
  OAI211_X1 U17784 ( .C1(n15901), .C2(n19915), .A(n15900), .B(n15899), .ZN(
        P1_U2972) );
  NAND3_X1 U17785 ( .A1(n15903), .A2(n15911), .A3(n15902), .ZN(n15904) );
  XNOR2_X1 U17786 ( .A(n15904), .B(n16042), .ZN(n16050) );
  NAND2_X1 U17787 ( .A1(n21390), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16044) );
  NAND2_X1 U17788 ( .A1(n19943), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15905) );
  OAI211_X1 U17789 ( .C1(n19952), .C2(n15906), .A(n16044), .B(n15905), .ZN(
        n15907) );
  AOI21_X1 U17790 ( .B1(n15908), .B2(n19948), .A(n15907), .ZN(n15909) );
  OAI21_X1 U17791 ( .B1(n21546), .B2(n16050), .A(n15909), .ZN(P1_U2973) );
  NAND2_X1 U17792 ( .A1(n16066), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15910) );
  OAI211_X1 U17793 ( .C1(n19883), .C2(n16066), .A(n15911), .B(n15910), .ZN(
        n15912) );
  AOI21_X1 U17794 ( .B1(n13580), .B2(n21404), .A(n15912), .ZN(n15913) );
  XNOR2_X1 U17795 ( .A(n15913), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16060) );
  NAND2_X1 U17796 ( .A1(n15914), .A2(n19948), .ZN(n15919) );
  NOR2_X1 U17797 ( .A1(n21401), .A2(n17152), .ZN(n16056) );
  NOR2_X1 U17798 ( .A1(n19901), .A2(n15915), .ZN(n15916) );
  AOI211_X1 U17799 ( .C1(n19927), .C2(n15917), .A(n16056), .B(n15916), .ZN(
        n15918) );
  OAI211_X1 U17800 ( .C1(n16060), .C2(n21546), .A(n15919), .B(n15918), .ZN(
        P1_U2974) );
  NAND3_X1 U17801 ( .A1(n13580), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n19883), .ZN(n15921) );
  NAND2_X1 U17802 ( .A1(n15921), .A2(n15920), .ZN(n15922) );
  XNOR2_X1 U17803 ( .A(n15922), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16069) );
  NOR2_X1 U17804 ( .A1(n21401), .A2(n17157), .ZN(n16064) );
  AOI21_X1 U17805 ( .B1(n19943), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16064), .ZN(n15923) );
  OAI21_X1 U17806 ( .B1(n19952), .B2(n15924), .A(n15923), .ZN(n15925) );
  AOI21_X1 U17807 ( .B1(n15926), .B2(n19948), .A(n15925), .ZN(n15927) );
  OAI21_X1 U17808 ( .B1(n16069), .B2(n21546), .A(n15927), .ZN(P1_U2975) );
  NAND2_X1 U17809 ( .A1(n21400), .A2(n19949), .ZN(n15930) );
  OAI22_X1 U17810 ( .A1(n19901), .A2(n21545), .B1(n21401), .B2(n21534), .ZN(
        n15928) );
  AOI21_X1 U17811 ( .B1(n19927), .B2(n21531), .A(n15928), .ZN(n15929) );
  OAI211_X1 U17812 ( .C1(n21538), .C2(n19915), .A(n15930), .B(n15929), .ZN(
        P1_U2976) );
  NOR2_X1 U17813 ( .A1(n17253), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15931) );
  AND3_X1 U17814 ( .A1(n15931), .A2(n19894), .A3(n21361), .ZN(n19940) );
  INV_X1 U17815 ( .A(n19940), .ZN(n15934) );
  AOI21_X1 U17816 ( .B1(n19936), .B2(n15934), .A(n15933), .ZN(n15935) );
  OAI21_X1 U17817 ( .B1(n15939), .B2(n19915), .A(n15938), .ZN(P1_U2978) );
  NAND2_X1 U17818 ( .A1(n19894), .A2(n15558), .ZN(n15940) );
  MUX2_X1 U17819 ( .A(n15558), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .S(
        n19883), .Z(n17252) );
  NAND2_X1 U17820 ( .A1(n17253), .A2(n17252), .ZN(n17251) );
  MUX2_X1 U17821 ( .A(n15941), .B(n15940), .S(n17251), .Z(n15942) );
  XOR2_X1 U17822 ( .A(n21361), .B(n15942), .Z(n21374) );
  NAND2_X1 U17823 ( .A1(n21374), .A2(n19949), .ZN(n15948) );
  INV_X1 U17824 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15943) );
  OAI22_X1 U17825 ( .A1(n19901), .A2(n15944), .B1(n21401), .B2(n15943), .ZN(
        n15945) );
  AOI21_X1 U17826 ( .B1(n19927), .B2(n15946), .A(n15945), .ZN(n15947) );
  OAI211_X1 U17827 ( .C1(n19915), .C2(n15949), .A(n15948), .B(n15947), .ZN(
        P1_U2980) );
  NOR2_X1 U17828 ( .A1(n15950), .A2(n15951), .ZN(n19912) );
  AOI21_X1 U17829 ( .B1(n19912), .B2(n15953), .A(n15952), .ZN(n15954) );
  MUX2_X1 U17830 ( .A(n15955), .B(n19894), .S(n15954), .Z(n15956) );
  XNOR2_X1 U17831 ( .A(n15956), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21344) );
  NAND2_X1 U17832 ( .A1(n21344), .A2(n19949), .ZN(n15961) );
  OAI22_X1 U17833 ( .A1(n19901), .A2(n15957), .B1(n21401), .B2(n19817), .ZN(
        n15958) );
  AOI21_X1 U17834 ( .B1(n19927), .B2(n15959), .A(n15958), .ZN(n15960) );
  OAI211_X1 U17835 ( .C1(n19915), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        P1_U2982) );
  INV_X1 U17836 ( .A(n15950), .ZN(n15964) );
  AOI21_X1 U17837 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n19894), .ZN(n19907) );
  OAI22_X1 U17838 ( .A1(n15964), .A2(n19907), .B1(n15963), .B2(n19945), .ZN(
        n19904) );
  INV_X1 U17839 ( .A(n15966), .ZN(n15965) );
  OAI21_X1 U17840 ( .B1(n19883), .B2(n21255), .A(n15965), .ZN(n19903) );
  NOR2_X1 U17841 ( .A1(n19904), .A2(n19903), .ZN(n19902) );
  NOR2_X1 U17842 ( .A1(n19902), .A2(n15966), .ZN(n15968) );
  XNOR2_X1 U17843 ( .A(n15968), .B(n15967), .ZN(n21246) );
  NAND2_X1 U17844 ( .A1(n21246), .A2(n19949), .ZN(n15974) );
  INV_X1 U17845 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15969) );
  OAI22_X1 U17846 ( .A1(n19901), .A2(n15970), .B1(n21401), .B2(n15969), .ZN(
        n15971) );
  AOI21_X1 U17847 ( .B1(n19927), .B2(n15972), .A(n15971), .ZN(n15973) );
  OAI211_X1 U17848 ( .C1(n19915), .C2(n15975), .A(n15974), .B(n15973), .ZN(
        P1_U2986) );
  NAND3_X1 U17849 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21343) );
  NOR2_X1 U17850 ( .A1(n15558), .A2(n21343), .ZN(n15978) );
  NOR2_X1 U17851 ( .A1(n21261), .A2(n21254), .ZN(n21331) );
  NAND2_X1 U17852 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21300) );
  NOR2_X1 U17853 ( .A1(n21300), .A2(n15976), .ZN(n21308) );
  AND2_X1 U17854 ( .A1(n21331), .A2(n21240), .ZN(n21329) );
  OAI221_X1 U17855 ( .B1(n21328), .B2(n15978), .C1(n21328), .C2(n21329), .A(
        n21327), .ZN(n21364) );
  NOR2_X1 U17856 ( .A1(n21364), .A2(n21337), .ZN(n16032) );
  NOR2_X1 U17857 ( .A1(n16032), .A2(n15988), .ZN(n15992) );
  NOR2_X1 U17858 ( .A1(n21378), .A2(n15977), .ZN(n15983) );
  OR2_X1 U17859 ( .A1(n21328), .A2(n15983), .ZN(n15981) );
  INV_X1 U17860 ( .A(n15978), .ZN(n21359) );
  NOR2_X1 U17861 ( .A1(n21300), .A2(n15979), .ZN(n21253) );
  NAND2_X1 U17862 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21253), .ZN(
        n21306) );
  NOR2_X1 U17863 ( .A1(n21255), .A2(n21306), .ZN(n21245) );
  NAND2_X1 U17864 ( .A1(n21331), .A2(n21245), .ZN(n21324) );
  NOR2_X1 U17865 ( .A1(n21359), .A2(n21324), .ZN(n21366) );
  NAND2_X1 U17866 ( .A1(n15983), .A2(n21366), .ZN(n15984) );
  AOI221_X1 U17867 ( .B1(n21404), .B2(n21325), .C1(n15984), .C2(n21325), .A(
        n21364), .ZN(n15980) );
  NAND2_X1 U17868 ( .A1(n15981), .A2(n15980), .ZN(n21405) );
  NOR2_X1 U17869 ( .A1(n21405), .A2(n16042), .ZN(n15982) );
  NAND2_X1 U17870 ( .A1(n21337), .A2(n16043), .ZN(n16053) );
  NAND2_X1 U17871 ( .A1(n15982), .A2(n16053), .ZN(n16047) );
  NOR2_X1 U17872 ( .A1(n16047), .A2(n16025), .ZN(n15997) );
  NAND2_X1 U17873 ( .A1(n21337), .A2(n16010), .ZN(n15998) );
  NAND3_X1 U17874 ( .A1(n15997), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15998), .ZN(n15991) );
  NAND2_X1 U17875 ( .A1(n21329), .A2(n21310), .ZN(n21332) );
  NOR2_X1 U17876 ( .A1(n21359), .A2(n21332), .ZN(n21360) );
  INV_X1 U17877 ( .A(n21360), .ZN(n15986) );
  INV_X1 U17878 ( .A(n15983), .ZN(n15985) );
  OAI22_X1 U17879 ( .A1(n15986), .A2(n15985), .B1(n15984), .B2(n21367), .ZN(
        n21403) );
  NAND3_X1 U17880 ( .A1(n21403), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15987), .ZN(n16024) );
  NOR3_X1 U17881 ( .A1(n16024), .A2(n16010), .A3(n16025), .ZN(n16003) );
  AND3_X1 U17882 ( .A1(n16003), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15988), .ZN(n15989) );
  AOI211_X1 U17883 ( .C1(n15992), .C2(n15991), .A(n15990), .B(n15989), .ZN(
        n15995) );
  NAND2_X1 U17884 ( .A1(n15993), .A2(n21409), .ZN(n15994) );
  OAI211_X1 U17885 ( .C1(n15996), .C2(n21335), .A(n15995), .B(n15994), .ZN(
        P1_U3000) );
  OR2_X1 U17886 ( .A1(n16032), .A2(n15997), .ZN(n16011) );
  AOI21_X1 U17887 ( .B1(n16011), .B2(n15998), .A(n16002), .ZN(n16001) );
  INV_X1 U17888 ( .A(n15999), .ZN(n16000) );
  AOI211_X1 U17889 ( .C1(n16003), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        n16006) );
  NAND2_X1 U17890 ( .A1(n16004), .A2(n21409), .ZN(n16005) );
  OAI211_X1 U17891 ( .C1(n16007), .C2(n21335), .A(n16006), .B(n16005), .ZN(
        P1_U3001) );
  INV_X1 U17892 ( .A(n16008), .ZN(n16014) );
  NOR3_X1 U17893 ( .A1(n16024), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16025), .ZN(n16013) );
  OAI21_X1 U17894 ( .B1(n16011), .B2(n16010), .A(n16009), .ZN(n16012) );
  AOI211_X1 U17895 ( .C1(n16014), .C2(n21409), .A(n16013), .B(n16012), .ZN(
        n16015) );
  OAI21_X1 U17896 ( .B1(n16016), .B2(n21335), .A(n16015), .ZN(P1_U3002) );
  INV_X1 U17897 ( .A(n16017), .ZN(n16029) );
  INV_X1 U17898 ( .A(n16018), .ZN(n16023) );
  NAND2_X1 U17899 ( .A1(n16047), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16021) );
  INV_X1 U17900 ( .A(n16019), .ZN(n16020) );
  OAI21_X1 U17901 ( .B1(n16032), .B2(n16021), .A(n16020), .ZN(n16022) );
  AOI21_X1 U17902 ( .B1(n16023), .B2(n21409), .A(n16022), .ZN(n16028) );
  INV_X1 U17903 ( .A(n16024), .ZN(n16039) );
  NAND3_X1 U17904 ( .A1(n16039), .A2(n16026), .A3(n16025), .ZN(n16027) );
  OAI211_X1 U17905 ( .C1(n16029), .C2(n21335), .A(n16028), .B(n16027), .ZN(
        P1_U3003) );
  INV_X1 U17906 ( .A(n16030), .ZN(n16041) );
  NAND2_X1 U17907 ( .A1(n16047), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16031) );
  NOR2_X1 U17908 ( .A1(n16032), .A2(n16031), .ZN(n16037) );
  INV_X1 U17909 ( .A(n16033), .ZN(n16034) );
  OAI21_X1 U17910 ( .B1(n16035), .B2(n21389), .A(n16034), .ZN(n16036) );
  AOI211_X1 U17911 ( .C1(n16039), .C2(n16038), .A(n16037), .B(n16036), .ZN(
        n16040) );
  OAI21_X1 U17912 ( .B1(n16041), .B2(n21335), .A(n16040), .ZN(P1_U3004) );
  INV_X1 U17913 ( .A(n21403), .ZN(n16051) );
  OAI21_X1 U17914 ( .B1(n16051), .B2(n16043), .A(n16042), .ZN(n16048) );
  OAI21_X1 U17915 ( .B1(n16045), .B2(n21389), .A(n16044), .ZN(n16046) );
  AOI21_X1 U17916 ( .B1(n16048), .B2(n16047), .A(n16046), .ZN(n16049) );
  OAI21_X1 U17917 ( .B1(n16050), .B2(n21335), .A(n16049), .ZN(P1_U3005) );
  NOR4_X1 U17918 ( .A1(n16051), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n16066), .A4(n21404), .ZN(n16058) );
  INV_X1 U17919 ( .A(n21405), .ZN(n16061) );
  AOI21_X1 U17920 ( .B1(n16061), .B2(n16053), .A(n16052), .ZN(n16057) );
  NOR2_X1 U17921 ( .A1(n16054), .A2(n21389), .ZN(n16055) );
  NOR4_X1 U17922 ( .A1(n16058), .A2(n16057), .A3(n16056), .A4(n16055), .ZN(
        n16059) );
  OAI21_X1 U17923 ( .B1(n16060), .B2(n21335), .A(n16059), .ZN(P1_U3006) );
  NAND2_X1 U17924 ( .A1(n21404), .A2(n21360), .ZN(n16062) );
  AOI21_X1 U17925 ( .B1(n16062), .B2(n16061), .A(n16066), .ZN(n16063) );
  AOI211_X1 U17926 ( .C1(n21409), .C2(n16065), .A(n16064), .B(n16063), .ZN(
        n16068) );
  NAND3_X1 U17927 ( .A1(n21403), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16066), .ZN(n16067) );
  OAI211_X1 U17928 ( .C1(n16069), .C2(n21335), .A(n16068), .B(n16067), .ZN(
        P1_U3007) );
  NAND2_X1 U17929 ( .A1(n16070), .A2(n21411), .ZN(n16082) );
  OR3_X1 U17930 ( .A1(n16076), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n21287), .ZN(n16081) );
  AOI21_X1 U17931 ( .B1(n21409), .B2(n16072), .A(n16071), .ZN(n16080) );
  NOR2_X1 U17932 ( .A1(n16073), .A2(n21328), .ZN(n16075) );
  AOI211_X1 U17933 ( .C1(n21325), .C2(n16076), .A(n16075), .B(n16074), .ZN(
        n21266) );
  NAND2_X1 U17934 ( .A1(n21265), .A2(n21310), .ZN(n16077) );
  AOI21_X1 U17935 ( .B1(n21266), .B2(n16077), .A(n14235), .ZN(n16078) );
  INV_X1 U17936 ( .A(n16078), .ZN(n16079) );
  NAND4_X1 U17937 ( .A1(n16082), .A2(n16081), .A3(n16080), .A4(n16079), .ZN(
        P1_U3025) );
  AND2_X1 U17938 ( .A1(n16084), .A2(n16083), .ZN(n21559) );
  AOI21_X1 U17939 ( .B1(n16086), .B2(n16085), .A(n21559), .ZN(n16087) );
  OAI21_X1 U17940 ( .B1(n13484), .B2(n21850), .A(n16087), .ZN(n16088) );
  MUX2_X1 U17941 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16088), .S(
        n17061), .Z(P1_U3478) );
  NOR3_X1 U17942 ( .A1(n16089), .A2(n16098), .A3(n16097), .ZN(n16092) );
  NOR2_X1 U17943 ( .A1(n13964), .A2(n16090), .ZN(n16091) );
  AOI211_X1 U17944 ( .C1(n17021), .C2(n16093), .A(n16092), .B(n16091), .ZN(
        n17025) );
  INV_X1 U17945 ( .A(n16094), .ZN(n16981) );
  INV_X1 U17946 ( .A(n16095), .ZN(n16101) );
  NOR3_X1 U17947 ( .A1(n16098), .A2(n16097), .A3(n16096), .ZN(n16099) );
  AOI21_X1 U17948 ( .B1(n16101), .B2(n16100), .A(n16099), .ZN(n16102) );
  OAI21_X1 U17949 ( .B1(n17025), .B2(n16981), .A(n16102), .ZN(n16103) );
  MUX2_X1 U17950 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16103), .S(
        n16984), .Z(P1_U3473) );
  INV_X1 U17951 ( .A(n16104), .ZN(n16245) );
  INV_X1 U17952 ( .A(n19110), .ZN(n16138) );
  AOI21_X1 U17953 ( .B1(n18565), .B2(n16132), .A(n16105), .ZN(n18561) );
  NOR2_X1 U17954 ( .A1(n16130), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16106) );
  OR2_X1 U17955 ( .A1(n16133), .A2(n16106), .ZN(n16412) );
  INV_X1 U17956 ( .A(n16412), .ZN(n16180) );
  INV_X1 U17957 ( .A(n16129), .ZN(n16107) );
  AOI21_X1 U17958 ( .B1(n18548), .B2(n16127), .A(n16107), .ZN(n18546) );
  AOI21_X1 U17959 ( .B1(n16457), .B2(n16124), .A(n16125), .ZN(n16455) );
  INV_X1 U17960 ( .A(n16122), .ZN(n16108) );
  AOI21_X1 U17961 ( .B1(n18514), .B2(n16120), .A(n16108), .ZN(n18524) );
  AOI21_X1 U17962 ( .B1(n16511), .B2(n16116), .A(n16118), .ZN(n18486) );
  INV_X1 U17963 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16109) );
  AOI21_X1 U17964 ( .B1(n16114), .B2(n16109), .A(n16117), .ZN(n18463) );
  NOR2_X1 U17965 ( .A1(n16110), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16111) );
  OR2_X1 U17966 ( .A1(n16113), .A2(n16111), .ZN(n16560) );
  INV_X1 U17967 ( .A(n16560), .ZN(n18438) );
  NAND2_X1 U17968 ( .A1(n16112), .A2(n16571), .ZN(n18437) );
  NOR2_X1 U17969 ( .A1(n18438), .A2(n18437), .ZN(n18449) );
  OR2_X1 U17970 ( .A1(n16113), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16115) );
  AND2_X1 U17971 ( .A1(n16115), .A2(n16114), .ZN(n18451) );
  INV_X1 U17972 ( .A(n18451), .ZN(n16543) );
  NAND2_X1 U17973 ( .A1(n18449), .A2(n16543), .ZN(n18461) );
  NOR2_X1 U17974 ( .A1(n18463), .A2(n18461), .ZN(n18473) );
  OAI21_X1 U17975 ( .B1(n16117), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16116), .ZN(n18474) );
  NAND2_X1 U17976 ( .A1(n18473), .A2(n18474), .ZN(n18484) );
  NOR2_X1 U17977 ( .A1(n18486), .A2(n18484), .ZN(n18504) );
  OR2_X1 U17978 ( .A1(n16118), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16119) );
  NAND2_X1 U17979 ( .A1(n16120), .A2(n16119), .ZN(n18508) );
  NAND2_X1 U17980 ( .A1(n18504), .A2(n18508), .ZN(n18503) );
  NOR2_X1 U17981 ( .A1(n18524), .A2(n18503), .ZN(n18534) );
  NAND2_X1 U17982 ( .A1(n16122), .A2(n16121), .ZN(n16123) );
  NAND2_X1 U17983 ( .A1(n16124), .A2(n16123), .ZN(n18533) );
  NAND2_X1 U17984 ( .A1(n18534), .A2(n18533), .ZN(n16214) );
  NOR2_X1 U17985 ( .A1(n16455), .A2(n16214), .ZN(n16206) );
  OR2_X1 U17986 ( .A1(n16125), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16126) );
  NAND2_X1 U17987 ( .A1(n16127), .A2(n16126), .ZN(n16446) );
  NAND2_X1 U17988 ( .A1(n16206), .A2(n16446), .ZN(n18543) );
  NOR2_X1 U17989 ( .A1(n18546), .A2(n18543), .ZN(n16192) );
  AND2_X1 U17990 ( .A1(n16129), .A2(n16128), .ZN(n16131) );
  OR2_X1 U17991 ( .A1(n16131), .A2(n16130), .ZN(n16428) );
  NAND2_X1 U17992 ( .A1(n16192), .A2(n16428), .ZN(n16177) );
  NOR2_X1 U17993 ( .A1(n16180), .A2(n16177), .ZN(n16157) );
  OAI21_X1 U17994 ( .B1(n16133), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16132), .ZN(n16404) );
  NAND2_X1 U17995 ( .A1(n16157), .A2(n16404), .ZN(n18556) );
  NOR2_X1 U17996 ( .A1(n18561), .A2(n18556), .ZN(n16143) );
  AND4_X1 U17997 ( .A1(n18558), .A2(n16143), .A3(n16144), .A4(n10997), .ZN(
        n16136) );
  OAI22_X1 U17998 ( .A1(n16247), .A2(n16134), .B1(n13416), .B2(n18562), .ZN(
        n16135) );
  AOI211_X1 U17999 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n18529), .A(
        n16136), .B(n16135), .ZN(n16137) );
  OAI21_X1 U18000 ( .B1(n16138), .B2(n18576), .A(n16137), .ZN(n16139) );
  AOI21_X1 U18001 ( .B1(n16245), .B2(n18570), .A(n16139), .ZN(n16140) );
  OAI21_X1 U18002 ( .B1(n16141), .B2(n18509), .A(n16140), .ZN(P2_U2824) );
  INV_X1 U18003 ( .A(n16142), .ZN(n16154) );
  NOR2_X1 U18004 ( .A1(n18535), .A2(n16143), .ZN(n16145) );
  XNOR2_X1 U18005 ( .A(n16145), .B(n16144), .ZN(n16146) );
  AOI22_X1 U18006 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18568), .B1(n18558), 
        .B2(n16146), .ZN(n16147) );
  OAI21_X1 U18007 ( .B1(n17386), .B2(n18562), .A(n16147), .ZN(n16151) );
  INV_X1 U18008 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16148) );
  OAI22_X1 U18009 ( .A1(n16149), .A2(n18576), .B1(n18564), .B2(n16148), .ZN(
        n16150) );
  AOI211_X1 U18010 ( .C1(n16152), .C2(n18570), .A(n16151), .B(n16150), .ZN(
        n16153) );
  OAI21_X1 U18011 ( .B1(n16154), .B2(n18509), .A(n16153), .ZN(P2_U2825) );
  AOI21_X1 U18012 ( .B1(n16156), .B2(n16170), .A(n16155), .ZN(n16646) );
  NOR2_X1 U18013 ( .A1(n18535), .A2(n16157), .ZN(n16158) );
  XNOR2_X1 U18014 ( .A(n16158), .B(n16404), .ZN(n16159) );
  AOI22_X1 U18015 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18568), .B1(n18558), 
        .B2(n16159), .ZN(n16160) );
  OAI21_X1 U18016 ( .B1(n17385), .B2(n18562), .A(n16160), .ZN(n16167) );
  NOR2_X1 U18017 ( .A1(n16162), .A2(n16161), .ZN(n16163) );
  INV_X1 U18018 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16165) );
  OAI22_X1 U18019 ( .A1(n16647), .A2(n18576), .B1(n18564), .B2(n16165), .ZN(
        n16166) );
  AOI211_X1 U18020 ( .C1(n16646), .C2(n18570), .A(n16167), .B(n16166), .ZN(
        n16168) );
  OAI21_X1 U18021 ( .B1(n16169), .B2(n18509), .A(n16168), .ZN(P2_U2827) );
  AOI21_X1 U18022 ( .B1(n16171), .B2(n16188), .A(n13160), .ZN(n16671) );
  XNOR2_X1 U18023 ( .A(n11020), .B(n16172), .ZN(n16659) );
  INV_X1 U18024 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16173) );
  OAI22_X1 U18025 ( .A1(n16173), .A2(n18564), .B1(n17384), .B2(n18562), .ZN(
        n16174) );
  AOI21_X1 U18026 ( .B1(n18568), .B2(P2_EBX_REG_27__SCAN_IN), .A(n16174), .ZN(
        n16175) );
  OAI21_X1 U18027 ( .B1(n16659), .B2(n18576), .A(n16175), .ZN(n16176) );
  AOI21_X1 U18028 ( .B1(n16671), .B2(n18570), .A(n16176), .ZN(n16183) );
  AND2_X1 U18029 ( .A1(n10997), .A2(n16177), .ZN(n16179) );
  OAI21_X1 U18030 ( .B1(n16180), .B2(n16179), .A(n18558), .ZN(n16178) );
  AOI21_X1 U18031 ( .B1(n16180), .B2(n16179), .A(n16178), .ZN(n16181) );
  INV_X1 U18032 ( .A(n16181), .ZN(n16182) );
  OAI211_X1 U18033 ( .C1(n18509), .C2(n16184), .A(n16183), .B(n16182), .ZN(
        P2_U2828) );
  INV_X1 U18034 ( .A(n16185), .ZN(n16200) );
  OR2_X1 U18035 ( .A1(n16273), .A2(n16186), .ZN(n16187) );
  NAND2_X1 U18036 ( .A1(n16188), .A2(n16187), .ZN(n16682) );
  INV_X1 U18037 ( .A(n16682), .ZN(n16198) );
  NAND2_X1 U18038 ( .A1(n16335), .A2(n16189), .ZN(n16190) );
  NAND2_X1 U18039 ( .A1(n11020), .A2(n16190), .ZN(n16677) );
  INV_X1 U18040 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16191) );
  OAI22_X1 U18041 ( .A1(n16677), .A2(n18576), .B1(n18516), .B2(n16191), .ZN(
        n16197) );
  NOR2_X1 U18042 ( .A1(n18535), .A2(n16192), .ZN(n16193) );
  XOR2_X1 U18043 ( .A(n16428), .B(n16193), .Z(n16195) );
  AOI22_X1 U18044 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18529), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18528), .ZN(n16194) );
  OAI21_X1 U18045 ( .B1(n18643), .B2(n16195), .A(n16194), .ZN(n16196) );
  AOI211_X1 U18046 ( .C1(n18570), .C2(n16198), .A(n16197), .B(n16196), .ZN(
        n16199) );
  OAI21_X1 U18047 ( .B1(n16200), .B2(n18509), .A(n16199), .ZN(P2_U2829) );
  NAND2_X1 U18048 ( .A1(n16218), .A2(n16201), .ZN(n16202) );
  NAND2_X1 U18049 ( .A1(n16274), .A2(n16202), .ZN(n16697) );
  AND2_X1 U18050 ( .A1(n16221), .A2(n16203), .ZN(n16204) );
  NOR2_X1 U18051 ( .A1(n16333), .A2(n16204), .ZN(n16699) );
  AOI22_X1 U18052 ( .A1(n16699), .A2(n18531), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n18568), .ZN(n16205) );
  OAI21_X1 U18053 ( .B1(n16697), .B2(n18511), .A(n16205), .ZN(n16211) );
  NOR2_X1 U18054 ( .A1(n18535), .A2(n16206), .ZN(n16207) );
  XOR2_X1 U18055 ( .A(n16446), .B(n16207), .Z(n16209) );
  AOI22_X1 U18056 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18529), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18528), .ZN(n16208) );
  OAI21_X1 U18057 ( .B1(n18643), .B2(n16209), .A(n16208), .ZN(n16210) );
  AOI211_X1 U18058 ( .C1(n18572), .C2(n16212), .A(n16211), .B(n16210), .ZN(
        n16213) );
  INV_X1 U18059 ( .A(n16213), .ZN(P2_U2831) );
  AND2_X1 U18060 ( .A1(n10997), .A2(n16214), .ZN(n16216) );
  OAI21_X1 U18061 ( .B1(n16455), .B2(n16216), .A(n18558), .ZN(n16215) );
  AOI21_X1 U18062 ( .B1(n16455), .B2(n16216), .A(n16215), .ZN(n16217) );
  INV_X1 U18063 ( .A(n16217), .ZN(n16229) );
  INV_X1 U18064 ( .A(n16218), .ZN(n16219) );
  AOI21_X1 U18065 ( .B1(n16220), .B2(n16291), .A(n16219), .ZN(n16719) );
  INV_X1 U18066 ( .A(n16221), .ZN(n16222) );
  AOI21_X1 U18067 ( .B1(n16223), .B2(n16723), .A(n16222), .ZN(n16712) );
  INV_X1 U18068 ( .A(n16712), .ZN(n16226) );
  OAI22_X1 U18069 ( .A1(n16457), .A2(n18564), .B1(n17380), .B2(n18562), .ZN(
        n16224) );
  AOI21_X1 U18070 ( .B1(n18568), .B2(P2_EBX_REG_23__SCAN_IN), .A(n16224), .ZN(
        n16225) );
  OAI21_X1 U18071 ( .B1(n16226), .B2(n18576), .A(n16225), .ZN(n16227) );
  AOI21_X1 U18072 ( .B1(n16719), .B2(n18570), .A(n16227), .ZN(n16228) );
  OAI211_X1 U18073 ( .C1(n18509), .C2(n16230), .A(n16229), .B(n16228), .ZN(
        P2_U2832) );
  AOI211_X1 U18074 ( .C1(n18348), .C2(n16232), .A(n18535), .B(n16231), .ZN(
        n16964) );
  NAND2_X1 U18075 ( .A1(n16964), .A2(n18558), .ZN(n16243) );
  INV_X1 U18076 ( .A(n16233), .ZN(n16239) );
  NAND2_X1 U18077 ( .A1(n18568), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n16238) );
  NAND2_X1 U18078 ( .A1(n18558), .A2(n18535), .ZN(n18507) );
  AOI22_X1 U18079 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18529), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18528), .ZN(n16234) );
  OAI21_X1 U18080 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18507), .A(
        n16234), .ZN(n16235) );
  AOI21_X1 U18081 ( .B1(n18531), .B2(n16236), .A(n16235), .ZN(n16237) );
  OAI211_X1 U18082 ( .C1(n18509), .C2(n16239), .A(n16238), .B(n16237), .ZN(
        n16240) );
  AOI21_X1 U18083 ( .B1(n18570), .B2(n16241), .A(n16240), .ZN(n16242) );
  OAI211_X1 U18084 ( .C1(n17320), .C2(n16244), .A(n16243), .B(n16242), .ZN(
        P2_U2854) );
  NAND2_X1 U18085 ( .A1(n16245), .A2(n16284), .ZN(n16246) );
  OAI21_X1 U18086 ( .B1(n16284), .B2(n16247), .A(n16246), .ZN(P2_U2856) );
  INV_X1 U18087 ( .A(n16248), .ZN(n16249) );
  NOR2_X1 U18088 ( .A1(n16250), .A2(n16249), .ZN(n16252) );
  XNOR2_X1 U18089 ( .A(n16252), .B(n16251), .ZN(n16315) );
  NOR2_X1 U18090 ( .A1(n18569), .A2(n14161), .ZN(n16253) );
  AOI21_X1 U18091 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n14161), .A(n16253), .ZN(
        n16254) );
  OAI21_X1 U18092 ( .B1(n16315), .B2(n16302), .A(n16254), .ZN(P2_U2858) );
  NAND2_X1 U18093 ( .A1(n11327), .A2(n16255), .ZN(n16257) );
  XNOR2_X1 U18094 ( .A(n16257), .B(n16256), .ZN(n16321) );
  NAND2_X1 U18095 ( .A1(n14161), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16259) );
  NAND2_X1 U18096 ( .A1(n16646), .A2(n16284), .ZN(n16258) );
  OAI211_X1 U18097 ( .C1(n16321), .C2(n16302), .A(n16259), .B(n16258), .ZN(
        P2_U2859) );
  NAND2_X1 U18098 ( .A1(n11327), .A2(n16260), .ZN(n16261) );
  XOR2_X1 U18099 ( .A(n16262), .B(n16261), .Z(n16326) );
  NAND2_X1 U18100 ( .A1(n14161), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16264) );
  NAND2_X1 U18101 ( .A1(n16671), .A2(n16284), .ZN(n16263) );
  OAI211_X1 U18102 ( .C1(n16326), .C2(n16302), .A(n16264), .B(n16263), .ZN(
        P2_U2860) );
  AOI21_X1 U18103 ( .B1(n16267), .B2(n16266), .A(n16265), .ZN(n16330) );
  NAND2_X1 U18104 ( .A1(n16330), .A2(n16307), .ZN(n16269) );
  NAND2_X1 U18105 ( .A1(n14161), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16268) );
  OAI211_X1 U18106 ( .C1(n16682), .C2(n14161), .A(n16269), .B(n16268), .ZN(
        P2_U2861) );
  OAI21_X1 U18107 ( .B1(n16272), .B2(n16271), .A(n16270), .ZN(n16341) );
  NAND2_X1 U18108 ( .A1(n14161), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16277) );
  AOI21_X1 U18109 ( .B1(n16275), .B2(n16274), .A(n16273), .ZN(n18552) );
  NAND2_X1 U18110 ( .A1(n18552), .A2(n16284), .ZN(n16276) );
  OAI211_X1 U18111 ( .C1(n16341), .C2(n16302), .A(n16277), .B(n16276), .ZN(
        P2_U2862) );
  OAI21_X1 U18112 ( .B1(n16280), .B2(n16279), .A(n16278), .ZN(n16351) );
  NOR2_X1 U18113 ( .A1(n16697), .A2(n14161), .ZN(n16281) );
  AOI21_X1 U18114 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14161), .A(n16281), .ZN(
        n16282) );
  OAI21_X1 U18115 ( .B1(n16351), .B2(n16302), .A(n16282), .ZN(P2_U2863) );
  XNOR2_X1 U18116 ( .A(n11005), .B(n16283), .ZN(n16359) );
  NAND2_X1 U18117 ( .A1(n14161), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16286) );
  NAND2_X1 U18118 ( .A1(n16719), .A2(n16284), .ZN(n16285) );
  OAI211_X1 U18119 ( .C1(n16359), .C2(n16302), .A(n16286), .B(n16285), .ZN(
        P2_U2864) );
  OAI21_X1 U18120 ( .B1(n16287), .B2(n16288), .A(n11005), .ZN(n19298) );
  OR2_X1 U18121 ( .A1(n16299), .A2(n16289), .ZN(n16290) );
  NAND2_X1 U18122 ( .A1(n16291), .A2(n16290), .ZN(n16730) );
  NOR2_X1 U18123 ( .A1(n16730), .A2(n14161), .ZN(n16292) );
  AOI21_X1 U18124 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n14161), .A(n16292), .ZN(
        n16293) );
  OAI21_X1 U18125 ( .B1(n19298), .B2(n16302), .A(n16293), .ZN(P2_U2865) );
  INV_X1 U18126 ( .A(n16287), .ZN(n16295) );
  OAI21_X1 U18127 ( .B1(n16294), .B2(n16296), .A(n16295), .ZN(n16360) );
  NOR2_X1 U18128 ( .A1(n16303), .A2(n16297), .ZN(n16298) );
  OR2_X1 U18129 ( .A1(n16299), .A2(n16298), .ZN(n18512) );
  NOR2_X1 U18130 ( .A1(n18512), .A2(n14161), .ZN(n16300) );
  AOI21_X1 U18131 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n14161), .A(n16300), .ZN(
        n16301) );
  OAI21_X1 U18132 ( .B1(n16360), .B2(n16302), .A(n16301), .ZN(P2_U2866) );
  AOI21_X1 U18133 ( .B1(n16304), .B2(n11018), .A(n16303), .ZN(n16769) );
  INV_X1 U18134 ( .A(n16769), .ZN(n18500) );
  AOI21_X1 U18135 ( .B1(n16306), .B2(n16305), .A(n16294), .ZN(n19396) );
  NAND2_X1 U18136 ( .A1(n19396), .A2(n16307), .ZN(n16309) );
  NAND2_X1 U18137 ( .A1(n14161), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16308) );
  OAI211_X1 U18138 ( .C1(n18500), .C2(n14161), .A(n16309), .B(n16308), .ZN(
        P2_U2867) );
  AOI22_X1 U18139 ( .A1(n19582), .A2(BUF2_REG_29__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16312) );
  AOI22_X1 U18140 ( .A1(n19583), .A2(BUF1_REG_29__SCAN_IN), .B1(n19581), .B2(
        n16310), .ZN(n16311) );
  OAI211_X1 U18141 ( .C1(n18577), .C2(n16373), .A(n16312), .B(n16311), .ZN(
        n16313) );
  INV_X1 U18142 ( .A(n16313), .ZN(n16314) );
  OAI21_X1 U18143 ( .B1(n16315), .B2(n19342), .A(n16314), .ZN(P2_U2890) );
  AOI22_X1 U18144 ( .A1(n19583), .A2(BUF1_REG_28__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U18145 ( .A1(n19582), .A2(BUF2_REG_28__SCAN_IN), .B1(n19581), .B2(
        n16316), .ZN(n16317) );
  OAI211_X1 U18146 ( .C1(n16647), .C2(n16373), .A(n16318), .B(n16317), .ZN(
        n16319) );
  INV_X1 U18147 ( .A(n16319), .ZN(n16320) );
  OAI21_X1 U18148 ( .B1(n16321), .B2(n19342), .A(n16320), .ZN(P2_U2891) );
  AOI22_X1 U18149 ( .A1(n19583), .A2(BUF1_REG_27__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16323) );
  AOI22_X1 U18150 ( .A1(n19582), .A2(BUF2_REG_27__SCAN_IN), .B1(n19581), .B2(
        n19113), .ZN(n16322) );
  OAI211_X1 U18151 ( .C1(n16659), .C2(n16373), .A(n16323), .B(n16322), .ZN(
        n16324) );
  INV_X1 U18152 ( .A(n16324), .ZN(n16325) );
  OAI21_X1 U18153 ( .B1(n16326), .B2(n19342), .A(n16325), .ZN(P2_U2892) );
  AOI22_X1 U18154 ( .A1(n19583), .A2(BUF1_REG_26__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16328) );
  AOI22_X1 U18155 ( .A1(n19582), .A2(BUF2_REG_26__SCAN_IN), .B1(n19581), .B2(
        n19116), .ZN(n16327) );
  OAI211_X1 U18156 ( .C1(n16677), .C2(n16373), .A(n16328), .B(n16327), .ZN(
        n16329) );
  AOI21_X1 U18157 ( .B1(n16330), .B2(n19586), .A(n16329), .ZN(n16331) );
  INV_X1 U18158 ( .A(n16331), .ZN(P2_U2893) );
  OR2_X1 U18159 ( .A1(n16333), .A2(n16332), .ZN(n16334) );
  NAND2_X1 U18160 ( .A1(n16335), .A2(n16334), .ZN(n18555) );
  AOI22_X1 U18161 ( .A1(n19582), .A2(BUF2_REG_25__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16338) );
  AOI22_X1 U18162 ( .A1(n19583), .A2(BUF1_REG_25__SCAN_IN), .B1(n19581), .B2(
        n16336), .ZN(n16337) );
  OAI211_X1 U18163 ( .C1(n18555), .C2(n16373), .A(n16338), .B(n16337), .ZN(
        n16339) );
  INV_X1 U18164 ( .A(n16339), .ZN(n16340) );
  OAI21_X1 U18165 ( .B1(n16341), .B2(n19342), .A(n16340), .ZN(P2_U2894) );
  INV_X1 U18166 ( .A(n19583), .ZN(n16355) );
  INV_X1 U18167 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16343) );
  OAI22_X1 U18168 ( .A1(n16355), .A2(n16343), .B1(n16342), .B2(n19496), .ZN(
        n16349) );
  INV_X1 U18169 ( .A(n19581), .ZN(n16346) );
  INV_X1 U18170 ( .A(n19582), .ZN(n16345) );
  INV_X1 U18171 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16344) );
  OAI22_X1 U18172 ( .A1(n16347), .A2(n16346), .B1(n16345), .B2(n16344), .ZN(
        n16348) );
  AOI211_X1 U18173 ( .C1(n16699), .C2(n19585), .A(n16349), .B(n16348), .ZN(
        n16350) );
  OAI21_X1 U18174 ( .B1(n16351), .B2(n19342), .A(n16350), .ZN(P2_U2895) );
  INV_X1 U18175 ( .A(n16352), .ZN(n16353) );
  AOI22_X1 U18176 ( .A1(n19582), .A2(BUF2_REG_23__SCAN_IN), .B1(n19581), .B2(
        n16353), .ZN(n16358) );
  OAI22_X1 U18177 ( .A1(n16355), .A2(n22135), .B1(n16354), .B2(n19496), .ZN(
        n16356) );
  AOI21_X1 U18178 ( .B1(n16712), .B2(n19585), .A(n16356), .ZN(n16357) );
  OAI211_X1 U18179 ( .C1(n16359), .C2(n19342), .A(n16358), .B(n16357), .ZN(
        P2_U2896) );
  OR2_X1 U18180 ( .A1(n16360), .A2(n19342), .ZN(n16369) );
  OR2_X1 U18181 ( .A1(n16768), .A2(n16361), .ZN(n16362) );
  NAND2_X1 U18182 ( .A1(n16725), .A2(n16362), .ZN(n18527) );
  OAI22_X1 U18183 ( .A1(n18527), .A2(n16373), .B1(n16363), .B2(n19496), .ZN(
        n16364) );
  INV_X1 U18184 ( .A(n16364), .ZN(n16368) );
  INV_X1 U18185 ( .A(n16365), .ZN(n19341) );
  AOI22_X1 U18186 ( .A1(n19583), .A2(BUF1_REG_21__SCAN_IN), .B1(n19581), .B2(
        n19341), .ZN(n16367) );
  NAND2_X1 U18187 ( .A1(n19582), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16366) );
  NAND4_X1 U18188 ( .A1(n16369), .A2(n16368), .A3(n16367), .A4(n16366), .ZN(
        P2_U2898) );
  AND2_X1 U18189 ( .A1(n16793), .A2(n16370), .ZN(n16371) );
  OR2_X1 U18190 ( .A1(n16371), .A2(n16766), .ZN(n18492) );
  OAI22_X1 U18191 ( .A1(n18492), .A2(n16373), .B1(n16372), .B2(n19496), .ZN(
        n16374) );
  AOI21_X1 U18192 ( .B1(n19582), .B2(BUF2_REG_19__SCAN_IN), .A(n16374), .ZN(
        n16377) );
  AOI22_X1 U18193 ( .A1(n19583), .A2(BUF1_REG_19__SCAN_IN), .B1(n19581), .B2(
        n16375), .ZN(n16376) );
  OAI211_X1 U18194 ( .C1(n16378), .C2(n19342), .A(n16377), .B(n16376), .ZN(
        P2_U2900) );
  OR2_X1 U18195 ( .A1(n16379), .A2(n19342), .ZN(n16387) );
  INV_X1 U18196 ( .A(n16381), .ZN(n16382) );
  XNOR2_X1 U18197 ( .A(n16380), .B(n16382), .ZN(n18468) );
  AOI22_X1 U18198 ( .A1(n19585), .A2(n18468), .B1(n19579), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16386) );
  AOI22_X1 U18199 ( .A1(n19583), .A2(BUF1_REG_17__SCAN_IN), .B1(n19581), .B2(
        n16383), .ZN(n16385) );
  NAND2_X1 U18200 ( .A1(n19582), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16384) );
  NAND4_X1 U18201 ( .A1(n16387), .A2(n16386), .A3(n16385), .A4(n16384), .ZN(
        P2_U2902) );
  OAI21_X1 U18202 ( .B1(n17268), .B2(n18565), .A(n16388), .ZN(n16389) );
  AOI21_X1 U18203 ( .B1(n17260), .B2(n18561), .A(n16389), .ZN(n16390) );
  OAI21_X1 U18204 ( .B1(n18569), .B2(n17296), .A(n16390), .ZN(n16391) );
  AOI21_X1 U18205 ( .B1(n16392), .B2(n17270), .A(n16391), .ZN(n16393) );
  OAI21_X1 U18206 ( .B1(n16394), .B2(n17295), .A(n16393), .ZN(P2_U2985) );
  INV_X1 U18207 ( .A(n16396), .ZN(n16397) );
  NAND2_X1 U18208 ( .A1(n16398), .A2(n16397), .ZN(n16407) );
  NOR2_X1 U18209 ( .A1(n16398), .A2(n16397), .ZN(n16409) );
  AOI21_X1 U18210 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16407), .A(
        n16409), .ZN(n16401) );
  XNOR2_X1 U18211 ( .A(n16399), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16400) );
  XNOR2_X1 U18212 ( .A(n16401), .B(n16400), .ZN(n16658) );
  XNOR2_X1 U18213 ( .A(n16414), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16656) );
  NAND2_X1 U18214 ( .A1(n16646), .A2(n17273), .ZN(n16403) );
  NOR2_X1 U18215 ( .A1(n18488), .A2(n17385), .ZN(n16649) );
  AOI21_X1 U18216 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16649), .ZN(n16402) );
  OAI211_X1 U18217 ( .C1(n17301), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        n16405) );
  AOI21_X1 U18218 ( .B1(n16656), .B2(n17270), .A(n16405), .ZN(n16406) );
  OAI21_X1 U18219 ( .B1(n16658), .B2(n17295), .A(n16406), .ZN(P2_U2986) );
  INV_X1 U18220 ( .A(n16407), .ZN(n16408) );
  NOR2_X1 U18221 ( .A1(n16409), .A2(n16408), .ZN(n16410) );
  XNOR2_X1 U18222 ( .A(n16410), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16673) );
  NOR2_X1 U18223 ( .A1(n18488), .A2(n17384), .ZN(n16663) );
  AOI21_X1 U18224 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16663), .ZN(n16411) );
  OAI21_X1 U18225 ( .B1(n17301), .B2(n16412), .A(n16411), .ZN(n16416) );
  NAND2_X1 U18226 ( .A1(n16424), .A2(n16666), .ZN(n16413) );
  NAND2_X1 U18227 ( .A1(n16414), .A2(n16413), .ZN(n16668) );
  NOR2_X1 U18228 ( .A1(n16668), .A2(n17294), .ZN(n16415) );
  OAI21_X1 U18229 ( .B1(n16673), .B2(n17295), .A(n16417), .ZN(P2_U2987) );
  INV_X1 U18230 ( .A(n16437), .ZN(n16418) );
  AOI21_X1 U18231 ( .B1(n16418), .B2(n16433), .A(n16434), .ZN(n16420) );
  MUX2_X1 U18232 ( .A(n16433), .B(n16420), .S(n16419), .Z(n16423) );
  INV_X1 U18233 ( .A(n16421), .ZN(n16422) );
  NAND2_X1 U18234 ( .A1(n16423), .A2(n16422), .ZN(n16686) );
  INV_X1 U18235 ( .A(n16424), .ZN(n16426) );
  AOI21_X1 U18236 ( .B1(n16441), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16425) );
  NOR2_X1 U18237 ( .A1(n16426), .A2(n16425), .ZN(n16684) );
  NOR2_X1 U18238 ( .A1(n16682), .A2(n17296), .ZN(n16430) );
  NAND2_X1 U18239 ( .A1(n18427), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16676) );
  NAND2_X1 U18240 ( .A1(n17286), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16427) );
  OAI211_X1 U18241 ( .C1(n17301), .C2(n16428), .A(n16676), .B(n16427), .ZN(
        n16429) );
  AOI211_X1 U18242 ( .C1(n16684), .C2(n17270), .A(n16430), .B(n16429), .ZN(
        n16431) );
  OAI21_X1 U18243 ( .B1(n16686), .B2(n17295), .A(n16431), .ZN(P2_U2988) );
  XNOR2_X1 U18244 ( .A(n16441), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16696) );
  NAND2_X1 U18245 ( .A1(n17260), .A2(n18546), .ZN(n16432) );
  NAND2_X1 U18246 ( .A1(n18427), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16687) );
  OAI211_X1 U18247 ( .C1(n17268), .C2(n18548), .A(n16432), .B(n16687), .ZN(
        n16439) );
  INV_X1 U18248 ( .A(n16433), .ZN(n16435) );
  NOR2_X1 U18249 ( .A1(n16435), .A2(n16434), .ZN(n16436) );
  NOR2_X1 U18250 ( .A1(n16692), .A2(n17295), .ZN(n16438) );
  AOI211_X1 U18251 ( .C1(n17273), .C2(n18552), .A(n16439), .B(n16438), .ZN(
        n16440) );
  OAI21_X1 U18252 ( .B1(n17294), .B2(n16696), .A(n16440), .ZN(P2_U2989) );
  INV_X1 U18253 ( .A(n16441), .ZN(n16442) );
  OAI21_X1 U18254 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16453), .A(
        n16442), .ZN(n16708) );
  XNOR2_X1 U18255 ( .A(n16443), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16444) );
  XNOR2_X1 U18256 ( .A(n16445), .B(n16444), .ZN(n16706) );
  INV_X1 U18257 ( .A(n16446), .ZN(n16449) );
  INV_X1 U18258 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16447) );
  NAND2_X1 U18259 ( .A1(n18427), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16700) );
  OAI21_X1 U18260 ( .B1(n17268), .B2(n16447), .A(n16700), .ZN(n16448) );
  AOI21_X1 U18261 ( .B1(n17260), .B2(n16449), .A(n16448), .ZN(n16450) );
  OAI21_X1 U18262 ( .B1(n16697), .B2(n17296), .A(n16450), .ZN(n16451) );
  AOI21_X1 U18263 ( .B1(n16706), .B2(n17274), .A(n16451), .ZN(n16452) );
  OAI21_X1 U18264 ( .B1(n16708), .B2(n17294), .A(n16452), .ZN(P2_U2990) );
  INV_X1 U18265 ( .A(n16453), .ZN(n16454) );
  OAI21_X1 U18266 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16470), .A(
        n16454), .ZN(n16721) );
  NAND2_X1 U18267 ( .A1(n17260), .A2(n16455), .ZN(n16456) );
  NAND2_X1 U18268 ( .A1(n18427), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16709) );
  OAI211_X1 U18269 ( .C1(n17268), .C2(n16457), .A(n16456), .B(n16709), .ZN(
        n16464) );
  INV_X1 U18270 ( .A(n16458), .ZN(n16460) );
  NOR2_X1 U18271 ( .A1(n16460), .A2(n16459), .ZN(n16461) );
  XNOR2_X1 U18272 ( .A(n16462), .B(n16461), .ZN(n16716) );
  NOR2_X1 U18273 ( .A1(n16716), .A2(n17295), .ZN(n16463) );
  AOI211_X1 U18274 ( .C1(n17273), .C2(n16719), .A(n16464), .B(n16463), .ZN(
        n16465) );
  OAI21_X1 U18275 ( .B1(n17294), .B2(n16721), .A(n16465), .ZN(P2_U2991) );
  XNOR2_X1 U18276 ( .A(n16467), .B(n16733), .ZN(n16468) );
  XNOR2_X1 U18277 ( .A(n16469), .B(n16468), .ZN(n16737) );
  AOI21_X1 U18278 ( .B1(n16733), .B2(n16492), .A(n16470), .ZN(n16722) );
  NAND2_X1 U18279 ( .A1(n16722), .A2(n17270), .ZN(n16474) );
  INV_X1 U18280 ( .A(n16730), .ZN(n18532) );
  NAND2_X1 U18281 ( .A1(n18427), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16727) );
  NAND2_X1 U18282 ( .A1(n17286), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16471) );
  OAI211_X1 U18283 ( .C1(n17301), .C2(n18533), .A(n16727), .B(n16471), .ZN(
        n16472) );
  AOI21_X1 U18284 ( .B1(n18532), .B2(n17273), .A(n16472), .ZN(n16473) );
  OAI211_X1 U18285 ( .C1(n16737), .C2(n17295), .A(n16474), .B(n16473), .ZN(
        P2_U2992) );
  INV_X1 U18286 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16864) );
  NAND2_X1 U18287 ( .A1(n16477), .A2(n16864), .ZN(n16587) );
  OAI21_X1 U18288 ( .B1(n16588), .B2(n16586), .A(n16587), .ZN(n16554) );
  NAND2_X1 U18289 ( .A1(n16554), .A2(n16478), .ZN(n16529) );
  INV_X1 U18290 ( .A(n16479), .ZN(n16480) );
  AOI21_X1 U18291 ( .B1(n16529), .B2(n16481), .A(n16480), .ZN(n16520) );
  INV_X1 U18292 ( .A(n16482), .ZN(n16483) );
  AOI21_X1 U18293 ( .B1(n16520), .B2(n16484), .A(n16483), .ZN(n16485) );
  XNOR2_X1 U18294 ( .A(n16485), .B(n16486), .ZN(n16503) );
  INV_X1 U18295 ( .A(n16503), .ZN(n16487) );
  AOI22_X1 U18296 ( .A1(n16487), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16486), .B2(n16485), .ZN(n16491) );
  NAND2_X1 U18297 ( .A1(n16489), .A2(n16488), .ZN(n16490) );
  XNOR2_X1 U18298 ( .A(n16491), .B(n16490), .ZN(n16748) );
  INV_X1 U18299 ( .A(n16492), .ZN(n16493) );
  AOI21_X1 U18300 ( .B1(n16494), .B2(n16499), .A(n16493), .ZN(n16746) );
  NOR2_X1 U18301 ( .A1(n18600), .A2(n18513), .ZN(n16740) );
  NOR2_X1 U18302 ( .A1(n17268), .A2(n18514), .ZN(n16495) );
  AOI211_X1 U18303 ( .C1(n18524), .C2(n17260), .A(n16740), .B(n16495), .ZN(
        n16496) );
  OAI21_X1 U18304 ( .B1(n18512), .B2(n17296), .A(n16496), .ZN(n16497) );
  AOI21_X1 U18305 ( .B1(n16746), .B2(n17270), .A(n16497), .ZN(n16498) );
  OAI21_X1 U18306 ( .B1(n16748), .B2(n17295), .A(n16498), .ZN(P2_U2993) );
  NAND2_X1 U18307 ( .A1(n16500), .A2(n16499), .ZN(n16776) );
  NAND2_X1 U18308 ( .A1(n18427), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16770) );
  NAND2_X1 U18309 ( .A1(n17286), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16501) );
  OAI211_X1 U18310 ( .C1(n17301), .C2(n18508), .A(n16770), .B(n16501), .ZN(
        n16502) );
  AOI21_X1 U18311 ( .B1(n16769), .B2(n17273), .A(n16502), .ZN(n16505) );
  XNOR2_X1 U18312 ( .A(n16503), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16774) );
  NAND2_X1 U18313 ( .A1(n16774), .A2(n17274), .ZN(n16504) );
  OAI211_X1 U18314 ( .C1(n16776), .C2(n17294), .A(n16505), .B(n16504), .ZN(
        P2_U2994) );
  XNOR2_X1 U18315 ( .A(n16517), .B(n16783), .ZN(n16788) );
  INV_X1 U18316 ( .A(n16519), .ZN(n16506) );
  AOI21_X1 U18317 ( .B1(n16520), .B2(n16518), .A(n16506), .ZN(n16510) );
  NAND2_X1 U18318 ( .A1(n16508), .A2(n16507), .ZN(n16509) );
  XNOR2_X1 U18319 ( .A(n16510), .B(n16509), .ZN(n16786) );
  NAND2_X1 U18320 ( .A1(n18427), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16778) );
  OAI21_X1 U18321 ( .B1(n17268), .B2(n16511), .A(n16778), .ZN(n16512) );
  AOI21_X1 U18322 ( .B1(n17260), .B2(n18486), .A(n16512), .ZN(n16513) );
  OAI21_X1 U18323 ( .B1(n18493), .B2(n17296), .A(n16513), .ZN(n16514) );
  AOI21_X1 U18324 ( .B1(n16786), .B2(n17274), .A(n16514), .ZN(n16515) );
  OAI21_X1 U18325 ( .B1(n16788), .B2(n17294), .A(n16515), .ZN(P2_U2995) );
  NAND2_X1 U18326 ( .A1(n16519), .A2(n16518), .ZN(n16521) );
  XOR2_X1 U18327 ( .A(n16521), .B(n16520), .Z(n16800) );
  NOR2_X1 U18328 ( .A1(n18600), .A2(n16522), .ZN(n16795) );
  NOR2_X1 U18329 ( .A1(n17301), .A2(n18474), .ZN(n16523) );
  AOI211_X1 U18330 ( .C1(n17286), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16795), .B(n16523), .ZN(n16524) );
  OAI21_X1 U18331 ( .B1(n18479), .B2(n17296), .A(n16524), .ZN(n16525) );
  AOI21_X1 U18332 ( .B1(n16800), .B2(n17274), .A(n16525), .ZN(n16526) );
  OAI21_X1 U18333 ( .B1(n16802), .B2(n17294), .A(n16526), .ZN(P2_U2996) );
  XNOR2_X1 U18334 ( .A(n16527), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16540) );
  AND2_X1 U18335 ( .A1(n16529), .A2(n16528), .ZN(n16545) );
  NAND2_X1 U18336 ( .A1(n16545), .A2(n16544), .ZN(n16546) );
  NAND2_X1 U18337 ( .A1(n16546), .A2(n16530), .ZN(n16534) );
  NAND2_X1 U18338 ( .A1(n16532), .A2(n16531), .ZN(n16533) );
  XNOR2_X1 U18339 ( .A(n16534), .B(n16533), .ZN(n16812) );
  NOR2_X1 U18340 ( .A1(n18600), .A2(n16535), .ZN(n16809) );
  AOI21_X1 U18341 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16809), .ZN(n16537) );
  NAND2_X1 U18342 ( .A1(n17260), .A2(n18463), .ZN(n16536) );
  OAI211_X1 U18343 ( .C1(n18467), .C2(n17296), .A(n16537), .B(n16536), .ZN(
        n16538) );
  AOI21_X1 U18344 ( .B1(n16812), .B2(n17274), .A(n16538), .ZN(n16539) );
  OAI21_X1 U18345 ( .B1(n16540), .B2(n17294), .A(n16539), .ZN(P2_U2997) );
  INV_X1 U18346 ( .A(n16820), .ZN(n16541) );
  OAI211_X1 U18347 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16541), .A(
        n11147), .B(n17270), .ZN(n16550) );
  NAND2_X1 U18348 ( .A1(n18427), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16824) );
  NAND2_X1 U18349 ( .A1(n17286), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16542) );
  OAI211_X1 U18350 ( .C1(n17301), .C2(n16543), .A(n16824), .B(n16542), .ZN(
        n16548) );
  NOR2_X1 U18351 ( .A1(n16545), .A2(n16544), .ZN(n16826) );
  INV_X1 U18352 ( .A(n16546), .ZN(n16825) );
  NOR3_X1 U18353 ( .A1(n16826), .A2(n16825), .A3(n17295), .ZN(n16547) );
  AOI211_X1 U18354 ( .C1(n17273), .C2(n18457), .A(n16548), .B(n16547), .ZN(
        n16549) );
  NAND2_X1 U18355 ( .A1(n16550), .A2(n16549), .ZN(P2_U2998) );
  OAI21_X1 U18356 ( .B1(n16551), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16820), .ZN(n16844) );
  NAND2_X1 U18357 ( .A1(n16553), .A2(n16552), .ZN(n16559) );
  INV_X1 U18358 ( .A(n16554), .ZN(n16581) );
  INV_X1 U18359 ( .A(n16578), .ZN(n16555) );
  OAI21_X1 U18360 ( .B1(n16581), .B2(n16555), .A(n16579), .ZN(n16569) );
  AND2_X1 U18361 ( .A1(n16557), .A2(n16556), .ZN(n16568) );
  NAND2_X1 U18362 ( .A1(n16569), .A2(n16568), .ZN(n16567) );
  NAND2_X1 U18363 ( .A1(n16567), .A2(n16557), .ZN(n16558) );
  XOR2_X1 U18364 ( .A(n16559), .B(n16558), .Z(n16842) );
  NOR2_X1 U18365 ( .A1(n18600), .A2(n18442), .ZN(n16833) );
  NOR2_X1 U18366 ( .A1(n17301), .A2(n16560), .ZN(n16561) );
  AOI211_X1 U18367 ( .C1(n17286), .C2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16833), .B(n16561), .ZN(n16562) );
  OAI21_X1 U18368 ( .B1(n18444), .B2(n17296), .A(n16562), .ZN(n16563) );
  AOI21_X1 U18369 ( .B1(n16842), .B2(n17274), .A(n16563), .ZN(n16564) );
  OAI21_X1 U18370 ( .B1(n16844), .B2(n17294), .A(n16564), .ZN(P2_U2999) );
  INV_X1 U18371 ( .A(n16577), .ZN(n16566) );
  INV_X1 U18372 ( .A(n16551), .ZN(n16565) );
  OAI21_X1 U18373 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16566), .A(
        n16565), .ZN(n16860) );
  OAI21_X1 U18374 ( .B1(n16569), .B2(n16568), .A(n16567), .ZN(n16857) );
  NOR2_X1 U18375 ( .A1(n18600), .A2(n16570), .ZN(n16848) );
  NOR2_X1 U18376 ( .A1(n17301), .A2(n16571), .ZN(n16572) );
  AOI211_X1 U18377 ( .C1(n17286), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16848), .B(n16572), .ZN(n16573) );
  OAI21_X1 U18378 ( .B1(n16851), .B2(n17296), .A(n16573), .ZN(n16574) );
  AOI21_X1 U18379 ( .B1(n16857), .B2(n17274), .A(n16574), .ZN(n16575) );
  OAI21_X1 U18380 ( .B1(n16860), .B2(n17294), .A(n16575), .ZN(P2_U3000) );
  OAI21_X1 U18381 ( .B1(n16576), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16577), .ZN(n16872) );
  NAND2_X1 U18382 ( .A1(n16579), .A2(n16578), .ZN(n16580) );
  XNOR2_X1 U18383 ( .A(n16581), .B(n16580), .ZN(n16869) );
  NAND2_X1 U18384 ( .A1(n18427), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16862) );
  OAI21_X1 U18385 ( .B1(n17268), .B2(n18425), .A(n16862), .ZN(n16582) );
  AOI21_X1 U18386 ( .B1(n17260), .B2(n18429), .A(n16582), .ZN(n16583) );
  OAI21_X1 U18387 ( .B1(n18431), .B2(n17296), .A(n16583), .ZN(n16584) );
  AOI21_X1 U18388 ( .B1(n16869), .B2(n17274), .A(n16584), .ZN(n16585) );
  OAI21_X1 U18389 ( .B1(n16872), .B2(n17294), .A(n16585), .ZN(P2_U3001) );
  NAND2_X1 U18390 ( .A1(n11233), .A2(n16587), .ZN(n16589) );
  XOR2_X1 U18391 ( .A(n16589), .B(n16588), .Z(n16885) );
  INV_X1 U18392 ( .A(n16576), .ZN(n16874) );
  NAND2_X1 U18393 ( .A1(n16596), .A2(n16864), .ZN(n16873) );
  NAND3_X1 U18394 ( .A1(n16874), .A2(n17270), .A3(n16873), .ZN(n16595) );
  NOR2_X1 U18395 ( .A1(n18600), .A2(n16590), .ZN(n16876) );
  AOI21_X1 U18396 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16876), .ZN(n16591) );
  OAI21_X1 U18397 ( .B1(n17301), .B2(n16592), .A(n16591), .ZN(n16593) );
  AOI21_X1 U18398 ( .B1(n16877), .B2(n17273), .A(n16593), .ZN(n16594) );
  OAI211_X1 U18399 ( .C1(n17295), .C2(n16885), .A(n16595), .B(n16594), .ZN(
        P2_U3002) );
  OAI21_X1 U18400 ( .B1(n16606), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16596), .ZN(n16904) );
  NOR2_X1 U18401 ( .A1(n18600), .A2(n16597), .ZN(n16896) );
  AOI21_X1 U18402 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16896), .ZN(n16598) );
  OAI21_X1 U18403 ( .B1(n18414), .B2(n17296), .A(n16598), .ZN(n16603) );
  INV_X1 U18404 ( .A(n16475), .ZN(n16599) );
  AOI21_X1 U18405 ( .B1(n16601), .B2(n16600), .A(n16599), .ZN(n16886) );
  NOR2_X1 U18406 ( .A1(n16886), .A2(n17295), .ZN(n16602) );
  AOI211_X1 U18407 ( .C1(n17260), .C2(n16604), .A(n16603), .B(n16602), .ZN(
        n16605) );
  OAI21_X1 U18408 ( .B1(n16904), .B2(n17294), .A(n16605), .ZN(P2_U3003) );
  INV_X1 U18409 ( .A(n16606), .ZN(n16607) );
  OAI21_X1 U18410 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16627), .A(
        n16607), .ZN(n16916) );
  NAND2_X1 U18411 ( .A1(n16608), .A2(n16635), .ZN(n17290) );
  INV_X1 U18412 ( .A(n16609), .ZN(n17288) );
  INV_X1 U18413 ( .A(n17287), .ZN(n16610) );
  AOI21_X1 U18414 ( .B1(n17290), .B2(n17288), .A(n16610), .ZN(n16624) );
  NAND2_X1 U18415 ( .A1(n16624), .A2(n16622), .ZN(n16626) );
  NAND2_X1 U18416 ( .A1(n16626), .A2(n16621), .ZN(n16614) );
  NAND2_X1 U18417 ( .A1(n16612), .A2(n16611), .ZN(n16613) );
  XNOR2_X1 U18418 ( .A(n16614), .B(n16613), .ZN(n16914) );
  NOR2_X1 U18419 ( .A1(n18600), .A2(n16615), .ZN(n16907) );
  NOR2_X1 U18420 ( .A1(n16911), .A2(n17296), .ZN(n16616) );
  AOI211_X1 U18421 ( .C1(n17286), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16907), .B(n16616), .ZN(n16617) );
  OAI21_X1 U18422 ( .B1(n17301), .B2(n16618), .A(n16617), .ZN(n16619) );
  AOI21_X1 U18423 ( .B1(n16914), .B2(n17274), .A(n16619), .ZN(n16620) );
  OAI21_X1 U18424 ( .B1(n16916), .B2(n17294), .A(n16620), .ZN(P2_U3004) );
  INV_X1 U18425 ( .A(n16621), .ZN(n16625) );
  AND2_X1 U18426 ( .A1(n16622), .A2(n16621), .ZN(n16623) );
  OAI22_X1 U18427 ( .A1(n16626), .A2(n16625), .B1(n16624), .B2(n16623), .ZN(
        n16927) );
  INV_X1 U18428 ( .A(n16628), .ZN(n16629) );
  NAND2_X1 U18429 ( .A1(n16629), .A2(n16888), .ZN(n16917) );
  NAND3_X1 U18430 ( .A1(n11291), .A2(n17270), .A3(n16917), .ZN(n16633) );
  INV_X1 U18431 ( .A(n16920), .ZN(n18404) );
  NOR2_X1 U18432 ( .A1(n18600), .A2(n18402), .ZN(n16919) );
  AOI21_X1 U18433 ( .B1(n17286), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16919), .ZN(n16630) );
  OAI21_X1 U18434 ( .B1(n18404), .B2(n17296), .A(n16630), .ZN(n16631) );
  AOI21_X1 U18435 ( .B1(n17260), .B2(n18397), .A(n16631), .ZN(n16632) );
  OAI211_X1 U18436 ( .C1(n17295), .C2(n16927), .A(n16633), .B(n16632), .ZN(
        P2_U3005) );
  NAND2_X1 U18437 ( .A1(n16635), .A2(n16634), .ZN(n16636) );
  XNOR2_X1 U18438 ( .A(n16637), .B(n16636), .ZN(n16941) );
  OR2_X1 U18439 ( .A1(n16639), .A2(n16638), .ZN(n16928) );
  NAND3_X1 U18440 ( .A1(n16928), .A2(n17270), .A3(n16640), .ZN(n16645) );
  NOR2_X1 U18441 ( .A1(n17296), .A2(n18391), .ZN(n16643) );
  OAI22_X1 U18442 ( .A1(n16641), .A2(n17268), .B1(n13095), .B2(n18488), .ZN(
        n16642) );
  AOI211_X1 U18443 ( .C1(n17260), .C2(n18386), .A(n16643), .B(n16642), .ZN(
        n16644) );
  OAI211_X1 U18444 ( .C1(n16941), .C2(n17295), .A(n16645), .B(n16644), .ZN(
        P2_U3007) );
  NAND2_X1 U18445 ( .A1(n16646), .A2(n18625), .ZN(n16652) );
  NOR2_X1 U18446 ( .A1(n16647), .A2(n18603), .ZN(n16648) );
  OAI211_X1 U18447 ( .C1(n16654), .C2(n16653), .A(n16652), .B(n16651), .ZN(
        n16655) );
  AOI21_X1 U18448 ( .B1(n16656), .B2(n18623), .A(n16655), .ZN(n16657) );
  OAI21_X1 U18449 ( .B1(n16658), .B2(n18614), .A(n16657), .ZN(P2_U3018) );
  INV_X1 U18450 ( .A(n16680), .ZN(n16667) );
  INV_X1 U18451 ( .A(n16659), .ZN(n16664) );
  INV_X1 U18452 ( .A(n16660), .ZN(n16661) );
  NOR3_X1 U18453 ( .A1(n16691), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16661), .ZN(n16662) );
  AOI211_X1 U18454 ( .C1(n16664), .C2(n18628), .A(n16663), .B(n16662), .ZN(
        n16665) );
  OAI21_X1 U18455 ( .B1(n16667), .B2(n16666), .A(n16665), .ZN(n16670) );
  NOR2_X1 U18456 ( .A1(n16668), .A2(n18608), .ZN(n16669) );
  AOI211_X1 U18457 ( .C1(n16671), .C2(n18625), .A(n16670), .B(n16669), .ZN(
        n16672) );
  OAI21_X1 U18458 ( .B1(n16673), .B2(n18614), .A(n16672), .ZN(P2_U3019) );
  OAI21_X1 U18459 ( .B1(n16691), .B2(n16675), .A(n16674), .ZN(n16679) );
  OAI21_X1 U18460 ( .B1(n16677), .B2(n18603), .A(n16676), .ZN(n16678) );
  AOI21_X1 U18461 ( .B1(n16680), .B2(n16679), .A(n16678), .ZN(n16681) );
  OAI21_X1 U18462 ( .B1(n16682), .B2(n18607), .A(n16681), .ZN(n16683) );
  AOI21_X1 U18463 ( .B1(n16684), .B2(n18623), .A(n16683), .ZN(n16685) );
  OAI21_X1 U18464 ( .B1(n16686), .B2(n18614), .A(n16685), .ZN(P2_U3020) );
  OAI21_X1 U18465 ( .B1(n18555), .B2(n18603), .A(n16687), .ZN(n16688) );
  AOI21_X1 U18466 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16689), .A(
        n16688), .ZN(n16690) );
  OAI21_X1 U18467 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16691), .A(
        n16690), .ZN(n16694) );
  NOR2_X1 U18468 ( .A1(n16692), .A2(n18614), .ZN(n16693) );
  AOI211_X1 U18469 ( .C1(n18552), .C2(n18625), .A(n16694), .B(n16693), .ZN(
        n16695) );
  NOR2_X1 U18470 ( .A1(n16697), .A2(n18607), .ZN(n16705) );
  INV_X1 U18471 ( .A(n16715), .ZN(n16734) );
  AOI21_X1 U18472 ( .B1(n16734), .B2(n16698), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16703) );
  NAND2_X1 U18473 ( .A1(n16699), .A2(n18628), .ZN(n16701) );
  OAI211_X1 U18474 ( .C1(n16703), .C2(n16702), .A(n16701), .B(n16700), .ZN(
        n16704) );
  AOI211_X1 U18475 ( .C1(n16706), .C2(n18627), .A(n16705), .B(n16704), .ZN(
        n16707) );
  OAI21_X1 U18476 ( .B1(n18608), .B2(n16708), .A(n16707), .ZN(P2_U3022) );
  XNOR2_X1 U18477 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16714) );
  OAI21_X1 U18478 ( .B1(n16729), .B2(n16710), .A(n16709), .ZN(n16711) );
  AOI21_X1 U18479 ( .B1(n16712), .B2(n18628), .A(n16711), .ZN(n16713) );
  OAI21_X1 U18480 ( .B1(n16715), .B2(n16714), .A(n16713), .ZN(n16718) );
  NOR2_X1 U18481 ( .A1(n16716), .A2(n18614), .ZN(n16717) );
  AOI211_X1 U18482 ( .C1(n16719), .C2(n18625), .A(n16718), .B(n16717), .ZN(
        n16720) );
  OAI21_X1 U18483 ( .B1(n18608), .B2(n16721), .A(n16720), .ZN(P2_U3023) );
  NAND2_X1 U18484 ( .A1(n16722), .A2(n18623), .ZN(n16736) );
  INV_X1 U18485 ( .A(n16723), .ZN(n16724) );
  AOI21_X1 U18486 ( .B1(n16726), .B2(n16725), .A(n16724), .ZN(n19299) );
  NAND2_X1 U18487 ( .A1(n19299), .A2(n18628), .ZN(n16728) );
  OAI211_X1 U18488 ( .C1(n16729), .C2(n16733), .A(n16728), .B(n16727), .ZN(
        n16732) );
  NOR2_X1 U18489 ( .A1(n16730), .A2(n18607), .ZN(n16731) );
  AOI211_X1 U18490 ( .C1(n16734), .C2(n16733), .A(n16732), .B(n16731), .ZN(
        n16735) );
  OAI211_X1 U18491 ( .C1(n16737), .C2(n18614), .A(n16736), .B(n16735), .ZN(
        P2_U3024) );
  INV_X1 U18492 ( .A(n18527), .ZN(n16741) );
  INV_X1 U18493 ( .A(n16738), .ZN(n16762) );
  NOR3_X1 U18494 ( .A1(n16762), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16763), .ZN(n16739) );
  AOI211_X1 U18495 ( .C1(n18628), .C2(n16741), .A(n16740), .B(n16739), .ZN(
        n16744) );
  NAND3_X1 U18496 ( .A1(n16742), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16887), .ZN(n16743) );
  OAI211_X1 U18497 ( .C1(n18512), .C2(n18607), .A(n16744), .B(n16743), .ZN(
        n16745) );
  AOI21_X1 U18498 ( .B1(n16746), .B2(n18623), .A(n16745), .ZN(n16747) );
  OAI21_X1 U18499 ( .B1(n16748), .B2(n18614), .A(n16747), .ZN(P2_U3025) );
  INV_X1 U18500 ( .A(n16813), .ZN(n16837) );
  NAND2_X1 U18501 ( .A1(n16837), .A2(n16754), .ZN(n16759) );
  NOR2_X1 U18502 ( .A1(n16759), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16789) );
  NOR2_X1 U18503 ( .A1(n18615), .A2(n16803), .ZN(n16749) );
  OR2_X1 U18504 ( .A1(n16750), .A2(n16749), .ZN(n16805) );
  INV_X1 U18505 ( .A(n16805), .ZN(n16758) );
  NOR2_X1 U18506 ( .A1(n16752), .A2(n16751), .ZN(n16753) );
  AOI22_X1 U18507 ( .A1(n16755), .A2(n16754), .B1(n16753), .B2(n16804), .ZN(
        n16756) );
  NAND2_X1 U18508 ( .A1(n16930), .A2(n16756), .ZN(n16757) );
  NAND2_X1 U18509 ( .A1(n16758), .A2(n16757), .ZN(n16796) );
  NOR2_X1 U18510 ( .A1(n16789), .A2(n16796), .ZN(n16784) );
  INV_X1 U18511 ( .A(n16759), .ZN(n16761) );
  NAND2_X1 U18512 ( .A1(n16761), .A2(n16760), .ZN(n16764) );
  AOI22_X1 U18513 ( .A1(n16784), .A2(n16764), .B1(n16763), .B2(n16762), .ZN(
        n16773) );
  NOR2_X1 U18514 ( .A1(n16766), .A2(n16765), .ZN(n16767) );
  OR2_X1 U18515 ( .A1(n16768), .A2(n16767), .ZN(n19394) );
  NAND2_X1 U18516 ( .A1(n16769), .A2(n18625), .ZN(n16771) );
  OAI211_X1 U18517 ( .C1(n18603), .C2(n19394), .A(n16771), .B(n16770), .ZN(
        n16772) );
  AOI211_X1 U18518 ( .C1(n16774), .C2(n18627), .A(n16773), .B(n16772), .ZN(
        n16775) );
  OAI21_X1 U18519 ( .B1(n16776), .B2(n18608), .A(n16775), .ZN(P2_U3026) );
  NAND3_X1 U18520 ( .A1(n16837), .A2(n16783), .A3(n16777), .ZN(n16779) );
  OAI211_X1 U18521 ( .C1(n18603), .C2(n18492), .A(n16779), .B(n16778), .ZN(
        n16780) );
  AOI21_X1 U18522 ( .B1(n16781), .B2(n18625), .A(n16780), .ZN(n16782) );
  OAI21_X1 U18523 ( .B1(n16784), .B2(n16783), .A(n16782), .ZN(n16785) );
  AOI21_X1 U18524 ( .B1(n16786), .B2(n18627), .A(n16785), .ZN(n16787) );
  OAI21_X1 U18525 ( .B1(n16788), .B2(n18608), .A(n16787), .ZN(P2_U3027) );
  INV_X1 U18526 ( .A(n16789), .ZN(n16798) );
  NAND2_X1 U18527 ( .A1(n16791), .A2(n16790), .ZN(n16792) );
  NAND2_X1 U18528 ( .A1(n16793), .A2(n16792), .ZN(n19481) );
  NOR2_X1 U18529 ( .A1(n18603), .A2(n19481), .ZN(n16794) );
  AOI211_X1 U18530 ( .C1(n16796), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16795), .B(n16794), .ZN(n16797) );
  OAI211_X1 U18531 ( .C1(n18479), .C2(n18607), .A(n16798), .B(n16797), .ZN(
        n16799) );
  AOI21_X1 U18532 ( .B1(n16800), .B2(n18627), .A(n16799), .ZN(n16801) );
  NAND2_X1 U18533 ( .A1(n18615), .A2(n18608), .ZN(n16819) );
  NAND3_X1 U18534 ( .A1(n16804), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16803), .ZN(n16806) );
  AOI21_X1 U18535 ( .B1(n16807), .B2(n16806), .A(n16805), .ZN(n16840) );
  OAI21_X1 U18536 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18593), .A(
        n16840), .ZN(n16808) );
  AOI21_X1 U18537 ( .B1(n11147), .B2(n16819), .A(n16808), .ZN(n16817) );
  AOI21_X1 U18538 ( .B1(n18628), .B2(n18468), .A(n16809), .ZN(n16810) );
  OAI21_X1 U18539 ( .B1(n18467), .B2(n18607), .A(n16810), .ZN(n16811) );
  AOI21_X1 U18540 ( .B1(n16812), .B2(n18627), .A(n16811), .ZN(n16815) );
  OAI22_X1 U18541 ( .A1(n16820), .A2(n18608), .B1(n16839), .B2(n16813), .ZN(
        n16821) );
  NAND3_X1 U18542 ( .A1(n16821), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16816), .ZN(n16814) );
  OAI211_X1 U18543 ( .C1(n16817), .C2(n16816), .A(n16815), .B(n16814), .ZN(
        P2_U3029) );
  INV_X1 U18544 ( .A(n16840), .ZN(n16818) );
  AOI21_X1 U18545 ( .B1(n16820), .B2(n16819), .A(n16818), .ZN(n16832) );
  NAND2_X1 U18546 ( .A1(n16821), .A2(n16831), .ZN(n16830) );
  NOR2_X1 U18547 ( .A1(n11062), .A2(n16822), .ZN(n16823) );
  OR2_X1 U18548 ( .A1(n16380), .A2(n16823), .ZN(n18456) );
  OAI21_X1 U18549 ( .B1(n18603), .B2(n18456), .A(n16824), .ZN(n16828) );
  NOR3_X1 U18550 ( .A1(n16826), .A2(n16825), .A3(n18614), .ZN(n16827) );
  AOI211_X1 U18551 ( .C1(n18625), .C2(n18457), .A(n16828), .B(n16827), .ZN(
        n16829) );
  OAI211_X1 U18552 ( .C1(n16832), .C2(n16831), .A(n16830), .B(n16829), .ZN(
        P2_U3030) );
  AOI21_X1 U18553 ( .B1(n18628), .B2(n16834), .A(n16833), .ZN(n16835) );
  OAI21_X1 U18554 ( .B1(n18444), .B2(n18607), .A(n16835), .ZN(n16836) );
  AOI21_X1 U18555 ( .B1(n16837), .B2(n16839), .A(n16836), .ZN(n16838) );
  OAI21_X1 U18556 ( .B1(n16840), .B2(n16839), .A(n16838), .ZN(n16841) );
  AOI21_X1 U18557 ( .B1(n16842), .B2(n18627), .A(n16841), .ZN(n16843) );
  OAI21_X1 U18558 ( .B1(n16844), .B2(n18608), .A(n16843), .ZN(P2_U3031) );
  NAND2_X1 U18559 ( .A1(n16890), .A2(n16845), .ZN(n16865) );
  INV_X1 U18560 ( .A(n16865), .ZN(n16846) );
  NAND2_X1 U18561 ( .A1(n16846), .A2(n16864), .ZN(n16879) );
  AOI21_X1 U18562 ( .B1(n16847), .B2(n16930), .A(n16924), .ZN(n16875) );
  NAND2_X1 U18563 ( .A1(n16879), .A2(n16875), .ZN(n16868) );
  AOI21_X1 U18564 ( .B1(n18628), .B2(n16849), .A(n16848), .ZN(n16850) );
  OAI21_X1 U18565 ( .B1(n16851), .B2(n18607), .A(n16850), .ZN(n16856) );
  AOI21_X1 U18566 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16854), .A(
        n16853), .ZN(n16852) );
  AOI211_X1 U18567 ( .C1(n16854), .C2(n16853), .A(n16852), .B(n16865), .ZN(
        n16855) );
  AOI211_X1 U18568 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16868), .A(
        n16856), .B(n16855), .ZN(n16859) );
  NAND2_X1 U18569 ( .A1(n16857), .A2(n18627), .ZN(n16858) );
  OAI211_X1 U18570 ( .C1(n16860), .C2(n18608), .A(n16859), .B(n16858), .ZN(
        P2_U3032) );
  INV_X1 U18571 ( .A(n18436), .ZN(n16861) );
  NAND2_X1 U18572 ( .A1(n18628), .A2(n16861), .ZN(n16863) );
  OAI211_X1 U18573 ( .C1(n18431), .C2(n18607), .A(n16863), .B(n16862), .ZN(
        n16867) );
  NOR3_X1 U18574 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n16864), .ZN(n16866) );
  AOI211_X1 U18575 ( .C1(n16868), .C2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16867), .B(n16866), .ZN(n16871) );
  NAND2_X1 U18576 ( .A1(n16869), .A2(n18627), .ZN(n16870) );
  OAI211_X1 U18577 ( .C1(n16872), .C2(n18608), .A(n16871), .B(n16870), .ZN(
        P2_U3033) );
  NAND3_X1 U18578 ( .A1(n16874), .A2(n18623), .A3(n16873), .ZN(n16884) );
  INV_X1 U18579 ( .A(n16875), .ZN(n16882) );
  AOI21_X1 U18580 ( .B1(n16877), .B2(n18625), .A(n16876), .ZN(n16878) );
  OAI211_X1 U18581 ( .C1(n18603), .C2(n16880), .A(n16879), .B(n16878), .ZN(
        n16881) );
  AOI21_X1 U18582 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16882), .A(
        n16881), .ZN(n16883) );
  OAI211_X1 U18583 ( .C1(n16885), .C2(n18614), .A(n16884), .B(n16883), .ZN(
        P2_U3034) );
  INV_X1 U18584 ( .A(n16886), .ZN(n16902) );
  OAI21_X1 U18585 ( .B1(n16924), .B2(n16888), .A(n16887), .ZN(n16906) );
  NOR2_X1 U18586 ( .A1(n16888), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16889) );
  NAND2_X1 U18587 ( .A1(n16890), .A2(n16889), .ZN(n16910) );
  AOI21_X1 U18588 ( .B1(n16906), .B2(n16910), .A(n16891), .ZN(n16901) );
  INV_X1 U18589 ( .A(n16890), .ZN(n16922) );
  NAND3_X1 U18590 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16891), .ZN(n16899) );
  INV_X1 U18591 ( .A(n18414), .ZN(n16897) );
  AND2_X1 U18592 ( .A1(n11070), .A2(n16892), .ZN(n16894) );
  OR2_X1 U18593 ( .A1(n16894), .A2(n16893), .ZN(n19115) );
  NOR2_X1 U18594 ( .A1(n18603), .A2(n19115), .ZN(n16895) );
  AOI211_X1 U18595 ( .C1(n16897), .C2(n18625), .A(n16896), .B(n16895), .ZN(
        n16898) );
  OAI21_X1 U18596 ( .B1(n16922), .B2(n16899), .A(n16898), .ZN(n16900) );
  AOI211_X1 U18597 ( .C1(n16902), .C2(n18627), .A(n16901), .B(n16900), .ZN(
        n16903) );
  OAI21_X1 U18598 ( .B1(n16904), .B2(n18608), .A(n16903), .ZN(P2_U3035) );
  NOR2_X1 U18599 ( .A1(n16906), .A2(n16905), .ZN(n16913) );
  AOI21_X1 U18600 ( .B1(n18628), .B2(n16908), .A(n16907), .ZN(n16909) );
  OAI211_X1 U18601 ( .C1(n18607), .C2(n16911), .A(n16910), .B(n16909), .ZN(
        n16912) );
  AOI211_X1 U18602 ( .C1(n16914), .C2(n18627), .A(n16913), .B(n16912), .ZN(
        n16915) );
  OAI21_X1 U18603 ( .B1(n16916), .B2(n18608), .A(n16915), .ZN(P2_U3036) );
  NAND3_X1 U18604 ( .A1(n11291), .A2(n18623), .A3(n16917), .ZN(n16926) );
  NOR2_X1 U18605 ( .A1(n18603), .A2(n18403), .ZN(n16918) );
  AOI211_X1 U18606 ( .C1(n16920), .C2(n18625), .A(n16919), .B(n16918), .ZN(
        n16921) );
  OAI21_X1 U18607 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16922), .A(
        n16921), .ZN(n16923) );
  AOI21_X1 U18608 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16924), .A(
        n16923), .ZN(n16925) );
  OAI211_X1 U18609 ( .C1(n16927), .C2(n18614), .A(n16926), .B(n16925), .ZN(
        P2_U3037) );
  NAND3_X1 U18610 ( .A1(n16928), .A2(n18623), .A3(n16640), .ZN(n16940) );
  NOR2_X1 U18611 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16931), .ZN(
        n16938) );
  AOI21_X1 U18612 ( .B1(n16931), .B2(n16930), .A(n16929), .ZN(n18599) );
  NOR2_X1 U18613 ( .A1(n13095), .A2(n18488), .ZN(n16933) );
  NOR2_X1 U18614 ( .A1(n18607), .A2(n18391), .ZN(n16932) );
  AOI211_X1 U18615 ( .C1(n16934), .C2(n18628), .A(n16933), .B(n16932), .ZN(
        n16935) );
  OAI21_X1 U18616 ( .B1(n18599), .B2(n18595), .A(n16935), .ZN(n16936) );
  AOI21_X1 U18617 ( .B1(n16938), .B2(n16937), .A(n16936), .ZN(n16939) );
  OAI211_X1 U18618 ( .C1(n16941), .C2(n18614), .A(n16940), .B(n16939), .ZN(
        P2_U3039) );
  XNOR2_X1 U18619 ( .A(n16943), .B(n16942), .ZN(n17281) );
  NOR2_X1 U18620 ( .A1(n16944), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17279) );
  INV_X1 U18621 ( .A(n17279), .ZN(n16946) );
  NAND3_X1 U18622 ( .A1(n16946), .A2(n18623), .A3(n16945), .ZN(n16955) );
  INV_X1 U18623 ( .A(n16947), .ZN(n16949) );
  NOR2_X1 U18624 ( .A1(n16949), .A2(n16948), .ZN(n18594) );
  INV_X1 U18625 ( .A(n17280), .ZN(n18380) );
  NOR2_X1 U18626 ( .A1(n18372), .A2(n18488), .ZN(n16951) );
  NOR2_X1 U18627 ( .A1(n18603), .A2(n18384), .ZN(n16950) );
  AOI211_X1 U18628 ( .C1(n18380), .C2(n18625), .A(n16951), .B(n16950), .ZN(
        n16952) );
  OAI21_X1 U18629 ( .B1(n18599), .B2(n18597), .A(n16952), .ZN(n16953) );
  AOI21_X1 U18630 ( .B1(n18594), .B2(n18597), .A(n16953), .ZN(n16954) );
  OAI211_X1 U18631 ( .C1(n17281), .C2(n18614), .A(n16955), .B(n16954), .ZN(
        P2_U3040) );
  NOR2_X1 U18632 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U18633 ( .A1(n18535), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18348), .B2(n10997), .ZN(n16963) );
  AOI222_X1 U18634 ( .A1(n16956), .A2(n16969), .B1(n19195), .B2(n18653), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n16963), .ZN(n16961) );
  OAI22_X1 U18635 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19262), .B1(n16957), 
        .B2(n18661), .ZN(n16958) );
  NAND2_X1 U18636 ( .A1(n18579), .A2(n16959), .ZN(n16960) );
  OAI21_X1 U18637 ( .B1(n16961), .B2(n18579), .A(n16960), .ZN(P2_U3601) );
  INV_X1 U18638 ( .A(n18653), .ZN(n16975) );
  NOR2_X1 U18639 ( .A1(n16963), .A2(n16962), .ZN(n16968) );
  AOI21_X1 U18640 ( .B1(n18535), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n16964), .ZN(n16971) );
  AOI22_X1 U18641 ( .A1(n16965), .A2(n16969), .B1(n16968), .B2(n16971), .ZN(
        n16966) );
  OAI21_X1 U18642 ( .B1(n17320), .B2(n16975), .A(n16966), .ZN(n16967) );
  MUX2_X1 U18643 ( .A(n16967), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n18579), .Z(P2_U3600) );
  INV_X1 U18644 ( .A(n16968), .ZN(n16972) );
  INV_X1 U18645 ( .A(n16969), .ZN(n18638) );
  OAI222_X1 U18646 ( .A1(n16975), .A2(n17309), .B1(n16972), .B2(n16971), .C1(
        n18638), .C2(n16970), .ZN(n16973) );
  MUX2_X1 U18647 ( .A(n16973), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n18579), .Z(P2_U3599) );
  OAI22_X1 U18648 ( .A1(n19162), .A2(n16975), .B1(n16974), .B2(n18638), .ZN(
        n16976) );
  MUX2_X1 U18649 ( .A(n16976), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n18579), .Z(P2_U3596) );
  NAND2_X1 U18650 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18712) );
  NOR2_X1 U18651 ( .A1(n20685), .A2(n21574), .ZN(n17849) );
  NOR2_X1 U18652 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17662), .ZN(n20004) );
  INV_X1 U18653 ( .A(n20004), .ZN(n17666) );
  NOR2_X1 U18654 ( .A1(n17849), .A2(n17666), .ZN(n16979) );
  INV_X1 U18655 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21166) );
  NAND2_X1 U18656 ( .A1(n21166), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18709) );
  NOR2_X1 U18657 ( .A1(n16977), .A2(n17735), .ZN(n17663) );
  NOR2_X1 U18658 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21210) );
  NAND2_X1 U18659 ( .A1(n20100), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20710) );
  OAI21_X1 U18660 ( .B1(n21210), .B2(n17662), .A(n20710), .ZN(n18693) );
  OAI211_X1 U18661 ( .C1(n17663), .C2(n21206), .A(n19011), .B(n16978), .ZN(
        n18231) );
  NAND2_X1 U18662 ( .A1(n18709), .A2(n18231), .ZN(n18232) );
  AOI221_X1 U18663 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18712), .C1(n16979), 
        .C2(n18712), .A(n18232), .ZN(n18229) );
  NAND3_X1 U18664 ( .A1(n21075), .A2(n21208), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18714) );
  INV_X1 U18665 ( .A(n18714), .ZN(n18732) );
  INV_X1 U18666 ( .A(n16979), .ZN(n16980) );
  OAI21_X1 U18667 ( .B1(n21166), .B2(n21208), .A(n16980), .ZN(n18230) );
  OAI221_X1 U18668 ( .B1(n18732), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18732), .C2(n18230), .A(n18231), .ZN(n18227) );
  AOI22_X1 U18669 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18229), .B1(
        n18227), .B2(n21174), .ZN(P3_U2865) );
  OR4_X1 U18670 ( .A1(n16982), .A2(n16981), .A3(n12382), .A4(n17039), .ZN(
        n16983) );
  OAI21_X1 U18671 ( .B1(n16984), .B2(n14443), .A(n16983), .ZN(P1_U3468) );
  INV_X1 U18672 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16985) );
  OAI21_X1 U18673 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21625), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18305) );
  NAND2_X1 U18674 ( .A1(n18326), .A2(n18305), .ZN(n16987) );
  INV_X1 U18675 ( .A(n21577), .ZN(n16986) );
  INV_X1 U18676 ( .A(BS16), .ZN(n17114) );
  NAND2_X1 U18677 ( .A1(n21622), .A2(n21625), .ZN(n21578) );
  AOI21_X1 U18678 ( .B1(n17114), .B2(n21578), .A(n16986), .ZN(n21573) );
  AOI21_X1 U18679 ( .B1(n16985), .B2(n16986), .A(n21573), .ZN(P3_U3280) );
  AND2_X1 U18680 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n16986), .ZN(P3_U3028) );
  AND2_X1 U18681 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n16986), .ZN(P3_U3027) );
  AND2_X1 U18682 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n16986), .ZN(P3_U3026) );
  AND2_X1 U18683 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n16986), .ZN(P3_U3025) );
  AND2_X1 U18684 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n16986), .ZN(P3_U3024) );
  AND2_X1 U18685 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n16986), .ZN(P3_U3023) );
  AND2_X1 U18686 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n16986), .ZN(P3_U3022) );
  AND2_X1 U18687 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n16986), .ZN(P3_U3021) );
  AND2_X1 U18688 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n16986), .ZN(
        P3_U3020) );
  AND2_X1 U18689 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n16986), .ZN(
        P3_U3019) );
  AND2_X1 U18690 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n16986), .ZN(
        P3_U3018) );
  AND2_X1 U18691 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n16986), .ZN(
        P3_U3017) );
  AND2_X1 U18692 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n16986), .ZN(
        P3_U3016) );
  AND2_X1 U18693 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n16987), .ZN(
        P3_U3015) );
  AND2_X1 U18694 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n16987), .ZN(
        P3_U3014) );
  AND2_X1 U18695 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n16987), .ZN(
        P3_U3013) );
  AND2_X1 U18696 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n16987), .ZN(
        P3_U3012) );
  AND2_X1 U18697 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n16987), .ZN(
        P3_U3011) );
  AND2_X1 U18698 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n16987), .ZN(
        P3_U3010) );
  AND2_X1 U18699 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n16987), .ZN(
        P3_U3009) );
  AND2_X1 U18700 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n16987), .ZN(
        P3_U3008) );
  AND2_X1 U18701 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n16987), .ZN(
        P3_U3007) );
  AND2_X1 U18702 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n16987), .ZN(
        P3_U3006) );
  AND2_X1 U18703 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n16987), .ZN(
        P3_U3005) );
  AND2_X1 U18704 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n16987), .ZN(
        P3_U3004) );
  AND2_X1 U18705 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n16987), .ZN(
        P3_U3003) );
  AND2_X1 U18706 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n16987), .ZN(
        P3_U3002) );
  AND2_X1 U18707 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n16986), .ZN(
        P3_U3001) );
  AND2_X1 U18708 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n16986), .ZN(
        P3_U3000) );
  AND2_X1 U18709 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n16987), .ZN(
        P3_U2999) );
  INV_X1 U18710 ( .A(n17849), .ZN(n18180) );
  AOI21_X1 U18711 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16989)
         );
  NOR4_X1 U18712 ( .A1(n20685), .A2(n20057), .A3(n21198), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21157) );
  AOI211_X1 U18713 ( .C1(n18180), .C2(n16989), .A(n16988), .B(n21157), .ZN(
        P3_U2998) );
  NOR2_X1 U18714 ( .A1(n21176), .A2(n18231), .ZN(P3_U2867) );
  NAND2_X1 U18715 ( .A1(n20057), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18222) );
  INV_X1 U18716 ( .A(n18222), .ZN(n17973) );
  NAND2_X1 U18717 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17973), .ZN(n20002) );
  INV_X2 U18718 ( .A(n20002), .ZN(n18302) );
  NOR2_X4 U18719 ( .A1(n18302), .A2(n18279), .ZN(n18293) );
  AND2_X1 U18720 ( .A1(n18293), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U18721 ( .A1(n21210), .A2(n21208), .ZN(n17824) );
  NAND2_X1 U18722 ( .A1(n17824), .A2(n20059), .ZN(n16994) );
  XOR2_X1 U18723 ( .A(n20738), .B(n20055), .Z(n20006) );
  OAI22_X1 U18724 ( .A1(P3_READREQUEST_REG_SCAN_IN), .A2(n16994), .B1(n20006), 
        .B2(n20059), .ZN(n16993) );
  INV_X1 U18725 ( .A(n16993), .ZN(P3_U3298) );
  NOR2_X1 U18726 ( .A1(n20495), .A2(n20059), .ZN(n20088) );
  NOR2_X1 U18727 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n16994), .ZN(n16995)
         );
  NOR2_X1 U18728 ( .A1(n20088), .A2(n16995), .ZN(P3_U3299) );
  NOR2_X1 U18729 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n16997), .ZN(n21601) );
  AOI21_X1 U18730 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21601), .A(n16996), 
        .ZN(n16998) );
  INV_X1 U18731 ( .A(n16998), .ZN(n21572) );
  INV_X1 U18732 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17014) );
  NAND2_X1 U18733 ( .A1(n21612), .A2(n16997), .ZN(n21596) );
  AOI21_X1 U18734 ( .B1(n17114), .B2(n21596), .A(n16999), .ZN(n21568) );
  AOI21_X1 U18735 ( .B1(n16999), .B2(n17014), .A(n21568), .ZN(P2_U3591) );
  AND2_X1 U18736 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n16999), .ZN(P2_U3208) );
  AND2_X1 U18737 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n16999), .ZN(P2_U3207) );
  AND2_X1 U18738 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n16999), .ZN(P2_U3206) );
  AND2_X1 U18739 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n16999), .ZN(P2_U3205) );
  AND2_X1 U18740 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n16999), .ZN(P2_U3204) );
  AND2_X1 U18741 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n16999), .ZN(P2_U3203) );
  AND2_X1 U18742 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n16999), .ZN(P2_U3202) );
  AND2_X1 U18743 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n16999), .ZN(P2_U3201) );
  AND2_X1 U18744 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n16999), .ZN(
        P2_U3200) );
  AND2_X1 U18745 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n16999), .ZN(
        P2_U3199) );
  AND2_X1 U18746 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n16999), .ZN(
        P2_U3198) );
  AND2_X1 U18747 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n16999), .ZN(
        P2_U3197) );
  AND2_X1 U18748 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n16999), .ZN(
        P2_U3196) );
  AND2_X1 U18749 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n16999), .ZN(
        P2_U3195) );
  AND2_X1 U18750 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n16998), .ZN(
        P2_U3194) );
  AND2_X1 U18751 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n16998), .ZN(
        P2_U3193) );
  AND2_X1 U18752 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n16998), .ZN(
        P2_U3192) );
  AND2_X1 U18753 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n16998), .ZN(
        P2_U3191) );
  AND2_X1 U18754 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n16998), .ZN(
        P2_U3190) );
  AND2_X1 U18755 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n16998), .ZN(
        P2_U3189) );
  AND2_X1 U18756 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n16998), .ZN(
        P2_U3188) );
  AND2_X1 U18757 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n16998), .ZN(
        P2_U3187) );
  AND2_X1 U18758 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n16998), .ZN(
        P2_U3186) );
  AND2_X1 U18759 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n16998), .ZN(
        P2_U3185) );
  AND2_X1 U18760 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n16998), .ZN(
        P2_U3184) );
  AND2_X1 U18761 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n16998), .ZN(
        P2_U3183) );
  AND2_X1 U18762 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n16999), .ZN(
        P2_U3182) );
  AND2_X1 U18763 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n16999), .ZN(
        P2_U3181) );
  AND2_X1 U18764 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n16999), .ZN(
        P2_U3180) );
  AND2_X1 U18765 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n16999), .ZN(
        P2_U3179) );
  NAND2_X1 U18766 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18655), .ZN(n18639) );
  AOI21_X1 U18767 ( .B1(n17000), .B2(n18340), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17002) );
  AOI221_X1 U18768 ( .B1(n18639), .B2(n17002), .C1(n16962), .C2(n17002), .A(
        n17001), .ZN(P2_U3178) );
  INV_X1 U18769 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18665) );
  OAI221_X1 U18770 ( .B1(n18665), .B2(n18647), .C1(n18645), .C2(n18647), .A(
        n19591), .ZN(n17316) );
  NOR2_X1 U18771 ( .A1(n17003), .A2(n17316), .ZN(P2_U3047) );
  AND2_X1 U18772 ( .A1(n17357), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18773 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17007) );
  NOR4_X1 U18774 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17006) );
  NOR4_X1 U18775 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17005) );
  NOR4_X1 U18776 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17004) );
  NAND4_X1 U18777 ( .A1(n17007), .A2(n17006), .A3(n17005), .A4(n17004), .ZN(
        n17013) );
  NOR4_X1 U18778 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17011) );
  AOI211_X1 U18779 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17010) );
  NOR4_X1 U18780 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17009) );
  NOR4_X1 U18781 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17008) );
  NAND4_X1 U18782 ( .A1(n17011), .A2(n17010), .A3(n17009), .A4(n17008), .ZN(
        n17012) );
  NOR2_X1 U18783 ( .A1(n17013), .A2(n17012), .ZN(n17333) );
  INV_X1 U18784 ( .A(n17333), .ZN(n17331) );
  NOR2_X1 U18785 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17331), .ZN(n17326) );
  INV_X1 U18786 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21571) );
  NAND3_X1 U18787 ( .A1(n12555), .A2(n21571), .A3(n17014), .ZN(n17330) );
  INV_X1 U18788 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U18789 ( .A1(n17326), .A2(n17330), .B1(n17331), .B2(n17015), .ZN(
        P2_U2821) );
  INV_X1 U18790 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U18791 ( .A1(n17326), .A2(n12555), .B1(n17331), .B2(n17016), .ZN(
        P2_U2820) );
  INV_X1 U18792 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17017) );
  NOR2_X2 U18793 ( .A1(n11627), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22246) );
  AND2_X1 U18794 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21580), .ZN(n17063) );
  NOR2_X1 U18795 ( .A1(n22246), .A2(n17063), .ZN(n21564) );
  OAI221_X1 U18796 ( .B1(n11627), .B2(BS16), .C1(n21585), .C2(BS16), .A(n21564), .ZN(n21563) );
  INV_X1 U18797 ( .A(n21563), .ZN(n21565) );
  AOI21_X1 U18798 ( .B1(n17017), .B2(n21566), .A(n21565), .ZN(P1_U3464) );
  AND2_X1 U18799 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21566), .ZN(P1_U3193) );
  AND2_X1 U18800 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21566), .ZN(P1_U3192) );
  AND2_X1 U18801 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21566), .ZN(P1_U3191) );
  AND2_X1 U18802 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21566), .ZN(P1_U3190) );
  AND2_X1 U18803 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21566), .ZN(P1_U3189) );
  AND2_X1 U18804 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21566), .ZN(P1_U3188) );
  AND2_X1 U18805 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21566), .ZN(P1_U3187) );
  AND2_X1 U18806 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21566), .ZN(P1_U3186) );
  AND2_X1 U18807 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21566), .ZN(
        P1_U3185) );
  AND2_X1 U18808 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21566), .ZN(
        P1_U3184) );
  AND2_X1 U18809 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21566), .ZN(
        P1_U3183) );
  AND2_X1 U18810 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21566), .ZN(
        P1_U3182) );
  AND2_X1 U18811 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21566), .ZN(
        P1_U3181) );
  AND2_X1 U18812 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21566), .ZN(
        P1_U3180) );
  AND2_X1 U18813 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21566), .ZN(
        P1_U3179) );
  AND2_X1 U18814 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21566), .ZN(
        P1_U3178) );
  AND2_X1 U18815 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21566), .ZN(
        P1_U3177) );
  AND2_X1 U18816 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21566), .ZN(
        P1_U3176) );
  AND2_X1 U18817 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21566), .ZN(
        P1_U3175) );
  AND2_X1 U18818 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21566), .ZN(
        P1_U3174) );
  AND2_X1 U18819 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21566), .ZN(
        P1_U3173) );
  AND2_X1 U18820 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21566), .ZN(
        P1_U3172) );
  AND2_X1 U18821 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21566), .ZN(
        P1_U3171) );
  AND2_X1 U18822 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21566), .ZN(
        P1_U3170) );
  AND2_X1 U18823 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21566), .ZN(
        P1_U3169) );
  AND2_X1 U18824 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21566), .ZN(
        P1_U3168) );
  AND2_X1 U18825 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21566), .ZN(
        P1_U3167) );
  AND2_X1 U18826 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21566), .ZN(
        P1_U3166) );
  AND2_X1 U18827 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21566), .ZN(
        P1_U3165) );
  AND2_X1 U18828 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21566), .ZN(
        P1_U3164) );
  MUX2_X1 U18829 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17018), .S(
        n17044), .Z(n17048) );
  MUX2_X1 U18830 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17019), .S(
        n17044), .Z(n17047) );
  MUX2_X1 U18831 ( .A(n17021), .B(n17020), .S(n11541), .Z(n17022) );
  NOR2_X1 U18832 ( .A1(n17022), .A2(n21810), .ZN(n17023) );
  AND2_X1 U18833 ( .A1(n17024), .A2(n17023), .ZN(n17028) );
  AOI21_X1 U18834 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17028), .A(
        n17025), .ZN(n17026) );
  NAND2_X1 U18835 ( .A1(n17026), .A2(n17044), .ZN(n17027) );
  OAI21_X1 U18836 ( .B1(n17028), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17027), .ZN(n17029) );
  AOI222_X1 U18837 ( .A1(n17048), .A2(n21824), .B1(n17048), .B2(n17029), .C1(
        n21824), .C2(n17029), .ZN(n17032) );
  NAND2_X1 U18838 ( .A1(n21825), .A2(n17047), .ZN(n17031) );
  INV_X1 U18839 ( .A(n17047), .ZN(n17030) );
  AOI221_X1 U18840 ( .B1(n17032), .B2(n17031), .C1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n17030), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17046) );
  INV_X1 U18841 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17228) );
  NAND2_X1 U18842 ( .A1(n21547), .A2(n17228), .ZN(n17033) );
  NAND2_X1 U18843 ( .A1(n17034), .A2(n17033), .ZN(n17038) );
  NOR2_X1 U18844 ( .A1(n17036), .A2(n17035), .ZN(n17037) );
  AND2_X1 U18845 ( .A1(n17038), .A2(n17037), .ZN(n17043) );
  INV_X1 U18846 ( .A(n17039), .ZN(n17041) );
  INV_X1 U18847 ( .A(n12382), .ZN(n17040) );
  NAND2_X1 U18848 ( .A1(n17041), .A2(n17040), .ZN(n17042) );
  OAI211_X1 U18849 ( .C1(n14443), .C2(n17044), .A(n17043), .B(n17042), .ZN(
        n17045) );
  AOI211_X1 U18850 ( .C1(n17048), .C2(n17047), .A(n17046), .B(n17045), .ZN(
        n21562) );
  OR2_X1 U18851 ( .A1(n21229), .A2(n17049), .ZN(n17054) );
  NOR3_X1 U18852 ( .A1(n17051), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n17050), 
        .ZN(n17052) );
  AOI21_X1 U18853 ( .B1(n17054), .B2(n17053), .A(n17052), .ZN(n17058) );
  OAI221_X1 U18854 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n21562), 
        .A(n17058), .ZN(n21553) );
  OAI211_X1 U18855 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21229), .A(n17055), 
        .B(n21553), .ZN(n21558) );
  NAND4_X1 U18856 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n11847), .A4(n21229), .ZN(n17056) );
  AND2_X1 U18857 ( .A1(n17057), .A2(n17056), .ZN(n21550) );
  AOI21_X1 U18858 ( .B1(n21550), .B2(n17059), .A(n17058), .ZN(n17060) );
  AOI21_X1 U18859 ( .B1(n21549), .B2(n21558), .A(n17060), .ZN(P1_U3162) );
  NOR2_X1 U18860 ( .A1(n17062), .A2(n17061), .ZN(P1_U3032) );
  AND2_X1 U18861 ( .A1(n19784), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U18862 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17122) );
  AOI21_X1 U18863 ( .B1(n17063), .B2(n17122), .A(n22246), .ZN(P1_U2802) );
  INV_X1 U18864 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n19821) );
  INV_X1 U18865 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21523) );
  OAI22_X1 U18866 ( .A1(n21523), .A2(keyinput_61), .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .ZN(n17064) );
  AOI221_X1 U18867 ( .B1(n21523), .B2(keyinput_61), .C1(keyinput_62), .C2(
        P1_REIP_REG_21__SCAN_IN), .A(n17064), .ZN(n17154) );
  INV_X1 U18868 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n17242) );
  INV_X1 U18869 ( .A(keyinput_57), .ZN(n17147) );
  INV_X1 U18870 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19855) );
  XOR2_X1 U18871 ( .A(n21547), .B(keyinput_46), .Z(n17136) );
  OAI22_X1 U18872 ( .A1(NA), .A2(keyinput_34), .B1(HOLD), .B2(keyinput_33), 
        .ZN(n17065) );
  AOI221_X1 U18873 ( .B1(NA), .B2(keyinput_34), .C1(keyinput_33), .C2(HOLD), 
        .A(n17065), .ZN(n17127) );
  XOR2_X1 U18874 ( .A(DATAI_0_), .B(keyinput_32), .Z(n17120) );
  INV_X1 U18875 ( .A(DATAI_5_), .ZN(n17068) );
  INV_X1 U18876 ( .A(DATAI_7_), .ZN(n17067) );
  OAI22_X1 U18877 ( .A1(n17068), .A2(keyinput_27), .B1(n17067), .B2(
        keyinput_25), .ZN(n17066) );
  AOI221_X1 U18878 ( .B1(n17068), .B2(keyinput_27), .C1(keyinput_25), .C2(
        n17067), .A(n17066), .ZN(n17112) );
  AOI22_X1 U18879 ( .A1(DATAI_10_), .A2(keyinput_22), .B1(DATAI_8_), .B2(
        keyinput_24), .ZN(n17069) );
  OAI221_X1 U18880 ( .B1(DATAI_10_), .B2(keyinput_22), .C1(DATAI_8_), .C2(
        keyinput_24), .A(n17069), .ZN(n17076) );
  INV_X1 U18881 ( .A(DATAI_2_), .ZN(n17205) );
  AOI22_X1 U18882 ( .A1(DATAI_6_), .A2(keyinput_26), .B1(n17205), .B2(
        keyinput_30), .ZN(n17070) );
  OAI221_X1 U18883 ( .B1(DATAI_6_), .B2(keyinput_26), .C1(n17205), .C2(
        keyinput_30), .A(n17070), .ZN(n17075) );
  INV_X1 U18884 ( .A(DATAI_4_), .ZN(n17197) );
  INV_X1 U18885 ( .A(DATAI_3_), .ZN(n17198) );
  AOI22_X1 U18886 ( .A1(n17197), .A2(keyinput_28), .B1(keyinput_29), .B2(
        n17198), .ZN(n17071) );
  OAI221_X1 U18887 ( .B1(n17197), .B2(keyinput_28), .C1(n17198), .C2(
        keyinput_29), .A(n17071), .ZN(n17074) );
  INV_X1 U18888 ( .A(DATAI_1_), .ZN(n17202) );
  AOI22_X1 U18889 ( .A1(keyinput_23), .A2(DATAI_9_), .B1(n17202), .B2(
        keyinput_31), .ZN(n17072) );
  OAI221_X1 U18890 ( .B1(keyinput_23), .B2(DATAI_9_), .C1(n17202), .C2(
        keyinput_31), .A(n17072), .ZN(n17073) );
  NOR4_X1 U18891 ( .A1(n17076), .A2(n17075), .A3(n17074), .A4(n17073), .ZN(
        n17111) );
  INV_X1 U18892 ( .A(DATAI_14_), .ZN(n17104) );
  INV_X1 U18893 ( .A(DATAI_16_), .ZN(n21676) );
  AOI22_X1 U18894 ( .A1(n21676), .A2(keyinput_16), .B1(keyinput_17), .B2(
        n13935), .ZN(n17077) );
  OAI221_X1 U18895 ( .B1(n21676), .B2(keyinput_16), .C1(n13935), .C2(
        keyinput_17), .A(n17077), .ZN(n17102) );
  INV_X1 U18896 ( .A(keyinput_15), .ZN(n17100) );
  INV_X1 U18897 ( .A(DATAI_18_), .ZN(n21904) );
  INV_X1 U18898 ( .A(keyinput_11), .ZN(n17094) );
  INV_X1 U18899 ( .A(DATAI_22_), .ZN(n22086) );
  INV_X1 U18900 ( .A(keyinput_10), .ZN(n17092) );
  INV_X1 U18901 ( .A(keyinput_9), .ZN(n17090) );
  INV_X1 U18902 ( .A(keyinput_8), .ZN(n17088) );
  INV_X1 U18903 ( .A(keyinput_7), .ZN(n17086) );
  XNOR2_X1 U18904 ( .A(n15830), .B(keyinput_6), .ZN(n17084) );
  AOI22_X1 U18905 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_0), .B1(
        DATAI_30_), .B2(keyinput_2), .ZN(n17078) );
  OAI221_X1 U18906 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .C1(
        DATAI_30_), .C2(keyinput_2), .A(n17078), .ZN(n17083) );
  AOI22_X1 U18907 ( .A1(DATAI_27_), .A2(keyinput_5), .B1(DATAI_31_), .B2(
        keyinput_1), .ZN(n17079) );
  OAI221_X1 U18908 ( .B1(DATAI_27_), .B2(keyinput_5), .C1(DATAI_31_), .C2(
        keyinput_1), .A(n17079), .ZN(n17082) );
  AOI22_X1 U18909 ( .A1(n15817), .A2(keyinput_4), .B1(n15810), .B2(keyinput_3), 
        .ZN(n17080) );
  OAI221_X1 U18910 ( .B1(n15817), .B2(keyinput_4), .C1(n15810), .C2(keyinput_3), .A(n17080), .ZN(n17081) );
  NOR4_X1 U18911 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17085) );
  AOI221_X1 U18912 ( .B1(DATAI_25_), .B2(n17086), .C1(n15835), .C2(keyinput_7), 
        .A(n17085), .ZN(n17087) );
  AOI221_X1 U18913 ( .B1(DATAI_24_), .B2(n17088), .C1(n21665), .C2(keyinput_8), 
        .A(n17087), .ZN(n17089) );
  AOI221_X1 U18914 ( .B1(DATAI_23_), .B2(keyinput_9), .C1(n15845), .C2(n17090), 
        .A(n17089), .ZN(n17091) );
  AOI221_X1 U18915 ( .B1(DATAI_22_), .B2(keyinput_10), .C1(n22086), .C2(n17092), .A(n17091), .ZN(n17093) );
  AOI221_X1 U18916 ( .B1(DATAI_21_), .B2(n17094), .C1(n15850), .C2(keyinput_11), .A(n17093), .ZN(n17098) );
  INV_X1 U18917 ( .A(DATAI_20_), .ZN(n21993) );
  OAI22_X1 U18918 ( .A1(n21993), .A2(keyinput_12), .B1(DATAI_19_), .B2(
        keyinput_13), .ZN(n17095) );
  AOI221_X1 U18919 ( .B1(n21993), .B2(keyinput_12), .C1(keyinput_13), .C2(
        DATAI_19_), .A(n17095), .ZN(n17096) );
  OAI21_X1 U18920 ( .B1(keyinput_14), .B2(n21904), .A(n17096), .ZN(n17097) );
  AOI211_X1 U18921 ( .C1(keyinput_14), .C2(n21904), .A(n17098), .B(n17097), 
        .ZN(n17099) );
  AOI221_X1 U18922 ( .B1(DATAI_17_), .B2(n17100), .C1(n15861), .C2(keyinput_15), .A(n17099), .ZN(n17101) );
  OAI22_X1 U18923 ( .A1(keyinput_18), .A2(n17104), .B1(n17102), .B2(n17101), 
        .ZN(n17103) );
  AOI21_X1 U18924 ( .B1(keyinput_18), .B2(n17104), .A(n17103), .ZN(n17108) );
  INV_X1 U18925 ( .A(DATAI_12_), .ZN(n17106) );
  AOI22_X1 U18926 ( .A1(DATAI_13_), .A2(keyinput_19), .B1(n17106), .B2(
        keyinput_20), .ZN(n17105) );
  OAI221_X1 U18927 ( .B1(DATAI_13_), .B2(keyinput_19), .C1(n17106), .C2(
        keyinput_20), .A(n17105), .ZN(n17107) );
  AOI211_X1 U18928 ( .C1(DATAI_11_), .C2(keyinput_21), .A(n17108), .B(n17107), 
        .ZN(n17109) );
  OAI21_X1 U18929 ( .B1(DATAI_11_), .B2(keyinput_21), .A(n17109), .ZN(n17110)
         );
  NAND3_X1 U18930 ( .A1(n17112), .A2(n17111), .A3(n17110), .ZN(n17119) );
  AOI22_X1 U18931 ( .A1(keyinput_37), .A2(READY2), .B1(n17114), .B2(
        keyinput_35), .ZN(n17113) );
  OAI221_X1 U18932 ( .B1(keyinput_37), .B2(READY2), .C1(n17114), .C2(
        keyinput_35), .A(n17113), .ZN(n17118) );
  INV_X1 U18933 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17116) );
  INV_X1 U18934 ( .A(READY1), .ZN(n17164) );
  AOI22_X1 U18935 ( .A1(n17116), .A2(keyinput_38), .B1(n17164), .B2(
        keyinput_36), .ZN(n17115) );
  OAI221_X1 U18936 ( .B1(n17116), .B2(keyinput_38), .C1(n17164), .C2(
        keyinput_36), .A(n17115), .ZN(n17117) );
  AOI211_X1 U18937 ( .C1(n17120), .C2(n17119), .A(n17118), .B(n17117), .ZN(
        n17126) );
  INV_X1 U18938 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n19957) );
  AOI22_X1 U18939 ( .A1(n19957), .A2(keyinput_42), .B1(keyinput_39), .B2(
        n17122), .ZN(n17121) );
  OAI221_X1 U18940 ( .B1(n19957), .B2(keyinput_42), .C1(n17122), .C2(
        keyinput_39), .A(n17121), .ZN(n17125) );
  AOI22_X1 U18941 ( .A1(keyinput_40), .A2(P1_CODEFETCH_REG_SCAN_IN), .B1(
        n22244), .B2(keyinput_41), .ZN(n17123) );
  OAI221_X1 U18942 ( .B1(keyinput_40), .B2(P1_CODEFETCH_REG_SCAN_IN), .C1(
        n22244), .C2(keyinput_41), .A(n17123), .ZN(n17124) );
  AOI211_X1 U18943 ( .C1(n17127), .C2(n17126), .A(n17125), .B(n17124), .ZN(
        n17134) );
  AOI22_X1 U18944 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_43), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_44), .ZN(n17128) );
  OAI221_X1 U18945 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_43), 
        .C1(P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_44), .A(n17128), .ZN(
        n17133) );
  OAI22_X1 U18946 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_47), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_48), .ZN(n17129) );
  AOI221_X1 U18947 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_47), .C1(
        keyinput_48), .C2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n17129), .ZN(
        n17132) );
  OAI22_X1 U18948 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_49), .B1(
        P1_MORE_REG_SCAN_IN), .B2(keyinput_45), .ZN(n17130) );
  AOI221_X1 U18949 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_49), .C1(
        keyinput_45), .C2(P1_MORE_REG_SCAN_IN), .A(n17130), .ZN(n17131) );
  OAI211_X1 U18950 ( .C1(n17134), .C2(n17133), .A(n17132), .B(n17131), .ZN(
        n17135) );
  OAI22_X1 U18951 ( .A1(keyinput_50), .A2(n19855), .B1(n17136), .B2(n17135), 
        .ZN(n17137) );
  AOI21_X1 U18952 ( .B1(keyinput_50), .B2(n19855), .A(n17137), .ZN(n17145) );
  AOI22_X1 U18953 ( .A1(n17139), .A2(keyinput_56), .B1(n15889), .B2(
        keyinput_55), .ZN(n17138) );
  OAI221_X1 U18954 ( .B1(n17139), .B2(keyinput_56), .C1(n15889), .C2(
        keyinput_55), .A(n17138), .ZN(n17144) );
  AOI22_X1 U18955 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_53), .B1(n19839), .B2(keyinput_52), .ZN(n17140) );
  OAI221_X1 U18956 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_53), .C1(
        n19839), .C2(keyinput_52), .A(n17140), .ZN(n17143) );
  INV_X1 U18957 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U18958 ( .A1(n19835), .A2(keyinput_54), .B1(keyinput_51), .B2(
        n17161), .ZN(n17141) );
  OAI221_X1 U18959 ( .B1(n19835), .B2(keyinput_54), .C1(n17161), .C2(
        keyinput_51), .A(n17141), .ZN(n17142) );
  NOR4_X1 U18960 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17146) );
  AOI221_X1 U18961 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .C1(
        n17242), .C2(n17147), .A(n17146), .ZN(n17150) );
  AOI22_X1 U18962 ( .A1(n21534), .A2(keyinput_60), .B1(n17157), .B2(
        keyinput_59), .ZN(n17148) );
  OAI221_X1 U18963 ( .B1(n21534), .B2(keyinput_60), .C1(n17157), .C2(
        keyinput_59), .A(n17148), .ZN(n17149) );
  AOI211_X1 U18964 ( .C1(n17152), .C2(keyinput_58), .A(n17150), .B(n17149), 
        .ZN(n17151) );
  OAI21_X1 U18965 ( .B1(n17152), .B2(keyinput_58), .A(n17151), .ZN(n17153) );
  OAI211_X1 U18966 ( .C1(n19821), .C2(keyinput_63), .A(n17154), .B(n17153), 
        .ZN(n17155) );
  AOI21_X1 U18967 ( .B1(n19821), .B2(keyinput_63), .A(n17155), .ZN(n17250) );
  XOR2_X1 U18968 ( .A(keyinput_126), .B(P1_REIP_REG_21__SCAN_IN), .Z(n17249)
         );
  OAI22_X1 U18969 ( .A1(n17157), .A2(keyinput_123), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_124), .ZN(n17156) );
  AOI221_X1 U18970 ( .B1(n17157), .B2(keyinput_123), .C1(keyinput_124), .C2(
        P1_REIP_REG_23__SCAN_IN), .A(n17156), .ZN(n17244) );
  INV_X1 U18971 ( .A(keyinput_121), .ZN(n17241) );
  OAI22_X1 U18972 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_118), .B1(
        keyinput_120), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n17158) );
  AOI221_X1 U18973 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_118), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_120), .A(n17158), .ZN(n17239)
         );
  OAI22_X1 U18974 ( .A1(n19839), .A2(keyinput_116), .B1(keyinput_117), .B2(
        P1_REIP_REG_30__SCAN_IN), .ZN(n17159) );
  AOI221_X1 U18975 ( .B1(n19839), .B2(keyinput_116), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_117), .A(n17159), .ZN(n17238)
         );
  OAI22_X1 U18976 ( .A1(n15889), .A2(keyinput_119), .B1(n17161), .B2(
        keyinput_115), .ZN(n17160) );
  AOI221_X1 U18977 ( .B1(n15889), .B2(keyinput_119), .C1(keyinput_115), .C2(
        n17161), .A(n17160), .ZN(n17237) );
  XOR2_X1 U18978 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_111), .Z(n17234) );
  OAI22_X1 U18979 ( .A1(n21829), .A2(keyinput_108), .B1(keyinput_107), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n17162) );
  AOI221_X1 U18980 ( .B1(n21829), .B2(keyinput_108), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_107), .A(n17162), .ZN(
        n17232) );
  INV_X1 U18981 ( .A(HOLD), .ZN(n21618) );
  AOI22_X1 U18982 ( .A1(n21618), .A2(keyinput_97), .B1(n17164), .B2(
        keyinput_100), .ZN(n17163) );
  OAI221_X1 U18983 ( .B1(n21618), .B2(keyinput_97), .C1(n17164), .C2(
        keyinput_100), .A(n17163), .ZN(n17225) );
  OAI22_X1 U18984 ( .A1(DATAI_13_), .A2(keyinput_83), .B1(DATAI_11_), .B2(
        keyinput_85), .ZN(n17165) );
  AOI221_X1 U18985 ( .B1(DATAI_13_), .B2(keyinput_83), .C1(keyinput_85), .C2(
        DATAI_11_), .A(n17165), .ZN(n17194) );
  OAI22_X1 U18986 ( .A1(n21676), .A2(keyinput_80), .B1(DATAI_15_), .B2(
        keyinput_81), .ZN(n17166) );
  AOI221_X1 U18987 ( .B1(n21676), .B2(keyinput_80), .C1(keyinput_81), .C2(
        DATAI_15_), .A(n17166), .ZN(n17191) );
  INV_X1 U18988 ( .A(keyinput_79), .ZN(n17189) );
  INV_X1 U18989 ( .A(keyinput_75), .ZN(n17183) );
  INV_X1 U18990 ( .A(keyinput_74), .ZN(n17181) );
  INV_X1 U18991 ( .A(keyinput_73), .ZN(n17179) );
  INV_X1 U18992 ( .A(keyinput_72), .ZN(n17177) );
  INV_X1 U18993 ( .A(keyinput_71), .ZN(n17175) );
  XNOR2_X1 U18994 ( .A(n15830), .B(keyinput_70), .ZN(n17173) );
  AOI22_X1 U18995 ( .A1(DATAI_30_), .A2(keyinput_66), .B1(DATAI_31_), .B2(
        keyinput_65), .ZN(n17167) );
  OAI221_X1 U18996 ( .B1(DATAI_30_), .B2(keyinput_66), .C1(DATAI_31_), .C2(
        keyinput_65), .A(n17167), .ZN(n17172) );
  AOI22_X1 U18997 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_64), .B1(
        DATAI_27_), .B2(keyinput_69), .ZN(n17168) );
  OAI221_X1 U18998 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_64), .C1(
        DATAI_27_), .C2(keyinput_69), .A(n17168), .ZN(n17171) );
  AOI22_X1 U18999 ( .A1(DATAI_29_), .A2(keyinput_67), .B1(n15817), .B2(
        keyinput_68), .ZN(n17169) );
  OAI221_X1 U19000 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(n15817), .C2(
        keyinput_68), .A(n17169), .ZN(n17170) );
  NOR4_X1 U19001 ( .A1(n17173), .A2(n17172), .A3(n17171), .A4(n17170), .ZN(
        n17174) );
  AOI221_X1 U19002 ( .B1(DATAI_25_), .B2(keyinput_71), .C1(n15835), .C2(n17175), .A(n17174), .ZN(n17176) );
  AOI221_X1 U19003 ( .B1(DATAI_24_), .B2(keyinput_72), .C1(n21665), .C2(n17177), .A(n17176), .ZN(n17178) );
  AOI221_X1 U19004 ( .B1(DATAI_23_), .B2(n17179), .C1(n15845), .C2(keyinput_73), .A(n17178), .ZN(n17180) );
  AOI221_X1 U19005 ( .B1(DATAI_22_), .B2(n17181), .C1(n22086), .C2(keyinput_74), .A(n17180), .ZN(n17182) );
  AOI221_X1 U19006 ( .B1(DATAI_21_), .B2(n17183), .C1(n15850), .C2(keyinput_75), .A(n17182), .ZN(n17186) );
  AOI22_X1 U19007 ( .A1(DATAI_19_), .A2(keyinput_77), .B1(n21904), .B2(
        keyinput_78), .ZN(n17184) );
  OAI221_X1 U19008 ( .B1(DATAI_19_), .B2(keyinput_77), .C1(n21904), .C2(
        keyinput_78), .A(n17184), .ZN(n17185) );
  AOI211_X1 U19009 ( .C1(DATAI_20_), .C2(keyinput_76), .A(n17186), .B(n17185), 
        .ZN(n17187) );
  OAI21_X1 U19010 ( .B1(DATAI_20_), .B2(keyinput_76), .A(n17187), .ZN(n17188)
         );
  OAI221_X1 U19011 ( .B1(DATAI_17_), .B2(n17189), .C1(n15861), .C2(keyinput_79), .A(n17188), .ZN(n17190) );
  AOI22_X1 U19012 ( .A1(n17191), .A2(n17190), .B1(keyinput_82), .B2(DATAI_14_), 
        .ZN(n17192) );
  OAI21_X1 U19013 ( .B1(keyinput_82), .B2(DATAI_14_), .A(n17192), .ZN(n17193)
         );
  OAI211_X1 U19014 ( .C1(DATAI_12_), .C2(keyinput_84), .A(n17194), .B(n17193), 
        .ZN(n17195) );
  AOI21_X1 U19015 ( .B1(DATAI_12_), .B2(keyinput_84), .A(n17195), .ZN(n17212)
         );
  AOI22_X1 U19016 ( .A1(n17198), .A2(keyinput_93), .B1(n17197), .B2(
        keyinput_92), .ZN(n17196) );
  OAI221_X1 U19017 ( .B1(n17198), .B2(keyinput_93), .C1(n17197), .C2(
        keyinput_92), .A(n17196), .ZN(n17211) );
  OAI22_X1 U19018 ( .A1(DATAI_7_), .A2(keyinput_89), .B1(keyinput_88), .B2(
        DATAI_8_), .ZN(n17199) );
  AOI221_X1 U19019 ( .B1(DATAI_7_), .B2(keyinput_89), .C1(DATAI_8_), .C2(
        keyinput_88), .A(n17199), .ZN(n17209) );
  OAI22_X1 U19020 ( .A1(DATAI_5_), .A2(keyinput_91), .B1(DATAI_9_), .B2(
        keyinput_87), .ZN(n17200) );
  AOI221_X1 U19021 ( .B1(DATAI_5_), .B2(keyinput_91), .C1(keyinput_87), .C2(
        DATAI_9_), .A(n17200), .ZN(n17208) );
  INV_X1 U19022 ( .A(DATAI_6_), .ZN(n17203) );
  OAI22_X1 U19023 ( .A1(n17203), .A2(keyinput_90), .B1(n17202), .B2(
        keyinput_95), .ZN(n17201) );
  AOI221_X1 U19024 ( .B1(n17203), .B2(keyinput_90), .C1(keyinput_95), .C2(
        n17202), .A(n17201), .ZN(n17207) );
  OAI22_X1 U19025 ( .A1(n17205), .A2(keyinput_94), .B1(keyinput_86), .B2(
        DATAI_10_), .ZN(n17204) );
  AOI221_X1 U19026 ( .B1(n17205), .B2(keyinput_94), .C1(DATAI_10_), .C2(
        keyinput_86), .A(n17204), .ZN(n17206) );
  NAND4_X1 U19027 ( .A1(n17209), .A2(n17208), .A3(n17207), .A4(n17206), .ZN(
        n17210) );
  NOR3_X1 U19028 ( .A1(n17212), .A2(n17211), .A3(n17210), .ZN(n17218) );
  XOR2_X1 U19029 ( .A(DATAI_0_), .B(keyinput_96), .Z(n17217) );
  OAI22_X1 U19030 ( .A1(READY2), .A2(keyinput_101), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_102), .ZN(n17213) );
  AOI221_X1 U19031 ( .B1(READY2), .B2(keyinput_101), .C1(keyinput_102), .C2(
        P1_READREQUEST_REG_SCAN_IN), .A(n17213), .ZN(n17216) );
  INV_X1 U19032 ( .A(NA), .ZN(n21607) );
  OAI22_X1 U19033 ( .A1(n21607), .A2(keyinput_98), .B1(keyinput_99), .B2(BS16), 
        .ZN(n17214) );
  AOI221_X1 U19034 ( .B1(n21607), .B2(keyinput_98), .C1(BS16), .C2(keyinput_99), .A(n17214), .ZN(n17215) );
  OAI211_X1 U19035 ( .C1(n17218), .C2(n17217), .A(n17216), .B(n17215), .ZN(
        n17224) );
  INV_X1 U19036 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17220) );
  OAI22_X1 U19037 ( .A1(n17220), .A2(keyinput_104), .B1(n22244), .B2(
        keyinput_105), .ZN(n17219) );
  AOI221_X1 U19038 ( .B1(n17220), .B2(keyinput_104), .C1(keyinput_105), .C2(
        n22244), .A(n17219), .ZN(n17223) );
  OAI22_X1 U19039 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_106), .B1(
        keyinput_103), .B2(P1_ADS_N_REG_SCAN_IN), .ZN(n17221) );
  AOI221_X1 U19040 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_106), .C1(
        P1_ADS_N_REG_SCAN_IN), .C2(keyinput_103), .A(n17221), .ZN(n17222) );
  OAI211_X1 U19041 ( .C1(n17225), .C2(n17224), .A(n17223), .B(n17222), .ZN(
        n17231) );
  INV_X1 U19042 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U19043 ( .A1(n21547), .A2(keyinput_110), .B1(keyinput_112), .B2(
        n19862), .ZN(n17226) );
  OAI221_X1 U19044 ( .B1(n21547), .B2(keyinput_110), .C1(n19862), .C2(
        keyinput_112), .A(n17226), .ZN(n17230) );
  INV_X1 U19045 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19046 ( .A1(n19859), .A2(keyinput_113), .B1(keyinput_109), .B2(
        n17228), .ZN(n17227) );
  OAI221_X1 U19047 ( .B1(n19859), .B2(keyinput_113), .C1(n17228), .C2(
        keyinput_109), .A(n17227), .ZN(n17229) );
  AOI211_X1 U19048 ( .C1(n17232), .C2(n17231), .A(n17230), .B(n17229), .ZN(
        n17233) );
  AOI22_X1 U19049 ( .A1(n17234), .A2(n17233), .B1(keyinput_114), .B2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n17235) );
  OAI21_X1 U19050 ( .B1(keyinput_114), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), .A(
        n17235), .ZN(n17236) );
  NAND4_X1 U19051 ( .A1(n17239), .A2(n17238), .A3(n17237), .A4(n17236), .ZN(
        n17240) );
  OAI221_X1 U19052 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_121), .C1(
        n17242), .C2(n17241), .A(n17240), .ZN(n17243) );
  OAI211_X1 U19053 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(keyinput_122), .A(
        n17244), .B(n17243), .ZN(n17245) );
  AOI21_X1 U19054 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_122), .A(n17245), .ZN(n17248) );
  AOI22_X1 U19055 ( .A1(n21523), .A2(keyinput_125), .B1(n19821), .B2(
        keyinput_127), .ZN(n17246) );
  OAI221_X1 U19056 ( .B1(n21523), .B2(keyinput_125), .C1(n19821), .C2(
        keyinput_127), .A(n17246), .ZN(n17247) );
  NOR4_X1 U19057 ( .A1(n17250), .A2(n17249), .A3(n17248), .A4(n17247), .ZN(
        n17258) );
  AOI22_X1 U19058 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n17256) );
  OAI21_X1 U19059 ( .B1(n17253), .B2(n17252), .A(n17251), .ZN(n17254) );
  INV_X1 U19060 ( .A(n17254), .ZN(n21339) );
  AOI22_X1 U19061 ( .A1(n21339), .A2(n19949), .B1(n19948), .B2(n21642), .ZN(
        n17255) );
  OAI211_X1 U19062 ( .C1(n19952), .C2(n21497), .A(n17256), .B(n17255), .ZN(
        n17257) );
  XOR2_X1 U19063 ( .A(n17258), .B(n17257), .Z(P1_U2981) );
  INV_X1 U19064 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17373) );
  OAI22_X1 U19065 ( .A1(n18341), .A2(n17373), .B1(n18638), .B2(n18646), .ZN(
        P2_U2816) );
  AOI22_X1 U19066 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n18427), .B1(n17260), 
        .B2(n17259), .ZN(n17267) );
  NOR3_X1 U19067 ( .A1(n17262), .A2(n17261), .A3(n17294), .ZN(n17265) );
  NOR2_X1 U19068 ( .A1(n17263), .A2(n17295), .ZN(n17264) );
  AOI211_X1 U19069 ( .C1(n17273), .C2(n14021), .A(n17265), .B(n17264), .ZN(
        n17266) );
  OAI211_X1 U19070 ( .C1(n17269), .C2(n17268), .A(n17267), .B(n17266), .ZN(
        P2_U3011) );
  AOI22_X1 U19071 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17286), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n18427), .ZN(n17277) );
  AOI222_X1 U19072 ( .A1(n17275), .A2(n17274), .B1(n17273), .B2(n17272), .C1(
        n17271), .C2(n17270), .ZN(n17276) );
  OAI211_X1 U19073 ( .C1(n17301), .C2(n17278), .A(n17277), .B(n17276), .ZN(
        P2_U3010) );
  AOI22_X1 U19074 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17286), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n18427), .ZN(n17285) );
  NOR2_X1 U19075 ( .A1(n17279), .A2(n17294), .ZN(n17283) );
  OAI22_X1 U19076 ( .A1(n17281), .A2(n17295), .B1(n17296), .B2(n17280), .ZN(
        n17282) );
  AOI21_X1 U19077 ( .B1(n17283), .B2(n16945), .A(n17282), .ZN(n17284) );
  OAI211_X1 U19078 ( .C1(n17301), .C2(n18378), .A(n17285), .B(n17284), .ZN(
        P2_U3008) );
  AOI22_X1 U19079 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17286), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18427), .ZN(n17299) );
  NAND2_X1 U19080 ( .A1(n17288), .A2(n17287), .ZN(n17289) );
  XNOR2_X1 U19081 ( .A(n17290), .B(n17289), .ZN(n18613) );
  OAI21_X1 U19082 ( .B1(n17293), .B2(n17292), .A(n17291), .ZN(n18609) );
  OAI222_X1 U19083 ( .A1(n18606), .A2(n17296), .B1(n18613), .B2(n17295), .C1(
        n18609), .C2(n17294), .ZN(n17297) );
  INV_X1 U19084 ( .A(n17297), .ZN(n17298) );
  OAI211_X1 U19085 ( .C1(n17301), .C2(n17300), .A(n17299), .B(n17298), .ZN(
        P2_U3006) );
  INV_X1 U19086 ( .A(n17316), .ZN(n17325) );
  INV_X1 U19087 ( .A(n17302), .ZN(n17304) );
  OAI22_X1 U19088 ( .A1(n17305), .A2(n18344), .B1(n17304), .B2(n17303), .ZN(
        n17306) );
  AOI21_X1 U19089 ( .B1(n19274), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17306), 
        .ZN(n17307) );
  OAI22_X1 U19090 ( .A1(n19274), .A2(n17316), .B1(n17325), .B2(n17307), .ZN(
        P2_U3605) );
  NOR2_X1 U19091 ( .A1(n17320), .A2(n21569), .ZN(n17308) );
  INV_X1 U19092 ( .A(n17308), .ZN(n19123) );
  NAND2_X1 U19093 ( .A1(n19123), .A2(n19282), .ZN(n17312) );
  NAND2_X1 U19094 ( .A1(n18638), .A2(n17312), .ZN(n17319) );
  NAND2_X1 U19095 ( .A1(n17309), .A2(n17308), .ZN(n19244) );
  INV_X1 U19096 ( .A(n19244), .ZN(n17310) );
  AOI222_X1 U19097 ( .A1(n19487), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19491), 
        .B2(n17319), .C1(n19282), .C2(n17310), .ZN(n17311) );
  AOI22_X1 U19098 ( .A1(n17325), .A2(n19172), .B1(n17311), .B2(n17316), .ZN(
        P2_U3603) );
  AOI21_X1 U19099 ( .B1(n17320), .B2(n21569), .A(n17312), .ZN(n17315) );
  OAI22_X1 U19100 ( .A1(n17320), .A2(n18638), .B1(n17313), .B2(n19262), .ZN(
        n17314) );
  NOR2_X1 U19101 ( .A1(n17315), .A2(n17314), .ZN(n17317) );
  AOI22_X1 U19102 ( .A1(n17325), .A2(n19272), .B1(n17317), .B2(n17316), .ZN(
        P2_U3604) );
  AOI22_X1 U19103 ( .A1(n19245), .A2(n17319), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n17318), .ZN(n17324) );
  AOI211_X1 U19104 ( .C1(n19185), .C2(n19212), .A(n19276), .B(n21569), .ZN(
        n17322) );
  NOR2_X1 U19105 ( .A1(n17325), .A2(n17322), .ZN(n17323) );
  AOI22_X1 U19106 ( .A1(n19154), .A2(n17325), .B1(n17324), .B2(n17323), .ZN(
        P2_U3602) );
  NAND2_X1 U19107 ( .A1(n17326), .A2(n21571), .ZN(n17329) );
  OAI21_X1 U19108 ( .B1(n12548), .B2(n12555), .A(n17333), .ZN(n17327) );
  OAI21_X1 U19109 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17333), .A(n17327), 
        .ZN(n17328) );
  OAI221_X1 U19110 ( .B1(n17329), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17329), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17328), .ZN(P2_U2822) );
  INV_X1 U19111 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17332) );
  OAI221_X1 U19112 ( .B1(n17333), .B2(n17332), .C1(n17331), .C2(n17330), .A(
        n17329), .ZN(P2_U2823) );
  OAI22_X1 U19113 ( .A1(n17390), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n21598), .ZN(n17334) );
  INV_X1 U19114 ( .A(n17334), .ZN(P2_U3611) );
  INV_X1 U19115 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17335) );
  AOI22_X1 U19116 ( .A1(n21598), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17335), 
        .B2(n17390), .ZN(P2_U3608) );
  AOI21_X1 U19117 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21572), .ZN(n17336) );
  INV_X1 U19118 ( .A(n17336), .ZN(P2_U2815) );
  INV_X1 U19119 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U19120 ( .A1(n17369), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17338) );
  OAI21_X1 U19121 ( .B1(n17339), .B2(n17371), .A(n17338), .ZN(P2_U2951) );
  INV_X1 U19122 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17341) );
  AOI22_X1 U19123 ( .A1(n17369), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17340) );
  OAI21_X1 U19124 ( .B1(n17341), .B2(n17371), .A(n17340), .ZN(P2_U2950) );
  INV_X1 U19125 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19495) );
  AOI22_X1 U19126 ( .A1(n17369), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17342) );
  OAI21_X1 U19127 ( .B1(n19495), .B2(n17371), .A(n17342), .ZN(P2_U2949) );
  INV_X1 U19128 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U19129 ( .A1(n17358), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17343) );
  OAI21_X1 U19130 ( .B1(n17344), .B2(n17371), .A(n17343), .ZN(P2_U2948) );
  INV_X1 U19131 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U19132 ( .A1(n17369), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17345) );
  OAI21_X1 U19133 ( .B1(n17346), .B2(n17371), .A(n17345), .ZN(P2_U2947) );
  INV_X1 U19134 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U19135 ( .A1(n17358), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17347) );
  OAI21_X1 U19136 ( .B1(n17348), .B2(n17371), .A(n17347), .ZN(P2_U2946) );
  AOI22_X1 U19137 ( .A1(n17358), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17349) );
  OAI21_X1 U19138 ( .B1(n17350), .B2(n17371), .A(n17349), .ZN(P2_U2945) );
  AOI22_X1 U19139 ( .A1(n17358), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17351) );
  OAI21_X1 U19140 ( .B1(n17352), .B2(n17371), .A(n17351), .ZN(P2_U2944) );
  AOI22_X1 U19141 ( .A1(n17358), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17353) );
  OAI21_X1 U19142 ( .B1(n17354), .B2(n17371), .A(n17353), .ZN(P2_U2943) );
  AOI22_X1 U19143 ( .A1(n17369), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17355) );
  OAI21_X1 U19144 ( .B1(n17356), .B2(n17371), .A(n17355), .ZN(P2_U2942) );
  AOI22_X1 U19145 ( .A1(n17358), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17359) );
  OAI21_X1 U19146 ( .B1(n17360), .B2(n17371), .A(n17359), .ZN(P2_U2941) );
  AOI22_X1 U19147 ( .A1(n17369), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U19148 ( .B1(n17362), .B2(n17371), .A(n17361), .ZN(P2_U2940) );
  AOI22_X1 U19149 ( .A1(n17369), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U19150 ( .B1(n17364), .B2(n17371), .A(n17363), .ZN(P2_U2939) );
  AOI22_X1 U19151 ( .A1(n17369), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U19152 ( .B1(n17366), .B2(n17371), .A(n17365), .ZN(P2_U2938) );
  AOI22_X1 U19153 ( .A1(n17369), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17367) );
  OAI21_X1 U19154 ( .B1(n17368), .B2(n17371), .A(n17367), .ZN(P2_U2937) );
  AOI22_X1 U19155 ( .A1(n17369), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17357), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17370) );
  OAI21_X1 U19156 ( .B1(n17372), .B2(n17371), .A(n17370), .ZN(P2_U2936) );
  AOI22_X1 U19157 ( .A1(n21598), .A2(n17373), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n17390), .ZN(n17374) );
  OAI21_X1 U19158 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21596), .A(n17374), 
        .ZN(P2_U2817) );
  INV_X1 U19159 ( .A(n17382), .ZN(n17387) );
  NOR2_X1 U19160 ( .A1(n21612), .A2(n17390), .ZN(n21600) );
  INV_X1 U19161 ( .A(n21600), .ZN(n21611) );
  OAI222_X1 U19162 ( .A1(n17387), .A2(n12577), .B1(n17375), .B2(n21598), .C1(
        n12548), .C2(n21611), .ZN(P2_U3212) );
  INV_X1 U19163 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19713) );
  OAI222_X1 U19164 ( .A1(n17387), .A2(n13263), .B1(n19713), .B2(n21598), .C1(
        n12577), .C2(n21611), .ZN(P2_U3213) );
  INV_X1 U19165 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19715) );
  OAI222_X1 U19166 ( .A1(n17387), .A2(n14618), .B1(n19715), .B2(n21598), .C1(
        n13263), .C2(n21611), .ZN(P2_U3214) );
  INV_X1 U19167 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19717) );
  OAI222_X1 U19168 ( .A1(n17387), .A2(n13225), .B1(n19717), .B2(n21598), .C1(
        n14618), .C2(n21611), .ZN(P2_U3215) );
  INV_X1 U19169 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19719) );
  OAI222_X1 U19170 ( .A1(n17387), .A2(n18372), .B1(n19719), .B2(n21598), .C1(
        n13225), .C2(n21611), .ZN(P2_U3216) );
  INV_X1 U19171 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19721) );
  OAI222_X1 U19172 ( .A1(n17387), .A2(n13095), .B1(n19721), .B2(n21598), .C1(
        n18372), .C2(n21611), .ZN(P2_U3217) );
  AOI222_X1 U19173 ( .A1(n17382), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n17390), .C1(P2_REIP_REG_7__SCAN_IN), 
        .C2(n21600), .ZN(n17376) );
  INV_X1 U19174 ( .A(n17376), .ZN(P2_U3218) );
  AOI222_X1 U19175 ( .A1(n17382), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n17390), .C1(P2_REIP_REG_8__SCAN_IN), 
        .C2(n21600), .ZN(n17377) );
  INV_X1 U19176 ( .A(n17377), .ZN(P2_U3219) );
  INV_X1 U19177 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19725) );
  OAI222_X1 U19178 ( .A1(n21611), .A2(n18402), .B1(n19725), .B2(n21598), .C1(
        n16615), .C2(n17387), .ZN(P2_U3220) );
  INV_X1 U19179 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19727) );
  OAI222_X1 U19180 ( .A1(n21611), .A2(n16615), .B1(n19727), .B2(n21598), .C1(
        n16597), .C2(n17387), .ZN(P2_U3221) );
  INV_X1 U19181 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19729) );
  OAI222_X1 U19182 ( .A1(n21611), .A2(n16597), .B1(n19729), .B2(n21598), .C1(
        n16590), .C2(n17387), .ZN(P2_U3222) );
  AOI222_X1 U19183 ( .A1(n21600), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n17390), .C1(P2_REIP_REG_13__SCAN_IN), 
        .C2(n17382), .ZN(n17378) );
  INV_X1 U19184 ( .A(n17378), .ZN(P2_U3223) );
  AOI222_X1 U19185 ( .A1(n21600), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n17390), .C1(P2_REIP_REG_14__SCAN_IN), 
        .C2(n17382), .ZN(n17379) );
  INV_X1 U19186 ( .A(n17379), .ZN(P2_U3224) );
  INV_X1 U19187 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19733) );
  OAI222_X1 U19188 ( .A1(n21611), .A2(n16570), .B1(n19733), .B2(n21598), .C1(
        n18442), .C2(n17387), .ZN(P2_U3225) );
  INV_X1 U19189 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19735) );
  OAI222_X1 U19190 ( .A1(n21611), .A2(n18442), .B1(n19735), .B2(n21598), .C1(
        n13124), .C2(n17387), .ZN(P2_U3226) );
  INV_X1 U19191 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19737) );
  OAI222_X1 U19192 ( .A1(n21611), .A2(n13124), .B1(n19737), .B2(n21598), .C1(
        n16535), .C2(n17387), .ZN(P2_U3227) );
  INV_X1 U19193 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19739) );
  OAI222_X1 U19194 ( .A1(n21611), .A2(n16535), .B1(n19739), .B2(n21598), .C1(
        n16522), .C2(n17387), .ZN(P2_U3228) );
  INV_X1 U19195 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19741) );
  OAI222_X1 U19196 ( .A1(n17387), .A2(n18490), .B1(n19741), .B2(n21598), .C1(
        n16522), .C2(n21611), .ZN(P2_U3229) );
  INV_X1 U19197 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19743) );
  OAI222_X1 U19198 ( .A1(n21611), .A2(n18490), .B1(n19743), .B2(n21598), .C1(
        n13136), .C2(n17387), .ZN(P2_U3230) );
  INV_X1 U19199 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19745) );
  OAI222_X1 U19200 ( .A1(n17387), .A2(n18513), .B1(n19745), .B2(n21598), .C1(
        n13136), .C2(n21611), .ZN(P2_U3231) );
  INV_X1 U19201 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19747) );
  OAI222_X1 U19202 ( .A1(n17387), .A2(n13143), .B1(n19747), .B2(n21598), .C1(
        n18513), .C2(n21611), .ZN(P2_U3232) );
  INV_X1 U19203 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19749) );
  OAI222_X1 U19204 ( .A1(n17387), .A2(n17380), .B1(n19749), .B2(n21598), .C1(
        n13143), .C2(n21611), .ZN(P2_U3233) );
  INV_X1 U19205 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19751) );
  OAI222_X1 U19206 ( .A1(n17387), .A2(n13149), .B1(n19751), .B2(n21598), .C1(
        n17380), .C2(n21611), .ZN(P2_U3234) );
  INV_X1 U19207 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19753) );
  OAI222_X1 U19208 ( .A1(n17387), .A2(n18547), .B1(n19753), .B2(n21598), .C1(
        n13149), .C2(n21611), .ZN(P2_U3235) );
  AOI222_X1 U19209 ( .A1(n21600), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(n17390), .C1(P2_REIP_REG_26__SCAN_IN), 
        .C2(n17382), .ZN(n17381) );
  INV_X1 U19210 ( .A(n17381), .ZN(P2_U3236) );
  AOI222_X1 U19211 ( .A1(n17382), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(n17390), .C1(P2_REIP_REG_26__SCAN_IN), 
        .C2(n21600), .ZN(n17383) );
  INV_X1 U19212 ( .A(n17383), .ZN(P2_U3237) );
  INV_X1 U19213 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19757) );
  OAI222_X1 U19214 ( .A1(n21611), .A2(n17384), .B1(n19757), .B2(n21598), .C1(
        n17385), .C2(n17387), .ZN(P2_U3238) );
  INV_X1 U19215 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19759) );
  OAI222_X1 U19216 ( .A1(n21611), .A2(n17385), .B1(n19759), .B2(n21598), .C1(
        n18563), .C2(n17387), .ZN(P2_U3239) );
  INV_X1 U19217 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19761) );
  OAI222_X1 U19218 ( .A1(n21611), .A2(n18563), .B1(n19761), .B2(n21598), .C1(
        n17386), .C2(n17387), .ZN(P2_U3240) );
  INV_X1 U19219 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19764) );
  OAI222_X1 U19220 ( .A1(n17387), .A2(n13416), .B1(n19764), .B2(n21598), .C1(
        n17386), .C2(n21611), .ZN(P2_U3241) );
  OAI22_X1 U19221 ( .A1(n17390), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n21598), .ZN(n17388) );
  INV_X1 U19222 ( .A(n17388), .ZN(P2_U3588) );
  OAI22_X1 U19223 ( .A1(n17390), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n21598), .ZN(n17389) );
  INV_X1 U19224 ( .A(n17389), .ZN(P2_U3587) );
  MUX2_X1 U19225 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n17390), .Z(P2_U3586) );
  OAI22_X1 U19226 ( .A1(n17390), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n21598), .ZN(n17391) );
  INV_X1 U19227 ( .A(n17391), .ZN(P2_U3585) );
  NAND2_X1 U19228 ( .A1(n17655), .A2(n17392), .ZN(n17411) );
  INV_X1 U19229 ( .A(n17411), .ZN(n17419) );
  NOR2_X1 U19230 ( .A1(n20592), .A2(n17657), .ZN(n17650) );
  AOI22_X1 U19231 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17654), .B1(n17393), .B2(
        n17650), .ZN(n17394) );
  OAI22_X1 U19232 ( .A1(n17419), .A2(n17394), .B1(n17725), .B2(n17654), .ZN(
        P3_U2699) );
  NAND4_X1 U19233 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(n17650), .ZN(n17398) );
  NAND3_X1 U19234 ( .A1(n17398), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17654), .ZN(
        n17395) );
  OAI221_X1 U19235 ( .B1(n17398), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17654), 
        .C2(n17396), .A(n17395), .ZN(P3_U2700) );
  INV_X1 U19236 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17699) );
  NAND2_X1 U19237 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17397) );
  INV_X1 U19238 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20078) );
  OAI21_X1 U19239 ( .B1(n17657), .B2(n17397), .A(n20078), .ZN(n17399) );
  NAND3_X1 U19240 ( .A1(n17654), .A2(n17399), .A3(n17398), .ZN(n17400) );
  OAI21_X1 U19241 ( .B1(n17654), .B2(n17699), .A(n17400), .ZN(P3_U2701) );
  AOI22_X1 U19242 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U19243 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17403) );
  AOI22_X1 U19244 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U19245 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17401) );
  NAND4_X1 U19246 ( .A1(n17404), .A2(n17403), .A3(n17402), .A4(n17401), .ZN(
        n17410) );
  AOI22_X1 U19247 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U19248 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17759), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U19249 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U19250 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17405) );
  NAND4_X1 U19251 ( .A1(n17408), .A2(n17407), .A3(n17406), .A4(n17405), .ZN(
        n17409) );
  NOR2_X1 U19252 ( .A1(n17410), .A2(n17409), .ZN(n20661) );
  NAND2_X1 U19253 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17422), .ZN(n17417) );
  NOR2_X1 U19254 ( .A1(n20146), .A2(n17417), .ZN(n17416) );
  NAND2_X1 U19255 ( .A1(n17412), .A2(n17422), .ZN(n17528) );
  OAI221_X1 U19256 ( .B1(n17416), .B2(P3_EBX_REG_8__SCAN_IN), .C1(n20671), 
        .C2(n17657), .A(n17528), .ZN(n17413) );
  OAI21_X1 U19257 ( .B1(n20661), .B2(n17654), .A(n17413), .ZN(P3_U2695) );
  NOR2_X1 U19258 ( .A1(n20592), .A2(n17417), .ZN(n17504) );
  AOI21_X1 U19259 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17654), .A(n17504), .ZN(
        n17415) );
  OAI22_X1 U19260 ( .A1(n17416), .A2(n17415), .B1(n17414), .B2(n17654), .ZN(
        P3_U2696) );
  OAI21_X1 U19261 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17422), .A(n17417), .ZN(
        n17418) );
  AOI22_X1 U19262 ( .A1(n17658), .A2(n17739), .B1(n17418), .B2(n17654), .ZN(
        P3_U2697) );
  OAI21_X1 U19263 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17419), .A(n17654), .ZN(
        n17421) );
  OAI22_X1 U19264 ( .A1(n17422), .A2(n17421), .B1(n17420), .B2(n17654), .ZN(
        P3_U2698) );
  AOI22_X1 U19265 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U19266 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U19267 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U19268 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17423) );
  NAND4_X1 U19269 ( .A1(n17426), .A2(n17425), .A3(n17424), .A4(n17423), .ZN(
        n17432) );
  AOI22_X1 U19270 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U19271 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U19272 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U19273 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17427) );
  NAND4_X1 U19274 ( .A1(n17430), .A2(n17429), .A3(n17428), .A4(n17427), .ZN(
        n17431) );
  NOR2_X1 U19275 ( .A1(n17432), .A2(n17431), .ZN(n20643) );
  INV_X1 U19276 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20260) );
  INV_X1 U19277 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20233) );
  NOR2_X1 U19278 ( .A1(n17433), .A2(n17528), .ZN(n17502) );
  NAND2_X1 U19279 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17478), .ZN(n17460) );
  NOR2_X1 U19280 ( .A1(n20233), .A2(n17460), .ZN(n17476) );
  NAND2_X1 U19281 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17476), .ZN(n17436) );
  NOR2_X1 U19282 ( .A1(n20260), .A2(n17436), .ZN(n17449) );
  NAND2_X1 U19283 ( .A1(n17449), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17434) );
  OAI221_X1 U19284 ( .B1(n17449), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n20671), 
        .C2(n17657), .A(n17434), .ZN(n17435) );
  OAI21_X1 U19285 ( .B1(n20643), .B2(n17654), .A(n17435), .ZN(P3_U2687) );
  NAND2_X1 U19286 ( .A1(n20260), .A2(n17436), .ZN(n17437) );
  NAND2_X1 U19287 ( .A1(n17437), .A2(n17654), .ZN(n17448) );
  AOI22_X1 U19288 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U19289 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U19290 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U19291 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17438) );
  NAND4_X1 U19292 ( .A1(n17441), .A2(n17440), .A3(n17439), .A4(n17438), .ZN(
        n17447) );
  AOI22_X1 U19293 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U19294 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U19295 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U19296 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17442) );
  NAND4_X1 U19297 ( .A1(n17445), .A2(n17444), .A3(n17443), .A4(n17442), .ZN(
        n17446) );
  NOR2_X1 U19298 ( .A1(n17447), .A2(n17446), .ZN(n20654) );
  OAI22_X1 U19299 ( .A1(n17449), .A2(n17448), .B1(n20654), .B2(n17654), .ZN(
        P3_U2688) );
  AOI22_X1 U19300 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U19301 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U19302 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U19303 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17450) );
  NAND4_X1 U19304 ( .A1(n17453), .A2(n17452), .A3(n17451), .A4(n17450), .ZN(
        n17459) );
  AOI22_X1 U19305 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U19306 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U19307 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U19308 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17454) );
  NAND4_X1 U19309 ( .A1(n17457), .A2(n17456), .A3(n17455), .A4(n17454), .ZN(
        n17458) );
  NOR2_X1 U19310 ( .A1(n17459), .A2(n17458), .ZN(n20507) );
  INV_X1 U19311 ( .A(n17460), .ZN(n17462) );
  NOR2_X1 U19312 ( .A1(n17658), .A2(n17476), .ZN(n17461) );
  OAI21_X1 U19313 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17462), .A(n17461), .ZN(
        n17463) );
  OAI21_X1 U19314 ( .B1(n20507), .B2(n17654), .A(n17463), .ZN(P3_U2690) );
  AOI22_X1 U19315 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U19316 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19317 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U19318 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17465) );
  NAND4_X1 U19319 ( .A1(n17468), .A2(n17467), .A3(n17466), .A4(n17465), .ZN(
        n17474) );
  AOI22_X1 U19320 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U19321 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19322 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U19323 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17469) );
  NAND4_X1 U19324 ( .A1(n17472), .A2(n17471), .A3(n17470), .A4(n17469), .ZN(
        n17473) );
  NOR2_X1 U19325 ( .A1(n17474), .A2(n17473), .ZN(n20648) );
  OAI22_X1 U19326 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20592), .B1(n17658), 
        .B2(n17476), .ZN(n17475) );
  OAI21_X1 U19327 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17476), .A(n17475), .ZN(
        n17477) );
  OAI21_X1 U19328 ( .B1(n20648), .B2(n17654), .A(n17477), .ZN(P3_U2689) );
  NAND2_X1 U19329 ( .A1(n20671), .A2(n17478), .ZN(n17490) );
  NOR2_X1 U19330 ( .A1(n17658), .A2(n17478), .ZN(n17501) );
  AOI22_X1 U19331 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U19332 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U19333 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17479) );
  OAI21_X1 U19334 ( .B1(n17518), .B2(n17725), .A(n17479), .ZN(n17485) );
  AOI22_X1 U19335 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U19336 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U19337 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U19338 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17480) );
  NAND4_X1 U19339 ( .A1(n17483), .A2(n17482), .A3(n17481), .A4(n17480), .ZN(
        n17484) );
  AOI211_X1 U19340 ( .C1(n10993), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17485), .B(n17484), .ZN(n17486) );
  NAND3_X1 U19341 ( .A1(n17488), .A2(n17487), .A3(n17486), .ZN(n20510) );
  AOI22_X1 U19342 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17501), .B1(n17658), 
        .B2(n20510), .ZN(n17489) );
  OAI21_X1 U19343 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17490), .A(n17489), .ZN(
        P3_U2691) );
  AOI22_X1 U19344 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U19345 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U19346 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U19347 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17491) );
  NAND4_X1 U19348 ( .A1(n17494), .A2(n17493), .A3(n17492), .A4(n17491), .ZN(
        n17500) );
  AOI22_X1 U19349 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U19350 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U19351 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U19352 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17495) );
  NAND4_X1 U19353 ( .A1(n17498), .A2(n17497), .A3(n17496), .A4(n17495), .ZN(
        n17499) );
  NOR2_X1 U19354 ( .A1(n17500), .A2(n17499), .ZN(n20514) );
  OAI21_X1 U19355 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17502), .A(n17501), .ZN(
        n17503) );
  OAI21_X1 U19356 ( .B1(n20514), .B2(n17654), .A(n17503), .ZN(P3_U2692) );
  NAND4_X1 U19357 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_7__SCAN_IN), .A4(n17504), .ZN(n17529) );
  AOI22_X1 U19358 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U19359 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U19360 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U19361 ( .B1(n17518), .B2(n17699), .A(n17505), .ZN(n17511) );
  AOI22_X1 U19362 ( .A1(n15054), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U19363 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U19364 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U19365 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17506) );
  NAND4_X1 U19366 ( .A1(n17509), .A2(n17508), .A3(n17507), .A4(n17506), .ZN(
        n17510) );
  AOI211_X1 U19367 ( .C1(n17759), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n17511), .B(n17510), .ZN(n17512) );
  NAND3_X1 U19368 ( .A1(n17514), .A2(n17513), .A3(n17512), .ZN(n20520) );
  INV_X1 U19369 ( .A(n20520), .ZN(n17516) );
  NAND3_X1 U19370 ( .A1(n17529), .A2(P3_EBX_REG_10__SCAN_IN), .A3(n17654), 
        .ZN(n17515) );
  OAI221_X1 U19371 ( .B1(n17529), .B2(P3_EBX_REG_10__SCAN_IN), .C1(n17654), 
        .C2(n17516), .A(n17515), .ZN(P3_U2693) );
  AOI22_X1 U19372 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10972), .ZN(n17527) );
  AOI22_X1 U19373 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17741), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U19374 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10976), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U19375 ( .B1(n17518), .B2(n17712), .A(n17517), .ZN(n17524) );
  AOI22_X1 U19376 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17722), .ZN(n17522) );
  AOI22_X1 U19377 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17521) );
  AOI22_X1 U19378 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17520) );
  AOI22_X1 U19379 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17687), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17737), .ZN(n17519) );
  NAND4_X1 U19380 ( .A1(n17522), .A2(n17521), .A3(n17520), .A4(n17519), .ZN(
        n17523) );
  AOI211_X1 U19381 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n10970), .A(
        n17524), .B(n17523), .ZN(n17525) );
  NAND3_X1 U19382 ( .A1(n17527), .A2(n17526), .A3(n17525), .ZN(n20523) );
  INV_X1 U19383 ( .A(n20523), .ZN(n17532) );
  INV_X1 U19384 ( .A(n17528), .ZN(n17530) );
  OAI211_X1 U19385 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17530), .A(n17529), .B(
        n17654), .ZN(n17531) );
  OAI21_X1 U19386 ( .B1(n17532), .B2(n17654), .A(n17531), .ZN(P3_U2694) );
  INV_X1 U19387 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20064) );
  OAI33_X1 U19388 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17534), .A3(n20592), 
        .B1(n20064), .B2(n17658), .B3(n17533), .ZN(P3_U2672) );
  OR2_X1 U19389 ( .A1(n20592), .A2(n17535), .ZN(n17547) );
  INV_X1 U19390 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20352) );
  NAND2_X1 U19391 ( .A1(n17654), .A2(n17535), .ZN(n17611) );
  AOI22_X1 U19392 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U19393 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U19394 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U19395 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17536) );
  NAND4_X1 U19396 ( .A1(n17539), .A2(n17538), .A3(n17537), .A4(n17536), .ZN(
        n17545) );
  AOI22_X1 U19397 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U19398 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U19399 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U19400 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17540) );
  NAND4_X1 U19401 ( .A1(n17543), .A2(n17542), .A3(n17541), .A4(n17540), .ZN(
        n17544) );
  NOR2_X1 U19402 ( .A1(n17545), .A2(n17544), .ZN(n20560) );
  OR2_X1 U19403 ( .A1(n20560), .A2(n17654), .ZN(n17546) );
  OAI221_X1 U19404 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17547), .C1(n20352), 
        .C2(n17611), .A(n17546), .ZN(P3_U2682) );
  INV_X1 U19405 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20370) );
  NOR2_X1 U19406 ( .A1(n20352), .A2(n17547), .ZN(n17585) );
  NAND2_X1 U19407 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17585), .ZN(n17578) );
  NOR2_X1 U19408 ( .A1(n20370), .A2(n17578), .ZN(n17584) );
  NAND2_X1 U19409 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17584), .ZN(n17564) );
  NAND3_X1 U19410 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17577), .ZN(n17548) );
  INV_X1 U19411 ( .A(n17548), .ZN(n17568) );
  NAND2_X1 U19412 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17568), .ZN(n17563) );
  INV_X1 U19413 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20426) );
  OAI21_X1 U19414 ( .B1(n20426), .B2(n17658), .A(n17548), .ZN(n17550) );
  AOI21_X1 U19415 ( .B1(n17549), .B2(n17565), .A(n17561), .ZN(n20619) );
  AOI22_X1 U19416 ( .A1(n17563), .A2(n17550), .B1(n20619), .B2(n17658), .ZN(
        n17551) );
  INV_X1 U19417 ( .A(n17551), .ZN(P3_U2676) );
  INV_X1 U19418 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20453) );
  NAND3_X1 U19419 ( .A1(n20453), .A2(n17552), .A3(n20671), .ZN(n17558) );
  INV_X1 U19420 ( .A(n17650), .ZN(n17660) );
  NAND2_X1 U19421 ( .A1(n17654), .A2(n17563), .ZN(n17553) );
  OAI21_X1 U19422 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17660), .A(n17553), .ZN(
        n17556) );
  AOI21_X1 U19423 ( .B1(n17555), .B2(n17559), .A(n17554), .ZN(n20609) );
  AOI22_X1 U19424 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17556), .B1(n20609), 
        .B2(n17658), .ZN(n17557) );
  NAND2_X1 U19425 ( .A1(n17558), .A2(n17557), .ZN(P3_U2674) );
  OAI21_X1 U19426 ( .B1(n17561), .B2(n17560), .A(n17559), .ZN(n20618) );
  NAND3_X1 U19427 ( .A1(n17563), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n17654), 
        .ZN(n17562) );
  OAI221_X1 U19428 ( .B1(n17563), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n17654), 
        .C2(n20618), .A(n17562), .ZN(P3_U2675) );
  INV_X1 U19429 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20397) );
  NOR2_X1 U19430 ( .A1(n20397), .A2(n17564), .ZN(n17573) );
  AOI21_X1 U19431 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17654), .A(n17573), .ZN(
        n17567) );
  OAI21_X1 U19432 ( .B1(n17569), .B2(n17566), .A(n17565), .ZN(n20601) );
  OAI22_X1 U19433 ( .A1(n17568), .A2(n17567), .B1(n20601), .B2(n17654), .ZN(
        P3_U2677) );
  AOI21_X1 U19434 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17654), .A(n17577), .ZN(
        n17572) );
  AOI21_X1 U19435 ( .B1(n17570), .B2(n17574), .A(n17569), .ZN(n20591) );
  INV_X1 U19436 ( .A(n20591), .ZN(n17571) );
  OAI22_X1 U19437 ( .A1(n17573), .A2(n17572), .B1(n17571), .B2(n17654), .ZN(
        P3_U2678) );
  AOI21_X1 U19438 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17654), .A(n17584), .ZN(
        n17576) );
  OAI21_X1 U19439 ( .B1(n17579), .B2(n17575), .A(n17574), .ZN(n20629) );
  OAI22_X1 U19440 ( .A1(n17577), .A2(n17576), .B1(n20629), .B2(n17654), .ZN(
        P3_U2679) );
  INV_X1 U19441 ( .A(n17578), .ZN(n17599) );
  AOI21_X1 U19442 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17654), .A(n17599), .ZN(
        n17583) );
  AOI21_X1 U19443 ( .B1(n17581), .B2(n17580), .A(n17579), .ZN(n20630) );
  INV_X1 U19444 ( .A(n20630), .ZN(n17582) );
  OAI22_X1 U19445 ( .A1(n17584), .A2(n17583), .B1(n17582), .B2(n17654), .ZN(
        P3_U2680) );
  AOI21_X1 U19446 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17654), .A(n17585), .ZN(
        n17598) );
  AOI22_X1 U19447 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19448 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U19449 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17586) );
  OAI21_X1 U19450 ( .B1(n17587), .B2(n17739), .A(n17586), .ZN(n17593) );
  AOI22_X1 U19451 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17759), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17591) );
  AOI22_X1 U19452 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17590) );
  AOI22_X1 U19453 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17589) );
  AOI22_X1 U19454 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17588) );
  NAND4_X1 U19455 ( .A1(n17591), .A2(n17590), .A3(n17589), .A4(n17588), .ZN(
        n17592) );
  AOI211_X1 U19456 ( .C1(n10977), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17593), .B(n17592), .ZN(n17594) );
  NAND3_X1 U19457 ( .A1(n17596), .A2(n17595), .A3(n17594), .ZN(n20573) );
  INV_X1 U19458 ( .A(n20573), .ZN(n17597) );
  OAI22_X1 U19459 ( .A1(n17599), .A2(n17598), .B1(n17597), .B2(n17654), .ZN(
        P3_U2681) );
  AOI22_X1 U19460 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17603) );
  AOI22_X1 U19461 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17602) );
  AOI22_X1 U19462 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17464), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17601) );
  AOI22_X1 U19463 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17600) );
  NAND4_X1 U19464 ( .A1(n17603), .A2(n17602), .A3(n17601), .A4(n17600), .ZN(
        n17609) );
  AOI22_X1 U19465 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U19466 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U19467 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17605) );
  AOI22_X1 U19468 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17604) );
  NAND4_X1 U19469 ( .A1(n17607), .A2(n17606), .A3(n17605), .A4(n17604), .ZN(
        n17608) );
  NOR2_X1 U19470 ( .A1(n17609), .A2(n17608), .ZN(n20567) );
  AND2_X1 U19471 ( .A1(n17610), .A2(n17650), .ZN(n17636) );
  AOI21_X1 U19472 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17636), .A(
        P3_EBX_REG_20__SCAN_IN), .ZN(n17612) );
  OAI22_X1 U19473 ( .A1(n20567), .A2(n17654), .B1(n17612), .B2(n17611), .ZN(
        P3_U2683) );
  AOI22_X1 U19474 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U19475 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17615) );
  AOI22_X1 U19476 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U19477 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17613) );
  NAND4_X1 U19478 ( .A1(n17616), .A2(n17615), .A3(n17614), .A4(n17613), .ZN(
        n17622) );
  AOI22_X1 U19479 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U19480 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17619) );
  AOI22_X1 U19481 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U19482 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17617) );
  NAND4_X1 U19483 ( .A1(n17620), .A2(n17619), .A3(n17618), .A4(n17617), .ZN(
        n17621) );
  NOR2_X1 U19484 ( .A1(n17622), .A2(n17621), .ZN(n20585) );
  OAI21_X1 U19485 ( .B1(n17649), .B2(n17660), .A(n20304), .ZN(n17624) );
  NOR2_X1 U19486 ( .A1(n17658), .A2(n17623), .ZN(n17637) );
  NAND2_X1 U19487 ( .A1(n17624), .A2(n17637), .ZN(n17625) );
  OAI21_X1 U19488 ( .B1(n20585), .B2(n17654), .A(n17625), .ZN(P3_U2685) );
  AOI22_X1 U19489 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17629) );
  AOI22_X1 U19490 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15091), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U19491 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U19492 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17626) );
  NAND4_X1 U19493 ( .A1(n17629), .A2(n17628), .A3(n17627), .A4(n17626), .ZN(
        n17635) );
  AOI22_X1 U19494 ( .A1(n17759), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U19495 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17632) );
  AOI22_X1 U19496 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17631) );
  AOI22_X1 U19497 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17630) );
  NAND4_X1 U19498 ( .A1(n17633), .A2(n17632), .A3(n17631), .A4(n17630), .ZN(
        n17634) );
  NOR2_X1 U19499 ( .A1(n17635), .A2(n17634), .ZN(n20581) );
  INV_X1 U19500 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20317) );
  AOI22_X1 U19501 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17637), .B1(n17636), 
        .B2(n20317), .ZN(n17638) );
  OAI21_X1 U19502 ( .B1(n20581), .B2(n17654), .A(n17638), .ZN(P3_U2684) );
  AOI22_X1 U19503 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17740), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U19504 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17641) );
  AOI22_X1 U19505 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17764), .ZN(n17640) );
  AOI22_X1 U19506 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17687), .ZN(n17639) );
  NAND4_X1 U19507 ( .A1(n17642), .A2(n17641), .A3(n17640), .A4(n17639), .ZN(
        n17648) );
  AOI22_X1 U19508 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17759), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n10993), .ZN(n17646) );
  AOI22_X1 U19509 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17741), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17735), .ZN(n17645) );
  AOI22_X1 U19510 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10972), .ZN(n17644) );
  AOI22_X1 U19511 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10970), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17643) );
  NAND4_X1 U19512 ( .A1(n17646), .A2(n17645), .A3(n17644), .A4(n17643), .ZN(
        n17647) );
  NOR2_X1 U19513 ( .A1(n17648), .A2(n17647), .ZN(n20590) );
  NAND2_X1 U19514 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17657), .ZN(n17653) );
  OAI211_X1 U19515 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17651), .A(n17650), .B(
        n17649), .ZN(n17652) );
  OAI211_X1 U19516 ( .C1(n20590), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        P3_U2686) );
  NOR2_X1 U19517 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20071) );
  AOI21_X1 U19518 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n20071), .ZN(n20060) );
  INV_X1 U19519 ( .A(n20060), .ZN(n17656) );
  INV_X1 U19520 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20065) );
  OAI222_X1 U19521 ( .A1(n17656), .A2(n17660), .B1(n20065), .B2(n17655), .C1(
        n17712), .C2(n17654), .ZN(P3_U2702) );
  AOI22_X1 U19522 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17658), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17657), .ZN(n17659) );
  OAI21_X1 U19523 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17660), .A(n17659), .ZN(
        P3_U2703) );
  OAI21_X1 U19524 ( .B1(n21158), .B2(n20013), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17661) );
  OAI21_X1 U19525 ( .B1(n17824), .B2(n20057), .A(n17661), .ZN(P3_U2634) );
  OAI21_X1 U19526 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17663), .A(n17662), .ZN(
        n17664) );
  INV_X1 U19527 ( .A(n17664), .ZN(n21213) );
  INV_X1 U19528 ( .A(n18709), .ZN(n18695) );
  OAI21_X1 U19529 ( .B1(n21213), .B2(n18695), .A(n18231), .ZN(n17665) );
  OAI221_X1 U19530 ( .B1(n21166), .B2(n17666), .C1(n21166), .C2(n18231), .A(
        n17665), .ZN(P3_U2863) );
  AOI22_X1 U19531 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17670) );
  AOI22_X1 U19532 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17669) );
  AOI22_X1 U19533 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U19534 ( .A1(n10970), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17667) );
  NAND4_X1 U19535 ( .A1(n17670), .A2(n17669), .A3(n17668), .A4(n17667), .ZN(
        n17676) );
  AOI22_X1 U19536 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U19537 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U19538 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17672) );
  AOI22_X1 U19539 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17671) );
  NAND4_X1 U19540 ( .A1(n17674), .A2(n17673), .A3(n17672), .A4(n17671), .ZN(
        n17675) );
  AOI22_X1 U19541 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U19542 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U19543 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U19544 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17677) );
  NAND4_X1 U19545 ( .A1(n17680), .A2(n17679), .A3(n17678), .A4(n17677), .ZN(
        n17686) );
  AOI22_X1 U19546 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17684) );
  AOI22_X1 U19547 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17683) );
  AOI22_X1 U19548 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10993), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U19549 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17681) );
  NAND4_X1 U19550 ( .A1(n17684), .A2(n17683), .A3(n17682), .A4(n17681), .ZN(
        n17685) );
  AOI22_X1 U19551 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U19552 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U19553 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17689) );
  AOI22_X1 U19554 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17688) );
  NAND4_X1 U19555 ( .A1(n17691), .A2(n17690), .A3(n17689), .A4(n17688), .ZN(
        n17697) );
  AOI22_X1 U19556 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17695) );
  AOI22_X1 U19557 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17694) );
  AOI22_X1 U19558 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U19559 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17692) );
  NAND4_X1 U19560 ( .A1(n17695), .A2(n17694), .A3(n17693), .A4(n17692), .ZN(
        n17696) );
  NOR2_X1 U19561 ( .A1(n17697), .A2(n17696), .ZN(n17791) );
  INV_X1 U19562 ( .A(n17791), .ZN(n20544) );
  AOI22_X1 U19563 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U19564 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17709) );
  AOI22_X1 U19565 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17698) );
  OAI21_X1 U19566 ( .B1(n11024), .B2(n17699), .A(n17698), .ZN(n17707) );
  AOI22_X1 U19567 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17705) );
  AOI22_X1 U19568 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U19569 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U19570 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17702) );
  NAND4_X1 U19571 ( .A1(n17705), .A2(n17704), .A3(n17703), .A4(n17702), .ZN(
        n17706) );
  AOI211_X1 U19572 ( .C1(n10994), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17707), .B(n17706), .ZN(n17708) );
  AOI22_X1 U19573 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17764), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17721) );
  AOI22_X1 U19574 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17735), .ZN(n17720) );
  AOI22_X1 U19575 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10969), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17737), .ZN(n17711) );
  OAI21_X1 U19576 ( .B1(n17712), .B2(n11024), .A(n17711), .ZN(n17718) );
  AOI22_X1 U19577 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U19578 ( .A1(n10984), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17722), .ZN(n17715) );
  AOI22_X1 U19579 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n15077), .ZN(n17714) );
  AOI22_X1 U19580 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17713) );
  NAND4_X1 U19581 ( .A1(n17716), .A2(n17715), .A3(n17714), .A4(n17713), .ZN(
        n17717) );
  AOI211_X1 U19582 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n10977), .A(
        n17718), .B(n17717), .ZN(n17719) );
  NAND3_X1 U19583 ( .A1(n17721), .A2(n17720), .A3(n17719), .ZN(n17790) );
  AOI22_X1 U19584 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U19585 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17733) );
  AOI22_X1 U19586 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17724) );
  OAI21_X1 U19587 ( .B1(n11024), .B2(n17725), .A(n17724), .ZN(n17731) );
  AOI22_X1 U19588 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17729) );
  AOI22_X1 U19589 ( .A1(n17764), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17728) );
  AOI22_X1 U19590 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17727) );
  AOI22_X1 U19591 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17726) );
  NAND4_X1 U19592 ( .A1(n17729), .A2(n17728), .A3(n17727), .A4(n17726), .ZN(
        n17730) );
  AOI211_X1 U19593 ( .C1(n17736), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n17731), .B(n17730), .ZN(n17732) );
  NAND3_X1 U19594 ( .A1(n17734), .A2(n17733), .A3(n17732), .ZN(n17804) );
  NAND2_X1 U19595 ( .A1(n17756), .A2(n17804), .ZN(n17755) );
  AOI22_X1 U19596 ( .A1(n17735), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U19597 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10993), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U19598 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17738) );
  OAI21_X1 U19599 ( .B1(n11024), .B2(n17739), .A(n17738), .ZN(n17748) );
  AOI22_X1 U19600 ( .A1(n17740), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U19601 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17741), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17745) );
  AOI22_X1 U19602 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17744) );
  AOI22_X1 U19603 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17743) );
  NAND4_X1 U19604 ( .A1(n17746), .A2(n17745), .A3(n17744), .A4(n17743), .ZN(
        n17747) );
  AOI211_X1 U19605 ( .C1(n15079), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17748), .B(n17747), .ZN(n17749) );
  NAND3_X1 U19606 ( .A1(n17751), .A2(n17750), .A3(n17749), .ZN(n17789) );
  AOI21_X1 U19607 ( .B1(n21021), .B2(n17752), .A(n18099), .ZN(n17780) );
  XOR2_X1 U19608 ( .A(n17789), .B(n17753), .Z(n17754) );
  NAND2_X1 U19609 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17754), .ZN(
        n17779) );
  XOR2_X1 U19610 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n17754), .Z(
        n18153) );
  INV_X1 U19611 ( .A(n20535), .ZN(n17793) );
  XNOR2_X1 U19612 ( .A(n17793), .B(n17755), .ZN(n17776) );
  XOR2_X1 U19613 ( .A(n17804), .B(n17756), .Z(n17757) );
  NAND2_X1 U19614 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17757), .ZN(
        n17775) );
  XOR2_X1 U19615 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n17757), .Z(
        n18174) );
  INV_X1 U19616 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20789) );
  OR2_X1 U19617 ( .A1(n20789), .A2(n17758), .ZN(n17772) );
  INV_X1 U19618 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20783) );
  AOI22_X1 U19619 ( .A1(n15079), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17763) );
  AOI22_X1 U19620 ( .A1(n17742), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17740), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17762) );
  AOI22_X1 U19621 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17735), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U19622 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17687), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17760) );
  NAND4_X1 U19623 ( .A1(n17763), .A2(n17762), .A3(n17761), .A4(n17760), .ZN(
        n17771) );
  AOI22_X1 U19624 ( .A1(n17736), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U19625 ( .A1(n10993), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10969), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17768) );
  AOI22_X1 U19626 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17764), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U19627 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17765), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17766) );
  NAND4_X1 U19628 ( .A1(n17769), .A2(n17768), .A3(n17767), .A4(n17766), .ZN(
        n17770) );
  NOR2_X1 U19629 ( .A1(n17771), .A2(n17770), .ZN(n20672) );
  INV_X1 U19630 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20862) );
  NOR2_X1 U19631 ( .A1(n20672), .A2(n20862), .ZN(n18220) );
  XNOR2_X1 U19632 ( .A(n17790), .B(n20783), .ZN(n18213) );
  INV_X1 U19633 ( .A(n18213), .ZN(n18211) );
  NAND2_X1 U19634 ( .A1(n18220), .A2(n18211), .ZN(n18210) );
  OAI21_X1 U19635 ( .B1(n20783), .B2(n17790), .A(n18210), .ZN(n18203) );
  NAND2_X1 U19636 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17773), .ZN(
        n17774) );
  INV_X1 U19637 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20795) );
  XNOR2_X1 U19638 ( .A(n20795), .B(n17773), .ZN(n18193) );
  XOR2_X1 U19639 ( .A(n20544), .B(n17796), .Z(n18192) );
  NAND2_X1 U19640 ( .A1(n18193), .A2(n18192), .ZN(n18191) );
  NAND2_X1 U19641 ( .A1(n17776), .A2(n17777), .ZN(n17778) );
  NAND2_X1 U19642 ( .A1(n17780), .A2(n17852), .ZN(n17781) );
  NAND2_X1 U19643 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18141), .ZN(
        n18140) );
  NAND2_X1 U19644 ( .A1(n20738), .A2(n17782), .ZN(n20689) );
  AOI21_X1 U19645 ( .B1(n17787), .B2(n17786), .A(n20741), .ZN(n21180) );
  NAND2_X2 U19646 ( .A1(n21224), .A2(n20738), .ZN(n18225) );
  NOR2_X4 U19647 ( .A1(n20749), .A2(n18225), .ZN(n18129) );
  INV_X1 U19648 ( .A(n17789), .ZN(n20531) );
  INV_X1 U19649 ( .A(n20672), .ZN(n17798) );
  NAND2_X1 U19650 ( .A1(n17790), .A2(n17798), .ZN(n17799) );
  NAND2_X1 U19651 ( .A1(n20550), .A2(n17799), .ZN(n17794) );
  NOR2_X1 U19652 ( .A1(n17791), .A2(n17795), .ZN(n17805) );
  NAND2_X1 U19653 ( .A1(n17792), .A2(n17793), .ZN(n17811) );
  NOR2_X1 U19654 ( .A1(n20531), .A2(n17811), .ZN(n17815) );
  NAND2_X1 U19655 ( .A1(n17815), .A2(n20749), .ZN(n17816) );
  XOR2_X1 U19656 ( .A(n17793), .B(n17792), .Z(n17809) );
  AND2_X1 U19657 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17809), .ZN(
        n17810) );
  XNOR2_X1 U19658 ( .A(n20544), .B(n17794), .ZN(n17802) );
  NOR2_X1 U19659 ( .A1(n20795), .A2(n17802), .ZN(n17803) );
  NOR2_X1 U19660 ( .A1(n17797), .A2(n20789), .ZN(n17801) );
  NAND2_X1 U19661 ( .A1(n20669), .A2(n20783), .ZN(n17800) );
  NOR2_X1 U19662 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17798), .ZN(
        n18219) );
  NAND2_X1 U19663 ( .A1(n18213), .A2(n18219), .ZN(n18212) );
  NAND3_X1 U19664 ( .A1(n17800), .A2(n17799), .A3(n18212), .ZN(n18200) );
  NOR2_X1 U19665 ( .A1(n17801), .A2(n18199), .ZN(n18190) );
  XOR2_X1 U19666 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n17802), .Z(
        n18189) );
  NOR2_X1 U19667 ( .A1(n18190), .A2(n18189), .ZN(n18188) );
  INV_X1 U19668 ( .A(n17804), .ZN(n20540) );
  XOR2_X1 U19669 ( .A(n20540), .B(n17805), .Z(n17807) );
  NOR2_X1 U19670 ( .A1(n17806), .A2(n17807), .ZN(n17808) );
  INV_X1 U19671 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20814) );
  INV_X1 U19672 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20823) );
  XOR2_X1 U19673 ( .A(n20823), .B(n17809), .Z(n18162) );
  NOR2_X1 U19674 ( .A1(n18163), .A2(n18162), .ZN(n18161) );
  NOR2_X1 U19675 ( .A1(n17810), .A2(n18161), .ZN(n17812) );
  XNOR2_X1 U19676 ( .A(n20531), .B(n17811), .ZN(n17813) );
  NOR2_X1 U19677 ( .A1(n17812), .A2(n17813), .ZN(n17814) );
  INV_X1 U19678 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20839) );
  XNOR2_X1 U19679 ( .A(n17813), .B(n17812), .ZN(n18156) );
  NOR2_X1 U19680 ( .A1(n20839), .A2(n18156), .ZN(n18155) );
  OR2_X2 U19681 ( .A1(n17814), .A2(n18155), .ZN(n17817) );
  XOR2_X1 U19682 ( .A(n20749), .B(n17815), .Z(n17818) );
  OR2_X2 U19683 ( .A1(n17817), .A2(n17818), .ZN(n18145) );
  NOR2_X1 U19684 ( .A1(n17816), .A2(n17820), .ZN(n17822) );
  INV_X1 U19685 ( .A(n17816), .ZN(n17821) );
  NAND2_X1 U19686 ( .A1(n17818), .A2(n17817), .ZN(n18146) );
  OAI21_X1 U19687 ( .B1(n17821), .B2(n17820), .A(n18146), .ZN(n17819) );
  AOI21_X1 U19688 ( .B1(n17821), .B2(n17820), .A(n17819), .ZN(n18131) );
  INV_X1 U19689 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20850) );
  NOR2_X2 U19690 ( .A1(n18131), .A2(n20850), .ZN(n18130) );
  AOI22_X2 U19691 ( .A1(n20750), .A2(n18129), .B1(n18214), .B2(n20859), .ZN(
        n18125) );
  INV_X1 U19692 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20903) );
  NOR2_X1 U19693 ( .A1(n21149), .A2(n18104), .ZN(n18083) );
  NAND3_X1 U19694 ( .A1(n18083), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20877) );
  NAND2_X1 U19695 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20876), .ZN(
        n20892) );
  NOR2_X1 U19696 ( .A1(n20903), .A2(n20892), .ZN(n20908) );
  INV_X1 U19697 ( .A(n20908), .ZN(n20911) );
  NOR2_X1 U19698 ( .A1(n20924), .A2(n20911), .ZN(n21083) );
  INV_X1 U19699 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21101) );
  NOR2_X1 U19700 ( .A1(n21109), .A2(n21101), .ZN(n21089) );
  INV_X1 U19701 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21095) );
  NAND2_X1 U19702 ( .A1(n21089), .A2(n21095), .ZN(n21100) );
  NAND2_X1 U19703 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18177) );
  NAND2_X1 U19704 ( .A1(n18181), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20103) );
  NAND3_X1 U19705 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18116) );
  NAND2_X1 U19706 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20265) );
  NOR2_X1 U19707 ( .A1(n17823), .A2(n20067), .ZN(n20288) );
  AOI21_X1 U19708 ( .B1(n17849), .B2(n17823), .A(n18195), .ZN(n18060) );
  OAI21_X1 U19709 ( .B1(n20288), .B2(n18222), .A(n18060), .ZN(n17840) );
  AOI21_X1 U19710 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17975), .A(
        n19012), .ZN(n18020) );
  NOR3_X1 U19711 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18020), .A3(
        n17823), .ZN(n17841) );
  INV_X1 U19712 ( .A(n20288), .ZN(n18055) );
  INV_X1 U19713 ( .A(n20312), .ZN(n17838) );
  NOR2_X1 U19714 ( .A1(n17838), .A2(n20067), .ZN(n17839) );
  AOI21_X1 U19715 ( .B1(n20305), .B2(n18055), .A(n17839), .ZN(n20302) );
  INV_X1 U19716 ( .A(n20302), .ZN(n20300) );
  OR2_X2 U19717 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17824), .ZN(n21129) );
  INV_X2 U19718 ( .A(n21129), .ZN(n21156) );
  NAND2_X1 U19719 ( .A1(n21156), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n21098) );
  OAI21_X1 U19720 ( .B1(n18003), .B2(n20300), .A(n21098), .ZN(n17825) );
  AOI211_X1 U19721 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17840), .A(
        n17841), .B(n17825), .ZN(n17834) );
  INV_X1 U19722 ( .A(n18129), .ZN(n18077) );
  NOR2_X1 U19723 ( .A1(n20863), .A2(n20892), .ZN(n18075) );
  NAND2_X1 U19724 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18075), .ZN(
        n20917) );
  OAI22_X1 U19725 ( .A1(n18077), .A2(n20915), .B1(n18226), .B2(n21084), .ZN(
        n17826) );
  INV_X1 U19726 ( .A(n17826), .ZN(n17869) );
  OAI21_X1 U19727 ( .B1(n21089), .B2(n17870), .A(n17869), .ZN(n18063) );
  NAND2_X1 U19728 ( .A1(n21034), .A2(n21095), .ZN(n17835) );
  AOI21_X1 U19729 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18099), .A(
        n17913), .ZN(n17832) );
  NAND2_X1 U19730 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21034), .ZN(
        n17827) );
  AOI22_X1 U19731 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21034), .B1(
        n18099), .B2(n20850), .ZN(n18128) );
  INV_X1 U19732 ( .A(n17828), .ZN(n18101) );
  INV_X1 U19733 ( .A(n21083), .ZN(n20755) );
  INV_X1 U19734 ( .A(n17830), .ZN(n17829) );
  NAND2_X1 U19735 ( .A1(n21149), .A2(n18104), .ZN(n18107) );
  NOR4_X1 U19736 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(n18107), .ZN(n18072) );
  NOR2_X1 U19737 ( .A1(n17831), .A2(n17830), .ZN(n17951) );
  INV_X1 U19738 ( .A(n17951), .ZN(n17862) );
  NAND2_X1 U19739 ( .A1(n21089), .A2(n17862), .ZN(n17836) );
  XNOR2_X1 U19740 ( .A(n17832), .B(n17891), .ZN(n21097) );
  AOI22_X1 U19741 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18063), .B1(
        n18122), .B2(n21097), .ZN(n17833) );
  OAI211_X1 U19742 ( .C1(n17870), .C2(n21100), .A(n17834), .B(n17833), .ZN(
        P3_U2812) );
  NAND2_X1 U19743 ( .A1(n21089), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17890) );
  INV_X1 U19744 ( .A(n17890), .ZN(n20752) );
  NAND2_X1 U19745 ( .A1(n20752), .A2(n18064), .ZN(n17915) );
  INV_X1 U19746 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17912) );
  NOR2_X1 U19747 ( .A1(n17890), .A2(n17912), .ZN(n20756) );
  NAND2_X1 U19748 ( .A1(n20915), .A2(n20756), .ZN(n21064) );
  NAND2_X1 U19749 ( .A1(n21084), .A2(n20756), .ZN(n21063) );
  AOI22_X1 U19750 ( .A1(n18129), .A2(n21064), .B1(n18214), .B2(n21063), .ZN(
        n17917) );
  NOR2_X1 U19751 ( .A1(n17835), .A2(n17891), .ZN(n17901) );
  NOR3_X1 U19752 ( .A1(n21034), .A2(n21095), .A3(n17836), .ZN(n17911) );
  NOR2_X1 U19753 ( .A1(n17901), .A2(n17911), .ZN(n17837) );
  XOR2_X1 U19754 ( .A(n17837), .B(n17912), .Z(n21071) );
  NOR3_X1 U19755 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18020), .A3(
        n17838), .ZN(n17844) );
  NAND2_X1 U19756 ( .A1(n20312), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17893) );
  INV_X1 U19757 ( .A(n17893), .ZN(n20330) );
  NAND2_X1 U19758 ( .A1(n20330), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17920) );
  OAI21_X1 U19759 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17839), .A(
        n17920), .ZN(n20314) );
  NAND2_X1 U19760 ( .A1(n21156), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21072) );
  OAI21_X1 U19761 ( .B1(n17841), .B2(n17840), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17842) );
  OAI211_X1 U19762 ( .C1(n18003), .C2(n20314), .A(n21072), .B(n17842), .ZN(
        n17843) );
  AOI211_X1 U19763 ( .C1(n18122), .C2(n21071), .A(n17844), .B(n17843), .ZN(
        n17845) );
  OAI221_X1 U19764 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17915), 
        .C1(n17912), .C2(n17917), .A(n17845), .ZN(P3_U2811) );
  NOR2_X1 U19765 ( .A1(n17846), .A2(n18226), .ZN(n17847) );
  AOI21_X1 U19766 ( .B1(n20908), .B2(n17847), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17860) );
  NOR2_X1 U19767 ( .A1(n18020), .A2(n17848), .ZN(n17864) );
  INV_X1 U19768 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17851) );
  NOR2_X1 U19769 ( .A1(n17848), .A2(n20067), .ZN(n18069) );
  AOI21_X1 U19770 ( .B1(n17849), .B2(n17848), .A(n18195), .ZN(n18081) );
  OAI21_X1 U19771 ( .B1(n18069), .B2(n18222), .A(n18081), .ZN(n17863) );
  INV_X1 U19772 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20280) );
  NAND2_X1 U19773 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18069), .ZN(
        n20268) );
  OAI21_X1 U19774 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18069), .A(
        n20268), .ZN(n20257) );
  OAI22_X1 U19775 ( .A1(n21129), .A2(n20280), .B1(n18003), .B2(n20257), .ZN(
        n17850) );
  AOI221_X1 U19776 ( .B1(n17864), .B2(n17851), .C1(n17863), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17850), .ZN(n17859) );
  INV_X1 U19777 ( .A(n20917), .ZN(n17857) );
  NOR2_X1 U19778 ( .A1(n20915), .A2(n18077), .ZN(n17856) );
  NAND4_X1 U19779 ( .A1(n18099), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n17852), .ZN(n18112) );
  NOR2_X1 U19780 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17853), .ZN(
        n18071) );
  NAND3_X1 U19781 ( .A1(n18072), .A2(n18071), .A3(n20903), .ZN(n17854) );
  OAI21_X1 U19782 ( .B1(n20911), .B2(n18112), .A(n17854), .ZN(n17855) );
  XOR2_X1 U19783 ( .A(n17855), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n20910) );
  AOI22_X1 U19784 ( .A1(n17857), .A2(n17856), .B1(n18122), .B2(n20910), .ZN(
        n17858) );
  OAI211_X1 U19785 ( .C1(n17869), .C2(n17860), .A(n17859), .B(n17858), .ZN(
        P3_U2815) );
  AOI22_X1 U19786 ( .A1(n18099), .A2(n21109), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21034), .ZN(n17861) );
  XOR2_X1 U19787 ( .A(n17862), .B(n17861), .Z(n21114) );
  INV_X1 U19788 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20281) );
  NOR2_X1 U19789 ( .A1(n21129), .A2(n20281), .ZN(n21113) );
  INV_X1 U19790 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20279) );
  AND2_X1 U19791 ( .A1(n18059), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18056) );
  AOI21_X1 U19792 ( .B1(n20279), .B2(n20268), .A(n18056), .ZN(n20275) );
  AOI22_X1 U19793 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17863), .B1(
        n18050), .B2(n20275), .ZN(n17866) );
  OAI211_X1 U19794 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17864), .B(n20265), .ZN(n17865) );
  NAND2_X1 U19795 ( .A1(n17866), .A2(n17865), .ZN(n17867) );
  AOI211_X1 U19796 ( .C1(n18122), .C2(n21114), .A(n21113), .B(n17867), .ZN(
        n17868) );
  OAI221_X1 U19797 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17870), 
        .C1(n21109), .C2(n17869), .A(n17868), .ZN(P3_U2814) );
  OAI22_X1 U19798 ( .A1(n20750), .A2(n18077), .B1(n18226), .B2(n20859), .ZN(
        n18089) );
  INV_X1 U19799 ( .A(n18089), .ZN(n18124) );
  OAI21_X1 U19800 ( .B1(n20876), .B2(n18125), .A(n18124), .ZN(n17887) );
  INV_X1 U19801 ( .A(n17887), .ZN(n17878) );
  INV_X1 U19802 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20889) );
  INV_X1 U19803 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20225) );
  NAND2_X1 U19804 ( .A1(n18067), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17872) );
  INV_X1 U19805 ( .A(n17872), .ZN(n18084) );
  NAND2_X1 U19806 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18084), .ZN(
        n20226) );
  INV_X1 U19807 ( .A(n20226), .ZN(n17883) );
  AOI21_X1 U19808 ( .B1(n20225), .B2(n17872), .A(n17883), .ZN(n20220) );
  NAND2_X1 U19809 ( .A1(n18067), .A2(n17976), .ZN(n17882) );
  OAI21_X1 U19810 ( .B1(n18067), .B2(n18180), .A(n18222), .ZN(n17871) );
  AOI21_X1 U19811 ( .B1(n17872), .B2(n17871), .A(n18195), .ZN(n17884) );
  NAND2_X1 U19812 ( .A1(n21156), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n20884) );
  OAI221_X1 U19813 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17882), .C1(
        n20225), .C2(n17884), .A(n20884), .ZN(n17873) );
  AOI21_X1 U19814 ( .B1(n18050), .B2(n20220), .A(n17873), .ZN(n17877) );
  INV_X1 U19815 ( .A(n18071), .ZN(n18113) );
  NOR3_X1 U19816 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18107), .A3(
        n18113), .ZN(n17879) );
  NAND2_X1 U19817 ( .A1(n18083), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20873) );
  NOR2_X1 U19818 ( .A1(n18112), .A2(n20873), .ZN(n17880) );
  NOR2_X1 U19819 ( .A1(n17879), .A2(n17880), .ZN(n17874) );
  XOR2_X1 U19820 ( .A(n17874), .B(n20889), .Z(n20883) );
  INV_X1 U19821 ( .A(n20873), .ZN(n20860) );
  NOR2_X1 U19822 ( .A1(n20876), .A2(n18125), .ZN(n17875) );
  AOI22_X1 U19823 ( .A1(n18122), .A2(n20883), .B1(n20860), .B2(n17875), .ZN(
        n17876) );
  OAI211_X1 U19824 ( .C1(n17878), .C2(n20889), .A(n17877), .B(n17876), .ZN(
        P3_U2818) );
  AOI22_X1 U19825 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17880), .B1(
        n17879), .B2(n20889), .ZN(n17881) );
  XOR2_X1 U19826 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17881), .Z(
        n21124) );
  INV_X1 U19827 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20230) );
  AOI221_X1 U19828 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C1(n20225), .C2(n20230), .A(
        n17882), .ZN(n17886) );
  NAND2_X1 U19829 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17883), .ZN(
        n20243) );
  OAI21_X1 U19830 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17883), .A(
        n20243), .ZN(n20228) );
  OAI22_X1 U19831 ( .A1(n17884), .A2(n20230), .B1(n18003), .B2(n20228), .ZN(
        n17885) );
  AOI211_X1 U19832 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n21156), .A(n17886), 
        .B(n17885), .ZN(n17889) );
  NOR2_X1 U19833 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20877), .ZN(
        n21117) );
  AOI22_X1 U19834 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17887), .B1(
        n21117), .B2(n18106), .ZN(n17888) );
  OAI211_X1 U19835 ( .C1(n21124), .C2(n18139), .A(n17889), .B(n17888), .ZN(
        P3_U2817) );
  INV_X1 U19836 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17916) );
  NOR2_X1 U19837 ( .A1(n17916), .A2(n17912), .ZN(n20762) );
  NAND2_X1 U19838 ( .A1(n20762), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n20987) );
  NOR2_X1 U19839 ( .A1(n17890), .A2(n20987), .ZN(n17950) );
  INV_X1 U19840 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21048) );
  NAND2_X1 U19841 ( .A1(n17950), .A2(n20915), .ZN(n21040) );
  NAND2_X1 U19842 ( .A1(n17950), .A2(n21084), .ZN(n21041) );
  AOI22_X1 U19843 ( .A1(n18129), .A2(n21040), .B1(n18214), .B2(n21041), .ZN(
        n17907) );
  NOR2_X1 U19844 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17902) );
  INV_X1 U19845 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20764) );
  NAND3_X1 U19846 ( .A1(n17913), .A2(n17902), .A3(n20764), .ZN(n17927) );
  INV_X1 U19847 ( .A(n20987), .ZN(n20927) );
  INV_X1 U19848 ( .A(n17952), .ZN(n17892) );
  AOI21_X1 U19849 ( .B1(n17927), .B2(n17955), .A(n17892), .ZN(n17928) );
  XOR2_X1 U19850 ( .A(n17928), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n20925) );
  INV_X1 U19851 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17897) );
  INV_X1 U19852 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20346) );
  NAND2_X1 U19853 ( .A1(n17922), .A2(n17976), .ZN(n17906) );
  AOI221_X1 U19854 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n17897), .C2(n20346), .A(
        n17906), .ZN(n17899) );
  AOI21_X1 U19855 ( .B1(n17973), .B2(n17920), .A(n18195), .ZN(n17894) );
  OAI21_X1 U19856 ( .B1(n17922), .B2(n18180), .A(n17894), .ZN(n17919) );
  AOI21_X1 U19857 ( .B1(n17975), .B2(n17921), .A(n17919), .ZN(n17905) );
  NAND3_X1 U19858 ( .A1(n17922), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17895) );
  NOR2_X1 U19859 ( .A1(n17936), .A2(n20067), .ZN(n17930) );
  AOI21_X1 U19860 ( .B1(n17897), .B2(n17895), .A(n17930), .ZN(n20358) );
  AOI22_X1 U19861 ( .A1(n21156), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18050), 
        .B2(n20358), .ZN(n17896) );
  OAI21_X1 U19862 ( .B1(n17905), .B2(n17897), .A(n17896), .ZN(n17898) );
  AOI211_X1 U19863 ( .C1(n20925), .C2(n18122), .A(n17899), .B(n17898), .ZN(
        n17900) );
  OAI221_X1 U19864 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18011), 
        .C1(n21048), .C2(n17907), .A(n17900), .ZN(P3_U2808) );
  AOI22_X1 U19865 ( .A1(n20762), .A2(n17911), .B1(n17902), .B2(n17901), .ZN(
        n17903) );
  XOR2_X1 U19866 ( .A(n17903), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n20754) );
  NAND2_X1 U19867 ( .A1(n17922), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17904) );
  XOR2_X1 U19868 ( .A(n20346), .B(n17904), .Z(n20343) );
  NAND2_X1 U19869 ( .A1(n21156), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n20768) );
  OAI221_X1 U19870 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17906), .C1(
        n20346), .C2(n17905), .A(n20768), .ZN(n17909) );
  NAND2_X1 U19871 ( .A1(n20762), .A2(n20764), .ZN(n20770) );
  OAI22_X1 U19872 ( .A1(n17907), .A2(n20764), .B1(n20770), .B2(n17915), .ZN(
        n17908) );
  AOI211_X1 U19873 ( .C1(n18050), .C2(n20343), .A(n17909), .B(n17908), .ZN(
        n17910) );
  OAI21_X1 U19874 ( .B1(n20754), .B2(n18139), .A(n17910), .ZN(P3_U2809) );
  OAI221_X1 U19875 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17913), 
        .C1(n17912), .C2(n17911), .A(n17952), .ZN(n17914) );
  XOR2_X1 U19876 ( .A(n17916), .B(n17914), .Z(n21074) );
  NAND2_X1 U19877 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17916), .ZN(
        n21082) );
  OAI22_X1 U19878 ( .A1(n17917), .A2(n17916), .B1(n17915), .B2(n21082), .ZN(
        n17918) );
  AOI21_X1 U19879 ( .B1(n18122), .B2(n21074), .A(n17918), .ZN(n17926) );
  NAND2_X1 U19880 ( .A1(n21156), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17925) );
  OAI221_X1 U19881 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20330), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19012), .A(n17919), .ZN(
        n17924) );
  AOI22_X1 U19882 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17922), .B1(
        n17921), .B2(n17920), .ZN(n20332) );
  OAI21_X1 U19883 ( .B1(n18050), .B2(n17975), .A(n20332), .ZN(n17923) );
  NAND4_X1 U19884 ( .A1(n17926), .A2(n17925), .A3(n17924), .A4(n17923), .ZN(
        P3_U2810) );
  NOR2_X1 U19885 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17927), .ZN(
        n17954) );
  OAI221_X1 U19886 ( .B1(n17954), .B2(n18099), .C1(n17954), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17928), .ZN(n17929) );
  XOR2_X1 U19887 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17929), .Z(
        n21053) );
  INV_X1 U19888 ( .A(n17930), .ZN(n17932) );
  OAI21_X1 U19889 ( .B1(n18021), .B2(n17932), .A(n17933), .ZN(n17938) );
  AOI221_X1 U19890 ( .B1(n17933), .B2(n17973), .C1(n17932), .C2(n17973), .A(
        n18195), .ZN(n17931) );
  OAI21_X1 U19891 ( .B1(n11059), .B2(n18965), .A(n17931), .ZN(n17963) );
  INV_X1 U19892 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20367) );
  NOR2_X1 U19893 ( .A1(n21129), .A2(n20367), .ZN(n21050) );
  OR2_X1 U19894 ( .A1(n18965), .A2(n11059), .ZN(n17935) );
  NAND2_X1 U19895 ( .A1(n11059), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17962) );
  NAND2_X1 U19896 ( .A1(n17933), .A2(n17932), .ZN(n17934) );
  NAND2_X1 U19897 ( .A1(n17962), .A2(n17934), .ZN(n20377) );
  OAI22_X1 U19898 ( .A1(n17936), .A2(n17935), .B1(n18003), .B2(n20377), .ZN(
        n17937) );
  AOI211_X1 U19899 ( .C1(n17938), .C2(n17963), .A(n21050), .B(n17937), .ZN(
        n17943) );
  NAND2_X1 U19900 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21054) );
  OAI21_X1 U19901 ( .B1(n21054), .B2(n21041), .A(n18214), .ZN(n17939) );
  OAI21_X1 U19902 ( .B1(n21054), .B2(n21040), .A(n18129), .ZN(n17940) );
  OAI22_X1 U19903 ( .A1(n21041), .A2(n17939), .B1(n21040), .B2(n17940), .ZN(
        n17941) );
  NAND2_X1 U19904 ( .A1(n17940), .A2(n17939), .ZN(n17969) );
  AOI22_X1 U19905 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17941), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17969), .ZN(n17942) );
  OAI211_X1 U19906 ( .C1(n18139), .C2(n21053), .A(n17943), .B(n17942), .ZN(
        P3_U2807) );
  INV_X1 U19907 ( .A(n21041), .ZN(n20759) );
  INV_X1 U19908 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17944) );
  NOR2_X1 U19909 ( .A1(n17944), .A2(n21054), .ZN(n20936) );
  NAND2_X1 U19910 ( .A1(n20759), .A2(n20936), .ZN(n17945) );
  XOR2_X1 U19911 ( .A(n17945), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n20947) );
  INV_X1 U19912 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20403) );
  NOR2_X1 U19913 ( .A1(n21129), .A2(n20403), .ZN(n20949) );
  NOR2_X1 U19914 ( .A1(n11317), .A2(n11318), .ZN(n17947) );
  OAI211_X1 U19915 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n11059), .B(n17976), .ZN(n17946) );
  NOR2_X1 U19916 ( .A1(n11318), .A2(n17962), .ZN(n17961) );
  OAI22_X1 U19917 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17961), .B1(
        n20067), .B2(n18006), .ZN(n20389) );
  OAI22_X1 U19918 ( .A1(n17947), .A2(n17946), .B1(n20389), .B2(n18003), .ZN(
        n17948) );
  AOI211_X1 U19919 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17963), .A(
        n20949), .B(n17948), .ZN(n17958) );
  INV_X1 U19920 ( .A(n21040), .ZN(n17980) );
  NAND2_X1 U19921 ( .A1(n17980), .A2(n20936), .ZN(n17949) );
  INV_X1 U19922 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20937) );
  XOR2_X1 U19923 ( .A(n17949), .B(n20937), .Z(n20944) );
  NAND2_X1 U19924 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17950), .ZN(
        n20938) );
  OAI21_X1 U19925 ( .B1(n17951), .B2(n20938), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17953) );
  OAI21_X1 U19926 ( .B1(n21034), .B2(n18009), .A(n11030), .ZN(n17956) );
  XOR2_X1 U19927 ( .A(n17956), .B(n20937), .Z(n20945) );
  AOI22_X1 U19928 ( .A1(n18129), .A2(n20944), .B1(n18122), .B2(n20945), .ZN(
        n17957) );
  OAI211_X1 U19929 ( .C1(n20947), .C2(n18226), .A(n17958), .B(n17957), .ZN(
        P3_U2805) );
  AOI21_X1 U19930 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17960), .A(
        n17959), .ZN(n21062) );
  AOI21_X1 U19931 ( .B1(n11318), .B2(n17962), .A(n17961), .ZN(n20379) );
  NAND2_X1 U19932 ( .A1(n11059), .A2(n17976), .ZN(n17966) );
  INV_X1 U19933 ( .A(n17963), .ZN(n17965) );
  NAND2_X1 U19934 ( .A1(n21156), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17964) );
  OAI221_X1 U19935 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17966), .C1(
        n11318), .C2(n17965), .A(n17964), .ZN(n17967) );
  AOI21_X1 U19936 ( .B1(n18050), .B2(n20379), .A(n17967), .ZN(n17971) );
  NOR2_X1 U19937 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21054), .ZN(
        n17968) );
  AOI22_X1 U19938 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17969), .B1(
        n17981), .B2(n17968), .ZN(n17970) );
  OAI211_X1 U19939 ( .C1(n21062), .C2(n18139), .A(n17971), .B(n17970), .ZN(
        P3_U2806) );
  INV_X1 U19940 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17977) );
  NAND2_X1 U19941 ( .A1(n17972), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17993) );
  NAND2_X1 U19942 ( .A1(n18053), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18044) );
  INV_X1 U19943 ( .A(n18044), .ZN(n18024) );
  AOI21_X1 U19944 ( .B1(n17977), .B2(n17993), .A(n18024), .ZN(n20436) );
  AND3_X1 U19945 ( .A1(n17977), .A2(n17976), .A3(n17972), .ZN(n17979) );
  OAI21_X1 U19946 ( .B1(n18006), .B2(n20067), .A(n17973), .ZN(n17974) );
  OAI211_X1 U19947 ( .C1(n17992), .C2(n18180), .A(n17974), .B(n18221), .ZN(
        n18008) );
  AOI21_X1 U19948 ( .B1(n17975), .B2(n20417), .A(n18008), .ZN(n18002) );
  INV_X1 U19949 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20423) );
  NAND3_X1 U19950 ( .A1(n17992), .A2(n20423), .A3(n17976), .ZN(n17995) );
  NAND2_X1 U19951 ( .A1(n21156), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21038) );
  OAI221_X1 U19952 ( .B1(n17977), .B2(n18002), .C1(n17977), .C2(n17995), .A(
        n21038), .ZN(n17978) );
  AOI211_X1 U19953 ( .C1(n18050), .C2(n20436), .A(n17979), .B(n17978), .ZN(
        n17989) );
  INV_X1 U19954 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20960) );
  NOR2_X1 U19955 ( .A1(n20960), .A2(n20937), .ZN(n17983) );
  AND2_X1 U19956 ( .A1(n20936), .A2(n17983), .ZN(n18018) );
  NAND2_X1 U19957 ( .A1(n20759), .A2(n18018), .ZN(n20954) );
  NAND2_X1 U19958 ( .A1(n18018), .A2(n17980), .ZN(n20956) );
  AOI22_X1 U19959 ( .A1(n18214), .A2(n20954), .B1(n18129), .B2(n20956), .ZN(
        n18012) );
  NAND2_X1 U19960 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18012), .ZN(
        n17998) );
  OAI211_X1 U19961 ( .C1(n18129), .C2(n18214), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17998), .ZN(n17988) );
  INV_X1 U19962 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21031) );
  NAND2_X1 U19963 ( .A1(n18018), .A2(n17981), .ZN(n18037) );
  NOR2_X1 U19964 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18099), .ZN(
        n18046) );
  AOI21_X1 U19965 ( .B1(n18099), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18046), .ZN(n21036) );
  AOI21_X1 U19966 ( .B1(n20960), .B2(n20937), .A(n18099), .ZN(n17982) );
  NAND2_X1 U19967 ( .A1(n17984), .A2(n21031), .ZN(n21037) );
  NAND2_X1 U19968 ( .A1(n21036), .A2(n17985), .ZN(n21018) );
  OAI211_X1 U19969 ( .C1(n21036), .C2(n17985), .A(n18122), .B(n21018), .ZN(
        n17986) );
  NAND4_X1 U19970 ( .A1(n17989), .A2(n17988), .A3(n17987), .A4(n17986), .ZN(
        P3_U2802) );
  OAI21_X1 U19971 ( .B1(n18099), .B2(n17991), .A(n17990), .ZN(n20973) );
  NAND2_X1 U19972 ( .A1(n17992), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18004) );
  INV_X1 U19973 ( .A(n17993), .ZN(n17994) );
  AOI21_X1 U19974 ( .B1(n20423), .B2(n18004), .A(n17994), .ZN(n20422) );
  INV_X1 U19975 ( .A(n20422), .ZN(n17996) );
  NAND2_X1 U19976 ( .A1(n21156), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n20974) );
  OAI211_X1 U19977 ( .C1(n18003), .C2(n17996), .A(n20974), .B(n17995), .ZN(
        n17997) );
  AOI21_X1 U19978 ( .B1(n18122), .B2(n20973), .A(n17997), .ZN(n18001) );
  INV_X1 U19979 ( .A(n18037), .ZN(n17999) );
  OAI21_X1 U19980 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17999), .A(
        n17998), .ZN(n18000) );
  OAI211_X1 U19981 ( .C1(n18002), .C2(n20423), .A(n18001), .B(n18000), .ZN(
        P3_U2803) );
  NOR2_X1 U19982 ( .A1(n18006), .A2(n20067), .ZN(n18005) );
  OAI21_X1 U19983 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18005), .A(
        n18004), .ZN(n20409) );
  OAI21_X1 U19984 ( .B1(n18006), .B2(n18965), .A(n20417), .ZN(n18007) );
  AOI22_X1 U19985 ( .A1(n21156), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18008), 
        .B2(n18007), .ZN(n18017) );
  OAI221_X1 U19986 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21034), 
        .C1(n20937), .C2(n18009), .A(n11030), .ZN(n18010) );
  XOR2_X1 U19987 ( .A(n20960), .B(n18010), .Z(n20952) );
  NAND2_X1 U19988 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n20936), .ZN(
        n20953) );
  NOR2_X1 U19989 ( .A1(n20953), .A2(n18011), .ZN(n18014) );
  INV_X1 U19990 ( .A(n18012), .ZN(n18013) );
  MUX2_X1 U19991 ( .A(n18014), .B(n18013), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n18015) );
  AOI21_X1 U19992 ( .B1(n18122), .B2(n20952), .A(n18015), .ZN(n18016) );
  OAI211_X1 U19993 ( .C1(n18205), .C2(n20409), .A(n18017), .B(n18016), .ZN(
        P3_U2804) );
  INV_X1 U19994 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20684) );
  NAND3_X1 U19995 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n18018), .ZN(n20986) );
  NOR2_X2 U19996 ( .A1(n21041), .A2(n20986), .ZN(n21027) );
  NAND3_X1 U19997 ( .A1(n21027), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n18019) );
  XNOR2_X1 U19998 ( .A(n20684), .B(n18019), .ZN(n21017) );
  INV_X1 U19999 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20485) );
  INV_X1 U20000 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20477) );
  NOR2_X1 U20001 ( .A1(n21129), .A2(n20477), .ZN(n21003) );
  OR2_X1 U20002 ( .A1(n18022), .A2(n18020), .ZN(n18036) );
  XNOR2_X1 U20003 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18025) );
  NOR2_X1 U20004 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18021), .ZN(
        n18051) );
  AOI21_X1 U20005 ( .B1(n19012), .B2(n18022), .A(n18195), .ZN(n18023) );
  OAI21_X1 U20006 ( .B1(n18024), .B2(n18222), .A(n18023), .ZN(n18052) );
  NOR2_X1 U20007 ( .A1(n18051), .A2(n18052), .ZN(n18035) );
  OAI22_X1 U20008 ( .A1(n18036), .A2(n18025), .B1(n18035), .B2(n20485), .ZN(
        n18026) );
  AOI211_X1 U20009 ( .C1(n20269), .C2(n18050), .A(n21003), .B(n18026), .ZN(
        n18031) );
  NAND3_X1 U20010 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n20995) );
  NOR2_X1 U20011 ( .A1(n20956), .A2(n20995), .ZN(n18038) );
  NAND2_X1 U20012 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18038), .ZN(
        n18027) );
  XOR2_X1 U20013 ( .A(n20684), .B(n18027), .Z(n21008) );
  NAND2_X1 U20014 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18099), .ZN(
        n18028) );
  NOR2_X1 U20015 ( .A1(n11033), .A2(n18028), .ZN(n21020) );
  NAND2_X1 U20016 ( .A1(n21020), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18032) );
  INV_X1 U20017 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21004) );
  NAND3_X1 U20018 ( .A1(n18046), .A2(n18045), .A3(n21004), .ZN(n18033) );
  INV_X1 U20019 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21005) );
  AOI22_X1 U20020 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18032), .B1(
        n18033), .B2(n21005), .ZN(n18029) );
  XNOR2_X1 U20021 ( .A(n20684), .B(n18029), .ZN(n21012) );
  AOI22_X1 U20022 ( .A1(n21008), .A2(n18129), .B1(n18122), .B2(n21012), .ZN(
        n18030) );
  OAI211_X1 U20023 ( .C1(n21017), .C2(n18226), .A(n18031), .B(n18030), .ZN(
        P3_U2799) );
  NAND2_X1 U20024 ( .A1(n18033), .A2(n18032), .ZN(n18034) );
  XOR2_X1 U20025 ( .A(n18034), .B(n21005), .Z(n21002) );
  XNOR2_X1 U20026 ( .A(n11315), .B(n11088), .ZN(n20475) );
  NAND2_X1 U20027 ( .A1(n21156), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21000) );
  OAI221_X1 U20028 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18036), .C1(
        n11315), .C2(n18035), .A(n21000), .ZN(n18042) );
  NOR2_X1 U20029 ( .A1(n20995), .A2(n18037), .ZN(n18040) );
  NAND2_X1 U20030 ( .A1(n21027), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n20983) );
  INV_X1 U20031 ( .A(n18038), .ZN(n20984) );
  AOI22_X1 U20032 ( .A1(n18214), .A2(n20983), .B1(n18129), .B2(n20984), .ZN(
        n18049) );
  INV_X1 U20033 ( .A(n18049), .ZN(n18039) );
  MUX2_X1 U20034 ( .A(n18040), .B(n18039), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n18041) );
  AOI211_X1 U20035 ( .C1(n18050), .C2(n20475), .A(n18042), .B(n18041), .ZN(
        n18043) );
  OAI21_X1 U20036 ( .B1(n21002), .B2(n18139), .A(n18043), .ZN(P3_U2800) );
  INV_X1 U20037 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20457) );
  AOI21_X1 U20038 ( .B1(n11314), .B2(n18044), .A(n11088), .ZN(n20446) );
  NOR2_X1 U20039 ( .A1(n20986), .A2(n21040), .ZN(n21025) );
  AOI211_X1 U20040 ( .C1(n21027), .C2(n18214), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n21025), .ZN(n18048) );
  AOI21_X1 U20041 ( .B1(n18046), .B2(n18045), .A(n21020), .ZN(n18047) );
  OAI221_X1 U20042 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18053), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19012), .A(n18052), .ZN(
        n18054) );
  OAI21_X1 U20043 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18056), .A(
        n18055), .ZN(n20292) );
  OAI21_X1 U20044 ( .B1(n18058), .B2(n21101), .A(n18057), .ZN(n21105) );
  AOI21_X1 U20045 ( .B1(n18059), .B2(n19012), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18061) );
  INV_X1 U20046 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21107) );
  OAI22_X1 U20047 ( .A1(n18061), .A2(n18060), .B1(n21129), .B2(n21107), .ZN(
        n18062) );
  AOI21_X1 U20048 ( .B1(n18122), .B2(n21105), .A(n18062), .ZN(n18066) );
  OAI221_X1 U20049 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18064), .A(n18063), .ZN(
        n18065) );
  OAI211_X1 U20050 ( .C1(n18205), .C2(n20292), .A(n18066), .B(n18065), .ZN(
        P3_U2813) );
  NOR2_X1 U20051 ( .A1(n20225), .A2(n20230), .ZN(n18068) );
  AND2_X1 U20052 ( .A1(n18067), .A2(n19012), .ZN(n18085) );
  AOI21_X1 U20053 ( .B1(n18068), .B2(n18085), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18082) );
  INV_X1 U20054 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18070) );
  AOI21_X1 U20055 ( .B1(n18070), .B2(n20243), .A(n18069), .ZN(n20245) );
  AOI22_X1 U20056 ( .A1(n21156), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n20245), 
        .B2(n18215), .ZN(n18080) );
  NAND2_X1 U20057 ( .A1(n18072), .A2(n18071), .ZN(n18073) );
  OAI21_X1 U20058 ( .B1(n20892), .B2(n18112), .A(n18073), .ZN(n18074) );
  XOR2_X1 U20059 ( .A(n18074), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n20887) );
  OAI21_X1 U20060 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18075), .A(
        n20917), .ZN(n20898) );
  OAI21_X1 U20061 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18076), .A(
        n20919), .ZN(n20897) );
  OAI22_X1 U20062 ( .A1(n18077), .A2(n20898), .B1(n18226), .B2(n20897), .ZN(
        n18078) );
  AOI21_X1 U20063 ( .B1(n18122), .B2(n20887), .A(n18078), .ZN(n18079) );
  OAI211_X1 U20064 ( .C1(n18082), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        P3_U2816) );
  INV_X1 U20065 ( .A(n18083), .ZN(n20865) );
  NOR2_X1 U20066 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n20865), .ZN(
        n20868) );
  AOI21_X1 U20067 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n20865), .A(
        n20868), .ZN(n18092) );
  AOI221_X1 U20068 ( .B1(n18093), .B2(n20217), .C1(n20067), .C2(n20217), .A(
        n18084), .ZN(n20201) );
  NOR3_X1 U20069 ( .A1(n18157), .A2(n20134), .A3(n18965), .ZN(n18143) );
  NAND2_X1 U20070 ( .A1(n20200), .A2(n18143), .ZN(n18098) );
  NAND2_X1 U20071 ( .A1(n18221), .A2(n18180), .ZN(n18216) );
  INV_X1 U20072 ( .A(n18216), .ZN(n18096) );
  AOI211_X1 U20073 ( .C1(n18098), .C2(n20217), .A(n18096), .B(n18085), .ZN(
        n18087) );
  INV_X1 U20074 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20871) );
  NOR2_X1 U20075 ( .A1(n21129), .A2(n20871), .ZN(n18086) );
  AOI211_X1 U20076 ( .C1(n20201), .C2(n18215), .A(n18087), .B(n18086), .ZN(
        n18091) );
  OAI22_X1 U20077 ( .A1(n20865), .A2(n18112), .B1(n18107), .B2(n18113), .ZN(
        n18088) );
  XOR2_X1 U20078 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18088), .Z(
        n20869) );
  AOI22_X1 U20079 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18089), .B1(
        n18122), .B2(n20869), .ZN(n18090) );
  OAI211_X1 U20080 ( .C1(n18125), .C2(n18092), .A(n18091), .B(n18090), .ZN(
        P3_U2819) );
  AND3_X1 U20081 ( .A1(n18148), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20162) );
  NAND2_X1 U20082 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20162), .ZN(
        n20170) );
  INV_X1 U20083 ( .A(n20170), .ZN(n18117) );
  NAND2_X1 U20084 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18117), .ZN(
        n20169) );
  NOR2_X1 U20085 ( .A1(n18093), .A2(n20067), .ZN(n18094) );
  AOI21_X1 U20086 ( .B1(n18095), .B2(n20169), .A(n18094), .ZN(n20183) );
  INV_X1 U20087 ( .A(n18143), .ZN(n18115) );
  OAI22_X1 U20088 ( .A1(n18096), .A2(n18095), .B1(n18116), .B2(n18115), .ZN(
        n18097) );
  AOI22_X1 U20089 ( .A1(n20183), .A2(n18215), .B1(n18098), .B2(n18097), .ZN(
        n18111) );
  OAI21_X1 U20090 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18099), .A(
        n18112), .ZN(n18100) );
  OAI21_X1 U20091 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18101), .A(
        n18100), .ZN(n18103) );
  OAI221_X1 U20092 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18113), .C1(
        n21149), .C2(n18112), .A(n18104), .ZN(n18102) );
  OAI21_X1 U20093 ( .B1(n18104), .B2(n18103), .A(n18102), .ZN(n21134) );
  OAI22_X1 U20094 ( .A1(n18104), .A2(n18124), .B1(n18139), .B2(n21134), .ZN(
        n18105) );
  INV_X1 U20095 ( .A(n18105), .ZN(n18110) );
  NAND2_X1 U20096 ( .A1(n21156), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18109) );
  NAND3_X1 U20097 ( .A1(n20865), .A2(n18107), .A3(n18106), .ZN(n18108) );
  NAND4_X1 U20098 ( .A1(n18111), .A2(n18110), .A3(n18109), .A4(n18108), .ZN(
        P3_U2820) );
  NAND2_X1 U20099 ( .A1(n18113), .A2(n18112), .ZN(n18114) );
  XOR2_X1 U20100 ( .A(n18114), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21151) );
  INV_X1 U20101 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21154) );
  NOR2_X1 U20102 ( .A1(n21129), .A2(n21154), .ZN(n18121) );
  NOR2_X1 U20103 ( .A1(n18116), .A2(n18115), .ZN(n18119) );
  INV_X1 U20104 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18134) );
  INV_X1 U20105 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20145) );
  NOR2_X1 U20106 ( .A1(n18134), .A2(n20145), .ZN(n18132) );
  AOI22_X1 U20107 ( .A1(n18132), .A2(n18143), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18216), .ZN(n18118) );
  OAI21_X1 U20108 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18117), .A(
        n20169), .ZN(n20172) );
  OAI22_X1 U20109 ( .A1(n18119), .A2(n18118), .B1(n18205), .B2(n20172), .ZN(
        n18120) );
  AOI211_X1 U20110 ( .C1(n18122), .C2(n21151), .A(n18121), .B(n18120), .ZN(
        n18123) );
  OAI221_X1 U20111 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18125), .C1(
        n21149), .C2(n18124), .A(n18123), .ZN(P3_U2821) );
  OAI21_X1 U20112 ( .B1(n18128), .B2(n18127), .A(n18126), .ZN(n20857) );
  OAI21_X1 U20113 ( .B1(n18148), .B2(n18180), .A(n18221), .ZN(n18144) );
  AOI22_X1 U20114 ( .A1(n18129), .A2(n20857), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18144), .ZN(n18138) );
  AOI21_X1 U20115 ( .B1(n18131), .B2(n20850), .A(n18130), .ZN(n20848) );
  NAND2_X1 U20116 ( .A1(n18148), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18133) );
  AOI211_X1 U20117 ( .C1(n18134), .C2(n18133), .A(n18132), .B(n18965), .ZN(
        n18136) );
  OAI21_X1 U20118 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20162), .A(
        n20170), .ZN(n20163) );
  NAND2_X1 U20119 ( .A1(n21156), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n20855) );
  OAI21_X1 U20120 ( .B1(n18205), .B2(n20163), .A(n20855), .ZN(n18135) );
  AOI211_X1 U20121 ( .C1(n20848), .C2(n18214), .A(n18136), .B(n18135), .ZN(
        n18137) );
  OAI211_X1 U20122 ( .C1(n18139), .C2(n20857), .A(n18138), .B(n18137), .ZN(
        P3_U2822) );
  INV_X1 U20123 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20835) );
  OAI21_X1 U20124 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18141), .A(
        n18140), .ZN(n20847) );
  OAI22_X1 U20125 ( .A1(n21129), .A2(n20835), .B1(n18225), .B2(n20847), .ZN(
        n18142) );
  AOI221_X1 U20126 ( .B1(n18144), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18143), .C2(n20145), .A(n18142), .ZN(n18150) );
  NAND2_X1 U20127 ( .A1(n18146), .A2(n18145), .ZN(n18147) );
  INV_X1 U20128 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20840) );
  XOR2_X1 U20129 ( .A(n18147), .B(n20840), .Z(n20837) );
  NAND2_X1 U20130 ( .A1(n18148), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20129) );
  AOI21_X1 U20131 ( .B1(n20145), .B2(n20129), .A(n20162), .ZN(n20150) );
  AOI22_X1 U20132 ( .A1(n18214), .A2(n20837), .B1(n20150), .B2(n18215), .ZN(
        n18149) );
  NAND2_X1 U20133 ( .A1(n18150), .A2(n18149), .ZN(P3_U2823) );
  OAI21_X1 U20134 ( .B1(n18153), .B2(n18152), .A(n18151), .ZN(n20834) );
  NOR2_X1 U20135 ( .A1(n18157), .A2(n18965), .ZN(n18154) );
  AOI22_X1 U20136 ( .A1(n21156), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18154), 
        .B2(n20134), .ZN(n18160) );
  AOI21_X1 U20137 ( .B1(n20839), .B2(n18156), .A(n18155), .ZN(n20831) );
  NOR2_X1 U20138 ( .A1(n18157), .A2(n20067), .ZN(n18164) );
  OAI21_X1 U20139 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18164), .A(
        n20129), .ZN(n20136) );
  OAI21_X1 U20140 ( .B1(n18965), .B2(n18157), .A(n18216), .ZN(n18170) );
  OAI22_X1 U20141 ( .A1(n18205), .A2(n20136), .B1(n20134), .B2(n18170), .ZN(
        n18158) );
  AOI21_X1 U20142 ( .B1(n18214), .B2(n20831), .A(n18158), .ZN(n18159) );
  OAI211_X1 U20143 ( .C1(n18225), .C2(n20834), .A(n18160), .B(n18159), .ZN(
        P3_U2824) );
  AOI21_X1 U20144 ( .B1(n11299), .B2(n18221), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18171) );
  AOI21_X1 U20145 ( .B1(n18163), .B2(n18162), .A(n18161), .ZN(n20821) );
  NOR2_X1 U20146 ( .A1(n21129), .A2(n20122), .ZN(n20820) );
  NOR2_X1 U20147 ( .A1(n20103), .A2(n20067), .ZN(n18182) );
  INV_X1 U20148 ( .A(n18164), .ZN(n18165) );
  OAI21_X1 U20149 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18182), .A(
        n18165), .ZN(n20116) );
  OAI21_X1 U20150 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18167), .A(
        n18166), .ZN(n20818) );
  OAI22_X1 U20151 ( .A1(n18205), .A2(n20116), .B1(n18225), .B2(n20818), .ZN(
        n18168) );
  AOI211_X1 U20152 ( .C1(n18214), .C2(n20821), .A(n20820), .B(n18168), .ZN(
        n18169) );
  OAI21_X1 U20153 ( .B1(n18171), .B2(n18170), .A(n18169), .ZN(P3_U2825) );
  OAI21_X1 U20154 ( .B1(n18174), .B2(n18173), .A(n18172), .ZN(n20809) );
  AOI21_X1 U20155 ( .B1(n20814), .B2(n18176), .A(n18175), .ZN(n20810) );
  NAND2_X1 U20156 ( .A1(n21156), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n20812) );
  INV_X1 U20157 ( .A(n20812), .ZN(n18179) );
  NOR3_X1 U20158 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18177), .A3(
        n18965), .ZN(n18178) );
  AOI211_X1 U20159 ( .C1(n18214), .C2(n20810), .A(n18179), .B(n18178), .ZN(
        n18185) );
  OAI21_X1 U20160 ( .B1(n18181), .B2(n18180), .A(n18221), .ZN(n18196) );
  INV_X1 U20161 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18183) );
  NAND2_X1 U20162 ( .A1(n18181), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18186) );
  AOI21_X1 U20163 ( .B1(n18183), .B2(n18186), .A(n18182), .ZN(n20108) );
  AOI22_X1 U20164 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18196), .B1(
        n20108), .B2(n18215), .ZN(n18184) );
  OAI211_X1 U20165 ( .C1(n18225), .C2(n20809), .A(n18185), .B(n18184), .ZN(
        P3_U2826) );
  INV_X1 U20166 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20082) );
  NOR2_X1 U20167 ( .A1(n20082), .A2(n20067), .ZN(n18187) );
  OAI21_X1 U20168 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18187), .A(
        n18186), .ZN(n20091) );
  AOI21_X1 U20169 ( .B1(n18190), .B2(n18189), .A(n18188), .ZN(n20798) );
  INV_X1 U20170 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20796) );
  OAI21_X1 U20171 ( .B1(n18193), .B2(n18192), .A(n18191), .ZN(n20805) );
  OAI22_X1 U20172 ( .A1(n21129), .A2(n20796), .B1(n18225), .B2(n20805), .ZN(
        n18194) );
  AOI21_X1 U20173 ( .B1(n18214), .B2(n20798), .A(n18194), .ZN(n18198) );
  NOR2_X1 U20174 ( .A1(n18195), .A2(n20082), .ZN(n18209) );
  OAI21_X1 U20175 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18209), .A(
        n18196), .ZN(n18197) );
  OAI211_X1 U20176 ( .C1(n18205), .C2(n20091), .A(n18198), .B(n18197), .ZN(
        P3_U2827) );
  AOI21_X1 U20177 ( .B1(n18201), .B2(n18200), .A(n18199), .ZN(n20791) );
  NAND2_X1 U20178 ( .A1(n21156), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n20792) );
  INV_X1 U20179 ( .A(n20792), .ZN(n18207) );
  AOI22_X1 U20180 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20067), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20082), .ZN(n20085) );
  OAI21_X1 U20181 ( .B1(n18204), .B2(n18203), .A(n18202), .ZN(n20785) );
  OAI22_X1 U20182 ( .A1(n18205), .A2(n20085), .B1(n18225), .B2(n20785), .ZN(
        n18206) );
  AOI211_X1 U20183 ( .C1(n18214), .C2(n20791), .A(n18207), .B(n18206), .ZN(
        n18208) );
  OAI221_X1 U20184 ( .B1(n18209), .B2(n20082), .C1(n18209), .C2(n18965), .A(
        n18208), .ZN(P3_U2828) );
  OAI21_X1 U20185 ( .B1(n18220), .B2(n18211), .A(n18210), .ZN(n20778) );
  OAI21_X1 U20186 ( .B1(n18213), .B2(n18219), .A(n18212), .ZN(n20776) );
  AOI22_X1 U20187 ( .A1(n21156), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18214), 
        .B2(n20776), .ZN(n18218) );
  AOI22_X1 U20188 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18216), .B1(
        n18215), .B2(n20067), .ZN(n18217) );
  OAI211_X1 U20189 ( .C1(n18225), .C2(n20778), .A(n18218), .B(n18217), .ZN(
        P3_U2829) );
  NOR2_X1 U20190 ( .A1(n18220), .A2(n18219), .ZN(n20775) );
  INV_X1 U20191 ( .A(n20775), .ZN(n20774) );
  NAND3_X1 U20192 ( .A1(n20685), .A2(n18222), .A3(n18221), .ZN(n18223) );
  AOI22_X1 U20193 ( .A1(n21156), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18223), .ZN(n18224) );
  OAI221_X1 U20194 ( .B1(n20775), .B2(n18226), .C1(n20774), .C2(n18225), .A(
        n18224), .ZN(P3_U2830) );
  INV_X1 U20195 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21175) );
  NAND2_X1 U20196 ( .A1(n21174), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18718) );
  INV_X1 U20197 ( .A(n18718), .ZN(n18719) );
  NOR2_X1 U20198 ( .A1(n21174), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18737) );
  NOR2_X1 U20199 ( .A1(n18719), .A2(n18737), .ZN(n18228) );
  OAI22_X1 U20200 ( .A1(n18229), .A2(n21175), .B1(n18228), .B2(n18227), .ZN(
        P3_U2866) );
  NAND2_X1 U20201 ( .A1(n18231), .A2(n18230), .ZN(n18234) );
  OAI21_X1 U20202 ( .B1(n18232), .B2(n18732), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18233) );
  OAI21_X1 U20203 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18234), .A(
        n18233), .ZN(P3_U2864) );
  NOR4_X1 U20204 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18238) );
  NOR4_X1 U20205 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18237) );
  NOR4_X1 U20206 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18236) );
  NOR4_X1 U20207 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18235) );
  NAND4_X1 U20208 ( .A1(n18238), .A2(n18237), .A3(n18236), .A4(n18235), .ZN(
        n18244) );
  NOR4_X1 U20209 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18242) );
  AOI211_X1 U20210 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18241) );
  NOR4_X1 U20211 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18240) );
  NOR4_X1 U20212 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18239) );
  NAND4_X1 U20213 ( .A1(n18242), .A2(n18241), .A3(n18240), .A4(n18239), .ZN(
        n18243) );
  NOR2_X1 U20214 ( .A1(n18244), .A2(n18243), .ZN(n18255) );
  INV_X1 U20215 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18246) );
  OAI21_X1 U20216 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18255), .ZN(n18245) );
  OAI21_X1 U20217 ( .B1(n18255), .B2(n18246), .A(n18245), .ZN(P3_U3293) );
  INV_X1 U20218 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18249) );
  AOI21_X1 U20219 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18247) );
  INV_X1 U20220 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20074) );
  OAI221_X1 U20221 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18247), .C1(n20074), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18255), .ZN(n18248) );
  OAI21_X1 U20222 ( .B1(n18255), .B2(n18249), .A(n18248), .ZN(P3_U3292) );
  INV_X1 U20223 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18251) );
  NOR3_X1 U20224 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18252) );
  OAI21_X1 U20225 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18252), .A(n18255), .ZN(
        n18250) );
  OAI21_X1 U20226 ( .B1(n18255), .B2(n18251), .A(n18250), .ZN(P3_U2638) );
  INV_X1 U20227 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18254) );
  INV_X1 U20228 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21576) );
  OAI211_X1 U20229 ( .C1(n18252), .C2(n20074), .A(n21576), .B(n18255), .ZN(
        n18253) );
  OAI21_X1 U20230 ( .B1(n18255), .B2(n18254), .A(n18253), .ZN(P3_U2639) );
  INV_X2 U20231 ( .A(n18326), .ZN(n21621) );
  OAI22_X1 U20232 ( .A1(n18326), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n21621), .ZN(n18256) );
  INV_X1 U20233 ( .A(n18256), .ZN(P3_U3297) );
  INV_X1 U20234 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18257) );
  AOI22_X1 U20235 ( .A1(n21621), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18257), 
        .B2(n18326), .ZN(P3_U3294) );
  INV_X1 U20236 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21614) );
  AOI21_X1 U20237 ( .B1(n21622), .B2(n21614), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18258) );
  AOI22_X1 U20238 ( .A1(n21621), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18258), 
        .B2(n18326), .ZN(P3_U2635) );
  INV_X1 U20239 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20500) );
  AOI22_X1 U20240 ( .A1(n18302), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18259) );
  OAI21_X1 U20241 ( .B1(n20500), .B2(n18278), .A(n18259), .ZN(P3_U2767) );
  AOI22_X1 U20242 ( .A1(n18302), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18260) );
  OAI21_X1 U20243 ( .B1(n20664), .B2(n18278), .A(n18260), .ZN(P3_U2766) );
  INV_X1 U20244 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20502) );
  AOI22_X1 U20245 ( .A1(n18302), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18261) );
  OAI21_X1 U20246 ( .B1(n20502), .B2(n18278), .A(n18261), .ZN(P3_U2765) );
  INV_X1 U20247 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20546) );
  AOI22_X1 U20248 ( .A1(n18302), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18262) );
  OAI21_X1 U20249 ( .B1(n20546), .B2(n18278), .A(n18262), .ZN(P3_U2764) );
  INV_X1 U20250 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18264) );
  AOI22_X1 U20251 ( .A1(n18302), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18263) );
  OAI21_X1 U20252 ( .B1(n18264), .B2(n18278), .A(n18263), .ZN(P3_U2763) );
  INV_X1 U20253 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18266) );
  AOI22_X1 U20254 ( .A1(n18302), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18265) );
  OAI21_X1 U20255 ( .B1(n18266), .B2(n18278), .A(n18265), .ZN(P3_U2762) );
  INV_X1 U20256 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20527) );
  AOI22_X1 U20257 ( .A1(n18302), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18267) );
  OAI21_X1 U20258 ( .B1(n20527), .B2(n18278), .A(n18267), .ZN(P3_U2761) );
  INV_X1 U20259 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20501) );
  AOI22_X1 U20260 ( .A1(n18302), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18268) );
  OAI21_X1 U20261 ( .B1(n20501), .B2(n18278), .A(n18268), .ZN(P3_U2760) );
  INV_X1 U20262 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U20263 ( .A1(n18302), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18269) );
  OAI21_X1 U20264 ( .B1(n20655), .B2(n18278), .A(n18269), .ZN(P3_U2759) );
  INV_X1 U20265 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20552) );
  AOI22_X1 U20266 ( .A1(n18302), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18270) );
  OAI21_X1 U20267 ( .B1(n20552), .B2(n18278), .A(n18270), .ZN(P3_U2758) );
  INV_X1 U20268 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20554) );
  AOI22_X1 U20269 ( .A1(n18302), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18271) );
  OAI21_X1 U20270 ( .B1(n20554), .B2(n18278), .A(n18271), .ZN(P3_U2757) );
  INV_X1 U20271 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20553) );
  AOI22_X1 U20272 ( .A1(n18302), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18272) );
  OAI21_X1 U20273 ( .B1(n20553), .B2(n18278), .A(n18272), .ZN(P3_U2756) );
  INV_X1 U20274 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U20275 ( .A1(n18302), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18273) );
  OAI21_X1 U20276 ( .B1(n20045), .B2(n18278), .A(n18273), .ZN(P3_U2755) );
  INV_X1 U20277 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U20278 ( .A1(n18302), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18274) );
  OAI21_X1 U20279 ( .B1(n18275), .B2(n18278), .A(n18274), .ZN(P3_U2754) );
  INV_X1 U20280 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20644) );
  AOI22_X1 U20281 ( .A1(n18302), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18276) );
  OAI21_X1 U20282 ( .B1(n20644), .B2(n18278), .A(n18276), .ZN(P3_U2753) );
  INV_X1 U20283 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U20284 ( .A1(n18302), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18277) );
  OAI21_X1 U20285 ( .B1(n20650), .B2(n18278), .A(n18277), .ZN(P3_U2752) );
  INV_X1 U20286 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U20287 ( .A1(n18302), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18280) );
  OAI21_X1 U20288 ( .B1(n18281), .B2(n18304), .A(n18280), .ZN(P3_U2751) );
  INV_X1 U20289 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20568) );
  AOI22_X1 U20290 ( .A1(n18302), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18282) );
  OAI21_X1 U20291 ( .B1(n20568), .B2(n18304), .A(n18282), .ZN(P3_U2750) );
  INV_X1 U20292 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U20293 ( .A1(n18302), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18283) );
  OAI21_X1 U20294 ( .B1(n18284), .B2(n18304), .A(n18283), .ZN(P3_U2749) );
  INV_X1 U20295 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20577) );
  AOI22_X1 U20296 ( .A1(n18302), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18285) );
  OAI21_X1 U20297 ( .B1(n20577), .B2(n18304), .A(n18285), .ZN(P3_U2748) );
  INV_X1 U20298 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18287) );
  AOI22_X1 U20299 ( .A1(n18302), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18286) );
  OAI21_X1 U20300 ( .B1(n18287), .B2(n18304), .A(n18286), .ZN(P3_U2747) );
  INV_X1 U20301 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18289) );
  AOI22_X1 U20302 ( .A1(n18302), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18288) );
  OAI21_X1 U20303 ( .B1(n18289), .B2(n18304), .A(n18288), .ZN(P3_U2746) );
  INV_X1 U20304 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20570) );
  AOI22_X1 U20305 ( .A1(n18302), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18290) );
  OAI21_X1 U20306 ( .B1(n20570), .B2(n18304), .A(n18290), .ZN(P3_U2745) );
  INV_X1 U20307 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U20308 ( .A1(n18302), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18291) );
  OAI21_X1 U20309 ( .B1(n18292), .B2(n18304), .A(n18291), .ZN(P3_U2744) );
  AOI22_X1 U20310 ( .A1(n18302), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18294) );
  OAI21_X1 U20311 ( .B1(n11276), .B2(n18304), .A(n18294), .ZN(P3_U2743) );
  INV_X1 U20312 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20024) );
  AOI22_X1 U20313 ( .A1(n18302), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18295) );
  OAI21_X1 U20314 ( .B1(n20024), .B2(n18304), .A(n18295), .ZN(P3_U2742) );
  INV_X1 U20315 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20597) );
  AOI22_X1 U20316 ( .A1(n18302), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18296) );
  OAI21_X1 U20317 ( .B1(n20597), .B2(n18304), .A(n18296), .ZN(P3_U2741) );
  INV_X1 U20318 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U20319 ( .A1(n18302), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18297) );
  OAI21_X1 U20320 ( .B1(n18298), .B2(n18304), .A(n18297), .ZN(P3_U2740) );
  INV_X1 U20321 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20614) );
  AOI22_X1 U20322 ( .A1(n18302), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18299) );
  OAI21_X1 U20323 ( .B1(n20614), .B2(n18304), .A(n18299), .ZN(P3_U2739) );
  INV_X1 U20324 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18301) );
  AOI22_X1 U20325 ( .A1(n18302), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18300) );
  OAI21_X1 U20326 ( .B1(n18301), .B2(n18304), .A(n18300), .ZN(P3_U2738) );
  INV_X1 U20327 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20030) );
  AOI22_X1 U20328 ( .A1(n18302), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18293), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18303) );
  OAI21_X1 U20329 ( .B1(n20030), .B2(n18304), .A(n18303), .ZN(P3_U2737) );
  NOR2_X1 U20330 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18305), .ZN(n18306) );
  NOR2_X1 U20331 ( .A1(n21621), .A2(n18306), .ZN(P3_U2633) );
  INV_X1 U20332 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20075) );
  NOR2_X1 U20333 ( .A1(n18326), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18320) );
  INV_X2 U20334 ( .A(n18320), .ZN(n18325) );
  AOI22_X1 U20335 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n18326), .ZN(n18307) );
  OAI21_X1 U20336 ( .B1(n20075), .B2(n18325), .A(n18307), .ZN(P3_U3032) );
  AOI22_X1 U20337 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n18326), .ZN(n18308) );
  OAI21_X1 U20338 ( .B1(n20796), .B2(n18325), .A(n18308), .ZN(P3_U3033) );
  INV_X1 U20339 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U20340 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n18326), .ZN(n18309) );
  OAI21_X1 U20341 ( .B1(n20110), .B2(n18325), .A(n18309), .ZN(P3_U3034) );
  AOI22_X1 U20342 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n18326), .ZN(n18310) );
  OAI21_X1 U20343 ( .B1(n20122), .B2(n18325), .A(n18310), .ZN(P3_U3035) );
  INV_X1 U20344 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U20345 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n18326), .ZN(n18311) );
  OAI21_X1 U20346 ( .B1(n20141), .B2(n18325), .A(n18311), .ZN(P3_U3036) );
  AOI22_X1 U20347 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n18326), .ZN(n18312) );
  OAI21_X1 U20348 ( .B1(n20835), .B2(n18325), .A(n18312), .ZN(P3_U3037) );
  AOI22_X1 U20349 ( .A1(n18320), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n18326), .ZN(n18313) );
  OAI21_X1 U20350 ( .B1(n18324), .B2(n20835), .A(n18313), .ZN(P3_U3038) );
  AOI22_X1 U20351 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n18326), .ZN(n18314) );
  OAI21_X1 U20352 ( .B1(n21154), .B2(n18325), .A(n18314), .ZN(P3_U3039) );
  INV_X1 U20353 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20204) );
  INV_X1 U20354 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19726) );
  OAI222_X1 U20355 ( .A1(n18325), .A2(n20204), .B1(n19726), .B2(n21621), .C1(
        n21154), .C2(n18324), .ZN(P3_U3040) );
  INV_X1 U20356 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19728) );
  OAI222_X1 U20357 ( .A1(n18325), .A2(n20871), .B1(n19728), .B2(n21621), .C1(
        n20204), .C2(n18324), .ZN(P3_U3041) );
  INV_X1 U20358 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19730) );
  INV_X1 U20359 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20222) );
  OAI222_X1 U20360 ( .A1(n20871), .A2(n18324), .B1(n19730), .B2(n21621), .C1(
        n20222), .C2(n18325), .ZN(P3_U3042) );
  AOI22_X1 U20361 ( .A1(n18320), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n18326), .ZN(n18315) );
  OAI21_X1 U20362 ( .B1(n18324), .B2(n20222), .A(n18315), .ZN(P3_U3043) );
  INV_X1 U20363 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U20364 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n18326), .ZN(n18316) );
  OAI21_X1 U20365 ( .B1(n18317), .B2(n18325), .A(n18316), .ZN(P3_U3044) );
  INV_X1 U20366 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19734) );
  OAI222_X1 U20367 ( .A1(n18317), .A2(n18324), .B1(n19734), .B2(n21621), .C1(
        n20280), .C2(n18325), .ZN(P3_U3045) );
  INV_X1 U20368 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19736) );
  OAI222_X1 U20369 ( .A1(n18325), .A2(n20281), .B1(n19736), .B2(n21621), .C1(
        n20280), .C2(n18324), .ZN(P3_U3046) );
  INV_X1 U20370 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19738) );
  OAI222_X1 U20371 ( .A1(n18325), .A2(n21107), .B1(n19738), .B2(n21621), .C1(
        n20281), .C2(n18324), .ZN(P3_U3047) );
  INV_X1 U20372 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20310) );
  INV_X1 U20373 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19740) );
  OAI222_X1 U20374 ( .A1(n18325), .A2(n20310), .B1(n19740), .B2(n21621), .C1(
        n21107), .C2(n18324), .ZN(P3_U3048) );
  INV_X1 U20375 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19742) );
  INV_X1 U20376 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20321) );
  OAI222_X1 U20377 ( .A1(n20310), .A2(n18324), .B1(n19742), .B2(n21621), .C1(
        n20321), .C2(n18325), .ZN(P3_U3049) );
  INV_X1 U20378 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20339) );
  INV_X1 U20379 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19744) );
  OAI222_X1 U20380 ( .A1(n18325), .A2(n20339), .B1(n19744), .B2(n21621), .C1(
        n20321), .C2(n18324), .ZN(P3_U3050) );
  INV_X1 U20381 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20354) );
  INV_X1 U20382 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19746) );
  OAI222_X1 U20383 ( .A1(n18325), .A2(n20354), .B1(n19746), .B2(n21621), .C1(
        n20339), .C2(n18324), .ZN(P3_U3051) );
  INV_X1 U20384 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20364) );
  INV_X1 U20385 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19748) );
  OAI222_X1 U20386 ( .A1(n18325), .A2(n20364), .B1(n19748), .B2(n21621), .C1(
        n20354), .C2(n18324), .ZN(P3_U3052) );
  INV_X1 U20387 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19750) );
  OAI222_X1 U20388 ( .A1(n18325), .A2(n20367), .B1(n19750), .B2(n21621), .C1(
        n20364), .C2(n18324), .ZN(P3_U3053) );
  INV_X1 U20389 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19752) );
  INV_X1 U20390 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20388) );
  OAI222_X1 U20391 ( .A1(n20367), .A2(n18324), .B1(n19752), .B2(n21621), .C1(
        n20388), .C2(n18325), .ZN(P3_U3054) );
  INV_X1 U20392 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19754) );
  OAI222_X1 U20393 ( .A1(n18325), .A2(n20403), .B1(n19754), .B2(n21621), .C1(
        n20388), .C2(n18324), .ZN(P3_U3055) );
  AOI22_X1 U20394 ( .A1(n18320), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n18326), .ZN(n18318) );
  OAI21_X1 U20395 ( .B1(n18324), .B2(n20403), .A(n18318), .ZN(P3_U3056) );
  INV_X1 U20396 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20430) );
  AOI22_X1 U20397 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n18326), .ZN(n18319) );
  OAI21_X1 U20398 ( .B1(n20430), .B2(n18325), .A(n18319), .ZN(P3_U3057) );
  AOI22_X1 U20399 ( .A1(n18320), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n18326), .ZN(n18321) );
  OAI21_X1 U20400 ( .B1(n18324), .B2(n20430), .A(n18321), .ZN(P3_U3058) );
  AOI22_X1 U20401 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18322), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n18326), .ZN(n18323) );
  OAI21_X1 U20402 ( .B1(n20457), .B2(n18325), .A(n18323), .ZN(P3_U3059) );
  INV_X1 U20403 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20470) );
  INV_X1 U20404 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19762) );
  OAI222_X1 U20405 ( .A1(n18325), .A2(n20470), .B1(n19762), .B2(n21621), .C1(
        n20457), .C2(n18324), .ZN(P3_U3060) );
  INV_X1 U20406 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19765) );
  OAI222_X1 U20407 ( .A1(n18325), .A2(n20477), .B1(n19765), .B2(n21621), .C1(
        n20470), .C2(n18324), .ZN(P3_U3061) );
  OAI22_X1 U20408 ( .A1(n18326), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n21621), .ZN(n18327) );
  INV_X1 U20409 ( .A(n18327), .ZN(P3_U3277) );
  OAI22_X1 U20410 ( .A1(n18326), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n21621), .ZN(n18328) );
  INV_X1 U20411 ( .A(n18328), .ZN(P3_U3276) );
  OAI22_X1 U20412 ( .A1(n18326), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n21621), .ZN(n18329) );
  INV_X1 U20413 ( .A(n18329), .ZN(P3_U3275) );
  OAI22_X1 U20414 ( .A1(n18326), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n21621), .ZN(n18330) );
  INV_X1 U20415 ( .A(n18330), .ZN(P3_U3274) );
  NOR4_X1 U20416 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18333)
         );
  INV_X1 U20417 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18331) );
  NOR4_X1 U20418 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18331), .ZN(n18332) );
  INV_X2 U20419 ( .A(n19008), .ZN(U215) );
  NAND3_X1 U20420 ( .A1(n18333), .A2(n18332), .A3(U215), .ZN(U213) );
  NOR2_X1 U20421 ( .A1(n21594), .A2(n19263), .ZN(n18339) );
  OAI21_X1 U20422 ( .B1(n21604), .B2(n21569), .A(n12525), .ZN(n18337) );
  NAND3_X1 U20423 ( .A1(n21604), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n18334), 
        .ZN(n18336) );
  MUX2_X1 U20424 ( .A(n18337), .B(n18336), .S(n18335), .Z(n18338) );
  OAI21_X1 U20425 ( .B1(n18339), .B2(n18656), .A(n18338), .ZN(n18347) );
  NAND4_X1 U20426 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n18340), .A4(n18655), .ZN(n18343) );
  INV_X1 U20427 ( .A(n18341), .ZN(n18342) );
  OAI211_X1 U20428 ( .C1(n18345), .C2(n18344), .A(n18343), .B(n18342), .ZN(
        n18346) );
  MUX2_X1 U20429 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n18347), .S(n18346), 
        .Z(P2_U3610) );
  INV_X1 U20430 ( .A(n18348), .ZN(n18361) );
  NAND2_X1 U20431 ( .A1(n18349), .A2(n18570), .ZN(n18355) );
  OAI22_X1 U20432 ( .A1(n18576), .A2(n18583), .B1(n12555), .B2(n18562), .ZN(
        n18350) );
  INV_X1 U20433 ( .A(n18350), .ZN(n18354) );
  NAND2_X1 U20434 ( .A1(n18568), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18353) );
  NAND2_X1 U20435 ( .A1(n18572), .A2(n18351), .ZN(n18352) );
  AND4_X1 U20436 ( .A1(n18355), .A2(n18354), .A3(n18353), .A4(n18352), .ZN(
        n18360) );
  NOR2_X1 U20437 ( .A1(n18564), .A2(n18356), .ZN(n18357) );
  AOI21_X1 U20438 ( .B1(n19195), .B2(n18358), .A(n18357), .ZN(n18359) );
  OAI211_X1 U20439 ( .C1(n18643), .C2(n18361), .A(n18360), .B(n18359), .ZN(
        P2_U2855) );
  OAI21_X1 U20440 ( .B1(n13225), .B2(n18562), .A(n18488), .ZN(n18364) );
  OAI22_X1 U20441 ( .A1(n18516), .A2(n12782), .B1(n18362), .B2(n18509), .ZN(
        n18363) );
  AOI211_X1 U20442 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18529), .A(
        n18364), .B(n18363), .ZN(n18371) );
  NAND2_X1 U20443 ( .A1(n10997), .A2(n18365), .ZN(n18366) );
  XNOR2_X1 U20444 ( .A(n18367), .B(n18366), .ZN(n18369) );
  AOI22_X1 U20445 ( .A1(n18369), .A2(n18558), .B1(n18368), .B2(n18570), .ZN(
        n18370) );
  OAI211_X1 U20446 ( .C1(n18576), .C2(n19347), .A(n18371), .B(n18370), .ZN(
        P2_U2850) );
  OAI21_X1 U20447 ( .B1(n18372), .B2(n18562), .A(n18488), .ZN(n18376) );
  INV_X1 U20448 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18374) );
  OAI22_X1 U20449 ( .A1(n18516), .A2(n18374), .B1(n18373), .B2(n18509), .ZN(
        n18375) );
  AOI211_X1 U20450 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18529), .A(
        n18376), .B(n18375), .ZN(n18383) );
  NOR2_X1 U20451 ( .A1(n18535), .A2(n18377), .ZN(n18379) );
  XNOR2_X1 U20452 ( .A(n18379), .B(n18378), .ZN(n18381) );
  AOI22_X1 U20453 ( .A1(n18381), .A2(n18558), .B1(n18380), .B2(n18570), .ZN(
        n18382) );
  OAI211_X1 U20454 ( .C1(n18576), .C2(n18384), .A(n18383), .B(n18382), .ZN(
        P2_U2849) );
  NAND2_X1 U20455 ( .A1(n10997), .A2(n18385), .ZN(n18387) );
  XOR2_X1 U20456 ( .A(n18387), .B(n18386), .Z(n18395) );
  AOI22_X1 U20457 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n18568), .B1(n18572), .B2(
        n18388), .ZN(n18389) );
  OAI211_X1 U20458 ( .C1(n13095), .C2(n18562), .A(n18389), .B(n18600), .ZN(
        n18393) );
  OAI22_X1 U20459 ( .A1(n18511), .A2(n18391), .B1(n18576), .B2(n18390), .ZN(
        n18392) );
  AOI211_X1 U20460 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18529), .A(
        n18393), .B(n18392), .ZN(n18394) );
  OAI21_X1 U20461 ( .B1(n18395), .B2(n18643), .A(n18394), .ZN(P2_U2848) );
  NAND2_X1 U20462 ( .A1(n10997), .A2(n18396), .ZN(n18399) );
  INV_X1 U20463 ( .A(n18397), .ZN(n18398) );
  XNOR2_X1 U20464 ( .A(n18399), .B(n18398), .ZN(n18408) );
  AOI22_X1 U20465 ( .A1(n18400), .A2(n18572), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18529), .ZN(n18401) );
  OAI211_X1 U20466 ( .C1(n18402), .C2(n18562), .A(n18401), .B(n18488), .ZN(
        n18406) );
  OAI22_X1 U20467 ( .A1(n18404), .A2(n18511), .B1(n18403), .B2(n18576), .ZN(
        n18405) );
  AOI211_X1 U20468 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18568), .A(n18406), .B(
        n18405), .ZN(n18407) );
  OAI21_X1 U20469 ( .B1(n18408), .B2(n18643), .A(n18407), .ZN(P2_U2846) );
  INV_X1 U20470 ( .A(n18409), .ZN(n18416) );
  INV_X1 U20471 ( .A(n19115), .ZN(n18412) );
  AOI22_X1 U20472 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18568), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18529), .ZN(n18410) );
  OAI211_X1 U20473 ( .C1(n16597), .C2(n18562), .A(n18600), .B(n18410), .ZN(
        n18411) );
  AOI21_X1 U20474 ( .B1(n18531), .B2(n18412), .A(n18411), .ZN(n18413) );
  OAI21_X1 U20475 ( .B1(n18414), .B2(n18511), .A(n18413), .ZN(n18415) );
  AOI21_X1 U20476 ( .B1(n18416), .B2(n18572), .A(n18415), .ZN(n18421) );
  INV_X1 U20477 ( .A(n18417), .ZN(n18419) );
  OAI21_X1 U20478 ( .B1(n18419), .B2(n18422), .A(n18418), .ZN(n18420) );
  OAI211_X1 U20479 ( .C1(n18507), .C2(n18422), .A(n18421), .B(n18420), .ZN(
        P2_U2844) );
  AOI22_X1 U20480 ( .A1(n18423), .A2(n18572), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n18568), .ZN(n18424) );
  OAI21_X1 U20481 ( .B1(n18425), .B2(n18564), .A(n18424), .ZN(n18426) );
  AOI211_X1 U20482 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18528), .A(n18427), 
        .B(n18426), .ZN(n18435) );
  NAND2_X1 U20483 ( .A1(n10997), .A2(n18428), .ZN(n18430) );
  XNOR2_X1 U20484 ( .A(n18430), .B(n18429), .ZN(n18433) );
  INV_X1 U20485 ( .A(n18431), .ZN(n18432) );
  AOI22_X1 U20486 ( .A1(n18433), .A2(n18558), .B1(n18432), .B2(n18570), .ZN(
        n18434) );
  OAI211_X1 U20487 ( .C1(n18436), .C2(n18576), .A(n18435), .B(n18434), .ZN(
        P2_U2842) );
  NAND2_X1 U20488 ( .A1(n10997), .A2(n18437), .ZN(n18439) );
  XOR2_X1 U20489 ( .A(n18439), .B(n18438), .Z(n18448) );
  AOI22_X1 U20490 ( .A1(n18440), .A2(n18572), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18529), .ZN(n18441) );
  OAI211_X1 U20491 ( .C1(n18442), .C2(n18562), .A(n18441), .B(n18488), .ZN(
        n18446) );
  OAI22_X1 U20492 ( .A1(n18444), .A2(n18511), .B1(n18443), .B2(n18576), .ZN(
        n18445) );
  AOI211_X1 U20493 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n18568), .A(n18446), .B(
        n18445), .ZN(n18447) );
  OAI21_X1 U20494 ( .B1(n18448), .B2(n18643), .A(n18447), .ZN(P2_U2840) );
  NOR2_X1 U20495 ( .A1(n18535), .A2(n18449), .ZN(n18450) );
  XNOR2_X1 U20496 ( .A(n18451), .B(n18450), .ZN(n18460) );
  INV_X1 U20497 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U20498 ( .A1(n18452), .A2(n18572), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18568), .ZN(n18453) );
  OAI21_X1 U20499 ( .B1(n18454), .B2(n18564), .A(n18453), .ZN(n18455) );
  AOI211_X1 U20500 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18528), .A(n18427), 
        .B(n18455), .ZN(n18459) );
  INV_X1 U20501 ( .A(n18456), .ZN(n19584) );
  AOI22_X1 U20502 ( .A1(n18457), .A2(n18570), .B1(n18531), .B2(n19584), .ZN(
        n18458) );
  OAI211_X1 U20503 ( .C1(n18643), .C2(n18460), .A(n18459), .B(n18458), .ZN(
        P2_U2839) );
  NAND2_X1 U20504 ( .A1(n10997), .A2(n18461), .ZN(n18462) );
  XOR2_X1 U20505 ( .A(n18463), .B(n18462), .Z(n18472) );
  AOI22_X1 U20506 ( .A1(n18464), .A2(n18572), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n18568), .ZN(n18465) );
  OAI211_X1 U20507 ( .C1(n16535), .C2(n18562), .A(n18465), .B(n18488), .ZN(
        n18466) );
  AOI21_X1 U20508 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18529), .A(
        n18466), .ZN(n18471) );
  INV_X1 U20509 ( .A(n18467), .ZN(n18469) );
  AOI22_X1 U20510 ( .A1(n18469), .A2(n18570), .B1(n18531), .B2(n18468), .ZN(
        n18470) );
  OAI211_X1 U20511 ( .C1(n18643), .C2(n18472), .A(n18471), .B(n18470), .ZN(
        P2_U2838) );
  NOR2_X1 U20512 ( .A1(n18535), .A2(n18473), .ZN(n18475) );
  XOR2_X1 U20513 ( .A(n18475), .B(n18474), .Z(n18483) );
  AOI22_X1 U20514 ( .A1(n18476), .A2(n18572), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18568), .ZN(n18477) );
  OAI211_X1 U20515 ( .C1(n16522), .C2(n18562), .A(n18477), .B(n18600), .ZN(
        n18478) );
  AOI21_X1 U20516 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18529), .A(
        n18478), .ZN(n18482) );
  OAI22_X1 U20517 ( .A1(n18479), .A2(n18511), .B1(n19481), .B2(n18576), .ZN(
        n18480) );
  INV_X1 U20518 ( .A(n18480), .ZN(n18481) );
  OAI211_X1 U20519 ( .C1(n18643), .C2(n18483), .A(n18482), .B(n18481), .ZN(
        P2_U2837) );
  NAND2_X1 U20520 ( .A1(n10997), .A2(n18484), .ZN(n18485) );
  XOR2_X1 U20521 ( .A(n18486), .B(n18485), .Z(n18497) );
  AOI22_X1 U20522 ( .A1(n18487), .A2(n18572), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n18568), .ZN(n18489) );
  OAI211_X1 U20523 ( .C1(n18490), .C2(n18562), .A(n18489), .B(n18488), .ZN(
        n18491) );
  AOI21_X1 U20524 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18529), .A(
        n18491), .ZN(n18496) );
  OAI22_X1 U20525 ( .A1(n18493), .A2(n18511), .B1(n18492), .B2(n18576), .ZN(
        n18494) );
  INV_X1 U20526 ( .A(n18494), .ZN(n18495) );
  OAI211_X1 U20527 ( .C1(n18643), .C2(n18497), .A(n18496), .B(n18495), .ZN(
        P2_U2836) );
  AOI22_X1 U20528 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18529), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18528), .ZN(n18498) );
  OAI21_X1 U20529 ( .B1(n18499), .B2(n18509), .A(n18498), .ZN(n18502) );
  OAI22_X1 U20530 ( .A1(n18500), .A2(n18511), .B1(n19394), .B2(n18576), .ZN(
        n18501) );
  AOI211_X1 U20531 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n18568), .A(n18502), .B(
        n18501), .ZN(n18506) );
  NAND2_X1 U20532 ( .A1(n10997), .A2(n18503), .ZN(n18521) );
  INV_X1 U20533 ( .A(n18521), .ZN(n18523) );
  OAI211_X1 U20534 ( .C1(n18504), .C2(n18508), .A(n18558), .B(n18523), .ZN(
        n18505) );
  OAI211_X1 U20535 ( .C1(n18508), .C2(n18507), .A(n18506), .B(n18505), .ZN(
        P2_U2835) );
  NOR2_X1 U20536 ( .A1(n18510), .A2(n18509), .ZN(n18520) );
  NOR2_X1 U20537 ( .A1(n18512), .A2(n18511), .ZN(n18519) );
  OAI22_X1 U20538 ( .A1(n18514), .A2(n18564), .B1(n18513), .B2(n18562), .ZN(
        n18518) );
  INV_X1 U20539 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n18515) );
  NOR2_X1 U20540 ( .A1(n18516), .A2(n18515), .ZN(n18517) );
  NOR4_X1 U20541 ( .A1(n18520), .A2(n18519), .A3(n18518), .A4(n18517), .ZN(
        n18526) );
  INV_X1 U20542 ( .A(n18524), .ZN(n18522) );
  OAI221_X1 U20543 ( .B1(n18524), .B2(n18523), .C1(n18522), .C2(n18521), .A(
        n18558), .ZN(n18525) );
  OAI211_X1 U20544 ( .C1(n18576), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        P2_U2834) );
  AOI22_X1 U20545 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18529), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18528), .ZN(n18542) );
  AOI22_X1 U20546 ( .A1(n18530), .A2(n18572), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n18568), .ZN(n18541) );
  AOI22_X1 U20547 ( .A1(n18532), .A2(n18570), .B1(n19299), .B2(n18531), .ZN(
        n18540) );
  INV_X1 U20548 ( .A(n18533), .ZN(n18538) );
  NOR2_X1 U20549 ( .A1(n18535), .A2(n18534), .ZN(n18537) );
  AOI21_X1 U20550 ( .B1(n18538), .B2(n18537), .A(n18643), .ZN(n18536) );
  OAI21_X1 U20551 ( .B1(n18538), .B2(n18537), .A(n18536), .ZN(n18539) );
  NAND4_X1 U20552 ( .A1(n18542), .A2(n18541), .A3(n18540), .A4(n18539), .ZN(
        P2_U2833) );
  AND2_X1 U20553 ( .A1(n10997), .A2(n18543), .ZN(n18545) );
  OAI21_X1 U20554 ( .B1(n18546), .B2(n18545), .A(n18558), .ZN(n18544) );
  AOI21_X1 U20555 ( .B1(n18546), .B2(n18545), .A(n18544), .ZN(n18550) );
  OAI22_X1 U20556 ( .A1(n18548), .A2(n18564), .B1(n18547), .B2(n18562), .ZN(
        n18549) );
  AOI211_X1 U20557 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n18568), .A(n18550), .B(
        n18549), .ZN(n18554) );
  AOI22_X1 U20558 ( .A1(n18552), .A2(n18570), .B1(n18551), .B2(n18572), .ZN(
        n18553) );
  OAI211_X1 U20559 ( .C1(n18555), .C2(n18576), .A(n18554), .B(n18553), .ZN(
        P2_U2830) );
  AND2_X1 U20560 ( .A1(n10997), .A2(n18556), .ZN(n18560) );
  OAI21_X1 U20561 ( .B1(n18561), .B2(n18560), .A(n18558), .ZN(n18559) );
  AOI21_X1 U20562 ( .B1(n18561), .B2(n18560), .A(n18559), .ZN(n18567) );
  OAI22_X1 U20563 ( .A1(n18565), .A2(n18564), .B1(n18563), .B2(n18562), .ZN(
        n18566) );
  AOI211_X1 U20564 ( .C1(P2_EBX_REG_29__SCAN_IN), .C2(n18568), .A(n18567), .B(
        n18566), .ZN(n18575) );
  INV_X1 U20565 ( .A(n18569), .ZN(n18571) );
  AOI22_X1 U20566 ( .A1(n18573), .A2(n18572), .B1(n18571), .B2(n18570), .ZN(
        n18574) );
  OAI211_X1 U20567 ( .C1(n18577), .C2(n18576), .A(n18575), .B(n18574), .ZN(
        P2_U2826) );
  INV_X1 U20568 ( .A(n18579), .ZN(n18582) );
  OR3_X1 U20569 ( .A1(n18579), .A2(n18638), .A3(n18578), .ZN(n18580) );
  OAI21_X1 U20570 ( .B1(n18582), .B2(n18581), .A(n18580), .ZN(P2_U3595) );
  OAI22_X1 U20571 ( .A1(n18584), .A2(n18614), .B1(n18603), .B2(n18583), .ZN(
        n18585) );
  INV_X1 U20572 ( .A(n18585), .ZN(n18592) );
  OAI22_X1 U20573 ( .A1(n18587), .A2(n18607), .B1(n18608), .B2(n18586), .ZN(
        n18588) );
  AOI211_X1 U20574 ( .C1(n18590), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18589), .B(n18588), .ZN(n18591) );
  OAI211_X1 U20575 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18593), .A(
        n18592), .B(n18591), .ZN(P2_U3046) );
  OAI221_X1 U20576 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n18598), .C2(n18595), .A(
        n18594), .ZN(n18596) );
  OAI22_X1 U20577 ( .A1(n18599), .A2(n18598), .B1(n18597), .B2(n18596), .ZN(
        n18605) );
  OAI22_X1 U20578 ( .A1(n18603), .A2(n18602), .B1(n18601), .B2(n18600), .ZN(
        n18604) );
  NOR2_X1 U20579 ( .A1(n18605), .A2(n18604), .ZN(n18612) );
  OAI22_X1 U20580 ( .A1(n18609), .A2(n18608), .B1(n18607), .B2(n18606), .ZN(
        n18610) );
  INV_X1 U20581 ( .A(n18610), .ZN(n18611) );
  OAI211_X1 U20582 ( .C1(n18614), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P2_U3038) );
  AOI21_X1 U20583 ( .B1(n18617), .B2(n18616), .A(n18615), .ZN(n18618) );
  AOI21_X1 U20584 ( .B1(n18620), .B2(n18619), .A(n18618), .ZN(n18634) );
  AOI21_X1 U20585 ( .B1(n18623), .B2(n18622), .A(n18621), .ZN(n18632) );
  NAND2_X1 U20586 ( .A1(n18625), .A2(n18624), .ZN(n18631) );
  NAND2_X1 U20587 ( .A1(n18627), .A2(n18626), .ZN(n18630) );
  NAND2_X1 U20588 ( .A1(n18628), .A2(n19487), .ZN(n18629) );
  AND4_X1 U20589 ( .A1(n18632), .A2(n18631), .A3(n18630), .A4(n18629), .ZN(
        n18633) );
  OAI211_X1 U20590 ( .C1(n18636), .C2(n18635), .A(n18634), .B(n18633), .ZN(
        P2_U3044) );
  NAND2_X1 U20591 ( .A1(n18652), .A2(n18637), .ZN(n18654) );
  OAI21_X1 U20592 ( .B1(n18639), .B2(n18638), .A(n18661), .ZN(n18642) );
  NAND2_X1 U20593 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21594), .ZN(n18640) );
  AOI21_X1 U20594 ( .B1(n18646), .B2(n18654), .A(n18640), .ZN(n18641) );
  AOI21_X1 U20595 ( .B1(n18654), .B2(n18642), .A(n18641), .ZN(n18644) );
  NAND2_X1 U20596 ( .A1(n18644), .A2(n18643), .ZN(P2_U3177) );
  INV_X1 U20597 ( .A(n18645), .ZN(n18648) );
  OAI22_X1 U20598 ( .A1(n18648), .A2(n18647), .B1(n18655), .B2(n18646), .ZN(
        n18650) );
  OR2_X1 U20599 ( .A1(n18650), .A2(n18649), .ZN(n18651) );
  AOI21_X1 U20600 ( .B1(n18652), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n18651), 
        .ZN(n18659) );
  NOR2_X1 U20601 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18653), .ZN(n18657) );
  OAI22_X1 U20602 ( .A1(n18657), .A2(n18656), .B1(n18655), .B2(n18654), .ZN(
        n18658) );
  OAI211_X1 U20603 ( .C1(n18660), .C2(n18661), .A(n18659), .B(n18658), .ZN(
        P2_U3176) );
  NOR2_X1 U20604 ( .A1(n18662), .A2(n18661), .ZN(n18666) );
  MUX2_X1 U20605 ( .A(P2_MORE_REG_SCAN_IN), .B(n18663), .S(n18666), .Z(
        P2_U3609) );
  OAI21_X1 U20606 ( .B1(n18666), .B2(n18665), .A(n18664), .ZN(P2_U2819) );
  INV_X1 U20607 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20000) );
  INV_X1 U20608 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18694) );
  AOI22_X1 U20609 ( .A1(n19008), .A2(n20000), .B1(n18694), .B2(U215), .ZN(U282) );
  OAI22_X1 U20610 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19008), .ZN(n18667) );
  INV_X1 U20611 ( .A(n18667), .ZN(U281) );
  OAI22_X1 U20612 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19008), .ZN(n18668) );
  INV_X1 U20613 ( .A(n18668), .ZN(U280) );
  OAI22_X1 U20614 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19008), .ZN(n18669) );
  INV_X1 U20615 ( .A(n18669), .ZN(U279) );
  OAI22_X1 U20616 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19008), .ZN(n18670) );
  INV_X1 U20617 ( .A(n18670), .ZN(U278) );
  OAI22_X1 U20618 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19008), .ZN(n18671) );
  INV_X1 U20619 ( .A(n18671), .ZN(U277) );
  OAI22_X1 U20620 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19008), .ZN(n18672) );
  INV_X1 U20621 ( .A(n18672), .ZN(U276) );
  OAI22_X1 U20622 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19008), .ZN(n18673) );
  INV_X1 U20623 ( .A(n18673), .ZN(U275) );
  OAI22_X1 U20624 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19008), .ZN(n18674) );
  INV_X1 U20625 ( .A(n18674), .ZN(U274) );
  OAI22_X1 U20626 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19008), .ZN(n18675) );
  INV_X1 U20627 ( .A(n18675), .ZN(U273) );
  OAI22_X1 U20628 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19008), .ZN(n18676) );
  INV_X1 U20629 ( .A(n18676), .ZN(U272) );
  OAI22_X1 U20630 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19008), .ZN(n18677) );
  INV_X1 U20631 ( .A(n18677), .ZN(U271) );
  OAI22_X1 U20632 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18690), .ZN(n18678) );
  INV_X1 U20633 ( .A(n18678), .ZN(U270) );
  OAI22_X1 U20634 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19008), .ZN(n18679) );
  INV_X1 U20635 ( .A(n18679), .ZN(U269) );
  OAI22_X1 U20636 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18690), .ZN(n18680) );
  INV_X1 U20637 ( .A(n18680), .ZN(U268) );
  OAI22_X1 U20638 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19008), .ZN(n18681) );
  INV_X1 U20639 ( .A(n18681), .ZN(U267) );
  OAI22_X1 U20640 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18690), .ZN(n18682) );
  INV_X1 U20641 ( .A(n18682), .ZN(U266) );
  OAI22_X1 U20642 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19008), .ZN(n18683) );
  INV_X1 U20643 ( .A(n18683), .ZN(U265) );
  OAI22_X1 U20644 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18690), .ZN(n18684) );
  INV_X1 U20645 ( .A(n18684), .ZN(U264) );
  OAI22_X1 U20646 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18690), .ZN(n18685) );
  INV_X1 U20647 ( .A(n18685), .ZN(U263) );
  OAI22_X1 U20648 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18690), .ZN(n18686) );
  INV_X1 U20649 ( .A(n18686), .ZN(U262) );
  OAI22_X1 U20650 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18690), .ZN(n18687) );
  INV_X1 U20651 ( .A(n18687), .ZN(U261) );
  OAI22_X1 U20652 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n18690), .ZN(n18688) );
  INV_X1 U20653 ( .A(n18688), .ZN(U260) );
  OAI22_X1 U20654 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18690), .ZN(n18689) );
  INV_X1 U20655 ( .A(n18689), .ZN(U259) );
  OAI22_X1 U20656 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18690), .ZN(n18691) );
  INV_X1 U20657 ( .A(n18691), .ZN(U258) );
  NOR2_X1 U20658 ( .A1(n21175), .A2(n18712), .ZN(n18755) );
  NAND2_X1 U20659 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18755), .ZN(
        n18913) );
  NAND2_X1 U20660 ( .A1(n18693), .A2(n18692), .ZN(n19014) );
  INV_X1 U20661 ( .A(n19014), .ZN(n18806) );
  NAND2_X1 U20662 ( .A1(n18806), .A2(n20592), .ZN(n18766) );
  NAND2_X1 U20663 ( .A1(n21075), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21199) );
  AND2_X1 U20664 ( .A1(n21199), .A2(n18755), .ZN(n19013) );
  INV_X1 U20665 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20529) );
  NOR2_X2 U20666 ( .A1(n20529), .A2(n19011), .ZN(n18758) );
  NOR3_X1 U20667 ( .A1(n21174), .A2(n21175), .A3(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18700) );
  NAND2_X1 U20668 ( .A1(n21166), .A2(n18700), .ZN(n18969) );
  INV_X1 U20669 ( .A(n18969), .ZN(n19029) );
  NOR2_X2 U20670 ( .A1(n18694), .A2(n18965), .ZN(n18759) );
  AOI22_X1 U20671 ( .A1(n19013), .A2(n18758), .B1(n19029), .B2(n18759), .ZN(
        n18697) );
  NOR2_X1 U20672 ( .A1(n18695), .A2(n19011), .ZN(n18729) );
  AOI22_X1 U20673 ( .A1(n19012), .A2(n18700), .B1(n18755), .B2(n18729), .ZN(
        n19015) );
  NAND2_X1 U20674 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18700), .ZN(
        n19109) );
  INV_X1 U20675 ( .A(n19109), .ZN(n19023) );
  NOR2_X2 U20676 ( .A1(n20636), .A2(n18965), .ZN(n18763) );
  AOI22_X1 U20677 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19015), .B1(
        n19023), .B2(n18763), .ZN(n18696) );
  OAI211_X1 U20678 ( .C1(n18913), .C2(n18766), .A(n18697), .B(n18696), .ZN(
        P3_U2995) );
  NAND2_X1 U20679 ( .A1(n18755), .A2(n21166), .ZN(n19098) );
  NAND2_X1 U20680 ( .A1(n19109), .A2(n19098), .ZN(n18762) );
  AND2_X1 U20681 ( .A1(n21199), .A2(n18762), .ZN(n19018) );
  NOR2_X1 U20682 ( .A1(n21169), .A2(n18718), .ZN(n18707) );
  NAND2_X1 U20683 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18707), .ZN(
        n19027) );
  INV_X1 U20684 ( .A(n19027), .ZN(n19035) );
  AOI22_X1 U20685 ( .A1(n18758), .A2(n19018), .B1(n18759), .B2(n19035), .ZN(
        n18699) );
  NAND2_X1 U20686 ( .A1(n18969), .A2(n19027), .ZN(n18703) );
  AOI21_X1 U20687 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19011), .ZN(n18761) );
  OAI221_X1 U20688 ( .B1(n18762), .B2(n18732), .C1(n18762), .C2(n18703), .A(
        n18761), .ZN(n19019) );
  AOI22_X1 U20689 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19019), .B1(
        n18763), .B2(n19029), .ZN(n18698) );
  OAI211_X1 U20690 ( .C1(n18766), .C2(n19098), .A(n18699), .B(n18698), .ZN(
        P3_U2987) );
  AND2_X1 U20691 ( .A1(n21199), .A2(n18700), .ZN(n19022) );
  NAND2_X1 U20692 ( .A1(n21166), .A2(n18707), .ZN(n18931) );
  INV_X1 U20693 ( .A(n18931), .ZN(n19040) );
  AOI22_X1 U20694 ( .A1(n18758), .A2(n19022), .B1(n18759), .B2(n19040), .ZN(
        n18702) );
  AOI22_X1 U20695 ( .A1(n19012), .A2(n18707), .B1(n18700), .B2(n18729), .ZN(
        n19024) );
  AOI22_X1 U20696 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19024), .B1(
        n18763), .B2(n19035), .ZN(n18701) );
  OAI211_X1 U20697 ( .C1(n19109), .C2(n18766), .A(n18702), .B(n18701), .ZN(
        P3_U2979) );
  AND2_X1 U20698 ( .A1(n21199), .A2(n18703), .ZN(n19028) );
  AOI22_X1 U20699 ( .A1(n18763), .A2(n19040), .B1(n18758), .B2(n19028), .ZN(
        n18706) );
  NAND2_X1 U20700 ( .A1(n21169), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18723) );
  NOR2_X2 U20701 ( .A1(n18718), .A2(n18723), .ZN(n19046) );
  NOR2_X1 U20702 ( .A1(n19040), .A2(n19046), .ZN(n18713) );
  INV_X1 U20703 ( .A(n18713), .ZN(n18704) );
  AOI22_X1 U20704 ( .A1(n19012), .A2(n18704), .B1(n18761), .B2(n18703), .ZN(
        n19030) );
  AOI22_X1 U20705 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19030), .B1(
        n18759), .B2(n19046), .ZN(n18705) );
  OAI211_X1 U20706 ( .C1(n18766), .C2(n18969), .A(n18706), .B(n18705), .ZN(
        P3_U2971) );
  INV_X1 U20707 ( .A(n21199), .ZN(n20058) );
  INV_X1 U20708 ( .A(n18707), .ZN(n18708) );
  NOR2_X1 U20709 ( .A1(n20058), .A2(n18708), .ZN(n19033) );
  NAND2_X1 U20710 ( .A1(n21169), .A2(n21166), .ZN(n21171) );
  NOR2_X2 U20711 ( .A1(n21171), .A2(n18718), .ZN(n19052) );
  AOI22_X1 U20712 ( .A1(n18758), .A2(n19033), .B1(n18759), .B2(n19052), .ZN(
        n18711) );
  AOI21_X1 U20713 ( .B1(n21169), .B2(n18714), .A(n19011), .ZN(n18744) );
  NAND3_X1 U20714 ( .A1(n18719), .A2(n18744), .A3(n18709), .ZN(n19034) );
  AOI22_X1 U20715 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19034), .B1(
        n18763), .B2(n19046), .ZN(n18710) );
  OAI211_X1 U20716 ( .C1(n18766), .C2(n19027), .A(n18711), .B(n18710), .ZN(
        P3_U2963) );
  NOR2_X1 U20717 ( .A1(n20058), .A2(n18713), .ZN(n19039) );
  AOI22_X1 U20718 ( .A1(n18763), .A2(n19052), .B1(n18758), .B2(n19039), .ZN(
        n18717) );
  INV_X1 U20719 ( .A(n19011), .ZN(n18966) );
  NOR2_X1 U20720 ( .A1(n18712), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18727) );
  NAND2_X1 U20721 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18727), .ZN(
        n19044) );
  NAND2_X1 U20722 ( .A1(n18980), .A2(n19044), .ZN(n18724) );
  INV_X1 U20723 ( .A(n18724), .ZN(n18722) );
  OAI21_X1 U20724 ( .B1(n18722), .B2(n18714), .A(n18713), .ZN(n18715) );
  OAI211_X1 U20725 ( .C1(n19040), .C2(n21208), .A(n18966), .B(n18715), .ZN(
        n19041) );
  AOI22_X1 U20726 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19041), .B1(
        n18759), .B2(n19058), .ZN(n18716) );
  OAI211_X1 U20727 ( .C1(n18766), .C2(n18931), .A(n18717), .B(n18716), .ZN(
        P3_U2955) );
  INV_X1 U20728 ( .A(n19046), .ZN(n19038) );
  NAND2_X1 U20729 ( .A1(n21169), .A2(n21199), .ZN(n18752) );
  NOR2_X1 U20730 ( .A1(n18718), .A2(n18752), .ZN(n19045) );
  AOI22_X1 U20731 ( .A1(n18763), .A2(n19058), .B1(n18758), .B2(n19045), .ZN(
        n18721) );
  AND2_X1 U20732 ( .A1(n21169), .A2(n18729), .ZN(n18754) );
  AOI22_X1 U20733 ( .A1(n19012), .A2(n18727), .B1(n18719), .B2(n18754), .ZN(
        n19047) );
  NAND2_X1 U20734 ( .A1(n21166), .A2(n18727), .ZN(n19050) );
  AOI22_X1 U20735 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19047), .B1(
        n18759), .B2(n19063), .ZN(n18720) );
  OAI211_X1 U20736 ( .C1(n18766), .C2(n19038), .A(n18721), .B(n18720), .ZN(
        P3_U2947) );
  NOR2_X1 U20737 ( .A1(n20058), .A2(n18722), .ZN(n19051) );
  INV_X1 U20738 ( .A(n18723), .ZN(n18740) );
  NAND2_X1 U20739 ( .A1(n18740), .A2(n18737), .ZN(n19061) );
  INV_X1 U20740 ( .A(n19061), .ZN(n19069) );
  AOI22_X1 U20741 ( .A1(n18758), .A2(n19051), .B1(n18759), .B2(n19069), .ZN(
        n18726) );
  NAND2_X1 U20742 ( .A1(n19050), .A2(n19061), .ZN(n18733) );
  AOI22_X1 U20743 ( .A1(n19012), .A2(n18733), .B1(n18761), .B2(n18724), .ZN(
        n19053) );
  AOI22_X1 U20744 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19053), .B1(
        n18763), .B2(n19063), .ZN(n18725) );
  OAI211_X1 U20745 ( .C1(n18766), .C2(n18980), .A(n18726), .B(n18725), .ZN(
        P3_U2939) );
  INV_X1 U20746 ( .A(n18727), .ZN(n18728) );
  NOR2_X1 U20747 ( .A1(n20058), .A2(n18728), .ZN(n19056) );
  INV_X1 U20748 ( .A(n18737), .ZN(n18736) );
  NOR2_X2 U20749 ( .A1(n21171), .A2(n18736), .ZN(n19074) );
  AOI22_X1 U20750 ( .A1(n18758), .A2(n19056), .B1(n18759), .B2(n19074), .ZN(
        n18731) );
  OAI211_X1 U20751 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18732), .A(
        n18729), .B(n18737), .ZN(n19057) );
  AOI22_X1 U20752 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19057), .B1(
        n18763), .B2(n19069), .ZN(n18730) );
  OAI211_X1 U20753 ( .C1(n18766), .C2(n19044), .A(n18731), .B(n18730), .ZN(
        P3_U2931) );
  AND2_X1 U20754 ( .A1(n21199), .A2(n18733), .ZN(n19062) );
  NAND2_X1 U20755 ( .A1(n21174), .A2(n21175), .ZN(n18751) );
  NOR2_X1 U20756 ( .A1(n21169), .A2(n18751), .ZN(n18745) );
  NAND2_X1 U20757 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18745), .ZN(
        n19067) );
  AOI22_X1 U20758 ( .A1(n18758), .A2(n19062), .B1(n18759), .B2(n19081), .ZN(
        n18735) );
  NAND2_X1 U20759 ( .A1(n18989), .A2(n19067), .ZN(n18741) );
  OAI221_X1 U20760 ( .B1(n18733), .B2(n18732), .C1(n18733), .C2(n18741), .A(
        n18761), .ZN(n19064) );
  AOI22_X1 U20761 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19064), .B1(
        n18763), .B2(n19074), .ZN(n18734) );
  OAI211_X1 U20762 ( .C1(n18766), .C2(n19050), .A(n18735), .B(n18734), .ZN(
        P3_U2923) );
  NOR2_X1 U20763 ( .A1(n18752), .A2(n18736), .ZN(n19068) );
  NAND2_X1 U20764 ( .A1(n21166), .A2(n18745), .ZN(n19078) );
  AOI22_X1 U20765 ( .A1(n18758), .A2(n19068), .B1(n18759), .B2(n19086), .ZN(
        n18739) );
  AOI22_X1 U20766 ( .A1(n19012), .A2(n18745), .B1(n18754), .B2(n18737), .ZN(
        n19070) );
  AOI22_X1 U20767 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19070), .B1(
        n18763), .B2(n19081), .ZN(n18738) );
  OAI211_X1 U20768 ( .C1(n18766), .C2(n19061), .A(n18739), .B(n18738), .ZN(
        P3_U2915) );
  AND2_X1 U20769 ( .A1(n21199), .A2(n18741), .ZN(n19073) );
  INV_X1 U20770 ( .A(n18751), .ZN(n18753) );
  NAND2_X1 U20771 ( .A1(n18740), .A2(n18753), .ZN(n18908) );
  AOI22_X1 U20772 ( .A1(n18758), .A2(n19073), .B1(n18759), .B2(n19094), .ZN(
        n18743) );
  NAND2_X1 U20773 ( .A1(n19078), .A2(n18908), .ZN(n18748) );
  AOI22_X1 U20774 ( .A1(n19012), .A2(n18748), .B1(n18761), .B2(n18741), .ZN(
        n19075) );
  AOI22_X1 U20775 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19075), .B1(
        n18763), .B2(n19086), .ZN(n18742) );
  OAI211_X1 U20776 ( .C1(n18766), .C2(n18989), .A(n18743), .B(n18742), .ZN(
        P3_U2907) );
  OAI211_X1 U20777 ( .C1(n19081), .C2(n21208), .A(n18753), .B(n18744), .ZN(
        n19080) );
  AND2_X1 U20778 ( .A1(n21199), .A2(n18745), .ZN(n19079) );
  AOI22_X1 U20779 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19080), .B1(
        n18758), .B2(n19079), .ZN(n18747) );
  NOR2_X2 U20780 ( .A1(n21171), .A2(n18751), .ZN(n19104) );
  AOI22_X1 U20781 ( .A1(n18763), .A2(n19094), .B1(n18759), .B2(n19104), .ZN(
        n18746) );
  OAI211_X1 U20782 ( .C1(n18766), .C2(n19067), .A(n18747), .B(n18746), .ZN(
        P3_U2899) );
  INV_X1 U20783 ( .A(n18913), .ZN(n19093) );
  AND2_X1 U20784 ( .A1(n21199), .A2(n18748), .ZN(n19084) );
  AOI22_X1 U20785 ( .A1(n19093), .A2(n18759), .B1(n18758), .B2(n19084), .ZN(
        n18750) );
  NAND2_X1 U20786 ( .A1(n18913), .A2(n19091), .ZN(n18760) );
  AOI22_X1 U20787 ( .A1(n19012), .A2(n18760), .B1(n18761), .B2(n18748), .ZN(
        n19087) );
  AOI22_X1 U20788 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19087), .B1(
        n18763), .B2(n19104), .ZN(n18749) );
  OAI211_X1 U20789 ( .C1(n18766), .C2(n19078), .A(n18750), .B(n18749), .ZN(
        P3_U2891) );
  NOR2_X1 U20790 ( .A1(n18752), .A2(n18751), .ZN(n19092) );
  AOI22_X1 U20791 ( .A1(n18763), .A2(n19093), .B1(n18758), .B2(n19092), .ZN(
        n18757) );
  AOI22_X1 U20792 ( .A1(n19012), .A2(n18755), .B1(n18754), .B2(n18753), .ZN(
        n19095) );
  INV_X1 U20793 ( .A(n19098), .ZN(n19102) );
  AOI22_X1 U20794 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19095), .B1(
        n18759), .B2(n19102), .ZN(n18756) );
  OAI211_X1 U20795 ( .C1(n18766), .C2(n18908), .A(n18757), .B(n18756), .ZN(
        P3_U2883) );
  AND2_X1 U20796 ( .A1(n21199), .A2(n18760), .ZN(n19100) );
  AOI22_X1 U20797 ( .A1(n19023), .A2(n18759), .B1(n18758), .B2(n19100), .ZN(
        n18765) );
  AOI22_X1 U20798 ( .A1(n19012), .A2(n18762), .B1(n18761), .B2(n18760), .ZN(
        n19105) );
  AOI22_X1 U20799 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19105), .B1(
        n18763), .B2(n19102), .ZN(n18764) );
  OAI211_X1 U20800 ( .C1(n18766), .C2(n19091), .A(n18765), .B(n18764), .ZN(
        P3_U2875) );
  OAI22_X1 U20801 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19008), .ZN(n18767) );
  INV_X1 U20802 ( .A(n18767), .ZN(U257) );
  NAND2_X1 U20803 ( .A1(n18806), .A2(n20558), .ZN(n18804) );
  AND2_X1 U20804 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19012), .ZN(n18800) );
  NOR2_X2 U20805 ( .A1(n20534), .A2(n19011), .ZN(n18799) );
  AOI22_X1 U20806 ( .A1(n19023), .A2(n18800), .B1(n19013), .B2(n18799), .ZN(
        n18770) );
  INV_X1 U20807 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18768) );
  NOR2_X2 U20808 ( .A1(n18768), .A2(n18965), .ZN(n18801) );
  AOI22_X1 U20809 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19015), .B1(
        n19029), .B2(n18801), .ZN(n18769) );
  OAI211_X1 U20810 ( .C1(n18913), .C2(n18804), .A(n18770), .B(n18769), .ZN(
        P3_U2994) );
  AOI22_X1 U20811 ( .A1(n19029), .A2(n18800), .B1(n19018), .B2(n18799), .ZN(
        n18772) );
  AOI22_X1 U20812 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19019), .B1(
        n19035), .B2(n18801), .ZN(n18771) );
  OAI211_X1 U20813 ( .C1(n19098), .C2(n18804), .A(n18772), .B(n18771), .ZN(
        P3_U2986) );
  AOI22_X1 U20814 ( .A1(n19040), .A2(n18801), .B1(n19022), .B2(n18799), .ZN(
        n18774) );
  AOI22_X1 U20815 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19024), .B1(
        n19035), .B2(n18800), .ZN(n18773) );
  OAI211_X1 U20816 ( .C1(n19109), .C2(n18804), .A(n18774), .B(n18773), .ZN(
        P3_U2978) );
  AOI22_X1 U20817 ( .A1(n19040), .A2(n18800), .B1(n19028), .B2(n18799), .ZN(
        n18776) );
  AOI22_X1 U20818 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19030), .B1(
        n19046), .B2(n18801), .ZN(n18775) );
  OAI211_X1 U20819 ( .C1(n18969), .C2(n18804), .A(n18776), .B(n18775), .ZN(
        P3_U2970) );
  AOI22_X1 U20820 ( .A1(n19052), .A2(n18801), .B1(n19033), .B2(n18799), .ZN(
        n18778) );
  AOI22_X1 U20821 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19034), .B1(
        n19046), .B2(n18800), .ZN(n18777) );
  OAI211_X1 U20822 ( .C1(n19027), .C2(n18804), .A(n18778), .B(n18777), .ZN(
        P3_U2962) );
  AOI22_X1 U20823 ( .A1(n19058), .A2(n18801), .B1(n19039), .B2(n18799), .ZN(
        n18780) );
  AOI22_X1 U20824 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19041), .B1(
        n19052), .B2(n18800), .ZN(n18779) );
  OAI211_X1 U20825 ( .C1(n18931), .C2(n18804), .A(n18780), .B(n18779), .ZN(
        P3_U2954) );
  AOI22_X1 U20826 ( .A1(n19063), .A2(n18801), .B1(n19045), .B2(n18799), .ZN(
        n18782) );
  AOI22_X1 U20827 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19047), .B1(
        n19058), .B2(n18800), .ZN(n18781) );
  OAI211_X1 U20828 ( .C1(n19038), .C2(n18804), .A(n18782), .B(n18781), .ZN(
        P3_U2946) );
  AOI22_X1 U20829 ( .A1(n19063), .A2(n18800), .B1(n19051), .B2(n18799), .ZN(
        n18784) );
  AOI22_X1 U20830 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19053), .B1(
        n19069), .B2(n18801), .ZN(n18783) );
  OAI211_X1 U20831 ( .C1(n18980), .C2(n18804), .A(n18784), .B(n18783), .ZN(
        P3_U2938) );
  AOI22_X1 U20832 ( .A1(n19069), .A2(n18800), .B1(n19056), .B2(n18799), .ZN(
        n18786) );
  AOI22_X1 U20833 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19057), .B1(
        n19074), .B2(n18801), .ZN(n18785) );
  OAI211_X1 U20834 ( .C1(n19044), .C2(n18804), .A(n18786), .B(n18785), .ZN(
        P3_U2930) );
  AOI22_X1 U20835 ( .A1(n19081), .A2(n18801), .B1(n19062), .B2(n18799), .ZN(
        n18788) );
  AOI22_X1 U20836 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19064), .B1(
        n19074), .B2(n18800), .ZN(n18787) );
  OAI211_X1 U20837 ( .C1(n19050), .C2(n18804), .A(n18788), .B(n18787), .ZN(
        P3_U2922) );
  AOI22_X1 U20838 ( .A1(n19081), .A2(n18800), .B1(n19068), .B2(n18799), .ZN(
        n18790) );
  AOI22_X1 U20839 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19070), .B1(
        n19086), .B2(n18801), .ZN(n18789) );
  OAI211_X1 U20840 ( .C1(n19061), .C2(n18804), .A(n18790), .B(n18789), .ZN(
        P3_U2914) );
  AOI22_X1 U20841 ( .A1(n19086), .A2(n18800), .B1(n19073), .B2(n18799), .ZN(
        n18792) );
  AOI22_X1 U20842 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19075), .B1(
        n19094), .B2(n18801), .ZN(n18791) );
  OAI211_X1 U20843 ( .C1(n18989), .C2(n18804), .A(n18792), .B(n18791), .ZN(
        P3_U2906) );
  AOI22_X1 U20844 ( .A1(n19104), .A2(n18801), .B1(n19079), .B2(n18799), .ZN(
        n18794) );
  AOI22_X1 U20845 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19080), .B1(
        n19094), .B2(n18800), .ZN(n18793) );
  OAI211_X1 U20846 ( .C1(n19067), .C2(n18804), .A(n18794), .B(n18793), .ZN(
        P3_U2898) );
  AOI22_X1 U20847 ( .A1(n19093), .A2(n18801), .B1(n19084), .B2(n18799), .ZN(
        n18796) );
  AOI22_X1 U20848 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19087), .B1(
        n19104), .B2(n18800), .ZN(n18795) );
  OAI211_X1 U20849 ( .C1(n19078), .C2(n18804), .A(n18796), .B(n18795), .ZN(
        P3_U2890) );
  AOI22_X1 U20850 ( .A1(n19102), .A2(n18801), .B1(n19092), .B2(n18799), .ZN(
        n18798) );
  AOI22_X1 U20851 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19095), .B1(
        n19093), .B2(n18800), .ZN(n18797) );
  OAI211_X1 U20852 ( .C1(n18908), .C2(n18804), .A(n18798), .B(n18797), .ZN(
        P3_U2882) );
  AOI22_X1 U20853 ( .A1(n19102), .A2(n18800), .B1(n19100), .B2(n18799), .ZN(
        n18803) );
  AOI22_X1 U20854 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19105), .B1(
        n19023), .B2(n18801), .ZN(n18802) );
  OAI211_X1 U20855 ( .C1(n19091), .C2(n18804), .A(n18803), .B(n18802), .ZN(
        P3_U2874) );
  OAI22_X1 U20856 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19008), .ZN(n18805) );
  INV_X1 U20857 ( .A(n18805), .ZN(U256) );
  NAND2_X1 U20858 ( .A1(n18806), .A2(n20557), .ZN(n18842) );
  INV_X1 U20859 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20538) );
  NOR2_X2 U20860 ( .A1(n20538), .A2(n19011), .ZN(n18837) );
  INV_X1 U20861 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n20613) );
  NOR2_X2 U20862 ( .A1(n20613), .A2(n18965), .ZN(n18839) );
  AOI22_X1 U20863 ( .A1(n19013), .A2(n18837), .B1(n19029), .B2(n18839), .ZN(
        n18808) );
  NOR2_X2 U20864 ( .A1(n20559), .A2(n18965), .ZN(n18838) );
  AOI22_X1 U20865 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19015), .B1(
        n19023), .B2(n18838), .ZN(n18807) );
  OAI211_X1 U20866 ( .C1(n18913), .C2(n18842), .A(n18808), .B(n18807), .ZN(
        P3_U2993) );
  AOI22_X1 U20867 ( .A1(n19029), .A2(n18838), .B1(n19018), .B2(n18837), .ZN(
        n18810) );
  AOI22_X1 U20868 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19019), .B1(
        n19035), .B2(n18839), .ZN(n18809) );
  OAI211_X1 U20869 ( .C1(n19098), .C2(n18842), .A(n18810), .B(n18809), .ZN(
        P3_U2985) );
  AOI22_X1 U20870 ( .A1(n19035), .A2(n18838), .B1(n19022), .B2(n18837), .ZN(
        n18812) );
  AOI22_X1 U20871 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19024), .B1(
        n19040), .B2(n18839), .ZN(n18811) );
  OAI211_X1 U20872 ( .C1(n19109), .C2(n18842), .A(n18812), .B(n18811), .ZN(
        P3_U2977) );
  AOI22_X1 U20873 ( .A1(n19040), .A2(n18838), .B1(n19028), .B2(n18837), .ZN(
        n18814) );
  AOI22_X1 U20874 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19030), .B1(
        n19046), .B2(n18839), .ZN(n18813) );
  OAI211_X1 U20875 ( .C1(n18969), .C2(n18842), .A(n18814), .B(n18813), .ZN(
        P3_U2969) );
  AOI22_X1 U20876 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19034), .B1(
        n19033), .B2(n18837), .ZN(n18816) );
  AOI22_X1 U20877 ( .A1(n19046), .A2(n18838), .B1(n19052), .B2(n18839), .ZN(
        n18815) );
  OAI211_X1 U20878 ( .C1(n19027), .C2(n18842), .A(n18816), .B(n18815), .ZN(
        P3_U2961) );
  AOI22_X1 U20879 ( .A1(n19052), .A2(n18838), .B1(n19039), .B2(n18837), .ZN(
        n18818) );
  AOI22_X1 U20880 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19041), .B1(
        n19058), .B2(n18839), .ZN(n18817) );
  OAI211_X1 U20881 ( .C1(n18931), .C2(n18842), .A(n18818), .B(n18817), .ZN(
        P3_U2953) );
  AOI22_X1 U20882 ( .A1(n19058), .A2(n18838), .B1(n19045), .B2(n18837), .ZN(
        n18820) );
  AOI22_X1 U20883 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19047), .B1(
        n19063), .B2(n18839), .ZN(n18819) );
  OAI211_X1 U20884 ( .C1(n19038), .C2(n18842), .A(n18820), .B(n18819), .ZN(
        P3_U2945) );
  AOI22_X1 U20885 ( .A1(n19063), .A2(n18838), .B1(n19051), .B2(n18837), .ZN(
        n18822) );
  AOI22_X1 U20886 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19053), .B1(
        n19069), .B2(n18839), .ZN(n18821) );
  OAI211_X1 U20887 ( .C1(n18980), .C2(n18842), .A(n18822), .B(n18821), .ZN(
        P3_U2937) );
  AOI22_X1 U20888 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n18837), .ZN(n18824) );
  AOI22_X1 U20889 ( .A1(n19069), .A2(n18838), .B1(n19074), .B2(n18839), .ZN(
        n18823) );
  OAI211_X1 U20890 ( .C1(n19044), .C2(n18842), .A(n18824), .B(n18823), .ZN(
        P3_U2929) );
  AOI22_X1 U20891 ( .A1(n19074), .A2(n18838), .B1(n19062), .B2(n18837), .ZN(
        n18826) );
  AOI22_X1 U20892 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19064), .B1(
        n19081), .B2(n18839), .ZN(n18825) );
  OAI211_X1 U20893 ( .C1(n19050), .C2(n18842), .A(n18826), .B(n18825), .ZN(
        P3_U2921) );
  AOI22_X1 U20894 ( .A1(n19081), .A2(n18838), .B1(n19068), .B2(n18837), .ZN(
        n18828) );
  AOI22_X1 U20895 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19070), .B1(
        n19086), .B2(n18839), .ZN(n18827) );
  OAI211_X1 U20896 ( .C1(n19061), .C2(n18842), .A(n18828), .B(n18827), .ZN(
        P3_U2913) );
  AOI22_X1 U20897 ( .A1(n19086), .A2(n18838), .B1(n19073), .B2(n18837), .ZN(
        n18830) );
  AOI22_X1 U20898 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19075), .B1(
        n19094), .B2(n18839), .ZN(n18829) );
  OAI211_X1 U20899 ( .C1(n18989), .C2(n18842), .A(n18830), .B(n18829), .ZN(
        P3_U2905) );
  AOI22_X1 U20900 ( .A1(n19094), .A2(n18838), .B1(n19079), .B2(n18837), .ZN(
        n18832) );
  AOI22_X1 U20901 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19080), .B1(
        n19104), .B2(n18839), .ZN(n18831) );
  OAI211_X1 U20902 ( .C1(n19067), .C2(n18842), .A(n18832), .B(n18831), .ZN(
        P3_U2897) );
  AOI22_X1 U20903 ( .A1(n19093), .A2(n18839), .B1(n19084), .B2(n18837), .ZN(
        n18834) );
  AOI22_X1 U20904 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19087), .B1(
        n19104), .B2(n18838), .ZN(n18833) );
  OAI211_X1 U20905 ( .C1(n19078), .C2(n18842), .A(n18834), .B(n18833), .ZN(
        P3_U2889) );
  AOI22_X1 U20906 ( .A1(n19102), .A2(n18839), .B1(n19092), .B2(n18837), .ZN(
        n18836) );
  AOI22_X1 U20907 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19095), .B1(
        n19093), .B2(n18838), .ZN(n18835) );
  OAI211_X1 U20908 ( .C1(n18908), .C2(n18842), .A(n18836), .B(n18835), .ZN(
        P3_U2881) );
  AOI22_X1 U20909 ( .A1(n19102), .A2(n18838), .B1(n19100), .B2(n18837), .ZN(
        n18841) );
  AOI22_X1 U20910 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19105), .B1(
        n19023), .B2(n18839), .ZN(n18840) );
  OAI211_X1 U20911 ( .C1(n19091), .C2(n18842), .A(n18841), .B(n18840), .ZN(
        P3_U2873) );
  OAI22_X1 U20912 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19008), .ZN(n18843) );
  INV_X1 U20913 ( .A(n18843), .ZN(U255) );
  NAND2_X1 U20914 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19012), .ZN(n18875) );
  NOR2_X2 U20915 ( .A1(n20543), .A2(n19011), .ZN(n18876) );
  NAND2_X1 U20916 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19012), .ZN(n18881) );
  INV_X1 U20917 ( .A(n18881), .ZN(n18872) );
  AOI22_X1 U20918 ( .A1(n19013), .A2(n18876), .B1(n19029), .B2(n18872), .ZN(
        n18845) );
  NOR2_X2 U20919 ( .A1(n20748), .A2(n19014), .ZN(n18878) );
  AOI22_X1 U20920 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19015), .B1(
        n19093), .B2(n18878), .ZN(n18844) );
  OAI211_X1 U20921 ( .C1(n19109), .C2(n18875), .A(n18845), .B(n18844), .ZN(
        P3_U2992) );
  AOI22_X1 U20922 ( .A1(n19035), .A2(n18872), .B1(n19018), .B2(n18876), .ZN(
        n18847) );
  AOI22_X1 U20923 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19019), .B1(
        n19102), .B2(n18878), .ZN(n18846) );
  OAI211_X1 U20924 ( .C1(n18969), .C2(n18875), .A(n18847), .B(n18846), .ZN(
        P3_U2984) );
  AOI22_X1 U20925 ( .A1(n19040), .A2(n18872), .B1(n19022), .B2(n18876), .ZN(
        n18849) );
  AOI22_X1 U20926 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18878), .ZN(n18848) );
  OAI211_X1 U20927 ( .C1(n19027), .C2(n18875), .A(n18849), .B(n18848), .ZN(
        P3_U2976) );
  INV_X1 U20928 ( .A(n18875), .ZN(n18877) );
  AOI22_X1 U20929 ( .A1(n19040), .A2(n18877), .B1(n19028), .B2(n18876), .ZN(
        n18851) );
  AOI22_X1 U20930 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18878), .ZN(n18850) );
  OAI211_X1 U20931 ( .C1(n19038), .C2(n18881), .A(n18851), .B(n18850), .ZN(
        P3_U2968) );
  AOI22_X1 U20932 ( .A1(n19046), .A2(n18877), .B1(n19033), .B2(n18876), .ZN(
        n18853) );
  AOI22_X1 U20933 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19034), .B1(
        n19035), .B2(n18878), .ZN(n18852) );
  OAI211_X1 U20934 ( .C1(n18980), .C2(n18881), .A(n18853), .B(n18852), .ZN(
        P3_U2960) );
  AOI22_X1 U20935 ( .A1(n19058), .A2(n18872), .B1(n19039), .B2(n18876), .ZN(
        n18855) );
  AOI22_X1 U20936 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19041), .B1(
        n19040), .B2(n18878), .ZN(n18854) );
  OAI211_X1 U20937 ( .C1(n18980), .C2(n18875), .A(n18855), .B(n18854), .ZN(
        P3_U2952) );
  AOI22_X1 U20938 ( .A1(n19058), .A2(n18877), .B1(n19045), .B2(n18876), .ZN(
        n18857) );
  AOI22_X1 U20939 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19047), .B1(
        n19046), .B2(n18878), .ZN(n18856) );
  OAI211_X1 U20940 ( .C1(n19050), .C2(n18881), .A(n18857), .B(n18856), .ZN(
        P3_U2944) );
  AOI22_X1 U20941 ( .A1(n19063), .A2(n18877), .B1(n19051), .B2(n18876), .ZN(
        n18859) );
  AOI22_X1 U20942 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19053), .B1(
        n19052), .B2(n18878), .ZN(n18858) );
  OAI211_X1 U20943 ( .C1(n19061), .C2(n18881), .A(n18859), .B(n18858), .ZN(
        P3_U2936) );
  AOI22_X1 U20944 ( .A1(n19069), .A2(n18877), .B1(n19056), .B2(n18876), .ZN(
        n18861) );
  AOI22_X1 U20945 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19057), .B1(
        n19058), .B2(n18878), .ZN(n18860) );
  OAI211_X1 U20946 ( .C1(n18989), .C2(n18881), .A(n18861), .B(n18860), .ZN(
        P3_U2928) );
  AOI22_X1 U20947 ( .A1(n19081), .A2(n18872), .B1(n19062), .B2(n18876), .ZN(
        n18863) );
  AOI22_X1 U20948 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19064), .B1(
        n19063), .B2(n18878), .ZN(n18862) );
  OAI211_X1 U20949 ( .C1(n18989), .C2(n18875), .A(n18863), .B(n18862), .ZN(
        P3_U2920) );
  AOI22_X1 U20950 ( .A1(n19081), .A2(n18877), .B1(n19068), .B2(n18876), .ZN(
        n18865) );
  AOI22_X1 U20951 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19070), .B1(
        n19069), .B2(n18878), .ZN(n18864) );
  OAI211_X1 U20952 ( .C1(n19078), .C2(n18881), .A(n18865), .B(n18864), .ZN(
        P3_U2912) );
  AOI22_X1 U20953 ( .A1(n19094), .A2(n18872), .B1(n19073), .B2(n18876), .ZN(
        n18867) );
  AOI22_X1 U20954 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19075), .B1(
        n19074), .B2(n18878), .ZN(n18866) );
  OAI211_X1 U20955 ( .C1(n19078), .C2(n18875), .A(n18867), .B(n18866), .ZN(
        P3_U2904) );
  AOI22_X1 U20956 ( .A1(n19094), .A2(n18877), .B1(n19079), .B2(n18876), .ZN(
        n18869) );
  AOI22_X1 U20957 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19080), .B1(
        n19081), .B2(n18878), .ZN(n18868) );
  OAI211_X1 U20958 ( .C1(n19091), .C2(n18881), .A(n18869), .B(n18868), .ZN(
        P3_U2896) );
  AOI22_X1 U20959 ( .A1(n19104), .A2(n18877), .B1(n19084), .B2(n18876), .ZN(
        n18871) );
  AOI22_X1 U20960 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19087), .B1(
        n19086), .B2(n18878), .ZN(n18870) );
  OAI211_X1 U20961 ( .C1(n18913), .C2(n18881), .A(n18871), .B(n18870), .ZN(
        P3_U2888) );
  AOI22_X1 U20962 ( .A1(n19102), .A2(n18872), .B1(n19092), .B2(n18876), .ZN(
        n18874) );
  AOI22_X1 U20963 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18878), .ZN(n18873) );
  OAI211_X1 U20964 ( .C1(n18913), .C2(n18875), .A(n18874), .B(n18873), .ZN(
        P3_U2880) );
  AOI22_X1 U20965 ( .A1(n19102), .A2(n18877), .B1(n19100), .B2(n18876), .ZN(
        n18880) );
  AOI22_X1 U20966 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n18878), .ZN(n18879) );
  OAI211_X1 U20967 ( .C1(n19109), .C2(n18881), .A(n18880), .B(n18879), .ZN(
        P3_U2872) );
  OAI22_X1 U20968 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19008), .ZN(n18882) );
  INV_X1 U20969 ( .A(n18882), .ZN(U254) );
  NAND2_X1 U20970 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19012), .ZN(n18923) );
  AND2_X1 U20971 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18966), .ZN(n18918) );
  NAND2_X1 U20972 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19012), .ZN(n18917) );
  INV_X1 U20973 ( .A(n18917), .ZN(n18919) );
  AOI22_X1 U20974 ( .A1(n19013), .A2(n18918), .B1(n19029), .B2(n18919), .ZN(
        n18885) );
  NOR2_X2 U20975 ( .A1(n18883), .A2(n19014), .ZN(n18920) );
  AOI22_X1 U20976 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19015), .B1(
        n19093), .B2(n18920), .ZN(n18884) );
  OAI211_X1 U20977 ( .C1(n19109), .C2(n18923), .A(n18885), .B(n18884), .ZN(
        P3_U2991) );
  AOI22_X1 U20978 ( .A1(n19035), .A2(n18919), .B1(n19018), .B2(n18918), .ZN(
        n18887) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19019), .B1(
        n19102), .B2(n18920), .ZN(n18886) );
  OAI211_X1 U20980 ( .C1(n18969), .C2(n18923), .A(n18887), .B(n18886), .ZN(
        P3_U2983) );
  AOI22_X1 U20981 ( .A1(n19035), .A2(n18914), .B1(n19022), .B2(n18918), .ZN(
        n18889) );
  AOI22_X1 U20982 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18920), .ZN(n18888) );
  OAI211_X1 U20983 ( .C1(n18931), .C2(n18917), .A(n18889), .B(n18888), .ZN(
        P3_U2975) );
  AOI22_X1 U20984 ( .A1(n19046), .A2(n18919), .B1(n19028), .B2(n18918), .ZN(
        n18891) );
  AOI22_X1 U20985 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18920), .ZN(n18890) );
  OAI211_X1 U20986 ( .C1(n18931), .C2(n18923), .A(n18891), .B(n18890), .ZN(
        P3_U2967) );
  AOI22_X1 U20987 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19034), .B1(
        n19033), .B2(n18918), .ZN(n18893) );
  AOI22_X1 U20988 ( .A1(n19035), .A2(n18920), .B1(n19046), .B2(n18914), .ZN(
        n18892) );
  OAI211_X1 U20989 ( .C1(n18980), .C2(n18917), .A(n18893), .B(n18892), .ZN(
        P3_U2959) );
  AOI22_X1 U20990 ( .A1(n19058), .A2(n18919), .B1(n19039), .B2(n18918), .ZN(
        n18895) );
  AOI22_X1 U20991 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19041), .B1(
        n19040), .B2(n18920), .ZN(n18894) );
  OAI211_X1 U20992 ( .C1(n18980), .C2(n18923), .A(n18895), .B(n18894), .ZN(
        P3_U2951) );
  AOI22_X1 U20993 ( .A1(n19063), .A2(n18919), .B1(n19045), .B2(n18918), .ZN(
        n18897) );
  AOI22_X1 U20994 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19047), .B1(
        n19046), .B2(n18920), .ZN(n18896) );
  OAI211_X1 U20995 ( .C1(n19044), .C2(n18923), .A(n18897), .B(n18896), .ZN(
        P3_U2943) );
  AOI22_X1 U20996 ( .A1(n19069), .A2(n18919), .B1(n19051), .B2(n18918), .ZN(
        n18899) );
  AOI22_X1 U20997 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19053), .B1(
        n19052), .B2(n18920), .ZN(n18898) );
  OAI211_X1 U20998 ( .C1(n19050), .C2(n18923), .A(n18899), .B(n18898), .ZN(
        P3_U2935) );
  AOI22_X1 U20999 ( .A1(n19069), .A2(n18914), .B1(n19056), .B2(n18918), .ZN(
        n18901) );
  AOI22_X1 U21000 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19057), .B1(
        n19058), .B2(n18920), .ZN(n18900) );
  OAI211_X1 U21001 ( .C1(n18989), .C2(n18917), .A(n18901), .B(n18900), .ZN(
        P3_U2927) );
  AOI22_X1 U21002 ( .A1(n19081), .A2(n18919), .B1(n19062), .B2(n18918), .ZN(
        n18903) );
  AOI22_X1 U21003 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19064), .B1(
        n19063), .B2(n18920), .ZN(n18902) );
  OAI211_X1 U21004 ( .C1(n18989), .C2(n18923), .A(n18903), .B(n18902), .ZN(
        P3_U2919) );
  AOI22_X1 U21005 ( .A1(n19081), .A2(n18914), .B1(n19068), .B2(n18918), .ZN(
        n18905) );
  AOI22_X1 U21006 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19070), .B1(
        n19069), .B2(n18920), .ZN(n18904) );
  OAI211_X1 U21007 ( .C1(n19078), .C2(n18917), .A(n18905), .B(n18904), .ZN(
        P3_U2911) );
  AOI22_X1 U21008 ( .A1(n19086), .A2(n18914), .B1(n19073), .B2(n18918), .ZN(
        n18907) );
  AOI22_X1 U21009 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19075), .B1(
        n19074), .B2(n18920), .ZN(n18906) );
  OAI211_X1 U21010 ( .C1(n18908), .C2(n18917), .A(n18907), .B(n18906), .ZN(
        P3_U2903) );
  AOI22_X1 U21011 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n18918), .ZN(n18910) );
  AOI22_X1 U21012 ( .A1(n19081), .A2(n18920), .B1(n19094), .B2(n18914), .ZN(
        n18909) );
  OAI211_X1 U21013 ( .C1(n19091), .C2(n18917), .A(n18910), .B(n18909), .ZN(
        P3_U2895) );
  AOI22_X1 U21014 ( .A1(n19104), .A2(n18914), .B1(n19084), .B2(n18918), .ZN(
        n18912) );
  AOI22_X1 U21015 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19087), .B1(
        n19086), .B2(n18920), .ZN(n18911) );
  OAI211_X1 U21016 ( .C1(n18913), .C2(n18917), .A(n18912), .B(n18911), .ZN(
        P3_U2887) );
  AOI22_X1 U21017 ( .A1(n19093), .A2(n18914), .B1(n19092), .B2(n18918), .ZN(
        n18916) );
  AOI22_X1 U21018 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18920), .ZN(n18915) );
  OAI211_X1 U21019 ( .C1(n19098), .C2(n18917), .A(n18916), .B(n18915), .ZN(
        P3_U2879) );
  AOI22_X1 U21020 ( .A1(n19023), .A2(n18919), .B1(n19100), .B2(n18918), .ZN(
        n18922) );
  AOI22_X1 U21021 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n18920), .ZN(n18921) );
  OAI211_X1 U21022 ( .C1(n19098), .C2(n18923), .A(n18922), .B(n18921), .ZN(
        P3_U2871) );
  OAI22_X1 U21023 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19008), .ZN(n18924) );
  INV_X1 U21024 ( .A(n18924), .ZN(U253) );
  NAND2_X1 U21025 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19012), .ZN(n18957) );
  NAND2_X1 U21026 ( .A1(n19012), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18963) );
  INV_X1 U21027 ( .A(n18963), .ZN(n18954) );
  INV_X1 U21028 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20551) );
  NOR2_X2 U21029 ( .A1(n19011), .A2(n20551), .ZN(n18958) );
  AOI22_X1 U21030 ( .A1(n19023), .A2(n18954), .B1(n19013), .B2(n18958), .ZN(
        n18926) );
  NOR2_X2 U21031 ( .A1(n20746), .A2(n19014), .ZN(n18960) );
  AOI22_X1 U21032 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19015), .B1(
        n19093), .B2(n18960), .ZN(n18925) );
  OAI211_X1 U21033 ( .C1(n18969), .C2(n18957), .A(n18926), .B(n18925), .ZN(
        P3_U2990) );
  AOI22_X1 U21034 ( .A1(n19035), .A2(n18959), .B1(n19018), .B2(n18958), .ZN(
        n18928) );
  AOI22_X1 U21035 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19019), .B1(
        n19102), .B2(n18960), .ZN(n18927) );
  OAI211_X1 U21036 ( .C1(n18969), .C2(n18963), .A(n18928), .B(n18927), .ZN(
        P3_U2982) );
  AOI22_X1 U21037 ( .A1(n19035), .A2(n18954), .B1(n19022), .B2(n18958), .ZN(
        n18930) );
  AOI22_X1 U21038 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n18960), .ZN(n18929) );
  OAI211_X1 U21039 ( .C1(n18931), .C2(n18957), .A(n18930), .B(n18929), .ZN(
        P3_U2974) );
  AOI22_X1 U21040 ( .A1(n19040), .A2(n18954), .B1(n19028), .B2(n18958), .ZN(
        n18933) );
  AOI22_X1 U21041 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18960), .ZN(n18932) );
  OAI211_X1 U21042 ( .C1(n19038), .C2(n18957), .A(n18933), .B(n18932), .ZN(
        P3_U2966) );
  AOI22_X1 U21043 ( .A1(n19052), .A2(n18959), .B1(n19033), .B2(n18958), .ZN(
        n18935) );
  AOI22_X1 U21044 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19034), .B1(
        n19035), .B2(n18960), .ZN(n18934) );
  OAI211_X1 U21045 ( .C1(n19038), .C2(n18963), .A(n18935), .B(n18934), .ZN(
        P3_U2958) );
  AOI22_X1 U21046 ( .A1(n19058), .A2(n18959), .B1(n19039), .B2(n18958), .ZN(
        n18937) );
  AOI22_X1 U21047 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19041), .B1(
        n19040), .B2(n18960), .ZN(n18936) );
  OAI211_X1 U21048 ( .C1(n18980), .C2(n18963), .A(n18937), .B(n18936), .ZN(
        P3_U2950) );
  AOI22_X1 U21049 ( .A1(n19063), .A2(n18959), .B1(n19045), .B2(n18958), .ZN(
        n18939) );
  AOI22_X1 U21050 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19047), .B1(
        n19046), .B2(n18960), .ZN(n18938) );
  OAI211_X1 U21051 ( .C1(n19044), .C2(n18963), .A(n18939), .B(n18938), .ZN(
        P3_U2942) );
  AOI22_X1 U21052 ( .A1(n19069), .A2(n18959), .B1(n19051), .B2(n18958), .ZN(
        n18941) );
  AOI22_X1 U21053 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19053), .B1(
        n19052), .B2(n18960), .ZN(n18940) );
  OAI211_X1 U21054 ( .C1(n19050), .C2(n18963), .A(n18941), .B(n18940), .ZN(
        P3_U2934) );
  AOI22_X1 U21055 ( .A1(n19074), .A2(n18959), .B1(n19056), .B2(n18958), .ZN(
        n18943) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19057), .B1(
        n19058), .B2(n18960), .ZN(n18942) );
  OAI211_X1 U21057 ( .C1(n19061), .C2(n18963), .A(n18943), .B(n18942), .ZN(
        P3_U2926) );
  AOI22_X1 U21058 ( .A1(n19074), .A2(n18954), .B1(n19062), .B2(n18958), .ZN(
        n18945) );
  AOI22_X1 U21059 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19064), .B1(
        n19063), .B2(n18960), .ZN(n18944) );
  OAI211_X1 U21060 ( .C1(n19067), .C2(n18957), .A(n18945), .B(n18944), .ZN(
        P3_U2918) );
  AOI22_X1 U21061 ( .A1(n19086), .A2(n18959), .B1(n19068), .B2(n18958), .ZN(
        n18947) );
  AOI22_X1 U21062 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19070), .B1(
        n19069), .B2(n18960), .ZN(n18946) );
  OAI211_X1 U21063 ( .C1(n19067), .C2(n18963), .A(n18947), .B(n18946), .ZN(
        P3_U2910) );
  AOI22_X1 U21064 ( .A1(n19094), .A2(n18959), .B1(n19073), .B2(n18958), .ZN(
        n18949) );
  AOI22_X1 U21065 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19075), .B1(
        n19074), .B2(n18960), .ZN(n18948) );
  OAI211_X1 U21066 ( .C1(n19078), .C2(n18963), .A(n18949), .B(n18948), .ZN(
        P3_U2902) );
  AOI22_X1 U21067 ( .A1(n19094), .A2(n18954), .B1(n19079), .B2(n18958), .ZN(
        n18951) );
  AOI22_X1 U21068 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19080), .B1(
        n19081), .B2(n18960), .ZN(n18950) );
  OAI211_X1 U21069 ( .C1(n19091), .C2(n18957), .A(n18951), .B(n18950), .ZN(
        P3_U2894) );
  AOI22_X1 U21070 ( .A1(n19093), .A2(n18959), .B1(n19084), .B2(n18958), .ZN(
        n18953) );
  AOI22_X1 U21071 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19087), .B1(
        n19086), .B2(n18960), .ZN(n18952) );
  OAI211_X1 U21072 ( .C1(n19091), .C2(n18963), .A(n18953), .B(n18952), .ZN(
        P3_U2886) );
  AOI22_X1 U21073 ( .A1(n19093), .A2(n18954), .B1(n19092), .B2(n18958), .ZN(
        n18956) );
  AOI22_X1 U21074 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18960), .ZN(n18955) );
  OAI211_X1 U21075 ( .C1(n19098), .C2(n18957), .A(n18956), .B(n18955), .ZN(
        P3_U2878) );
  AOI22_X1 U21076 ( .A1(n19023), .A2(n18959), .B1(n19100), .B2(n18958), .ZN(
        n18962) );
  AOI22_X1 U21077 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n18960), .ZN(n18961) );
  OAI211_X1 U21078 ( .C1(n19098), .C2(n18963), .A(n18962), .B(n18961), .ZN(
        P3_U2870) );
  OAI22_X1 U21079 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19008), .ZN(n18964) );
  INV_X1 U21080 ( .A(n18964), .ZN(U252) );
  INV_X1 U21081 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n20596) );
  NOR2_X1 U21082 ( .A1(n20596), .A2(n18965), .ZN(n19003) );
  NAND2_X1 U21083 ( .A1(n19012), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19007) );
  INV_X1 U21084 ( .A(n19007), .ZN(n18998) );
  AND2_X1 U21085 ( .A1(n18966), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19002) );
  AOI22_X1 U21086 ( .A1(n19023), .A2(n18998), .B1(n19013), .B2(n19002), .ZN(
        n18968) );
  NOR2_X2 U21087 ( .A1(n20063), .A2(n19014), .ZN(n19004) );
  AOI22_X1 U21088 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19015), .B1(
        n19093), .B2(n19004), .ZN(n18967) );
  OAI211_X1 U21089 ( .C1(n18969), .C2(n19001), .A(n18968), .B(n18967), .ZN(
        P3_U2989) );
  AOI22_X1 U21090 ( .A1(n19029), .A2(n18998), .B1(n19018), .B2(n19002), .ZN(
        n18971) );
  AOI22_X1 U21091 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19019), .B1(
        n19102), .B2(n19004), .ZN(n18970) );
  OAI211_X1 U21092 ( .C1(n19027), .C2(n19001), .A(n18971), .B(n18970), .ZN(
        P3_U2981) );
  AOI22_X1 U21093 ( .A1(n19040), .A2(n19003), .B1(n19022), .B2(n19002), .ZN(
        n18973) );
  AOI22_X1 U21094 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n19004), .ZN(n18972) );
  OAI211_X1 U21095 ( .C1(n19027), .C2(n19007), .A(n18973), .B(n18972), .ZN(
        P3_U2973) );
  AOI22_X1 U21096 ( .A1(n19040), .A2(n18998), .B1(n19028), .B2(n19002), .ZN(
        n18975) );
  AOI22_X1 U21097 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n19004), .ZN(n18974) );
  OAI211_X1 U21098 ( .C1(n19038), .C2(n19001), .A(n18975), .B(n18974), .ZN(
        P3_U2965) );
  AOI22_X1 U21099 ( .A1(n19046), .A2(n18998), .B1(n19033), .B2(n19002), .ZN(
        n18977) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19034), .B1(
        n19035), .B2(n19004), .ZN(n18976) );
  OAI211_X1 U21101 ( .C1(n18980), .C2(n19001), .A(n18977), .B(n18976), .ZN(
        P3_U2957) );
  AOI22_X1 U21102 ( .A1(n19058), .A2(n19003), .B1(n19039), .B2(n19002), .ZN(
        n18979) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19041), .B1(
        n19040), .B2(n19004), .ZN(n18978) );
  OAI211_X1 U21104 ( .C1(n18980), .C2(n19007), .A(n18979), .B(n18978), .ZN(
        P3_U2949) );
  AOI22_X1 U21105 ( .A1(n19063), .A2(n19003), .B1(n19045), .B2(n19002), .ZN(
        n18982) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19047), .B1(
        n19046), .B2(n19004), .ZN(n18981) );
  OAI211_X1 U21107 ( .C1(n19044), .C2(n19007), .A(n18982), .B(n18981), .ZN(
        P3_U2941) );
  AOI22_X1 U21108 ( .A1(n19069), .A2(n19003), .B1(n19051), .B2(n19002), .ZN(
        n18984) );
  AOI22_X1 U21109 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19053), .B1(
        n19052), .B2(n19004), .ZN(n18983) );
  OAI211_X1 U21110 ( .C1(n19050), .C2(n19007), .A(n18984), .B(n18983), .ZN(
        P3_U2933) );
  AOI22_X1 U21111 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n19002), .ZN(n18986) );
  AOI22_X1 U21112 ( .A1(n19058), .A2(n19004), .B1(n19069), .B2(n18998), .ZN(
        n18985) );
  OAI211_X1 U21113 ( .C1(n18989), .C2(n19001), .A(n18986), .B(n18985), .ZN(
        P3_U2925) );
  AOI22_X1 U21114 ( .A1(n19081), .A2(n19003), .B1(n19062), .B2(n19002), .ZN(
        n18988) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19064), .B1(
        n19063), .B2(n19004), .ZN(n18987) );
  OAI211_X1 U21116 ( .C1(n18989), .C2(n19007), .A(n18988), .B(n18987), .ZN(
        P3_U2917) );
  AOI22_X1 U21117 ( .A1(n19081), .A2(n18998), .B1(n19068), .B2(n19002), .ZN(
        n18991) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19070), .B1(
        n19069), .B2(n19004), .ZN(n18990) );
  OAI211_X1 U21119 ( .C1(n19078), .C2(n19001), .A(n18991), .B(n18990), .ZN(
        P3_U2909) );
  AOI22_X1 U21120 ( .A1(n19094), .A2(n19003), .B1(n19073), .B2(n19002), .ZN(
        n18993) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19075), .B1(
        n19074), .B2(n19004), .ZN(n18992) );
  OAI211_X1 U21122 ( .C1(n19078), .C2(n19007), .A(n18993), .B(n18992), .ZN(
        P3_U2901) );
  AOI22_X1 U21123 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n19002), .ZN(n18995) );
  AOI22_X1 U21124 ( .A1(n19081), .A2(n19004), .B1(n19094), .B2(n18998), .ZN(
        n18994) );
  OAI211_X1 U21125 ( .C1(n19091), .C2(n19001), .A(n18995), .B(n18994), .ZN(
        P3_U2893) );
  AOI22_X1 U21126 ( .A1(n19093), .A2(n19003), .B1(n19084), .B2(n19002), .ZN(
        n18997) );
  AOI22_X1 U21127 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19087), .B1(
        n19086), .B2(n19004), .ZN(n18996) );
  OAI211_X1 U21128 ( .C1(n19091), .C2(n19007), .A(n18997), .B(n18996), .ZN(
        P3_U2885) );
  AOI22_X1 U21129 ( .A1(n19093), .A2(n18998), .B1(n19092), .B2(n19002), .ZN(
        n19000) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19004), .ZN(n18999) );
  OAI211_X1 U21131 ( .C1(n19098), .C2(n19001), .A(n19000), .B(n18999), .ZN(
        P3_U2877) );
  AOI22_X1 U21132 ( .A1(n19023), .A2(n19003), .B1(n19100), .B2(n19002), .ZN(
        n19006) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19004), .ZN(n19005) );
  OAI211_X1 U21134 ( .C1(n19098), .C2(n19007), .A(n19006), .B(n19005), .ZN(
        P3_U2869) );
  OAI22_X1 U21135 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19008), .ZN(n19010) );
  INV_X1 U21136 ( .A(n19010), .ZN(U251) );
  NAND2_X1 U21137 ( .A1(n19012), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19090) );
  INV_X1 U21138 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n20677) );
  NOR2_X2 U21139 ( .A1(n19011), .A2(n20677), .ZN(n19099) );
  NAND2_X1 U21140 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19012), .ZN(n19108) );
  INV_X1 U21141 ( .A(n19108), .ZN(n19085) );
  AOI22_X1 U21142 ( .A1(n19013), .A2(n19099), .B1(n19029), .B2(n19085), .ZN(
        n19017) );
  NOR2_X2 U21143 ( .A1(n20055), .A2(n19014), .ZN(n19103) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19015), .B1(
        n19093), .B2(n19103), .ZN(n19016) );
  OAI211_X1 U21145 ( .C1(n19109), .C2(n19090), .A(n19017), .B(n19016), .ZN(
        P3_U2988) );
  INV_X1 U21146 ( .A(n19090), .ZN(n19101) );
  AOI22_X1 U21147 ( .A1(n19029), .A2(n19101), .B1(n19018), .B2(n19099), .ZN(
        n19021) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19019), .B1(
        n19102), .B2(n19103), .ZN(n19020) );
  OAI211_X1 U21149 ( .C1(n19027), .C2(n19108), .A(n19021), .B(n19020), .ZN(
        P3_U2980) );
  AOI22_X1 U21150 ( .A1(n19040), .A2(n19085), .B1(n19022), .B2(n19099), .ZN(
        n19026) );
  AOI22_X1 U21151 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19024), .B1(
        n19023), .B2(n19103), .ZN(n19025) );
  OAI211_X1 U21152 ( .C1(n19027), .C2(n19090), .A(n19026), .B(n19025), .ZN(
        P3_U2972) );
  AOI22_X1 U21153 ( .A1(n19040), .A2(n19101), .B1(n19028), .B2(n19099), .ZN(
        n19032) );
  AOI22_X1 U21154 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n19103), .ZN(n19031) );
  OAI211_X1 U21155 ( .C1(n19038), .C2(n19108), .A(n19032), .B(n19031), .ZN(
        P3_U2964) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19034), .B1(
        n19033), .B2(n19099), .ZN(n19037) );
  AOI22_X1 U21157 ( .A1(n19035), .A2(n19103), .B1(n19052), .B2(n19085), .ZN(
        n19036) );
  OAI211_X1 U21158 ( .C1(n19038), .C2(n19090), .A(n19037), .B(n19036), .ZN(
        P3_U2956) );
  AOI22_X1 U21159 ( .A1(n19052), .A2(n19101), .B1(n19039), .B2(n19099), .ZN(
        n19043) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19041), .B1(
        n19040), .B2(n19103), .ZN(n19042) );
  OAI211_X1 U21161 ( .C1(n19044), .C2(n19108), .A(n19043), .B(n19042), .ZN(
        P3_U2948) );
  AOI22_X1 U21162 ( .A1(n19058), .A2(n19101), .B1(n19045), .B2(n19099), .ZN(
        n19049) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19047), .B1(
        n19046), .B2(n19103), .ZN(n19048) );
  OAI211_X1 U21164 ( .C1(n19050), .C2(n19108), .A(n19049), .B(n19048), .ZN(
        P3_U2940) );
  AOI22_X1 U21165 ( .A1(n19063), .A2(n19101), .B1(n19051), .B2(n19099), .ZN(
        n19055) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19053), .B1(
        n19052), .B2(n19103), .ZN(n19054) );
  OAI211_X1 U21167 ( .C1(n19061), .C2(n19108), .A(n19055), .B(n19054), .ZN(
        P3_U2932) );
  AOI22_X1 U21168 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n19099), .ZN(n19060) );
  AOI22_X1 U21169 ( .A1(n19058), .A2(n19103), .B1(n19074), .B2(n19085), .ZN(
        n19059) );
  OAI211_X1 U21170 ( .C1(n19061), .C2(n19090), .A(n19060), .B(n19059), .ZN(
        P3_U2924) );
  AOI22_X1 U21171 ( .A1(n19074), .A2(n19101), .B1(n19062), .B2(n19099), .ZN(
        n19066) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19064), .B1(
        n19063), .B2(n19103), .ZN(n19065) );
  OAI211_X1 U21173 ( .C1(n19067), .C2(n19108), .A(n19066), .B(n19065), .ZN(
        P3_U2916) );
  AOI22_X1 U21174 ( .A1(n19081), .A2(n19101), .B1(n19068), .B2(n19099), .ZN(
        n19072) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19070), .B1(
        n19069), .B2(n19103), .ZN(n19071) );
  OAI211_X1 U21176 ( .C1(n19078), .C2(n19108), .A(n19072), .B(n19071), .ZN(
        P3_U2908) );
  AOI22_X1 U21177 ( .A1(n19094), .A2(n19085), .B1(n19073), .B2(n19099), .ZN(
        n19077) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19075), .B1(
        n19074), .B2(n19103), .ZN(n19076) );
  OAI211_X1 U21179 ( .C1(n19078), .C2(n19090), .A(n19077), .B(n19076), .ZN(
        P3_U2900) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n19099), .ZN(n19083) );
  AOI22_X1 U21181 ( .A1(n19081), .A2(n19103), .B1(n19094), .B2(n19101), .ZN(
        n19082) );
  OAI211_X1 U21182 ( .C1(n19091), .C2(n19108), .A(n19083), .B(n19082), .ZN(
        P3_U2892) );
  AOI22_X1 U21183 ( .A1(n19093), .A2(n19085), .B1(n19084), .B2(n19099), .ZN(
        n19089) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19087), .B1(
        n19086), .B2(n19103), .ZN(n19088) );
  OAI211_X1 U21185 ( .C1(n19091), .C2(n19090), .A(n19089), .B(n19088), .ZN(
        P3_U2884) );
  AOI22_X1 U21186 ( .A1(n19093), .A2(n19101), .B1(n19092), .B2(n19099), .ZN(
        n19097) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19103), .ZN(n19096) );
  OAI211_X1 U21188 ( .C1(n19098), .C2(n19108), .A(n19097), .B(n19096), .ZN(
        P3_U2876) );
  AOI22_X1 U21189 ( .A1(n19102), .A2(n19101), .B1(n19100), .B2(n19099), .ZN(
        n19107) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19103), .ZN(n19106) );
  OAI211_X1 U21191 ( .C1(n19109), .C2(n19108), .A(n19107), .B(n19106), .ZN(
        P3_U2868) );
  AOI22_X1 U21192 ( .A1(n19110), .A2(n19585), .B1(n19582), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19112) );
  AOI22_X1 U21193 ( .A1(n19583), .A2(BUF1_REG_31__SCAN_IN), .B1(n19579), .B2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n19111) );
  NAND2_X1 U21194 ( .A1(n19112), .A2(n19111), .ZN(P2_U2888) );
  AOI22_X1 U21195 ( .A1(n19489), .A2(n19113), .B1(n19579), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n19114) );
  OAI21_X1 U21196 ( .B1(n19348), .B2(n19115), .A(n19114), .ZN(P2_U2908) );
  AOI22_X1 U21197 ( .A1(n19489), .A2(n19116), .B1(n19579), .B2(
        P2_EAX_REG_10__SCAN_IN), .ZN(n19117) );
  OAI21_X1 U21198 ( .B1(n19348), .B2(n19118), .A(n19117), .ZN(P2_U2909) );
  NAND3_X1 U21199 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19131) );
  OAI21_X1 U21200 ( .B1(n19121), .B2(n19595), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19122) );
  OAI21_X1 U21201 ( .B1(n19131), .B2(n19276), .A(n19122), .ZN(n19596) );
  INV_X1 U21202 ( .A(n19226), .ZN(n19291) );
  AOI22_X1 U21203 ( .A1(n19596), .A2(n14780), .B1(n19595), .B2(n19291), .ZN(
        n19130) );
  OAI21_X1 U21204 ( .B1(n19124), .B2(n19123), .A(n19131), .ZN(n19128) );
  OAI21_X1 U21205 ( .B1(n19282), .B2(n19595), .A(n19281), .ZN(n19125) );
  OAI21_X1 U21206 ( .B1(n19126), .B2(n19284), .A(n19125), .ZN(n19127) );
  NAND2_X1 U21207 ( .A1(n19128), .A2(n19127), .ZN(n19599) );
  AOI22_X1 U21208 ( .A1(n19705), .A2(n19292), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19129) );
  OAI211_X1 U21209 ( .C1(n19271), .C2(n19544), .A(n19130), .B(n19129), .ZN(
        P2_U3175) );
  INV_X1 U21210 ( .A(n19292), .ZN(n19290) );
  NOR2_X1 U21211 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19131), .ZN(
        n19603) );
  AOI22_X1 U21212 ( .A1(n19500), .A2(n19293), .B1(n19291), .B2(n19603), .ZN(
        n19142) );
  NAND2_X1 U21213 ( .A1(n19544), .A2(n19614), .ZN(n19132) );
  AOI21_X1 U21214 ( .B1(n19132), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19276), 
        .ZN(n19137) );
  AOI21_X1 U21215 ( .B1(n19138), .B2(n19133), .A(n19231), .ZN(n19134) );
  AOI21_X1 U21216 ( .B1(n19137), .B2(n19135), .A(n19134), .ZN(n19136) );
  AOI21_X1 U21217 ( .B1(n19603), .B2(n19281), .A(n19136), .ZN(n19606) );
  OAI21_X1 U21218 ( .B1(n19603), .B2(n19609), .A(n19137), .ZN(n19140) );
  OAI21_X1 U21219 ( .B1(n19138), .B2(n19603), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19139) );
  NAND2_X1 U21220 ( .A1(n19140), .A2(n19139), .ZN(n19605) );
  AOI22_X1 U21221 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19606), .B1(
        n14780), .B2(n19605), .ZN(n19141) );
  OAI211_X1 U21222 ( .C1(n19290), .C2(n19544), .A(n19142), .B(n19141), .ZN(
        P2_U3167) );
  INV_X1 U21223 ( .A(n19223), .ZN(n19143) );
  INV_X1 U21224 ( .A(n19144), .ZN(n19151) );
  INV_X1 U21225 ( .A(n19145), .ZN(n19147) );
  NAND2_X1 U21226 ( .A1(n19147), .A2(n19146), .ZN(n19229) );
  NOR2_X1 U21227 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19148), .ZN(
        n19615) );
  OAI21_X1 U21228 ( .B1(n19149), .B2(n19615), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19150) );
  OAI21_X1 U21229 ( .B1(n19151), .B2(n19229), .A(n19150), .ZN(n19616) );
  AOI22_X1 U21230 ( .A1(n19616), .A2(n14780), .B1(n19291), .B2(n19615), .ZN(
        n19159) );
  INV_X1 U21231 ( .A(n19615), .ZN(n19152) );
  AOI21_X1 U21232 ( .B1(n19152), .B2(n19276), .A(n19591), .ZN(n19157) );
  NOR2_X1 U21233 ( .A1(n12711), .A2(n19284), .ZN(n19156) );
  OAI21_X1 U21234 ( .B1(n19625), .B2(n19617), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19153) );
  OAI21_X1 U21235 ( .B1(n19229), .B2(n19154), .A(n19153), .ZN(n19155) );
  AOI22_X1 U21236 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19292), .B2(n19617), .ZN(n19158) );
  OAI211_X1 U21237 ( .C1(n19271), .C2(n19621), .A(n19159), .B(n19158), .ZN(
        P2_U3151) );
  NAND3_X1 U21238 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19172), .ZN(n19169) );
  NOR2_X1 U21239 ( .A1(n19274), .A2(n19169), .ZN(n19622) );
  OAI21_X1 U21240 ( .B1(n19160), .B2(n19622), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19161) );
  OAI21_X1 U21241 ( .B1(n19169), .B2(n19276), .A(n19161), .ZN(n19623) );
  AOI22_X1 U21242 ( .A1(n19623), .A2(n14780), .B1(n19291), .B2(n19622), .ZN(
        n19168) );
  OAI21_X1 U21243 ( .B1(n19162), .B2(n19244), .A(n19169), .ZN(n19166) );
  OAI21_X1 U21244 ( .B1(n19282), .B2(n19622), .A(n19281), .ZN(n19163) );
  OAI21_X1 U21245 ( .B1(n19164), .B2(n19284), .A(n19163), .ZN(n19165) );
  NAND2_X1 U21246 ( .A1(n19166), .A2(n19165), .ZN(n19624) );
  AOI22_X1 U21247 ( .A1(n19625), .A2(n19292), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n19624), .ZN(n19167) );
  OAI211_X1 U21248 ( .C1(n19271), .C2(n19628), .A(n19168), .B(n19167), .ZN(
        P2_U3143) );
  NOR2_X1 U21249 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19169), .ZN(
        n19629) );
  INV_X1 U21250 ( .A(n19629), .ZN(n19359) );
  OAI22_X1 U21251 ( .A1(n19628), .A2(n19290), .B1(n19226), .B2(n19359), .ZN(
        n19170) );
  INV_X1 U21252 ( .A(n19170), .ZN(n19181) );
  OAI21_X1 U21253 ( .B1(n19630), .B2(n19553), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19171) );
  NAND2_X1 U21254 ( .A1(n19171), .A2(n19282), .ZN(n19179) );
  NAND3_X1 U21255 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19272), .A3(
        n19172), .ZN(n19197) );
  NOR2_X1 U21256 ( .A1(n19274), .A2(n19197), .ZN(n19635) );
  NOR2_X1 U21257 ( .A1(n19635), .A2(n19629), .ZN(n19178) );
  INV_X1 U21258 ( .A(n19178), .ZN(n19176) );
  AOI21_X1 U21259 ( .B1(n12615), .B2(n19262), .A(n19629), .ZN(n19174) );
  NOR2_X1 U21260 ( .A1(n19174), .A2(n19591), .ZN(n19175) );
  OAI22_X1 U21261 ( .A1(n19179), .A2(n19176), .B1(n19231), .B2(n19175), .ZN(
        n19632) );
  OAI21_X1 U21262 ( .B1(n12615), .B2(n19629), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19177) );
  AOI22_X1 U21263 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19632), .B1(
        n14780), .B2(n19631), .ZN(n19180) );
  OAI211_X1 U21264 ( .C1(n19271), .C2(n19641), .A(n19181), .B(n19180), .ZN(
        P2_U3135) );
  INV_X1 U21265 ( .A(n19182), .ZN(n19183) );
  AOI22_X1 U21266 ( .A1(n19636), .A2(n19293), .B1(n19291), .B2(n19635), .ZN(
        n19194) );
  OAI21_X1 U21267 ( .B1(n19185), .B2(n19278), .A(n19282), .ZN(n19192) );
  INV_X1 U21268 ( .A(n19197), .ZN(n19189) );
  AOI21_X1 U21269 ( .B1(n19635), .B2(n19281), .A(n19231), .ZN(n19186) );
  OAI21_X1 U21270 ( .B1(n19187), .B2(n19284), .A(n19186), .ZN(n19188) );
  OAI21_X1 U21271 ( .B1(n19192), .B2(n19189), .A(n19188), .ZN(n19638) );
  OAI21_X1 U21272 ( .B1(n19190), .B2(n19635), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19191) );
  OAI21_X1 U21273 ( .B1(n19192), .B2(n19197), .A(n19191), .ZN(n19637) );
  AOI22_X1 U21274 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19638), .B1(
        n14780), .B2(n19637), .ZN(n19193) );
  OAI211_X1 U21275 ( .C1(n19290), .C2(n19641), .A(n19194), .B(n19193), .ZN(
        P2_U3127) );
  INV_X1 U21276 ( .A(n19212), .ZN(n19196) );
  NOR2_X1 U21277 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19197), .ZN(
        n19513) );
  INV_X1 U21278 ( .A(n19513), .ZN(n19643) );
  OAI22_X1 U21279 ( .A1(n19655), .A2(n19271), .B1(n19226), .B2(n19643), .ZN(
        n19198) );
  INV_X1 U21280 ( .A(n19198), .ZN(n19207) );
  AOI21_X1 U21281 ( .B1(n19655), .B2(n19649), .A(n21569), .ZN(n19199) );
  NOR2_X1 U21282 ( .A1(n19199), .A2(n19276), .ZN(n19202) );
  OAI21_X1 U21283 ( .B1(n19203), .B2(n19263), .A(n19262), .ZN(n19200) );
  AOI21_X1 U21284 ( .B1(n19202), .B2(n19209), .A(n19200), .ZN(n19201) );
  OAI21_X1 U21285 ( .B1(n19513), .B2(n19201), .A(n19281), .ZN(n19646) );
  INV_X1 U21286 ( .A(n19209), .ZN(n19650) );
  OAI21_X1 U21287 ( .B1(n19650), .B2(n19513), .A(n19202), .ZN(n19205) );
  OAI21_X1 U21288 ( .B1(n19203), .B2(n19513), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19204) );
  NAND2_X1 U21289 ( .A1(n19205), .A2(n19204), .ZN(n19645) );
  AOI22_X1 U21290 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n14780), .ZN(n19206) );
  OAI211_X1 U21291 ( .C1(n19290), .C2(n19649), .A(n19207), .B(n19206), .ZN(
        P2_U3119) );
  NOR2_X1 U21292 ( .A1(n19208), .A2(n19650), .ZN(n19210) );
  OAI22_X1 U21293 ( .A1(n19210), .A2(n19263), .B1(n19211), .B2(n19276), .ZN(
        n19651) );
  AOI22_X1 U21294 ( .A1(n19651), .A2(n14780), .B1(n19650), .B2(n19291), .ZN(
        n19216) );
  OAI22_X1 U21295 ( .A1(n19210), .A2(n19284), .B1(n19591), .B2(n19209), .ZN(
        n19214) );
  OAI21_X1 U21296 ( .B1(n21569), .B2(n19212), .A(n19211), .ZN(n19213) );
  OAI21_X1 U21297 ( .B1(n19231), .B2(n19214), .A(n19213), .ZN(n19652) );
  AOI22_X1 U21298 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19293), .ZN(n19215) );
  OAI211_X1 U21299 ( .C1(n19290), .C2(n19655), .A(n19216), .B(n19215), .ZN(
        P2_U3111) );
  INV_X1 U21300 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U21301 ( .A1(n19657), .A2(n14780), .B1(n19656), .B2(n19291), .ZN(
        n19218) );
  AOI22_X1 U21302 ( .A1(n19659), .A2(n19293), .B1(n19658), .B2(n19292), .ZN(
        n19217) );
  OAI211_X1 U21303 ( .C1(n19663), .C2(n19219), .A(n19218), .B(n19217), .ZN(
        P2_U3103) );
  AOI22_X1 U21304 ( .A1(n19671), .A2(n19293), .B1(n19664), .B2(n19291), .ZN(
        n19221) );
  AOI22_X1 U21305 ( .A1(n14780), .A2(n19665), .B1(n19659), .B2(n19292), .ZN(
        n19220) );
  OAI211_X1 U21306 ( .C1(n19524), .C2(n19222), .A(n19221), .B(n19220), .ZN(
        P2_U3095) );
  NAND2_X1 U21307 ( .A1(n19225), .A2(n19224), .ZN(n19375) );
  OAI22_X1 U21308 ( .A1(n19564), .A2(n19290), .B1(n19226), .B2(n19375), .ZN(
        n19227) );
  INV_X1 U21309 ( .A(n19227), .ZN(n19241) );
  OAI21_X1 U21310 ( .B1(n19678), .B2(n19671), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19228) );
  NAND2_X1 U21311 ( .A1(n19228), .A2(n19282), .ZN(n19239) );
  NOR2_X1 U21312 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19229), .ZN(
        n19235) );
  INV_X1 U21313 ( .A(n19236), .ZN(n19230) );
  NOR2_X1 U21314 ( .A1(n19230), .A2(n19284), .ZN(n19234) );
  INV_X1 U21315 ( .A(n19231), .ZN(n19232) );
  OAI21_X1 U21316 ( .B1(n19591), .B2(n19375), .A(n19232), .ZN(n19233) );
  INV_X1 U21317 ( .A(n19235), .ZN(n19238) );
  INV_X1 U21318 ( .A(n19375), .ZN(n19670) );
  OAI21_X1 U21319 ( .B1(n19236), .B2(n19670), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19237) );
  AOI22_X1 U21320 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19673), .B1(
        n14780), .B2(n19672), .ZN(n19240) );
  OAI211_X1 U21321 ( .C1(n19271), .C2(n19676), .A(n19241), .B(n19240), .ZN(
        P2_U3087) );
  AND2_X1 U21322 ( .A1(n19243), .A2(n19273), .ZN(n19677) );
  AOI22_X1 U21323 ( .A1(n19686), .A2(n19293), .B1(n19291), .B2(n19677), .ZN(
        n19255) );
  NOR2_X1 U21324 ( .A1(n19245), .A2(n19244), .ZN(n19253) );
  NAND2_X1 U21325 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19273), .ZN(
        n19258) );
  INV_X1 U21326 ( .A(n19258), .ZN(n19249) );
  INV_X1 U21327 ( .A(n19250), .ZN(n19247) );
  OAI21_X1 U21328 ( .B1(n19282), .B2(n19677), .A(n19281), .ZN(n19246) );
  OAI21_X1 U21329 ( .B1(n19247), .B2(n19284), .A(n19246), .ZN(n19248) );
  OAI21_X1 U21330 ( .B1(n19253), .B2(n19249), .A(n19248), .ZN(n19680) );
  NAND2_X1 U21331 ( .A1(n19282), .A2(n19249), .ZN(n19252) );
  OAI21_X1 U21332 ( .B1(n19250), .B2(n19677), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19251) );
  OAI21_X1 U21333 ( .B1(n19253), .B2(n19252), .A(n19251), .ZN(n19679) );
  AOI22_X1 U21334 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n14780), .ZN(n19254) );
  OAI211_X1 U21335 ( .C1(n19290), .C2(n19676), .A(n19255), .B(n19254), .ZN(
        P2_U3079) );
  NOR2_X1 U21336 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19258), .ZN(
        n19684) );
  OAI21_X1 U21337 ( .B1(n19264), .B2(n19684), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19260) );
  NAND3_X1 U21338 ( .A1(n19259), .A2(n19282), .A3(n19273), .ZN(n19261) );
  NAND2_X1 U21339 ( .A1(n19260), .A2(n19261), .ZN(n19685) );
  AOI22_X1 U21340 ( .A1(n19685), .A2(n14780), .B1(n19291), .B2(n19684), .ZN(
        n19270) );
  OAI221_X1 U21341 ( .B1(n21569), .B2(n19696), .C1(n21569), .C2(n19683), .A(
        n19261), .ZN(n19268) );
  OAI21_X1 U21342 ( .B1(n19264), .B2(n19263), .A(n19262), .ZN(n19266) );
  INV_X1 U21343 ( .A(n19684), .ZN(n19265) );
  AOI21_X1 U21344 ( .B1(n19266), .B2(n19265), .A(n19591), .ZN(n19267) );
  AOI22_X1 U21345 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19292), .ZN(n19269) );
  OAI211_X1 U21346 ( .C1(n19271), .C2(n19696), .A(n19270), .B(n19269), .ZN(
        P2_U3071) );
  NAND2_X1 U21347 ( .A1(n19273), .A2(n19272), .ZN(n19277) );
  NOR2_X1 U21348 ( .A1(n19274), .A2(n19277), .ZN(n19691) );
  OAI21_X1 U21349 ( .B1(n19280), .B2(n19691), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19275) );
  OAI21_X1 U21350 ( .B1(n19277), .B2(n19276), .A(n19275), .ZN(n19692) );
  AOI22_X1 U21351 ( .A1(n19692), .A2(n14780), .B1(n19291), .B2(n19691), .ZN(
        n19289) );
  OAI21_X1 U21352 ( .B1(n19279), .B2(n19278), .A(n19277), .ZN(n19287) );
  INV_X1 U21353 ( .A(n19280), .ZN(n19285) );
  OAI21_X1 U21354 ( .B1(n19282), .B2(n19691), .A(n19281), .ZN(n19283) );
  OAI21_X1 U21355 ( .B1(n19285), .B2(n19284), .A(n19283), .ZN(n19286) );
  NAND2_X1 U21356 ( .A1(n19287), .A2(n19286), .ZN(n19693) );
  AOI22_X1 U21357 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19293), .ZN(n19288) );
  OAI211_X1 U21358 ( .C1(n19290), .C2(n19696), .A(n19289), .B(n19288), .ZN(
        P2_U3063) );
  AOI22_X1 U21359 ( .A1(n19701), .A2(n19292), .B1(n19699), .B2(n19291), .ZN(
        n19295) );
  AOI22_X1 U21360 ( .A1(n14780), .A2(n19703), .B1(n19705), .B2(n19293), .ZN(
        n19294) );
  OAI211_X1 U21361 ( .C1(n19709), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        P2_U3055) );
  AOI22_X1 U21362 ( .A1(n19581), .A2(n19297), .B1(n19579), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n19303) );
  AOI22_X1 U21363 ( .A1(n19583), .A2(BUF1_REG_22__SCAN_IN), .B1(n19582), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n19302) );
  INV_X1 U21364 ( .A(n19298), .ZN(n19300) );
  AOI22_X1 U21365 ( .A1(n19300), .A2(n19586), .B1(n19585), .B2(n19299), .ZN(
        n19301) );
  NAND3_X1 U21366 ( .A1(n19303), .A2(n19302), .A3(n19301), .ZN(P2_U2897) );
  AOI22_X1 U21367 ( .A1(n19596), .A2(n14755), .B1(n19335), .B2(n19595), .ZN(
        n19305) );
  INV_X1 U21368 ( .A(n19544), .ZN(n19604) );
  AOI22_X1 U21369 ( .A1(n19604), .A2(n19336), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n19304) );
  OAI211_X1 U21370 ( .C1(n19334), .C2(n19602), .A(n19305), .B(n19304), .ZN(
        P2_U3174) );
  AOI22_X1 U21371 ( .A1(n19604), .A2(n19337), .B1(n19335), .B2(n19603), .ZN(
        n19307) );
  AOI22_X1 U21372 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19606), .B1(
        n14755), .B2(n19605), .ZN(n19306) );
  OAI211_X1 U21373 ( .C1(n19331), .C2(n19614), .A(n19307), .B(n19306), .ZN(
        P2_U3166) );
  AOI22_X1 U21374 ( .A1(n19616), .A2(n14755), .B1(n19335), .B2(n19615), .ZN(
        n19309) );
  AOI22_X1 U21375 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n19617), .B2(n19337), .ZN(n19308) );
  OAI211_X1 U21376 ( .C1(n19331), .C2(n19621), .A(n19309), .B(n19308), .ZN(
        P2_U3150) );
  AOI22_X1 U21377 ( .A1(n19623), .A2(n14755), .B1(n19335), .B2(n19622), .ZN(
        n19311) );
  AOI22_X1 U21378 ( .A1(n19625), .A2(n19337), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n19624), .ZN(n19310) );
  OAI211_X1 U21379 ( .C1(n19331), .C2(n19628), .A(n19311), .B(n19310), .ZN(
        P2_U3142) );
  AOI22_X1 U21380 ( .A1(n19630), .A2(n19337), .B1(n19335), .B2(n19629), .ZN(
        n19313) );
  AOI22_X1 U21381 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19632), .B1(
        n14755), .B2(n19631), .ZN(n19312) );
  OAI211_X1 U21382 ( .C1(n19331), .C2(n19641), .A(n19313), .B(n19312), .ZN(
        P2_U3134) );
  AOI22_X1 U21383 ( .A1(n19636), .A2(n19336), .B1(n19335), .B2(n19635), .ZN(
        n19315) );
  AOI22_X1 U21384 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19638), .B1(
        n14755), .B2(n19637), .ZN(n19314) );
  OAI211_X1 U21385 ( .C1(n19334), .C2(n19641), .A(n19315), .B(n19314), .ZN(
        P2_U3126) );
  OAI22_X1 U21386 ( .A1(n19655), .A2(n19331), .B1(n19316), .B2(n19643), .ZN(
        n19317) );
  INV_X1 U21387 ( .A(n19317), .ZN(n19319) );
  AOI22_X1 U21388 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n14755), .ZN(n19318) );
  OAI211_X1 U21389 ( .C1(n19334), .C2(n19649), .A(n19319), .B(n19318), .ZN(
        P2_U3118) );
  AOI22_X1 U21390 ( .A1(n19651), .A2(n14755), .B1(n19650), .B2(n19335), .ZN(
        n19321) );
  AOI22_X1 U21391 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19336), .ZN(n19320) );
  OAI211_X1 U21392 ( .C1(n19334), .C2(n19655), .A(n19321), .B(n19320), .ZN(
        P2_U3110) );
  INV_X1 U21393 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n19324) );
  AOI22_X1 U21394 ( .A1(n19671), .A2(n19336), .B1(n19335), .B2(n19664), .ZN(
        n19323) );
  AOI22_X1 U21395 ( .A1(n14755), .A2(n19665), .B1(n19659), .B2(n19337), .ZN(
        n19322) );
  OAI211_X1 U21396 ( .C1(n19524), .C2(n19324), .A(n19323), .B(n19322), .ZN(
        P2_U3094) );
  AOI22_X1 U21397 ( .A1(n19671), .A2(n19337), .B1(n19335), .B2(n19670), .ZN(
        n19326) );
  AOI22_X1 U21398 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19673), .B1(
        n14755), .B2(n19672), .ZN(n19325) );
  OAI211_X1 U21399 ( .C1(n19331), .C2(n19676), .A(n19326), .B(n19325), .ZN(
        P2_U3086) );
  AOI22_X1 U21400 ( .A1(n19686), .A2(n19336), .B1(n19335), .B2(n19677), .ZN(
        n19328) );
  AOI22_X1 U21401 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n14755), .ZN(n19327) );
  OAI211_X1 U21402 ( .C1(n19334), .C2(n19676), .A(n19328), .B(n19327), .ZN(
        P2_U3078) );
  AOI22_X1 U21403 ( .A1(n19685), .A2(n14755), .B1(n19335), .B2(n19684), .ZN(
        n19330) );
  AOI22_X1 U21404 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19337), .ZN(n19329) );
  OAI211_X1 U21405 ( .C1(n19331), .C2(n19696), .A(n19330), .B(n19329), .ZN(
        P2_U3070) );
  AOI22_X1 U21406 ( .A1(n19692), .A2(n14755), .B1(n19335), .B2(n19691), .ZN(
        n19333) );
  AOI22_X1 U21407 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19336), .ZN(n19332) );
  OAI211_X1 U21408 ( .C1(n19334), .C2(n19696), .A(n19333), .B(n19332), .ZN(
        P2_U3062) );
  AOI22_X1 U21409 ( .A1(n19705), .A2(n19336), .B1(n19335), .B2(n19699), .ZN(
        n19339) );
  AOI22_X1 U21410 ( .A1(n19701), .A2(n19337), .B1(n19703), .B2(n14755), .ZN(
        n19338) );
  OAI211_X1 U21411 ( .C1(n19709), .C2(n19340), .A(n19339), .B(n19338), .ZN(
        P2_U3054) );
  AOI22_X1 U21412 ( .A1(n19489), .A2(n19341), .B1(n19579), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n19346) );
  OR3_X1 U21413 ( .A1(n19344), .A2(n19343), .A3(n19342), .ZN(n19345) );
  OAI211_X1 U21414 ( .C1(n19348), .C2(n19347), .A(n19346), .B(n19345), .ZN(
        P2_U2914) );
  AOI22_X1 U21415 ( .A1(n19596), .A2(n14600), .B1(n19595), .B2(n19388), .ZN(
        n19350) );
  AOI22_X1 U21416 ( .A1(n19604), .A2(n19389), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n19349) );
  OAI211_X1 U21417 ( .C1(n19392), .C2(n19602), .A(n19350), .B(n19349), .ZN(
        P2_U3173) );
  AOI22_X1 U21418 ( .A1(n19500), .A2(n19389), .B1(n19388), .B2(n19603), .ZN(
        n19352) );
  AOI22_X1 U21419 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19606), .B1(
        n14600), .B2(n19605), .ZN(n19351) );
  OAI211_X1 U21420 ( .C1(n19392), .C2(n19544), .A(n19352), .B(n19351), .ZN(
        P2_U3165) );
  AOI22_X1 U21421 ( .A1(n19610), .A2(n14600), .B1(n19388), .B2(n19609), .ZN(
        n19354) );
  AOI22_X1 U21422 ( .A1(n19611), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n19617), .B2(n19389), .ZN(n19353) );
  OAI211_X1 U21423 ( .C1(n19392), .C2(n19614), .A(n19354), .B(n19353), .ZN(
        P2_U3157) );
  AOI22_X1 U21424 ( .A1(n19616), .A2(n14600), .B1(n19388), .B2(n19615), .ZN(
        n19356) );
  AOI22_X1 U21425 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n19617), .B2(n19384), .ZN(n19355) );
  OAI211_X1 U21426 ( .C1(n19387), .C2(n19621), .A(n19356), .B(n19355), .ZN(
        P2_U3149) );
  AOI22_X1 U21427 ( .A1(n19623), .A2(n14600), .B1(n19388), .B2(n19622), .ZN(
        n19358) );
  AOI22_X1 U21428 ( .A1(n19630), .A2(n19389), .B1(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n19624), .ZN(n19357) );
  OAI211_X1 U21429 ( .C1(n19392), .C2(n19621), .A(n19358), .B(n19357), .ZN(
        P2_U3141) );
  OAI22_X1 U21430 ( .A1(n19628), .A2(n19392), .B1(n19380), .B2(n19359), .ZN(
        n19360) );
  INV_X1 U21431 ( .A(n19360), .ZN(n19362) );
  AOI22_X1 U21432 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19632), .B1(
        n14600), .B2(n19631), .ZN(n19361) );
  OAI211_X1 U21433 ( .C1(n19387), .C2(n19641), .A(n19362), .B(n19361), .ZN(
        P2_U3133) );
  INV_X1 U21434 ( .A(n19635), .ZN(n19363) );
  OAI22_X1 U21435 ( .A1(n19641), .A2(n19392), .B1(n19380), .B2(n19363), .ZN(
        n19364) );
  INV_X1 U21436 ( .A(n19364), .ZN(n19366) );
  AOI22_X1 U21437 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19638), .B1(
        n14600), .B2(n19637), .ZN(n19365) );
  OAI211_X1 U21438 ( .C1(n19387), .C2(n19649), .A(n19366), .B(n19365), .ZN(
        P2_U3125) );
  OAI22_X1 U21439 ( .A1(n19655), .A2(n19387), .B1(n19380), .B2(n19643), .ZN(
        n19367) );
  INV_X1 U21440 ( .A(n19367), .ZN(n19369) );
  AOI22_X1 U21441 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n14600), .ZN(n19368) );
  OAI211_X1 U21442 ( .C1(n19392), .C2(n19649), .A(n19369), .B(n19368), .ZN(
        P2_U3117) );
  AOI22_X1 U21443 ( .A1(n19651), .A2(n14600), .B1(n19650), .B2(n19388), .ZN(
        n19371) );
  AOI22_X1 U21444 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19389), .ZN(n19370) );
  OAI211_X1 U21445 ( .C1(n19392), .C2(n19655), .A(n19371), .B(n19370), .ZN(
        P2_U3109) );
  INV_X1 U21446 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n19374) );
  AOI22_X1 U21447 ( .A1(n19657), .A2(n14600), .B1(n19656), .B2(n19388), .ZN(
        n19373) );
  AOI22_X1 U21448 ( .A1(n19659), .A2(n19389), .B1(n19658), .B2(n19384), .ZN(
        n19372) );
  OAI211_X1 U21449 ( .C1(n19663), .C2(n19374), .A(n19373), .B(n19372), .ZN(
        P2_U3101) );
  OAI22_X1 U21450 ( .A1(n19564), .A2(n19392), .B1(n19380), .B2(n19375), .ZN(
        n19376) );
  INV_X1 U21451 ( .A(n19376), .ZN(n19378) );
  AOI22_X1 U21452 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19673), .B1(
        n14600), .B2(n19672), .ZN(n19377) );
  OAI211_X1 U21453 ( .C1(n19387), .C2(n19676), .A(n19378), .B(n19377), .ZN(
        P2_U3085) );
  INV_X1 U21454 ( .A(n19677), .ZN(n19379) );
  OAI22_X1 U21455 ( .A1(n19676), .A2(n19392), .B1(n19380), .B2(n19379), .ZN(
        n19381) );
  INV_X1 U21456 ( .A(n19381), .ZN(n19383) );
  AOI22_X1 U21457 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n14600), .ZN(n19382) );
  OAI211_X1 U21458 ( .C1(n19387), .C2(n19683), .A(n19383), .B(n19382), .ZN(
        P2_U3077) );
  AOI22_X1 U21459 ( .A1(n19685), .A2(n14600), .B1(n19388), .B2(n19684), .ZN(
        n19386) );
  AOI22_X1 U21460 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19384), .ZN(n19385) );
  OAI211_X1 U21461 ( .C1(n19387), .C2(n19696), .A(n19386), .B(n19385), .ZN(
        P2_U3069) );
  AOI22_X1 U21462 ( .A1(n19692), .A2(n14600), .B1(n19388), .B2(n19691), .ZN(
        n19391) );
  AOI22_X1 U21463 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19389), .ZN(n19390) );
  OAI211_X1 U21464 ( .C1(n19392), .C2(n19696), .A(n19391), .B(n19390), .ZN(
        P2_U3061) );
  AOI22_X1 U21465 ( .A1(n19581), .A2(n19393), .B1(n19579), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n19399) );
  AOI22_X1 U21466 ( .A1(n19583), .A2(BUF1_REG_20__SCAN_IN), .B1(n19582), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n19398) );
  INV_X1 U21467 ( .A(n19394), .ZN(n19395) );
  AOI22_X1 U21468 ( .A1(n19396), .A2(n19586), .B1(n19585), .B2(n19395), .ZN(
        n19397) );
  NAND3_X1 U21469 ( .A1(n19399), .A2(n19398), .A3(n19397), .ZN(P2_U2899) );
  AOI22_X1 U21470 ( .A1(n19596), .A2(n14749), .B1(n19431), .B2(n19595), .ZN(
        n19401) );
  AOI22_X1 U21471 ( .A1(n19705), .A2(n19427), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19400) );
  OAI211_X1 U21472 ( .C1(n19430), .C2(n19544), .A(n19401), .B(n19400), .ZN(
        P2_U3172) );
  AOI22_X1 U21473 ( .A1(n19500), .A2(n19432), .B1(n19431), .B2(n19603), .ZN(
        n19403) );
  AOI22_X1 U21474 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19606), .B1(
        n14749), .B2(n19605), .ZN(n19402) );
  OAI211_X1 U21475 ( .C1(n19435), .C2(n19544), .A(n19403), .B(n19402), .ZN(
        P2_U3164) );
  AOI22_X1 U21476 ( .A1(n19610), .A2(n14749), .B1(n19431), .B2(n19609), .ZN(
        n19405) );
  AOI22_X1 U21477 ( .A1(n19611), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n19617), .B2(n19432), .ZN(n19404) );
  OAI211_X1 U21478 ( .C1(n19435), .C2(n19614), .A(n19405), .B(n19404), .ZN(
        P2_U3156) );
  AOI22_X1 U21479 ( .A1(n19616), .A2(n14749), .B1(n19431), .B2(n19615), .ZN(
        n19407) );
  AOI22_X1 U21480 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n19617), .B2(n19427), .ZN(n19406) );
  OAI211_X1 U21481 ( .C1(n19430), .C2(n19621), .A(n19407), .B(n19406), .ZN(
        P2_U3148) );
  AOI22_X1 U21482 ( .A1(n19623), .A2(n14749), .B1(n19431), .B2(n19622), .ZN(
        n19409) );
  AOI22_X1 U21483 ( .A1(n19630), .A2(n19432), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n19624), .ZN(n19408) );
  OAI211_X1 U21484 ( .C1(n19435), .C2(n19621), .A(n19409), .B(n19408), .ZN(
        P2_U3140) );
  AOI22_X1 U21485 ( .A1(n19630), .A2(n19427), .B1(n19431), .B2(n19629), .ZN(
        n19411) );
  AOI22_X1 U21486 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19632), .B1(
        n14749), .B2(n19631), .ZN(n19410) );
  OAI211_X1 U21487 ( .C1(n19430), .C2(n19641), .A(n19411), .B(n19410), .ZN(
        P2_U3132) );
  AOI22_X1 U21488 ( .A1(n19636), .A2(n19432), .B1(n19431), .B2(n19635), .ZN(
        n19413) );
  AOI22_X1 U21489 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19638), .B1(
        n14749), .B2(n19637), .ZN(n19412) );
  OAI211_X1 U21490 ( .C1(n19435), .C2(n19641), .A(n19413), .B(n19412), .ZN(
        P2_U3124) );
  INV_X1 U21491 ( .A(n19431), .ZN(n19414) );
  OAI22_X1 U21492 ( .A1(n19655), .A2(n19430), .B1(n19414), .B2(n19643), .ZN(
        n19415) );
  INV_X1 U21493 ( .A(n19415), .ZN(n19417) );
  AOI22_X1 U21494 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n14749), .ZN(n19416) );
  OAI211_X1 U21495 ( .C1(n19435), .C2(n19649), .A(n19417), .B(n19416), .ZN(
        P2_U3116) );
  AOI22_X1 U21496 ( .A1(n19651), .A2(n14749), .B1(n19650), .B2(n19431), .ZN(
        n19419) );
  AOI22_X1 U21497 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19432), .ZN(n19418) );
  OAI211_X1 U21498 ( .C1(n19435), .C2(n19655), .A(n19419), .B(n19418), .ZN(
        P2_U3108) );
  INV_X1 U21499 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19422) );
  AOI22_X1 U21500 ( .A1(n19671), .A2(n19432), .B1(n19431), .B2(n19664), .ZN(
        n19421) );
  AOI22_X1 U21501 ( .A1(n14749), .A2(n19665), .B1(n19659), .B2(n19427), .ZN(
        n19420) );
  OAI211_X1 U21502 ( .C1(n19524), .C2(n19422), .A(n19421), .B(n19420), .ZN(
        P2_U3092) );
  AOI22_X1 U21503 ( .A1(n19671), .A2(n19427), .B1(n19431), .B2(n19670), .ZN(
        n19424) );
  AOI22_X1 U21504 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19673), .B1(
        n14749), .B2(n19672), .ZN(n19423) );
  OAI211_X1 U21505 ( .C1(n19430), .C2(n19676), .A(n19424), .B(n19423), .ZN(
        P2_U3084) );
  AOI22_X1 U21506 ( .A1(n19686), .A2(n19432), .B1(n19431), .B2(n19677), .ZN(
        n19426) );
  AOI22_X1 U21507 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n14749), .ZN(n19425) );
  OAI211_X1 U21508 ( .C1(n19435), .C2(n19676), .A(n19426), .B(n19425), .ZN(
        P2_U3076) );
  AOI22_X1 U21509 ( .A1(n19685), .A2(n14749), .B1(n19431), .B2(n19684), .ZN(
        n19429) );
  AOI22_X1 U21510 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19427), .ZN(n19428) );
  OAI211_X1 U21511 ( .C1(n19430), .C2(n19696), .A(n19429), .B(n19428), .ZN(
        P2_U3068) );
  AOI22_X1 U21512 ( .A1(n19692), .A2(n14749), .B1(n19431), .B2(n19691), .ZN(
        n19434) );
  AOI22_X1 U21513 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19432), .ZN(n19433) );
  OAI211_X1 U21514 ( .C1(n19435), .C2(n19696), .A(n19434), .B(n19433), .ZN(
        P2_U3060) );
  NOR2_X2 U21515 ( .A1(n19436), .A2(n19591), .ZN(n19476) );
  NAND2_X1 U21516 ( .A1(n19437), .A2(n19593), .ZN(n19452) );
  AOI22_X1 U21517 ( .A1(n19596), .A2(n19476), .B1(n19595), .B2(n19474), .ZN(
        n19439) );
  AOI22_X1 U21518 ( .A1(n19604), .A2(n19477), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n19438) );
  OAI211_X1 U21519 ( .C1(n19473), .C2(n19602), .A(n19439), .B(n19438), .ZN(
        P2_U3171) );
  AOI22_X1 U21520 ( .A1(n19604), .A2(n19475), .B1(n19474), .B2(n19603), .ZN(
        n19441) );
  AOI22_X1 U21521 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19606), .B1(
        n19476), .B2(n19605), .ZN(n19440) );
  OAI211_X1 U21522 ( .C1(n19470), .C2(n19614), .A(n19441), .B(n19440), .ZN(
        P2_U3163) );
  AOI22_X1 U21523 ( .A1(n19610), .A2(n19476), .B1(n19609), .B2(n19474), .ZN(
        n19443) );
  AOI22_X1 U21524 ( .A1(n19611), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n19617), .B2(n19477), .ZN(n19442) );
  OAI211_X1 U21525 ( .C1(n19473), .C2(n19614), .A(n19443), .B(n19442), .ZN(
        P2_U3155) );
  AOI22_X1 U21526 ( .A1(n19616), .A2(n19476), .B1(n19474), .B2(n19615), .ZN(
        n19445) );
  AOI22_X1 U21527 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n19617), .B2(n19475), .ZN(n19444) );
  OAI211_X1 U21528 ( .C1(n19470), .C2(n19621), .A(n19445), .B(n19444), .ZN(
        P2_U3147) );
  AOI22_X1 U21529 ( .A1(n19623), .A2(n19476), .B1(n19474), .B2(n19622), .ZN(
        n19447) );
  AOI22_X1 U21530 ( .A1(n19630), .A2(n19477), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n19624), .ZN(n19446) );
  OAI211_X1 U21531 ( .C1(n19473), .C2(n19621), .A(n19447), .B(n19446), .ZN(
        P2_U3139) );
  AOI22_X1 U21532 ( .A1(n19553), .A2(n19477), .B1(n19474), .B2(n19629), .ZN(
        n19449) );
  AOI22_X1 U21533 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19632), .B1(
        n19476), .B2(n19631), .ZN(n19448) );
  OAI211_X1 U21534 ( .C1(n19473), .C2(n19628), .A(n19449), .B(n19448), .ZN(
        P2_U3131) );
  AOI22_X1 U21535 ( .A1(n19636), .A2(n19477), .B1(n19474), .B2(n19635), .ZN(
        n19451) );
  AOI22_X1 U21536 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19638), .B1(
        n19476), .B2(n19637), .ZN(n19450) );
  OAI211_X1 U21537 ( .C1(n19473), .C2(n19641), .A(n19451), .B(n19450), .ZN(
        P2_U3123) );
  OAI22_X1 U21538 ( .A1(n19655), .A2(n19470), .B1(n19643), .B2(n19452), .ZN(
        n19453) );
  INV_X1 U21539 ( .A(n19453), .ZN(n19455) );
  AOI22_X1 U21540 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19476), .ZN(n19454) );
  OAI211_X1 U21541 ( .C1(n19473), .C2(n19649), .A(n19455), .B(n19454), .ZN(
        P2_U3115) );
  AOI22_X1 U21542 ( .A1(n19651), .A2(n19476), .B1(n19650), .B2(n19474), .ZN(
        n19457) );
  AOI22_X1 U21543 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19477), .ZN(n19456) );
  OAI211_X1 U21544 ( .C1(n19473), .C2(n19655), .A(n19457), .B(n19456), .ZN(
        P2_U3107) );
  INV_X1 U21545 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n19460) );
  AOI22_X1 U21546 ( .A1(n19657), .A2(n19476), .B1(n19656), .B2(n19474), .ZN(
        n19459) );
  AOI22_X1 U21547 ( .A1(n19659), .A2(n19477), .B1(n19658), .B2(n19475), .ZN(
        n19458) );
  OAI211_X1 U21548 ( .C1(n19663), .C2(n19460), .A(n19459), .B(n19458), .ZN(
        P2_U3099) );
  INV_X1 U21549 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n19463) );
  AOI22_X1 U21550 ( .A1(n19671), .A2(n19477), .B1(n19664), .B2(n19474), .ZN(
        n19462) );
  AOI22_X1 U21551 ( .A1(n19476), .A2(n19665), .B1(n19659), .B2(n19475), .ZN(
        n19461) );
  OAI211_X1 U21552 ( .C1(n19524), .C2(n19463), .A(n19462), .B(n19461), .ZN(
        P2_U3091) );
  AOI22_X1 U21553 ( .A1(n19671), .A2(n19475), .B1(n19474), .B2(n19670), .ZN(
        n19465) );
  AOI22_X1 U21554 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19673), .B1(
        n19476), .B2(n19672), .ZN(n19464) );
  OAI211_X1 U21555 ( .C1(n19470), .C2(n19676), .A(n19465), .B(n19464), .ZN(
        P2_U3083) );
  AOI22_X1 U21556 ( .A1(n19678), .A2(n19475), .B1(n19474), .B2(n19677), .ZN(
        n19467) );
  AOI22_X1 U21557 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n19476), .ZN(n19466) );
  OAI211_X1 U21558 ( .C1(n19470), .C2(n19683), .A(n19467), .B(n19466), .ZN(
        P2_U3075) );
  AOI22_X1 U21559 ( .A1(n19685), .A2(n19476), .B1(n19474), .B2(n19684), .ZN(
        n19469) );
  AOI22_X1 U21560 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19475), .ZN(n19468) );
  OAI211_X1 U21561 ( .C1(n19470), .C2(n19696), .A(n19469), .B(n19468), .ZN(
        P2_U3067) );
  AOI22_X1 U21562 ( .A1(n19692), .A2(n19476), .B1(n19474), .B2(n19691), .ZN(
        n19472) );
  AOI22_X1 U21563 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19477), .ZN(n19471) );
  OAI211_X1 U21564 ( .C1(n19473), .C2(n19696), .A(n19472), .B(n19471), .ZN(
        P2_U3059) );
  AOI22_X1 U21565 ( .A1(n19701), .A2(n19475), .B1(n19699), .B2(n19474), .ZN(
        n19479) );
  AOI22_X1 U21566 ( .A1(n19705), .A2(n19477), .B1(n19703), .B2(n19476), .ZN(
        n19478) );
  OAI211_X1 U21567 ( .C1(n19709), .C2(n19480), .A(n19479), .B(n19478), .ZN(
        P2_U3051) );
  INV_X1 U21568 ( .A(n19497), .ZN(n19488) );
  AOI22_X1 U21569 ( .A1(n19581), .A2(n19488), .B1(n19579), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n19486) );
  AOI22_X1 U21570 ( .A1(n19583), .A2(BUF1_REG_18__SCAN_IN), .B1(n19582), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n19485) );
  INV_X1 U21571 ( .A(n19481), .ZN(n19482) );
  AOI22_X1 U21572 ( .A1(n19483), .A2(n19586), .B1(n19585), .B2(n19482), .ZN(
        n19484) );
  NAND3_X1 U21573 ( .A1(n19486), .A2(n19485), .A3(n19484), .ZN(P2_U2901) );
  AOI22_X1 U21574 ( .A1(n19489), .A2(n19488), .B1(n19585), .B2(n19487), .ZN(
        n19494) );
  OAI211_X1 U21575 ( .C1(n19492), .C2(n19491), .A(n19490), .B(n19586), .ZN(
        n19493) );
  OAI211_X1 U21576 ( .C1(n19496), .C2(n19495), .A(n19494), .B(n19493), .ZN(
        P2_U2917) );
  NOR2_X2 U21577 ( .A1(n19497), .A2(n19591), .ZN(n19537) );
  AOI22_X1 U21578 ( .A1(n19596), .A2(n19537), .B1(n19595), .B2(n19535), .ZN(
        n19499) );
  AOI22_X1 U21579 ( .A1(n19604), .A2(n19536), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19498) );
  OAI211_X1 U21580 ( .C1(n19534), .C2(n19602), .A(n19499), .B(n19498), .ZN(
        P2_U3170) );
  AOI22_X1 U21581 ( .A1(n19500), .A2(n19536), .B1(n19535), .B2(n19603), .ZN(
        n19502) );
  AOI22_X1 U21582 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19606), .B1(
        n19537), .B2(n19605), .ZN(n19501) );
  OAI211_X1 U21583 ( .C1(n19534), .C2(n19544), .A(n19502), .B(n19501), .ZN(
        P2_U3162) );
  AOI22_X1 U21584 ( .A1(n19610), .A2(n19537), .B1(n19609), .B2(n19535), .ZN(
        n19504) );
  AOI22_X1 U21585 ( .A1(n19611), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n19617), .B2(n19536), .ZN(n19503) );
  OAI211_X1 U21586 ( .C1(n19534), .C2(n19614), .A(n19504), .B(n19503), .ZN(
        P2_U3154) );
  AOI22_X1 U21587 ( .A1(n19616), .A2(n19537), .B1(n19535), .B2(n19615), .ZN(
        n19506) );
  AOI22_X1 U21588 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n19617), .B2(n19538), .ZN(n19505) );
  OAI211_X1 U21589 ( .C1(n19531), .C2(n19621), .A(n19506), .B(n19505), .ZN(
        P2_U3146) );
  AOI22_X1 U21590 ( .A1(n19623), .A2(n19537), .B1(n19535), .B2(n19622), .ZN(
        n19508) );
  AOI22_X1 U21591 ( .A1(n19630), .A2(n19536), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n19624), .ZN(n19507) );
  OAI211_X1 U21592 ( .C1(n19534), .C2(n19621), .A(n19508), .B(n19507), .ZN(
        P2_U3138) );
  AOI22_X1 U21593 ( .A1(n19630), .A2(n19538), .B1(n19629), .B2(n19535), .ZN(
        n19510) );
  AOI22_X1 U21594 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19632), .B1(
        n19537), .B2(n19631), .ZN(n19509) );
  OAI211_X1 U21595 ( .C1(n19531), .C2(n19641), .A(n19510), .B(n19509), .ZN(
        P2_U3130) );
  AOI22_X1 U21596 ( .A1(n19553), .A2(n19538), .B1(n19635), .B2(n19535), .ZN(
        n19512) );
  AOI22_X1 U21597 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19638), .B1(
        n19537), .B2(n19637), .ZN(n19511) );
  OAI211_X1 U21598 ( .C1(n19531), .C2(n19649), .A(n19512), .B(n19511), .ZN(
        P2_U3122) );
  AOI22_X1 U21599 ( .A1(n19636), .A2(n19538), .B1(n19513), .B2(n19535), .ZN(
        n19515) );
  AOI22_X1 U21600 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19537), .ZN(n19514) );
  OAI211_X1 U21601 ( .C1(n19531), .C2(n19655), .A(n19515), .B(n19514), .ZN(
        P2_U3114) );
  AOI22_X1 U21602 ( .A1(n19651), .A2(n19537), .B1(n19650), .B2(n19535), .ZN(
        n19517) );
  AOI22_X1 U21603 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19536), .ZN(n19516) );
  OAI211_X1 U21604 ( .C1(n19534), .C2(n19655), .A(n19517), .B(n19516), .ZN(
        P2_U3106) );
  INV_X1 U21605 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n19520) );
  AOI22_X1 U21606 ( .A1(n19657), .A2(n19537), .B1(n19656), .B2(n19535), .ZN(
        n19519) );
  AOI22_X1 U21607 ( .A1(n19658), .A2(n19538), .B1(n19659), .B2(n19536), .ZN(
        n19518) );
  OAI211_X1 U21608 ( .C1(n19663), .C2(n19520), .A(n19519), .B(n19518), .ZN(
        P2_U3098) );
  INV_X1 U21609 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19523) );
  AOI22_X1 U21610 ( .A1(n19671), .A2(n19536), .B1(n19664), .B2(n19535), .ZN(
        n19522) );
  AOI22_X1 U21611 ( .A1(n19537), .A2(n19665), .B1(n19659), .B2(n19538), .ZN(
        n19521) );
  OAI211_X1 U21612 ( .C1(n19524), .C2(n19523), .A(n19522), .B(n19521), .ZN(
        P2_U3090) );
  AOI22_X1 U21613 ( .A1(n19671), .A2(n19538), .B1(n19535), .B2(n19670), .ZN(
        n19526) );
  AOI22_X1 U21614 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19673), .B1(
        n19537), .B2(n19672), .ZN(n19525) );
  OAI211_X1 U21615 ( .C1(n19531), .C2(n19676), .A(n19526), .B(n19525), .ZN(
        P2_U3082) );
  AOI22_X1 U21616 ( .A1(n19686), .A2(n19536), .B1(n19677), .B2(n19535), .ZN(
        n19528) );
  AOI22_X1 U21617 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n19537), .ZN(n19527) );
  OAI211_X1 U21618 ( .C1(n19534), .C2(n19676), .A(n19528), .B(n19527), .ZN(
        P2_U3074) );
  AOI22_X1 U21619 ( .A1(n19685), .A2(n19537), .B1(n19535), .B2(n19684), .ZN(
        n19530) );
  AOI22_X1 U21620 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19538), .ZN(n19529) );
  OAI211_X1 U21621 ( .C1(n19531), .C2(n19696), .A(n19530), .B(n19529), .ZN(
        P2_U3066) );
  AOI22_X1 U21622 ( .A1(n19692), .A2(n19537), .B1(n19535), .B2(n19691), .ZN(
        n19533) );
  AOI22_X1 U21623 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19536), .ZN(n19532) );
  OAI211_X1 U21624 ( .C1(n19534), .C2(n19696), .A(n19533), .B(n19532), .ZN(
        P2_U3058) );
  INV_X1 U21625 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19541) );
  AOI22_X1 U21626 ( .A1(n19705), .A2(n19536), .B1(n19699), .B2(n19535), .ZN(
        n19540) );
  AOI22_X1 U21627 ( .A1(n19701), .A2(n19538), .B1(n19703), .B2(n19537), .ZN(
        n19539) );
  OAI211_X1 U21628 ( .C1(n19709), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3050) );
  AOI22_X1 U21629 ( .A1(n19596), .A2(n19574), .B1(n19573), .B2(n19595), .ZN(
        n19543) );
  AOI22_X1 U21630 ( .A1(n19705), .A2(n19569), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19542) );
  OAI211_X1 U21631 ( .C1(n19572), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        P2_U3169) );
  AOI22_X1 U21632 ( .A1(n19604), .A2(n19569), .B1(n19573), .B2(n19603), .ZN(
        n19546) );
  AOI22_X1 U21633 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19606), .B1(
        n19574), .B2(n19605), .ZN(n19545) );
  OAI211_X1 U21634 ( .C1(n19572), .C2(n19614), .A(n19546), .B(n19545), .ZN(
        P2_U3161) );
  AOI22_X1 U21635 ( .A1(n19616), .A2(n19574), .B1(n19573), .B2(n19615), .ZN(
        n19548) );
  AOI22_X1 U21636 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n19617), .B2(n19569), .ZN(n19547) );
  OAI211_X1 U21637 ( .C1(n19572), .C2(n19621), .A(n19548), .B(n19547), .ZN(
        P2_U3145) );
  AOI22_X1 U21638 ( .A1(n19623), .A2(n19574), .B1(n19573), .B2(n19622), .ZN(
        n19550) );
  AOI22_X1 U21639 ( .A1(n19630), .A2(n19575), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n19624), .ZN(n19549) );
  OAI211_X1 U21640 ( .C1(n19578), .C2(n19621), .A(n19550), .B(n19549), .ZN(
        P2_U3137) );
  AOI22_X1 U21641 ( .A1(n19553), .A2(n19575), .B1(n19573), .B2(n19629), .ZN(
        n19552) );
  AOI22_X1 U21642 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19632), .B1(
        n19574), .B2(n19631), .ZN(n19551) );
  OAI211_X1 U21643 ( .C1(n19578), .C2(n19628), .A(n19552), .B(n19551), .ZN(
        P2_U3129) );
  AOI22_X1 U21644 ( .A1(n19553), .A2(n19569), .B1(n19573), .B2(n19635), .ZN(
        n19555) );
  AOI22_X1 U21645 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19638), .B1(
        n19574), .B2(n19637), .ZN(n19554) );
  OAI211_X1 U21646 ( .C1(n19572), .C2(n19649), .A(n19555), .B(n19554), .ZN(
        P2_U3121) );
  OAI22_X1 U21647 ( .A1(n19655), .A2(n19572), .B1(n19556), .B2(n19643), .ZN(
        n19557) );
  INV_X1 U21648 ( .A(n19557), .ZN(n19559) );
  AOI22_X1 U21649 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19574), .ZN(n19558) );
  OAI211_X1 U21650 ( .C1(n19578), .C2(n19649), .A(n19559), .B(n19558), .ZN(
        P2_U3113) );
  AOI22_X1 U21651 ( .A1(n19651), .A2(n19574), .B1(n19650), .B2(n19573), .ZN(
        n19561) );
  AOI22_X1 U21652 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19575), .ZN(n19560) );
  OAI211_X1 U21653 ( .C1(n19578), .C2(n19655), .A(n19561), .B(n19560), .ZN(
        P2_U3105) );
  AOI22_X1 U21654 ( .A1(n19659), .A2(n19569), .B1(n19573), .B2(n19664), .ZN(
        n19563) );
  AOI22_X1 U21655 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19666), .B1(
        n19574), .B2(n19665), .ZN(n19562) );
  OAI211_X1 U21656 ( .C1(n19572), .C2(n19564), .A(n19563), .B(n19562), .ZN(
        P2_U3089) );
  AOI22_X1 U21657 ( .A1(n19671), .A2(n19569), .B1(n19573), .B2(n19670), .ZN(
        n19566) );
  AOI22_X1 U21658 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19673), .B1(
        n19574), .B2(n19672), .ZN(n19565) );
  OAI211_X1 U21659 ( .C1(n19572), .C2(n19676), .A(n19566), .B(n19565), .ZN(
        P2_U3081) );
  AOI22_X1 U21660 ( .A1(n19678), .A2(n19569), .B1(n19573), .B2(n19677), .ZN(
        n19568) );
  AOI22_X1 U21661 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n19574), .ZN(n19567) );
  OAI211_X1 U21662 ( .C1(n19572), .C2(n19683), .A(n19568), .B(n19567), .ZN(
        P2_U3073) );
  AOI22_X1 U21663 ( .A1(n19685), .A2(n19574), .B1(n19573), .B2(n19684), .ZN(
        n19571) );
  AOI22_X1 U21664 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19569), .ZN(n19570) );
  OAI211_X1 U21665 ( .C1(n19572), .C2(n19696), .A(n19571), .B(n19570), .ZN(
        P2_U3065) );
  AOI22_X1 U21666 ( .A1(n19692), .A2(n19574), .B1(n19573), .B2(n19691), .ZN(
        n19577) );
  AOI22_X1 U21667 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19575), .ZN(n19576) );
  OAI211_X1 U21668 ( .C1(n19578), .C2(n19696), .A(n19577), .B(n19576), .ZN(
        P2_U3057) );
  AOI22_X1 U21669 ( .A1(n19581), .A2(n19580), .B1(n19579), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19590) );
  AOI22_X1 U21670 ( .A1(n19583), .A2(BUF1_REG_16__SCAN_IN), .B1(n19582), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19589) );
  AOI22_X1 U21671 ( .A1(n19587), .A2(n19586), .B1(n19585), .B2(n19584), .ZN(
        n19588) );
  NAND3_X1 U21672 ( .A1(n19590), .A2(n19589), .A3(n19588), .ZN(P2_U2903) );
  NOR2_X2 U21673 ( .A1(n19592), .A2(n19591), .ZN(n19702) );
  NAND2_X1 U21674 ( .A1(n19594), .A2(n19593), .ZN(n19642) );
  AOI22_X1 U21675 ( .A1(n19596), .A2(n19702), .B1(n19595), .B2(n19698), .ZN(
        n19601) );
  AOI22_X1 U21676 ( .A1(n19604), .A2(n19704), .B1(n19599), .B2(
        P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19600) );
  OAI211_X1 U21677 ( .C1(n19697), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        P2_U3168) );
  AOI22_X1 U21678 ( .A1(n19604), .A2(n19700), .B1(n19698), .B2(n19603), .ZN(
        n19608) );
  AOI22_X1 U21679 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19606), .B1(
        n19702), .B2(n19605), .ZN(n19607) );
  OAI211_X1 U21680 ( .C1(n19690), .C2(n19614), .A(n19608), .B(n19607), .ZN(
        P2_U3160) );
  AOI22_X1 U21681 ( .A1(n19610), .A2(n19702), .B1(n19609), .B2(n19698), .ZN(
        n19613) );
  AOI22_X1 U21682 ( .A1(n19611), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n19617), .B2(n19704), .ZN(n19612) );
  OAI211_X1 U21683 ( .C1(n19697), .C2(n19614), .A(n19613), .B(n19612), .ZN(
        P2_U3152) );
  AOI22_X1 U21684 ( .A1(n19616), .A2(n19702), .B1(n19698), .B2(n19615), .ZN(
        n19620) );
  AOI22_X1 U21685 ( .A1(n19618), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n19617), .B2(n19700), .ZN(n19619) );
  OAI211_X1 U21686 ( .C1(n19690), .C2(n19621), .A(n19620), .B(n19619), .ZN(
        P2_U3144) );
  AOI22_X1 U21687 ( .A1(n19623), .A2(n19702), .B1(n19698), .B2(n19622), .ZN(
        n19627) );
  AOI22_X1 U21688 ( .A1(n19625), .A2(n19700), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n19624), .ZN(n19626) );
  OAI211_X1 U21689 ( .C1(n19690), .C2(n19628), .A(n19627), .B(n19626), .ZN(
        P2_U3136) );
  AOI22_X1 U21690 ( .A1(n19630), .A2(n19700), .B1(n19698), .B2(n19629), .ZN(
        n19634) );
  AOI22_X1 U21691 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19632), .B1(
        n19702), .B2(n19631), .ZN(n19633) );
  OAI211_X1 U21692 ( .C1(n19690), .C2(n19641), .A(n19634), .B(n19633), .ZN(
        P2_U3128) );
  AOI22_X1 U21693 ( .A1(n19636), .A2(n19704), .B1(n19698), .B2(n19635), .ZN(
        n19640) );
  AOI22_X1 U21694 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19638), .B1(
        n19702), .B2(n19637), .ZN(n19639) );
  OAI211_X1 U21695 ( .C1(n19697), .C2(n19641), .A(n19640), .B(n19639), .ZN(
        P2_U3120) );
  OAI22_X1 U21696 ( .A1(n19655), .A2(n19690), .B1(n19643), .B2(n19642), .ZN(
        n19644) );
  INV_X1 U21697 ( .A(n19644), .ZN(n19648) );
  AOI22_X1 U21698 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19646), .B1(
        n19645), .B2(n19702), .ZN(n19647) );
  OAI211_X1 U21699 ( .C1(n19697), .C2(n19649), .A(n19648), .B(n19647), .ZN(
        P2_U3112) );
  AOI22_X1 U21700 ( .A1(n19651), .A2(n19702), .B1(n19650), .B2(n19698), .ZN(
        n19654) );
  AOI22_X1 U21701 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19652), .B1(
        n19658), .B2(n19704), .ZN(n19653) );
  OAI211_X1 U21702 ( .C1(n19697), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3104) );
  INV_X1 U21703 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U21704 ( .A1(n19657), .A2(n19702), .B1(n19656), .B2(n19698), .ZN(
        n19661) );
  AOI22_X1 U21705 ( .A1(n19659), .A2(n19704), .B1(n19658), .B2(n19700), .ZN(
        n19660) );
  OAI211_X1 U21706 ( .C1(n19663), .C2(n19662), .A(n19661), .B(n19660), .ZN(
        P2_U3096) );
  AOI22_X1 U21707 ( .A1(n19671), .A2(n19704), .B1(n19664), .B2(n19698), .ZN(
        n19668) );
  AOI22_X1 U21708 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19666), .B1(
        n19702), .B2(n19665), .ZN(n19667) );
  OAI211_X1 U21709 ( .C1(n19697), .C2(n19669), .A(n19668), .B(n19667), .ZN(
        P2_U3088) );
  AOI22_X1 U21710 ( .A1(n19671), .A2(n19700), .B1(n19698), .B2(n19670), .ZN(
        n19675) );
  AOI22_X1 U21711 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19673), .B1(
        n19702), .B2(n19672), .ZN(n19674) );
  OAI211_X1 U21712 ( .C1(n19690), .C2(n19676), .A(n19675), .B(n19674), .ZN(
        P2_U3080) );
  AOI22_X1 U21713 ( .A1(n19678), .A2(n19700), .B1(n19698), .B2(n19677), .ZN(
        n19682) );
  AOI22_X1 U21714 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19680), .B1(
        n19679), .B2(n19702), .ZN(n19681) );
  OAI211_X1 U21715 ( .C1(n19690), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        P2_U3072) );
  AOI22_X1 U21716 ( .A1(n19685), .A2(n19702), .B1(n19698), .B2(n19684), .ZN(
        n19689) );
  AOI22_X1 U21717 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19700), .ZN(n19688) );
  OAI211_X1 U21718 ( .C1(n19690), .C2(n19696), .A(n19689), .B(n19688), .ZN(
        P2_U3064) );
  AOI22_X1 U21719 ( .A1(n19692), .A2(n19702), .B1(n19698), .B2(n19691), .ZN(
        n19695) );
  AOI22_X1 U21720 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19693), .B1(
        n19701), .B2(n19704), .ZN(n19694) );
  OAI211_X1 U21721 ( .C1(n19697), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        P2_U3056) );
  AOI22_X1 U21722 ( .A1(n19701), .A2(n19700), .B1(n19699), .B2(n19698), .ZN(
        n19707) );
  AOI22_X1 U21723 ( .A1(n19705), .A2(n19704), .B1(n19703), .B2(n19702), .ZN(
        n19706) );
  OAI211_X1 U21724 ( .C1(n19709), .C2(n19708), .A(n19707), .B(n19706), .ZN(
        P2_U3048) );
  INV_X1 U21725 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n19998) );
  INV_X1 U21726 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19710) );
  AOI222_X1 U21727 ( .A1(n19998), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20000), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19710), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19711) );
  OAI22_X1 U21728 ( .A1(n19763), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n19766), .ZN(n19712) );
  INV_X1 U21729 ( .A(n19712), .ZN(U376) );
  INV_X2 U21730 ( .A(n19763), .ZN(n19766) );
  INV_X1 U21731 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19714) );
  AOI22_X1 U21732 ( .A1(n19766), .A2(n19714), .B1(n19713), .B2(n19763), .ZN(
        U365) );
  INV_X1 U21733 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19716) );
  AOI22_X1 U21734 ( .A1(n19766), .A2(n19716), .B1(n19715), .B2(n19763), .ZN(
        U354) );
  INV_X1 U21735 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19718) );
  AOI22_X1 U21736 ( .A1(n19766), .A2(n19718), .B1(n19717), .B2(n19763), .ZN(
        U353) );
  INV_X1 U21737 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U21738 ( .A1(n19766), .A2(n19720), .B1(n19719), .B2(n19763), .ZN(
        U352) );
  INV_X1 U21739 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19722) );
  AOI22_X1 U21740 ( .A1(n19766), .A2(n19722), .B1(n19721), .B2(n19763), .ZN(
        U351) );
  OAI22_X1 U21741 ( .A1(n19763), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n19766), .ZN(n19723) );
  INV_X1 U21742 ( .A(n19723), .ZN(U350) );
  OAI22_X1 U21743 ( .A1(n19763), .A2(P3_ADDRESS_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n19766), .ZN(n19724) );
  INV_X1 U21744 ( .A(n19724), .ZN(U349) );
  AOI22_X1 U21745 ( .A1(n19766), .A2(n19726), .B1(n19725), .B2(n19763), .ZN(
        U348) );
  AOI22_X1 U21746 ( .A1(n19766), .A2(n19728), .B1(n19727), .B2(n19763), .ZN(
        U347) );
  AOI22_X1 U21747 ( .A1(n19766), .A2(n19730), .B1(n19729), .B2(n19763), .ZN(
        U375) );
  OAI22_X1 U21748 ( .A1(n19763), .A2(P3_ADDRESS_REG_11__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n19766), .ZN(n19731) );
  INV_X1 U21749 ( .A(n19731), .ZN(U374) );
  OAI22_X1 U21750 ( .A1(n19763), .A2(P3_ADDRESS_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n19766), .ZN(n19732) );
  INV_X1 U21751 ( .A(n19732), .ZN(U373) );
  AOI22_X1 U21752 ( .A1(n19766), .A2(n19734), .B1(n19733), .B2(n19763), .ZN(
        U372) );
  AOI22_X1 U21753 ( .A1(n19766), .A2(n19736), .B1(n19735), .B2(n19763), .ZN(
        U371) );
  AOI22_X1 U21754 ( .A1(n19766), .A2(n19738), .B1(n19737), .B2(n19763), .ZN(
        U370) );
  AOI22_X1 U21755 ( .A1(n19766), .A2(n19740), .B1(n19739), .B2(n19763), .ZN(
        U369) );
  AOI22_X1 U21756 ( .A1(n19766), .A2(n19742), .B1(n19741), .B2(n19763), .ZN(
        U368) );
  AOI22_X1 U21757 ( .A1(n19766), .A2(n19744), .B1(n19743), .B2(n19763), .ZN(
        U367) );
  AOI22_X1 U21758 ( .A1(n19766), .A2(n19746), .B1(n19745), .B2(n19763), .ZN(
        U366) );
  AOI22_X1 U21759 ( .A1(n19766), .A2(n19748), .B1(n19747), .B2(n19763), .ZN(
        U364) );
  AOI22_X1 U21760 ( .A1(n19766), .A2(n19750), .B1(n19749), .B2(n19763), .ZN(
        U363) );
  AOI22_X1 U21761 ( .A1(n19766), .A2(n19752), .B1(n19751), .B2(n19763), .ZN(
        U362) );
  AOI22_X1 U21762 ( .A1(n19766), .A2(n19754), .B1(n19753), .B2(n19763), .ZN(
        U361) );
  OAI22_X1 U21763 ( .A1(n19763), .A2(P3_ADDRESS_REG_24__SCAN_IN), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(n19766), .ZN(n19755) );
  INV_X1 U21764 ( .A(n19755), .ZN(U360) );
  OAI22_X1 U21765 ( .A1(n19763), .A2(P3_ADDRESS_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(n19766), .ZN(n19756) );
  INV_X1 U21766 ( .A(n19756), .ZN(U359) );
  INV_X1 U21767 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U21768 ( .A1(n19766), .A2(n19758), .B1(n19757), .B2(n19763), .ZN(
        U358) );
  INV_X1 U21769 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U21770 ( .A1(n19766), .A2(n19760), .B1(n19759), .B2(n19763), .ZN(
        U357) );
  AOI22_X1 U21771 ( .A1(n19766), .A2(n19762), .B1(n19761), .B2(n19763), .ZN(
        U356) );
  AOI22_X1 U21772 ( .A1(n19766), .A2(n19765), .B1(n19764), .B2(n19763), .ZN(
        U355) );
  AOI22_X1 U21773 ( .A1(n21230), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19768) );
  OAI21_X1 U21774 ( .B1(n11848), .B2(n19794), .A(n19768), .ZN(P1_U2936) );
  AOI22_X1 U21775 ( .A1(n19780), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19769) );
  OAI21_X1 U21776 ( .B1(n11838), .B2(n19794), .A(n19769), .ZN(P1_U2935) );
  AOI22_X1 U21777 ( .A1(n19780), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19770) );
  OAI21_X1 U21778 ( .B1(n19771), .B2(n19794), .A(n19770), .ZN(P1_U2934) );
  AOI22_X1 U21779 ( .A1(n19780), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19772) );
  OAI21_X1 U21780 ( .B1(n11864), .B2(n19794), .A(n19772), .ZN(P1_U2933) );
  AOI22_X1 U21781 ( .A1(n19780), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19773) );
  OAI21_X1 U21782 ( .B1(n19774), .B2(n19794), .A(n19773), .ZN(P1_U2932) );
  AOI22_X1 U21783 ( .A1(n19780), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19775) );
  OAI21_X1 U21784 ( .B1(n19776), .B2(n19794), .A(n19775), .ZN(P1_U2931) );
  AOI22_X1 U21785 ( .A1(n19780), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19777) );
  OAI21_X1 U21786 ( .B1(n19778), .B2(n19794), .A(n19777), .ZN(P1_U2930) );
  AOI22_X1 U21787 ( .A1(n21230), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19779) );
  OAI21_X1 U21788 ( .B1(n11828), .B2(n19794), .A(n19779), .ZN(P1_U2929) );
  AOI22_X1 U21789 ( .A1(n19780), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19781) );
  OAI21_X1 U21790 ( .B1(n14502), .B2(n19794), .A(n19781), .ZN(P1_U2928) );
  AOI22_X1 U21791 ( .A1(n21230), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19782) );
  OAI21_X1 U21792 ( .B1(n19783), .B2(n19794), .A(n19782), .ZN(P1_U2927) );
  AOI22_X1 U21793 ( .A1(n21230), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19785) );
  OAI21_X1 U21794 ( .B1(n19786), .B2(n19794), .A(n19785), .ZN(P1_U2926) );
  AOI22_X1 U21795 ( .A1(n21230), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19787) );
  OAI21_X1 U21796 ( .B1(n19788), .B2(n19794), .A(n19787), .ZN(P1_U2925) );
  AOI22_X1 U21797 ( .A1(n21230), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19789) );
  OAI21_X1 U21798 ( .B1(n15026), .B2(n19794), .A(n19789), .ZN(P1_U2924) );
  AOI22_X1 U21799 ( .A1(n21230), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19790) );
  OAI21_X1 U21800 ( .B1(n15001), .B2(n19794), .A(n19790), .ZN(P1_U2923) );
  AOI22_X1 U21801 ( .A1(n21230), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19791) );
  OAI21_X1 U21802 ( .B1(n19792), .B2(n19794), .A(n19791), .ZN(P1_U2922) );
  AOI22_X1 U21803 ( .A1(n21230), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19784), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19793) );
  OAI21_X1 U21804 ( .B1(n19795), .B2(n19794), .A(n19793), .ZN(P1_U2921) );
  INV_X2 U21805 ( .A(n22246), .ZN(n19831) );
  NOR2_X2 U21806 ( .A1(n21585), .A2(n19831), .ZN(n19836) );
  INV_X1 U21807 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19798) );
  NOR2_X2 U21808 ( .A1(n19831), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n19830) );
  OAI222_X1 U21809 ( .A1(n19834), .A2(n13941), .B1(n19796), .B2(n22246), .C1(
        n19798), .C2(n19838), .ZN(P1_U3197) );
  AOI22_X1 U21810 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n19831), .ZN(n19797) );
  OAI21_X1 U21811 ( .B1(n19798), .B2(n19834), .A(n19797), .ZN(P1_U3198) );
  AOI22_X1 U21812 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n19831), .ZN(n19799) );
  OAI21_X1 U21813 ( .B1(n19801), .B2(n19838), .A(n19799), .ZN(P1_U3199) );
  AOI22_X1 U21814 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n19831), .ZN(n19800) );
  OAI21_X1 U21815 ( .B1(n19801), .B2(n19834), .A(n19800), .ZN(P1_U3200) );
  AOI22_X1 U21816 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n19831), .ZN(n19802) );
  OAI21_X1 U21817 ( .B1(n21426), .B2(n19838), .A(n19802), .ZN(P1_U3201) );
  AOI22_X1 U21818 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n19831), .ZN(n19803) );
  OAI21_X1 U21819 ( .B1(n21426), .B2(n19834), .A(n19803), .ZN(P1_U3202) );
  AOI22_X1 U21820 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n19831), .ZN(n19804) );
  OAI21_X1 U21821 ( .B1(n19806), .B2(n19838), .A(n19804), .ZN(P1_U3203) );
  AOI22_X1 U21822 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n19831), .ZN(n19805) );
  OAI21_X1 U21823 ( .B1(n19806), .B2(n19834), .A(n19805), .ZN(P1_U3204) );
  AOI22_X1 U21824 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n19831), .ZN(n19807) );
  OAI21_X1 U21825 ( .B1(n21297), .B2(n19838), .A(n19807), .ZN(P1_U3205) );
  AOI22_X1 U21826 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n19831), .ZN(n19808) );
  OAI21_X1 U21827 ( .B1(n21297), .B2(n19834), .A(n19808), .ZN(P1_U3206) );
  AOI22_X1 U21828 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n19831), .ZN(n19809) );
  OAI21_X1 U21829 ( .B1(n21305), .B2(n19838), .A(n19809), .ZN(P1_U3207) );
  AOI22_X1 U21830 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n19831), .ZN(n19810) );
  OAI21_X1 U21831 ( .B1(n21305), .B2(n19834), .A(n19810), .ZN(P1_U3208) );
  INV_X1 U21832 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21469) );
  AOI22_X1 U21833 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n19831), .ZN(n19811) );
  OAI21_X1 U21834 ( .B1(n21469), .B2(n19838), .A(n19811), .ZN(P1_U3209) );
  AOI22_X1 U21835 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n19831), .ZN(n19812) );
  OAI21_X1 U21836 ( .B1(n21469), .B2(n19834), .A(n19812), .ZN(P1_U3210) );
  INV_X1 U21837 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U21838 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n19831), .ZN(n19813) );
  OAI21_X1 U21839 ( .B1(n19814), .B2(n19838), .A(n19813), .ZN(P1_U3211) );
  AOI222_X1 U21840 ( .A1(n19830), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n19836), .ZN(n19815) );
  INV_X1 U21841 ( .A(n19815), .ZN(P1_U3212) );
  AOI22_X1 U21842 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n19831), .ZN(n19816) );
  OAI21_X1 U21843 ( .B1(n19817), .B2(n19834), .A(n19816), .ZN(P1_U3213) );
  INV_X1 U21844 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U21845 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n19831), .ZN(n19818) );
  OAI21_X1 U21846 ( .B1(n19819), .B2(n19834), .A(n19818), .ZN(P1_U3214) );
  AOI22_X1 U21847 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n19831), .ZN(n19820) );
  OAI21_X1 U21848 ( .B1(n19821), .B2(n19838), .A(n19820), .ZN(P1_U3215) );
  AOI222_X1 U21849 ( .A1(n19836), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n19830), .ZN(n19822) );
  INV_X1 U21850 ( .A(n19822), .ZN(P1_U3216) );
  AOI222_X1 U21851 ( .A1(n19830), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n19836), .ZN(n19823) );
  INV_X1 U21852 ( .A(n19823), .ZN(P1_U3217) );
  AOI222_X1 U21853 ( .A1(n19830), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n19836), .ZN(n19824) );
  INV_X1 U21854 ( .A(n19824), .ZN(P1_U3218) );
  AOI222_X1 U21855 ( .A1(n19836), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n19830), .ZN(n19825) );
  INV_X1 U21856 ( .A(n19825), .ZN(P1_U3219) );
  AOI222_X1 U21857 ( .A1(n19830), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n19836), .ZN(n19826) );
  INV_X1 U21858 ( .A(n19826), .ZN(P1_U3220) );
  AOI222_X1 U21859 ( .A1(n19836), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n19830), .ZN(n19827) );
  INV_X1 U21860 ( .A(n19827), .ZN(P1_U3221) );
  AOI222_X1 U21861 ( .A1(n19830), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n19836), .ZN(n19828) );
  INV_X1 U21862 ( .A(n19828), .ZN(P1_U3222) );
  AOI222_X1 U21863 ( .A1(n19836), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n19830), .ZN(n19829) );
  INV_X1 U21864 ( .A(n19829), .ZN(P1_U3223) );
  AOI222_X1 U21865 ( .A1(n19836), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n19831), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n19830), .ZN(n19832) );
  INV_X1 U21866 ( .A(n19832), .ZN(P1_U3224) );
  AOI22_X1 U21867 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n19830), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n19831), .ZN(n19833) );
  OAI21_X1 U21868 ( .B1(n19835), .B2(n19834), .A(n19833), .ZN(P1_U3225) );
  AOI22_X1 U21869 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n19836), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n19831), .ZN(n19837) );
  OAI21_X1 U21870 ( .B1(n19839), .B2(n19838), .A(n19837), .ZN(P1_U3226) );
  OAI22_X1 U21871 ( .A1(n19831), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22246), .ZN(n19840) );
  INV_X1 U21872 ( .A(n19840), .ZN(P1_U3458) );
  AOI221_X1 U21873 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19851) );
  NOR4_X1 U21874 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19844) );
  NOR4_X1 U21875 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19843) );
  NOR4_X1 U21876 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19842) );
  NOR4_X1 U21877 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19841) );
  NAND4_X1 U21878 ( .A1(n19844), .A2(n19843), .A3(n19842), .A4(n19841), .ZN(
        n19850) );
  NOR4_X1 U21879 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19848) );
  AOI211_X1 U21880 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19847) );
  NOR4_X1 U21881 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19846) );
  NOR4_X1 U21882 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19845) );
  NAND4_X1 U21883 ( .A1(n19848), .A2(n19847), .A3(n19846), .A4(n19845), .ZN(
        n19849) );
  NOR2_X1 U21884 ( .A1(n19850), .A2(n19849), .ZN(n19863) );
  MUX2_X1 U21885 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n19851), .S(n19863), 
        .Z(P1_U2808) );
  OAI22_X1 U21886 ( .A1(n19831), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22246), .ZN(n19852) );
  INV_X1 U21887 ( .A(n19852), .ZN(P1_U3459) );
  AOI21_X1 U21888 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19853) );
  OAI221_X1 U21889 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19853), .C1(n13941), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n19863), .ZN(n19854) );
  OAI21_X1 U21890 ( .B1(n19863), .B2(n19855), .A(n19854), .ZN(P1_U3481) );
  OAI22_X1 U21891 ( .A1(n19831), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22246), .ZN(n19856) );
  INV_X1 U21892 ( .A(n19856), .ZN(P1_U3460) );
  NOR3_X1 U21893 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19857) );
  OAI21_X1 U21894 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19857), .A(n19863), .ZN(
        n19858) );
  OAI21_X1 U21895 ( .B1(n19863), .B2(n19859), .A(n19858), .ZN(P1_U2807) );
  OAI22_X1 U21896 ( .A1(n19831), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22246), .ZN(n19860) );
  INV_X1 U21897 ( .A(n19860), .ZN(P1_U3461) );
  OAI21_X1 U21898 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n19863), .ZN(n19861) );
  OAI21_X1 U21899 ( .B1(n19863), .B2(n19862), .A(n19861), .ZN(P1_U3482) );
  AOI22_X1 U21900 ( .A1(n19867), .A2(n19866), .B1(n19865), .B2(n19864), .ZN(
        n19868) );
  OAI21_X1 U21901 ( .B1(n19870), .B2(n19869), .A(n19868), .ZN(P1_U2869) );
  XNOR2_X1 U21902 ( .A(n19872), .B(n19871), .ZN(n21264) );
  OAI22_X1 U21903 ( .A1(n19874), .A2(n19915), .B1(n19873), .B2(n19952), .ZN(
        n19875) );
  AOI21_X1 U21904 ( .B1(n21264), .B2(n19949), .A(n19875), .ZN(n19876) );
  NAND2_X1 U21905 ( .A1(n21390), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n21270) );
  OAI211_X1 U21906 ( .C1(n19901), .C2(n19877), .A(n19876), .B(n21270), .ZN(
        P1_U2994) );
  INV_X1 U21907 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19882) );
  XOR2_X1 U21908 ( .A(n19879), .B(n19878), .Z(n21275) );
  INV_X1 U21909 ( .A(n21435), .ZN(n19880) );
  AOI222_X1 U21910 ( .A1(n21275), .A2(n19949), .B1(n19948), .B2(n21440), .C1(
        n19880), .C2(n19927), .ZN(n19881) );
  NAND2_X1 U21911 ( .A1(n21390), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n21274) );
  OAI211_X1 U21912 ( .C1(n19901), .C2(n19882), .A(n19881), .B(n21274), .ZN(
        P1_U2992) );
  MUX2_X1 U21913 ( .A(n15950), .B(n19884), .S(n19883), .Z(n19886) );
  INV_X1 U21914 ( .A(n19886), .ZN(n19888) );
  NOR2_X1 U21915 ( .A1(n19886), .A2(n19885), .ZN(n19896) );
  INV_X1 U21916 ( .A(n19896), .ZN(n19887) );
  OAI21_X1 U21917 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19888), .A(
        n19887), .ZN(n21304) );
  AOI22_X1 U21918 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n19893) );
  INV_X1 U21919 ( .A(n19889), .ZN(n19890) );
  AOI22_X1 U21920 ( .A1(n19891), .A2(n19948), .B1(n19890), .B2(n19927), .ZN(
        n19892) );
  OAI211_X1 U21921 ( .C1(n21546), .C2(n21304), .A(n19893), .B(n19892), .ZN(
        P1_U2989) );
  INV_X1 U21922 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19900) );
  NOR2_X1 U21923 ( .A1(n19896), .A2(n15950), .ZN(n19895) );
  MUX2_X1 U21924 ( .A(n19896), .B(n19895), .S(n19894), .Z(n19897) );
  XOR2_X1 U21925 ( .A(n21309), .B(n19897), .Z(n21318) );
  OAI22_X1 U21926 ( .A1(n21318), .A2(n21546), .B1(n19952), .B2(n21446), .ZN(
        n19898) );
  AOI21_X1 U21927 ( .B1(n19948), .B2(n21448), .A(n19898), .ZN(n19899) );
  NAND2_X1 U21928 ( .A1(n21390), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n21322) );
  OAI211_X1 U21929 ( .C1(n19901), .C2(n19900), .A(n19899), .B(n21322), .ZN(
        P1_U2988) );
  AOI21_X1 U21930 ( .B1(n19904), .B2(n19903), .A(n19902), .ZN(n21317) );
  AOI22_X1 U21931 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U21932 ( .A1(n19927), .A2(n21457), .B1(n19948), .B2(n21456), .ZN(
        n19905) );
  OAI211_X1 U21933 ( .C1(n21317), .C2(n21546), .A(n19906), .B(n19905), .ZN(
        P1_U2987) );
  INV_X1 U21934 ( .A(n19907), .ZN(n19909) );
  NAND2_X1 U21935 ( .A1(n19909), .A2(n19908), .ZN(n19911) );
  OAI21_X1 U21936 ( .B1(n19912), .B2(n19911), .A(n19910), .ZN(n19914) );
  XNOR2_X1 U21937 ( .A(n19945), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n19913) );
  XNOR2_X1 U21938 ( .A(n19914), .B(n19913), .ZN(n21256) );
  AOI22_X1 U21939 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n19917) );
  INV_X1 U21940 ( .A(n19948), .ZN(n19915) );
  AOI22_X1 U21941 ( .A1(n21468), .A2(n21664), .B1(n19927), .B2(n21467), .ZN(
        n19916) );
  OAI211_X1 U21942 ( .C1(n21256), .C2(n21546), .A(n19917), .B(n19916), .ZN(
        P1_U2985) );
  INV_X1 U21943 ( .A(n19918), .ZN(n19920) );
  AOI21_X1 U21944 ( .B1(n15950), .B2(n19920), .A(n19919), .ZN(n19923) );
  INV_X1 U21945 ( .A(n19923), .ZN(n19926) );
  OAI21_X1 U21946 ( .B1(n13569), .B2(n19945), .A(n19930), .ZN(n19925) );
  INV_X1 U21947 ( .A(n19921), .ZN(n19922) );
  NAND3_X1 U21948 ( .A1(n19923), .A2(n19922), .A3(n19930), .ZN(n19931) );
  INV_X1 U21949 ( .A(n19931), .ZN(n19924) );
  AOI21_X1 U21950 ( .B1(n19926), .B2(n19925), .A(n19924), .ZN(n21336) );
  AOI22_X1 U21951 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U21952 ( .A1(n21480), .A2(n21664), .B1(n19927), .B2(n21478), .ZN(
        n19928) );
  OAI211_X1 U21953 ( .C1(n21336), .C2(n21546), .A(n19929), .B(n19928), .ZN(
        P1_U2984) );
  AOI22_X1 U21954 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n19935) );
  NAND2_X1 U21955 ( .A1(n19931), .A2(n19930), .ZN(n19933) );
  XNOR2_X1 U21956 ( .A(n19933), .B(n19932), .ZN(n21354) );
  AOI22_X1 U21957 ( .A1(n21354), .A2(n19949), .B1(n19948), .B2(n21638), .ZN(
        n19934) );
  OAI211_X1 U21958 ( .C1(n19952), .C2(n21487), .A(n19935), .B(n19934), .ZN(
        P1_U2983) );
  AOI22_X1 U21959 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n19942) );
  OAI21_X1 U21960 ( .B1(n19937), .B2(n19940), .A(n19936), .ZN(n19938) );
  OAI21_X1 U21961 ( .B1(n19940), .B2(n19939), .A(n19938), .ZN(n21369) );
  AOI22_X1 U21962 ( .A1(n21369), .A2(n19949), .B1(n19948), .B2(n21646), .ZN(
        n19941) );
  OAI211_X1 U21963 ( .C1(n19952), .C2(n21507), .A(n19942), .B(n19941), .ZN(
        P1_U2979) );
  AOI22_X1 U21964 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19943), .B1(
        n21390), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n19951) );
  OAI21_X1 U21965 ( .B1(n19946), .B2(n19945), .A(n19944), .ZN(n19947) );
  XNOR2_X1 U21966 ( .A(n19947), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21381) );
  AOI22_X1 U21967 ( .A1(n21381), .A2(n19949), .B1(n19948), .B2(n21654), .ZN(
        n19950) );
  OAI211_X1 U21968 ( .C1(n19952), .C2(n21520), .A(n19951), .B(n19950), .ZN(
        P1_U2977) );
  OAI21_X1 U21969 ( .B1(n19953), .B2(n21561), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19954) );
  OAI21_X1 U21970 ( .B1(n19955), .B2(n11213), .A(n19954), .ZN(P1_U2803) );
  INV_X1 U21971 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21591) );
  OAI21_X1 U21972 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21585), .A(n21591), 
        .ZN(n19956) );
  AOI22_X1 U21973 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22246), .B1(n19957), 
        .B2(n19956), .ZN(P1_U2804) );
  AOI22_X1 U21974 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10979), .ZN(n19959) );
  OAI21_X1 U21975 ( .B1(n13914), .B2(n19999), .A(n19959), .ZN(U247) );
  AOI22_X1 U21976 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10979), .ZN(n19960) );
  OAI21_X1 U21977 ( .B1(n13892), .B2(n19999), .A(n19960), .ZN(U246) );
  AOI22_X1 U21978 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10979), .ZN(n19961) );
  OAI21_X1 U21979 ( .B1(n13862), .B2(n19999), .A(n19961), .ZN(U245) );
  AOI22_X1 U21980 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10979), .ZN(n19962) );
  OAI21_X1 U21981 ( .B1(n13899), .B2(n19999), .A(n19962), .ZN(U244) );
  AOI22_X1 U21982 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10979), .ZN(n19963) );
  OAI21_X1 U21983 ( .B1(n19964), .B2(n19999), .A(n19963), .ZN(U243) );
  AOI22_X1 U21984 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10979), .ZN(n19965) );
  OAI21_X1 U21985 ( .B1(n13675), .B2(n19999), .A(n19965), .ZN(U242) );
  AOI22_X1 U21986 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10979), .ZN(n19966) );
  OAI21_X1 U21987 ( .B1(n19967), .B2(n19999), .A(n19966), .ZN(U241) );
  AOI22_X1 U21988 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10979), .ZN(n19968) );
  OAI21_X1 U21989 ( .B1(n13687), .B2(n19999), .A(n19968), .ZN(U240) );
  AOI22_X1 U21990 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10979), .ZN(n19969) );
  OAI21_X1 U21991 ( .B1(n13666), .B2(n19999), .A(n19969), .ZN(U239) );
  AOI22_X1 U21992 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10979), .ZN(n19970) );
  OAI21_X1 U21993 ( .B1(n13661), .B2(n19999), .A(n19970), .ZN(U238) );
  AOI22_X1 U21994 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10979), .ZN(n19971) );
  OAI21_X1 U21995 ( .B1(n19972), .B2(n19999), .A(n19971), .ZN(U237) );
  AOI22_X1 U21996 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10979), .ZN(n19973) );
  OAI21_X1 U21997 ( .B1(n19974), .B2(n19999), .A(n19973), .ZN(U236) );
  AOI22_X1 U21998 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10979), .ZN(n19975) );
  OAI21_X1 U21999 ( .B1(n19976), .B2(n19999), .A(n19975), .ZN(U235) );
  AOI22_X1 U22000 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10979), .ZN(n19977) );
  OAI21_X1 U22001 ( .B1(n13680), .B2(n19999), .A(n19977), .ZN(U234) );
  AOI22_X1 U22002 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10979), .ZN(n19978) );
  OAI21_X1 U22003 ( .B1(n19979), .B2(n19999), .A(n19978), .ZN(U233) );
  INV_X1 U22004 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22005 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10979), .ZN(n19980) );
  OAI21_X1 U22006 ( .B1(n19981), .B2(n19999), .A(n19980), .ZN(U232) );
  INV_X1 U22007 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n21675) );
  AOI22_X1 U22008 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10979), .ZN(n19982) );
  OAI21_X1 U22009 ( .B1(n21675), .B2(n19999), .A(n19982), .ZN(U231) );
  INV_X1 U22010 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n21860) );
  AOI22_X1 U22011 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10979), .ZN(n19983) );
  OAI21_X1 U22012 ( .B1(n21860), .B2(n19999), .A(n19983), .ZN(U230) );
  INV_X1 U22013 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21903) );
  AOI22_X1 U22014 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10979), .ZN(n19984) );
  OAI21_X1 U22015 ( .B1(n21903), .B2(n19999), .A(n19984), .ZN(U229) );
  INV_X1 U22016 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n21947) );
  AOI22_X1 U22017 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10979), .ZN(n19985) );
  OAI21_X1 U22018 ( .B1(n21947), .B2(n19999), .A(n19985), .ZN(U228) );
  INV_X1 U22019 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21992) );
  AOI22_X1 U22020 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10979), .ZN(n19986) );
  OAI21_X1 U22021 ( .B1(n21992), .B2(n19999), .A(n19986), .ZN(U227) );
  AOI22_X1 U22022 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10979), .ZN(n19987) );
  OAI21_X1 U22023 ( .B1(n22039), .B2(n19999), .A(n19987), .ZN(U226) );
  INV_X1 U22024 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n22085) );
  AOI22_X1 U22025 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10979), .ZN(n19988) );
  OAI21_X1 U22026 ( .B1(n22085), .B2(n19999), .A(n19988), .ZN(U225) );
  AOI22_X1 U22027 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10979), .ZN(n19989) );
  OAI21_X1 U22028 ( .B1(n22135), .B2(n19999), .A(n19989), .ZN(U224) );
  AOI22_X1 U22029 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10979), .ZN(n19990) );
  OAI21_X1 U22030 ( .B1(n16343), .B2(n19999), .A(n19990), .ZN(U223) );
  INV_X1 U22031 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n21858) );
  AOI22_X1 U22032 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10979), .ZN(n19991) );
  OAI21_X1 U22033 ( .B1(n21858), .B2(n19999), .A(n19991), .ZN(U222) );
  INV_X1 U22034 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21901) );
  AOI22_X1 U22035 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10979), .ZN(n19992) );
  OAI21_X1 U22036 ( .B1(n21901), .B2(n19999), .A(n19992), .ZN(U221) );
  INV_X1 U22037 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n21945) );
  AOI22_X1 U22038 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10979), .ZN(n19994) );
  OAI21_X1 U22039 ( .B1(n21945), .B2(n19999), .A(n19994), .ZN(U220) );
  INV_X1 U22040 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n21990) );
  AOI22_X1 U22041 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10979), .ZN(n19995) );
  OAI21_X1 U22042 ( .B1(n21990), .B2(n19999), .A(n19995), .ZN(U219) );
  INV_X1 U22043 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n22036) );
  AOI22_X1 U22044 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10979), .ZN(n19996) );
  OAI21_X1 U22045 ( .B1(n22036), .B2(n19999), .A(n19996), .ZN(U218) );
  INV_X1 U22046 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n22084) );
  AOI22_X1 U22047 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n19993), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10979), .ZN(n19997) );
  OAI21_X1 U22048 ( .B1(n22084), .B2(n19999), .A(n19997), .ZN(U217) );
  INV_X1 U22049 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n22130) );
  OAI222_X1 U22050 ( .A1(U212), .A2(n20000), .B1(n19999), .B2(n22130), .C1(
        U214), .C2(n19998), .ZN(U216) );
  INV_X1 U22051 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20001) );
  AOI22_X1 U22052 ( .A1(n22246), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20001), 
        .B2(n19831), .ZN(P1_U3483) );
  OAI21_X1 U22053 ( .B1(n21628), .B2(n20002), .A(n20059), .ZN(n20003) );
  AOI21_X1 U22054 ( .B1(n20004), .B2(n21218), .A(n20003), .ZN(n20011) );
  INV_X1 U22055 ( .A(n20739), .ZN(n20005) );
  AOI21_X1 U22056 ( .B1(n20063), .B2(n21574), .A(n20005), .ZN(n20007) );
  OAI211_X1 U22057 ( .C1(n20007), .C2(n20006), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n21198), .ZN(n20008) );
  AOI21_X1 U22058 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20008), .A(n21210), 
        .ZN(n20010) );
  NAND2_X1 U22059 ( .A1(n20011), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20009) );
  OAI21_X1 U22060 ( .B1(n20011), .B2(n20010), .A(n20009), .ZN(P3_U3296) );
  AOI22_X1 U22061 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20050), .ZN(n20014) );
  OAI21_X1 U22062 ( .B1(n20677), .B2(n20048), .A(n20014), .ZN(P3_U2768) );
  AOI22_X1 U22063 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20051), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20050), .ZN(n20015) );
  OAI21_X1 U22064 ( .B1(n20568), .B2(n20053), .A(n20015), .ZN(P3_U2769) );
  AOI22_X1 U22065 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20050), .ZN(n20016) );
  OAI21_X1 U22066 ( .B1(n20551), .B2(n20048), .A(n20016), .ZN(P3_U2770) );
  AOI22_X1 U22067 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20051), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20050), .ZN(n20017) );
  OAI21_X1 U22068 ( .B1(n20577), .B2(n20053), .A(n20017), .ZN(P3_U2771) );
  AOI22_X1 U22069 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20050), .ZN(n20018) );
  OAI21_X1 U22070 ( .B1(n20543), .B2(n20048), .A(n20018), .ZN(P3_U2772) );
  AOI22_X1 U22071 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20043), .ZN(n20019) );
  OAI21_X1 U22072 ( .B1(n20538), .B2(n20048), .A(n20019), .ZN(P3_U2773) );
  AOI22_X1 U22073 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20043), .ZN(n20020) );
  OAI21_X1 U22074 ( .B1(n20534), .B2(n20048), .A(n20020), .ZN(P3_U2774) );
  AOI22_X1 U22075 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20043), .ZN(n20021) );
  OAI21_X1 U22076 ( .B1(n20529), .B2(n20048), .A(n20021), .ZN(P3_U2775) );
  AOI22_X1 U22077 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20051), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20043), .ZN(n20022) );
  OAI21_X1 U22078 ( .B1(n11276), .B2(n20053), .A(n20022), .ZN(P3_U2776) );
  AOI22_X1 U22079 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20051), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20043), .ZN(n20023) );
  OAI21_X1 U22080 ( .B1(n20024), .B2(n20053), .A(n20023), .ZN(P3_U2777) );
  INV_X1 U22081 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20522) );
  AOI22_X1 U22082 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20043), .ZN(n20025) );
  OAI21_X1 U22083 ( .B1(n20522), .B2(n20048), .A(n20025), .ZN(P3_U2778) );
  INV_X1 U22084 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20517) );
  AOI22_X1 U22085 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20043), .ZN(n20026) );
  OAI21_X1 U22086 ( .B1(n20517), .B2(n20048), .A(n20026), .ZN(P3_U2779) );
  AOI22_X1 U22087 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20051), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20050), .ZN(n20027) );
  OAI21_X1 U22088 ( .B1(n20614), .B2(n20053), .A(n20027), .ZN(P3_U2780) );
  INV_X1 U22089 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n20509) );
  AOI22_X1 U22090 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n20046), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20050), .ZN(n20028) );
  OAI21_X1 U22091 ( .B1(n20509), .B2(n20048), .A(n20028), .ZN(P3_U2781) );
  AOI22_X1 U22092 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20051), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20050), .ZN(n20029) );
  OAI21_X1 U22093 ( .B1(n20030), .B2(n20053), .A(n20029), .ZN(P3_U2782) );
  AOI22_X1 U22094 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20050), .ZN(n20031) );
  OAI21_X1 U22095 ( .B1(n20677), .B2(n20048), .A(n20031), .ZN(P3_U2783) );
  AOI22_X1 U22096 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20050), .ZN(n20032) );
  OAI21_X1 U22097 ( .B1(n20664), .B2(n20053), .A(n20032), .ZN(P3_U2784) );
  AOI22_X1 U22098 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20050), .ZN(n20033) );
  OAI21_X1 U22099 ( .B1(n20551), .B2(n20048), .A(n20033), .ZN(P3_U2785) );
  AOI22_X1 U22100 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20050), .ZN(n20034) );
  OAI21_X1 U22101 ( .B1(n20546), .B2(n20053), .A(n20034), .ZN(P3_U2786) );
  AOI22_X1 U22102 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20050), .ZN(n20035) );
  OAI21_X1 U22103 ( .B1(n20543), .B2(n20048), .A(n20035), .ZN(P3_U2787) );
  AOI22_X1 U22104 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20050), .ZN(n20036) );
  OAI21_X1 U22105 ( .B1(n20538), .B2(n20048), .A(n20036), .ZN(P3_U2788) );
  AOI22_X1 U22106 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20050), .ZN(n20037) );
  OAI21_X1 U22107 ( .B1(n20534), .B2(n20048), .A(n20037), .ZN(P3_U2789) );
  AOI22_X1 U22108 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20050), .ZN(n20038) );
  OAI21_X1 U22109 ( .B1(n20529), .B2(n20048), .A(n20038), .ZN(P3_U2790) );
  AOI22_X1 U22110 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20050), .ZN(n20039) );
  OAI21_X1 U22111 ( .B1(n20655), .B2(n20053), .A(n20039), .ZN(P3_U2791) );
  AOI22_X1 U22112 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20043), .ZN(n20040) );
  OAI21_X1 U22113 ( .B1(n20552), .B2(n20053), .A(n20040), .ZN(P3_U2792) );
  AOI22_X1 U22114 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20043), .ZN(n20041) );
  OAI21_X1 U22115 ( .B1(n20522), .B2(n20048), .A(n20041), .ZN(P3_U2793) );
  AOI22_X1 U22116 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20043), .ZN(n20042) );
  OAI21_X1 U22117 ( .B1(n20517), .B2(n20048), .A(n20042), .ZN(P3_U2794) );
  AOI22_X1 U22118 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20043), .ZN(n20044) );
  OAI21_X1 U22119 ( .B1(n20045), .B2(n20053), .A(n20044), .ZN(P3_U2795) );
  AOI22_X1 U22120 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20046), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20050), .ZN(n20047) );
  OAI21_X1 U22121 ( .B1(n20509), .B2(n20048), .A(n20047), .ZN(P3_U2796) );
  AOI22_X1 U22122 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20050), .ZN(n20049) );
  OAI21_X1 U22123 ( .B1(n20644), .B2(n20053), .A(n20049), .ZN(P3_U2797) );
  AOI22_X1 U22124 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20051), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20050), .ZN(n20052) );
  OAI21_X1 U22125 ( .B1(n20650), .B2(n20053), .A(n20052), .ZN(P3_U2798) );
  NAND2_X1 U22126 ( .A1(n20054), .A2(n20713), .ZN(n20683) );
  INV_X1 U22127 ( .A(n20088), .ZN(n20493) );
  NOR2_X1 U22128 ( .A1(n20064), .A2(n20063), .ZN(n20056) );
  OAI211_X2 U22129 ( .C1(n21628), .C2(P3_STATEBS16_REG_SCAN_IN), .A(n20062), 
        .B(n20056), .ZN(n20486) );
  NAND4_X1 U22130 ( .A1(n20057), .A2(n21075), .A3(n21574), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n21205) );
  NAND2_X1 U22131 ( .A1(n21201), .A2(n20058), .ZN(n21216) );
  AOI22_X1 U22132 ( .A1(n20451), .A2(n20060), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n20407), .ZN(n20070) );
  INV_X1 U22133 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20289) );
  NOR2_X1 U22134 ( .A1(n20458), .A2(n21205), .ZN(n20081) );
  INV_X1 U22135 ( .A(n20081), .ZN(n20473) );
  OAI21_X1 U22136 ( .B1(n20289), .B2(n20473), .A(n20484), .ZN(n20068) );
  AOI21_X1 U22137 ( .B1(n20269), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21205), .ZN(n20133) );
  OAI211_X1 U22138 ( .C1(n20738), .C2(n20739), .A(n21198), .B(n21574), .ZN(
        n21197) );
  INV_X1 U22139 ( .A(n21197), .ZN(n20061) );
  OAI211_X2 U22140 ( .C1(n20064), .C2(n20063), .A(n21197), .B(n20062), .ZN(
        n20487) );
  OAI22_X1 U22141 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20419), .B1(n20487), 
        .B2(n20065), .ZN(n20066) );
  AOI221_X1 U22142 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20068), .C1(
        n20067), .C2(n20133), .A(n20066), .ZN(n20069) );
  OAI211_X1 U22143 ( .C1(n20683), .C2(n20493), .A(n20070), .B(n20069), .ZN(
        P3_U2670) );
  INV_X1 U22144 ( .A(n21205), .ZN(n20463) );
  NAND2_X1 U22145 ( .A1(n20463), .A2(n20458), .ZN(n20291) );
  INV_X1 U22146 ( .A(n20071), .ZN(n20072) );
  NOR3_X1 U22147 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20095) );
  AOI211_X1 U22148 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20072), .A(n20095), .B(
        n20486), .ZN(n20080) );
  OAI21_X1 U22149 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20704), .A(
        n20721), .ZN(n20699) );
  OAI22_X1 U22150 ( .A1(n20075), .A2(n20490), .B1(n20699), .B2(n20493), .ZN(
        n20073) );
  INV_X1 U22151 ( .A(n20073), .ZN(n20077) );
  NOR2_X1 U22152 ( .A1(n20075), .A2(n20074), .ZN(n20090) );
  INV_X1 U22153 ( .A(n20090), .ZN(n20086) );
  OAI211_X1 U22154 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20404), .B(n20086), .ZN(n20076) );
  OAI211_X1 U22155 ( .C1(n20078), .C2(n20487), .A(n20077), .B(n20076), .ZN(
        n20079) );
  AOI211_X1 U22156 ( .C1(n20432), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20080), .B(n20079), .ZN(n20084) );
  NAND2_X1 U22157 ( .A1(n20289), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20102) );
  INV_X1 U22158 ( .A(n20102), .ZN(n20311) );
  OAI221_X1 U22159 ( .B1(n20311), .B2(n20085), .C1(n20102), .C2(n20082), .A(
        n20081), .ZN(n20083) );
  OAI211_X1 U22160 ( .C1(n20291), .C2(n20085), .A(n20084), .B(n20083), .ZN(
        P3_U2669) );
  AOI22_X1 U22161 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20432), .B1(
        n20472), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n20099) );
  NOR2_X1 U22162 ( .A1(n20796), .A2(n20086), .ZN(n20117) );
  NOR2_X1 U22163 ( .A1(n20117), .A2(n20419), .ZN(n20089) );
  NAND2_X1 U22164 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20721), .ZN(
        n20087) );
  NAND2_X1 U22165 ( .A1(n11511), .A2(n20087), .ZN(n20729) );
  AOI22_X1 U22166 ( .A1(n20090), .A2(n20089), .B1(n20088), .B2(n20729), .ZN(
        n20098) );
  AOI21_X1 U22167 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20311), .A(
        n20458), .ZN(n20092) );
  XNOR2_X1 U22168 ( .A(n20092), .B(n20091), .ZN(n20093) );
  OAI21_X1 U22169 ( .B1(n20117), .B2(n20419), .A(n20490), .ZN(n20109) );
  AOI22_X1 U22170 ( .A1(n20463), .A2(n20093), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n20109), .ZN(n20097) );
  INV_X1 U22171 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20094) );
  NAND2_X1 U22172 ( .A1(n20095), .A2(n20094), .ZN(n20104) );
  OAI211_X1 U22173 ( .C1(n20095), .C2(n20094), .A(n20451), .B(n20104), .ZN(
        n20096) );
  NAND4_X1 U22174 ( .A1(n20099), .A2(n20098), .A3(n20097), .A4(n20096), .ZN(
        P3_U2668) );
  AOI21_X1 U22175 ( .B1(n11024), .B2(n20100), .A(n20493), .ZN(n20101) );
  AOI211_X1 U22176 ( .C1(n20472), .C2(P3_EBX_REG_4__SCAN_IN), .A(n21156), .B(
        n20101), .ZN(n20114) );
  OAI21_X1 U22177 ( .B1(n20103), .B2(n20102), .A(n20269), .ZN(n20115) );
  NOR3_X1 U22178 ( .A1(n20108), .A2(n21205), .A3(n20115), .ZN(n20106) );
  NOR2_X1 U22179 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20104), .ZN(n20126) );
  AOI211_X1 U22180 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20104), .A(n20126), .B(
        n20486), .ZN(n20105) );
  AOI211_X1 U22181 ( .C1(n20432), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20106), .B(n20105), .ZN(n20113) );
  INV_X1 U22182 ( .A(n20133), .ZN(n20267) );
  AOI21_X1 U22183 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20291), .A(
        n20267), .ZN(n20107) );
  AOI22_X1 U22184 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20109), .B1(n20108), 
        .B2(n20107), .ZN(n20112) );
  NAND3_X1 U22185 ( .A1(n20404), .A2(n20117), .A3(n20110), .ZN(n20111) );
  NAND4_X1 U22186 ( .A1(n20114), .A2(n20113), .A3(n20112), .A4(n20111), .ZN(
        P3_U2667) );
  XOR2_X1 U22187 ( .A(n20116), .B(n20115), .Z(n20124) );
  NAND2_X1 U22188 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20117), .ZN(n20118) );
  NOR2_X1 U22189 ( .A1(n20122), .A2(n20118), .ZN(n20144) );
  NOR2_X1 U22190 ( .A1(n20144), .A2(n20419), .ZN(n20119) );
  NOR2_X1 U22191 ( .A1(n20407), .A2(n20119), .ZN(n20143) );
  INV_X1 U22192 ( .A(n20118), .ZN(n20120) );
  AOI22_X1 U22193 ( .A1(n20472), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n20120), .B2(
        n20119), .ZN(n20121) );
  OAI211_X1 U22194 ( .C1(n20143), .C2(n20122), .A(n20121), .B(n21129), .ZN(
        n20123) );
  AOI21_X1 U22195 ( .B1(n20463), .B2(n20124), .A(n20123), .ZN(n20128) );
  NAND2_X1 U22196 ( .A1(n20126), .A2(n20125), .ZN(n20132) );
  OAI211_X1 U22197 ( .C1(n20126), .C2(n20125), .A(n20451), .B(n20132), .ZN(
        n20127) );
  OAI211_X1 U22198 ( .C1(n20484), .C2(n11302), .A(n20128), .B(n20127), .ZN(
        P3_U2666) );
  NOR2_X1 U22199 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20129), .ZN(
        n20199) );
  NOR2_X1 U22200 ( .A1(n20199), .A2(n20458), .ZN(n20130) );
  NAND2_X1 U22201 ( .A1(n20463), .A2(n20130), .ZN(n20149) );
  INV_X1 U22202 ( .A(n20149), .ZN(n20131) );
  AOI22_X1 U22203 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20432), .B1(
        n20131), .B2(n20136), .ZN(n20140) );
  NOR2_X1 U22204 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20132), .ZN(n20147) );
  AOI211_X1 U22205 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20132), .A(n20147), .B(
        n20486), .ZN(n20138) );
  OAI21_X1 U22206 ( .B1(n20458), .B2(n20134), .A(n20133), .ZN(n20135) );
  NAND3_X1 U22207 ( .A1(n20404), .A2(n20144), .A3(n20141), .ZN(n20142) );
  OAI211_X1 U22208 ( .C1(n20136), .C2(n20135), .A(n21129), .B(n20142), .ZN(
        n20137) );
  AOI211_X1 U22209 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20472), .A(n20138), .B(
        n20137), .ZN(n20139) );
  OAI211_X1 U22210 ( .C1(n20143), .C2(n20141), .A(n20140), .B(n20139), .ZN(
        P3_U2665) );
  OAI21_X1 U22211 ( .B1(n20199), .B2(n20458), .A(n20150), .ZN(n20156) );
  AOI21_X1 U22212 ( .B1(n20143), .B2(n20142), .A(n20835), .ZN(n20154) );
  NAND2_X1 U22213 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20144), .ZN(n20157) );
  NOR3_X1 U22214 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20419), .A3(n20157), .ZN(
        n20153) );
  OAI22_X1 U22215 ( .A1(n20145), .A2(n20484), .B1(n20487), .B2(n20146), .ZN(
        n20152) );
  NAND2_X1 U22216 ( .A1(n20147), .A2(n20146), .ZN(n20160) );
  OAI211_X1 U22217 ( .C1(n20147), .C2(n20146), .A(n20451), .B(n20160), .ZN(
        n20148) );
  OAI21_X1 U22218 ( .B1(n20150), .B2(n20149), .A(n20148), .ZN(n20151) );
  NOR4_X1 U22219 ( .A1(n20154), .A2(n20153), .A3(n20152), .A4(n20151), .ZN(
        n20155) );
  OAI211_X1 U22220 ( .C1(n21205), .C2(n20156), .A(n20155), .B(n21129), .ZN(
        P3_U2664) );
  NOR2_X1 U22221 ( .A1(n20835), .A2(n20157), .ZN(n20159) );
  NAND2_X1 U22222 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20159), .ZN(n20173) );
  NOR2_X1 U22223 ( .A1(n20192), .A2(n20419), .ZN(n20158) );
  AOI22_X1 U22224 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20432), .B1(
        n20159), .B2(n20158), .ZN(n20168) );
  NOR2_X1 U22225 ( .A1(n20187), .A2(n20486), .ZN(n20178) );
  NAND2_X1 U22226 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20160), .ZN(n20161) );
  AOI22_X1 U22227 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20472), .B1(n20178), .B2(
        n20161), .ZN(n20167) );
  AOI21_X1 U22228 ( .B1(n20162), .B2(n20289), .A(n20458), .ZN(n20164) );
  XNOR2_X1 U22229 ( .A(n20164), .B(n20163), .ZN(n20165) );
  OAI21_X1 U22230 ( .B1(n20419), .B2(n20192), .A(n20490), .ZN(n20174) );
  AOI22_X1 U22231 ( .A1(n20463), .A2(n20165), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n20174), .ZN(n20166) );
  NAND4_X1 U22232 ( .A1(n20168), .A2(n20167), .A3(n20166), .A4(n21129), .ZN(
        P3_U2663) );
  INV_X1 U22233 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20181) );
  NOR2_X1 U22234 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20169), .ZN(
        n20185) );
  NOR2_X1 U22235 ( .A1(n20185), .A2(n20473), .ZN(n20182) );
  AOI211_X1 U22236 ( .C1(n20269), .C2(n20170), .A(n20267), .B(n20172), .ZN(
        n20171) );
  AOI211_X1 U22237 ( .C1(n20182), .C2(n20172), .A(n21156), .B(n20171), .ZN(
        n20180) );
  INV_X1 U22238 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20186) );
  NOR3_X1 U22239 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20419), .A3(n20173), .ZN(
        n20177) );
  INV_X1 U22240 ( .A(n20174), .ZN(n20191) );
  AOI21_X1 U22241 ( .B1(n20451), .B2(n20187), .A(n20472), .ZN(n20175) );
  OAI22_X1 U22242 ( .A1(n20191), .A2(n21154), .B1(n20186), .B2(n20175), .ZN(
        n20176) );
  AOI211_X1 U22243 ( .C1(n20178), .C2(n20186), .A(n20177), .B(n20176), .ZN(
        n20179) );
  OAI211_X1 U22244 ( .C1(n20181), .C2(n20484), .A(n20180), .B(n20179), .ZN(
        P3_U2662) );
  AOI21_X1 U22245 ( .B1(n20183), .B2(n20463), .A(n20182), .ZN(n20198) );
  INV_X1 U22246 ( .A(n20183), .ZN(n20184) );
  NOR3_X1 U22247 ( .A1(n20185), .A2(n20184), .A3(n20458), .ZN(n20197) );
  NAND2_X1 U22248 ( .A1(n20187), .A2(n20186), .ZN(n20188) );
  AOI211_X1 U22249 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20188), .A(n20207), .B(
        n20486), .ZN(n20189) );
  AOI211_X1 U22250 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n20432), .A(
        n21156), .B(n20189), .ZN(n20196) );
  NAND2_X1 U22251 ( .A1(n20404), .A2(n21154), .ZN(n20190) );
  AOI21_X1 U22252 ( .B1(n20191), .B2(n20190), .A(n20204), .ZN(n20194) );
  NAND2_X1 U22253 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20192), .ZN(n20203) );
  NOR3_X1 U22254 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20419), .A3(n20203), 
        .ZN(n20193) );
  AOI211_X1 U22255 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20472), .A(n20194), .B(
        n20193), .ZN(n20195) );
  OAI211_X1 U22256 ( .C1(n20198), .C2(n20197), .A(n20196), .B(n20195), .ZN(
        P3_U2661) );
  NAND2_X1 U22257 ( .A1(n20200), .A2(n20199), .ZN(n20216) );
  NAND2_X1 U22258 ( .A1(n20269), .A2(n20216), .ZN(n20202) );
  XOR2_X1 U22259 ( .A(n20202), .B(n20201), .Z(n20212) );
  OR2_X1 U22260 ( .A1(n20204), .A2(n20203), .ZN(n20215) );
  NOR2_X1 U22261 ( .A1(n20419), .A2(n20215), .ZN(n20205) );
  NAND2_X1 U22262 ( .A1(n20419), .A2(n20490), .ZN(n20488) );
  NOR2_X1 U22263 ( .A1(n20871), .A2(n20215), .ZN(n20284) );
  NAND2_X1 U22264 ( .A1(n20284), .A2(n20490), .ZN(n20242) );
  AND2_X1 U22265 ( .A1(n20488), .A2(n20242), .ZN(n20232) );
  OAI21_X1 U22266 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n20205), .A(n20232), 
        .ZN(n20209) );
  INV_X1 U22267 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20206) );
  NAND2_X1 U22268 ( .A1(n20207), .A2(n20206), .ZN(n20213) );
  OAI211_X1 U22269 ( .C1(n20207), .C2(n20206), .A(n20451), .B(n20213), .ZN(
        n20208) );
  OAI211_X1 U22270 ( .C1(n20484), .C2(n20217), .A(n20209), .B(n20208), .ZN(
        n20210) );
  AOI211_X1 U22271 ( .C1(n20472), .C2(P3_EBX_REG_11__SCAN_IN), .A(n21156), .B(
        n20210), .ZN(n20211) );
  OAI21_X1 U22272 ( .B1(n20212), .B2(n21205), .A(n20211), .ZN(P3_U2660) );
  AOI211_X1 U22273 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20213), .A(n20234), .B(
        n20486), .ZN(n20214) );
  AOI211_X1 U22274 ( .C1(n20472), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21156), .B(
        n20214), .ZN(n20224) );
  NOR2_X1 U22275 ( .A1(n20217), .A2(n20216), .ZN(n20254) );
  NOR2_X1 U22276 ( .A1(n20254), .A2(n20458), .ZN(n20219) );
  OAI21_X1 U22277 ( .B1(n20220), .B2(n20219), .A(n20463), .ZN(n20218) );
  AOI21_X1 U22278 ( .B1(n20220), .B2(n20219), .A(n20218), .ZN(n20221) );
  AOI221_X1 U22279 ( .B1(n20232), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n20253), 
        .C2(n20222), .A(n20221), .ZN(n20223) );
  OAI211_X1 U22280 ( .C1(n20225), .C2(n20484), .A(n20224), .B(n20223), .ZN(
        P3_U2659) );
  AOI211_X1 U22281 ( .C1(n20226), .C2(n20291), .A(n20267), .B(n20228), .ZN(
        n20227) );
  AOI21_X1 U22282 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n20472), .A(n20227), .ZN(
        n20238) );
  OAI21_X1 U22283 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20243), .A(
        n20228), .ZN(n20229) );
  OAI22_X1 U22284 ( .A1(n20230), .A2(n20484), .B1(n20473), .B2(n20229), .ZN(
        n20231) );
  AOI211_X1 U22285 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n20232), .A(n21156), 
        .B(n20231), .ZN(n20237) );
  NAND2_X1 U22286 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20240) );
  OAI211_X1 U22287 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(P3_REIP_REG_12__SCAN_IN), .A(n20253), .B(n20240), .ZN(n20236) );
  NAND2_X1 U22288 ( .A1(n20234), .A2(n20233), .ZN(n20239) );
  OAI211_X1 U22289 ( .C1(n20234), .C2(n20233), .A(n20451), .B(n20239), .ZN(
        n20235) );
  NAND4_X1 U22290 ( .A1(n20238), .A2(n20237), .A3(n20236), .A4(n20235), .ZN(
        P3_U2658) );
  INV_X1 U22291 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20251) );
  AOI211_X1 U22292 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20239), .A(n20258), .B(
        n20486), .ZN(n20249) );
  INV_X1 U22293 ( .A(n20240), .ZN(n20241) );
  AOI21_X1 U22294 ( .B1(n20241), .B2(n20253), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n20247) );
  NAND2_X1 U22295 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n20241), .ZN(n20252) );
  OAI21_X1 U22296 ( .B1(n20252), .B2(n20242), .A(n20488), .ZN(n20271) );
  OAI21_X1 U22297 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20243), .A(
        n20269), .ZN(n20244) );
  XOR2_X1 U22298 ( .A(n20245), .B(n20244), .Z(n20246) );
  OAI22_X1 U22299 ( .A1(n20247), .A2(n20271), .B1(n21205), .B2(n20246), .ZN(
        n20248) );
  AOI211_X1 U22300 ( .C1(n20432), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20249), .B(n20248), .ZN(n20250) );
  OAI211_X1 U22301 ( .C1(n20487), .C2(n20251), .A(n20250), .B(n21129), .ZN(
        P3_U2657) );
  INV_X1 U22302 ( .A(n20252), .ZN(n20283) );
  NAND2_X1 U22303 ( .A1(n20283), .A2(n20253), .ZN(n20282) );
  NAND4_X1 U22304 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A4(n20254), .ZN(n20264) );
  NAND2_X1 U22305 ( .A1(n20269), .A2(n20264), .ZN(n20256) );
  OAI21_X1 U22306 ( .B1(n20257), .B2(n20256), .A(n20463), .ZN(n20255) );
  AOI21_X1 U22307 ( .B1(n20257), .B2(n20256), .A(n20255), .ZN(n20262) );
  NAND2_X1 U22308 ( .A1(n20258), .A2(n20260), .ZN(n20270) );
  OAI211_X1 U22309 ( .C1(n20258), .C2(n20260), .A(n20451), .B(n20270), .ZN(
        n20259) );
  OAI211_X1 U22310 ( .C1(n20487), .C2(n20260), .A(n21129), .B(n20259), .ZN(
        n20261) );
  AOI211_X1 U22311 ( .C1(n20432), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20262), .B(n20261), .ZN(n20263) );
  OAI221_X1 U22312 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n20282), .C1(n20280), 
        .C2(n20271), .A(n20263), .ZN(P3_U2656) );
  NOR2_X1 U22313 ( .A1(n20265), .A2(n20264), .ZN(n20329) );
  NOR3_X1 U22314 ( .A1(n20329), .A2(n20275), .A3(n20473), .ZN(n20266) );
  AOI211_X1 U22315 ( .C1(n20472), .C2(P3_EBX_REG_16__SCAN_IN), .A(n21156), .B(
        n20266), .ZN(n20278) );
  AOI21_X1 U22316 ( .B1(n20269), .B2(n20268), .A(n20267), .ZN(n20276) );
  NOR2_X1 U22317 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20270), .ZN(n20285) );
  AOI211_X1 U22318 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20270), .A(n20285), .B(
        n20486), .ZN(n20274) );
  XOR2_X1 U22319 ( .A(P3_REIP_REG_16__SCAN_IN), .B(n20280), .Z(n20272) );
  OAI22_X1 U22320 ( .A1(n20282), .A2(n20272), .B1(n20281), .B2(n20271), .ZN(
        n20273) );
  AOI211_X1 U22321 ( .C1(n20276), .C2(n20275), .A(n20274), .B(n20273), .ZN(
        n20277) );
  OAI211_X1 U22322 ( .C1(n20279), .C2(n20484), .A(n20278), .B(n20277), .ZN(
        P3_U2655) );
  NOR2_X1 U22323 ( .A1(n20281), .A2(n20280), .ZN(n20298) );
  INV_X1 U22324 ( .A(n20282), .ZN(n20297) );
  AOI21_X1 U22325 ( .B1(n20298), .B2(n20297), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n20296) );
  NAND4_X1 U22326 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20284), .A3(n20283), 
        .A4(n20298), .ZN(n20326) );
  AOI21_X1 U22327 ( .B1(n20404), .B2(n20326), .A(n20407), .ZN(n20320) );
  INV_X1 U22328 ( .A(n20285), .ZN(n20286) );
  AOI21_X1 U22329 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n20286), .A(n20486), .ZN(
        n20287) );
  AOI22_X1 U22330 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20432), .B1(
        n20287), .B2(n20303), .ZN(n20295) );
  AOI21_X1 U22331 ( .B1(n20289), .B2(n20288), .A(n20458), .ZN(n20301) );
  INV_X1 U22332 ( .A(n20301), .ZN(n20299) );
  OAI21_X1 U22333 ( .B1(n20329), .B2(n20292), .A(n20463), .ZN(n20290) );
  AOI22_X1 U22334 ( .A1(n20292), .A2(n20299), .B1(n20291), .B2(n20290), .ZN(
        n20293) );
  AOI211_X1 U22335 ( .C1(n20472), .C2(P3_EBX_REG_17__SCAN_IN), .A(n21156), .B(
        n20293), .ZN(n20294) );
  OAI211_X1 U22336 ( .C1(n20296), .C2(n20320), .A(n20295), .B(n20294), .ZN(
        P3_U2654) );
  NAND3_X1 U22337 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20298), .A3(n20297), 
        .ZN(n20319) );
  AOI221_X1 U22338 ( .B1(n20302), .B2(n20301), .C1(n20300), .C2(n20299), .A(
        n21205), .ZN(n20308) );
  AOI211_X1 U22339 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20303), .A(n20315), .B(
        n20486), .ZN(n20307) );
  OAI22_X1 U22340 ( .A1(n20305), .A2(n20484), .B1(n20487), .B2(n20304), .ZN(
        n20306) );
  NOR4_X1 U22341 ( .A1(n21156), .A2(n20308), .A3(n20307), .A4(n20306), .ZN(
        n20309) );
  OAI221_X1 U22342 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n20319), .C1(n20310), 
        .C2(n20320), .A(n20309), .ZN(P3_U2653) );
  AOI21_X1 U22343 ( .B1(n20312), .B2(n20311), .A(n20458), .ZN(n20313) );
  XOR2_X1 U22344 ( .A(n20314), .B(n20313), .Z(n20325) );
  NAND2_X1 U22345 ( .A1(n20315), .A2(n20317), .ZN(n20328) );
  OAI211_X1 U22346 ( .C1(n20315), .C2(n20317), .A(n20451), .B(n20328), .ZN(
        n20316) );
  OAI211_X1 U22347 ( .C1(n20487), .C2(n20317), .A(n21129), .B(n20316), .ZN(
        n20323) );
  NAND2_X1 U22348 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n20327) );
  OAI21_X1 U22349 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), 
        .A(n20327), .ZN(n20318) );
  OAI22_X1 U22350 ( .A1(n20321), .A2(n20320), .B1(n20319), .B2(n20318), .ZN(
        n20322) );
  AOI211_X1 U22351 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n20432), .A(
        n20323), .B(n20322), .ZN(n20324) );
  OAI21_X1 U22352 ( .B1(n21205), .B2(n20325), .A(n20324), .ZN(P3_U2652) );
  NOR2_X1 U22353 ( .A1(n20327), .A2(n20326), .ZN(n20336) );
  NAND2_X1 U22354 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20336), .ZN(n20353) );
  AOI21_X1 U22355 ( .B1(n20353), .B2(n20404), .A(n20407), .ZN(n20340) );
  AOI22_X1 U22356 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20432), .B1(
        n20472), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n20338) );
  NOR2_X1 U22357 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20419), .ZN(n20335) );
  AOI211_X1 U22358 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20328), .A(n20344), .B(
        n20486), .ZN(n20334) );
  AOI21_X1 U22359 ( .B1(n20330), .B2(n20329), .A(n20458), .ZN(n20331) );
  NOR2_X1 U22360 ( .A1(n20332), .A2(n20331), .ZN(n20341) );
  AOI211_X1 U22361 ( .C1(n20332), .C2(n20331), .A(n20341), .B(n21205), .ZN(
        n20333) );
  AOI211_X1 U22362 ( .C1(n20336), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        n20337) );
  OAI211_X1 U22363 ( .C1(n20339), .C2(n20340), .A(n20338), .B(n20337), .ZN(
        P3_U2651) );
  INV_X1 U22364 ( .A(n20340), .ZN(n20349) );
  NOR2_X1 U22365 ( .A1(n20341), .A2(n20458), .ZN(n20342) );
  AOI211_X1 U22366 ( .C1(n20343), .C2(n20342), .A(n20356), .B(n21205), .ZN(
        n20348) );
  NAND2_X1 U22367 ( .A1(n20344), .A2(n20352), .ZN(n20355) );
  OAI211_X1 U22368 ( .C1(n20344), .C2(n20352), .A(n20451), .B(n20355), .ZN(
        n20345) );
  OAI21_X1 U22369 ( .B1(n20484), .B2(n20346), .A(n20345), .ZN(n20347) );
  AOI211_X1 U22370 ( .C1(n20349), .C2(P3_REIP_REG_21__SCAN_IN), .A(n20348), 
        .B(n20347), .ZN(n20351) );
  OR3_X1 U22371 ( .A1(n20419), .A2(n20353), .A3(P3_REIP_REG_21__SCAN_IN), .ZN(
        n20350) );
  OAI211_X1 U22372 ( .C1(n20352), .C2(n20487), .A(n20351), .B(n20350), .ZN(
        P3_U2650) );
  AOI221_X1 U22373 ( .B1(n20354), .B2(n20404), .C1(n20353), .C2(n20404), .A(
        n20407), .ZN(n20365) );
  AOI22_X1 U22374 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20432), .B1(
        n20472), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n20363) );
  NOR2_X1 U22375 ( .A1(n20354), .A2(n20353), .ZN(n20366) );
  NOR2_X1 U22376 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20419), .ZN(n20361) );
  AOI211_X1 U22377 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20355), .A(n20371), .B(
        n20486), .ZN(n20360) );
  AOI211_X1 U22378 ( .C1(n20358), .C2(n20357), .A(n11089), .B(n21205), .ZN(
        n20359) );
  AOI211_X1 U22379 ( .C1(n20366), .C2(n20361), .A(n20360), .B(n20359), .ZN(
        n20362) );
  OAI211_X1 U22380 ( .C1(n20365), .C2(n20364), .A(n20363), .B(n20362), .ZN(
        P3_U2649) );
  AOI22_X1 U22381 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20432), .B1(
        n20472), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n20376) );
  NAND2_X1 U22382 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20366), .ZN(n20372) );
  NOR2_X1 U22383 ( .A1(n20367), .A2(n20372), .ZN(n20393) );
  OAI21_X1 U22384 ( .B1(n20393), .B2(n20419), .A(n20490), .ZN(n20387) );
  NOR2_X1 U22385 ( .A1(n11089), .A2(n20458), .ZN(n20368) );
  XNOR2_X1 U22386 ( .A(n20368), .B(n20377), .ZN(n20369) );
  AOI22_X1 U22387 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20387), .B1(n20463), 
        .B2(n20369), .ZN(n20375) );
  NAND2_X1 U22388 ( .A1(n20371), .A2(n20370), .ZN(n20380) );
  OAI211_X1 U22389 ( .C1(n20371), .C2(n20370), .A(n20451), .B(n20380), .ZN(
        n20374) );
  OR3_X1 U22390 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20419), .A3(n20372), .ZN(
        n20373) );
  NAND4_X1 U22391 ( .A1(n20376), .A2(n20375), .A3(n20374), .A4(n20373), .ZN(
        P3_U2648) );
  INV_X1 U22392 ( .A(n20387), .ZN(n20386) );
  AOI22_X1 U22393 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20432), .B1(
        n20472), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n20385) );
  NOR2_X1 U22394 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20419), .ZN(n20383) );
  NOR2_X1 U22395 ( .A1(n20379), .A2(n20378), .ZN(n20390) );
  AOI211_X1 U22396 ( .C1(n20379), .C2(n20378), .A(n20390), .B(n21205), .ZN(
        n20382) );
  AOI211_X1 U22397 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20380), .A(n20398), .B(
        n20486), .ZN(n20381) );
  AOI211_X1 U22398 ( .C1(n20383), .C2(n20393), .A(n20382), .B(n20381), .ZN(
        n20384) );
  OAI211_X1 U22399 ( .C1(n20388), .C2(n20386), .A(n20385), .B(n20384), .ZN(
        P3_U2647) );
  AOI21_X1 U22400 ( .B1(n20404), .B2(n20388), .A(n20387), .ZN(n20401) );
  INV_X1 U22401 ( .A(n20389), .ZN(n20392) );
  NOR2_X1 U22402 ( .A1(n20390), .A2(n20458), .ZN(n20391) );
  NOR2_X1 U22403 ( .A1(n20392), .A2(n20391), .ZN(n20410) );
  AOI211_X1 U22404 ( .C1(n20392), .C2(n20391), .A(n20410), .B(n21205), .ZN(
        n20396) );
  NAND2_X1 U22405 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20393), .ZN(n20402) );
  NOR3_X1 U22406 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20419), .A3(n20402), 
        .ZN(n20395) );
  OAI22_X1 U22407 ( .A1(n11317), .A2(n20484), .B1(n20487), .B2(n20397), .ZN(
        n20394) );
  NOR3_X1 U22408 ( .A1(n20396), .A2(n20395), .A3(n20394), .ZN(n20400) );
  NAND2_X1 U22409 ( .A1(n20398), .A2(n20397), .ZN(n20408) );
  OAI211_X1 U22410 ( .C1(n20398), .C2(n20397), .A(n20451), .B(n20408), .ZN(
        n20399) );
  OAI211_X1 U22411 ( .C1(n20401), .C2(n20403), .A(n20400), .B(n20399), .ZN(
        P3_U2646) );
  NOR2_X1 U22412 ( .A1(n20403), .A2(n20402), .ZN(n20405) );
  NAND2_X1 U22413 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n20405), .ZN(n20418) );
  AND2_X1 U22414 ( .A1(n20404), .A2(n20418), .ZN(n20406) );
  AOI22_X1 U22415 ( .A1(n20472), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n20405), 
        .B2(n20406), .ZN(n20416) );
  NOR2_X1 U22416 ( .A1(n20407), .A2(n20406), .ZN(n20431) );
  INV_X1 U22417 ( .A(n20431), .ZN(n20442) );
  NOR2_X1 U22418 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20408), .ZN(n20427) );
  AOI211_X1 U22419 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20408), .A(n20427), .B(
        n20486), .ZN(n20414) );
  INV_X1 U22420 ( .A(n20409), .ZN(n20412) );
  NOR2_X1 U22421 ( .A1(n20410), .A2(n20458), .ZN(n20411) );
  NOR2_X1 U22422 ( .A1(n20412), .A2(n20411), .ZN(n20420) );
  AOI211_X1 U22423 ( .C1(n20412), .C2(n20411), .A(n20420), .B(n21205), .ZN(
        n20413) );
  AOI211_X1 U22424 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n20442), .A(n20414), 
        .B(n20413), .ZN(n20415) );
  OAI211_X1 U22425 ( .C1(n20417), .C2(n20484), .A(n20416), .B(n20415), .ZN(
        P3_U2645) );
  NOR2_X1 U22426 ( .A1(n20419), .A2(n20418), .ZN(n20460) );
  NOR2_X1 U22427 ( .A1(n20420), .A2(n20458), .ZN(n20421) );
  NOR2_X1 U22428 ( .A1(n20422), .A2(n20421), .ZN(n20434) );
  AOI211_X1 U22429 ( .C1(n20422), .C2(n20421), .A(n20434), .B(n21205), .ZN(
        n20425) );
  OAI22_X1 U22430 ( .A1(n20423), .A2(n20484), .B1(n20487), .B2(n20426), .ZN(
        n20424) );
  AOI211_X1 U22431 ( .C1(n20460), .C2(n20430), .A(n20425), .B(n20424), .ZN(
        n20429) );
  NAND2_X1 U22432 ( .A1(n20427), .A2(n20426), .ZN(n20433) );
  OAI211_X1 U22433 ( .C1(n20427), .C2(n20426), .A(n20451), .B(n20433), .ZN(
        n20428) );
  OAI211_X1 U22434 ( .C1(n20431), .C2(n20430), .A(n20429), .B(n20428), .ZN(
        P3_U2644) );
  AOI22_X1 U22435 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20432), .B1(
        n20472), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20441) );
  NOR2_X1 U22436 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20433), .ZN(n20454) );
  AOI211_X1 U22437 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20433), .A(n20454), .B(
        n20486), .ZN(n20438) );
  NOR2_X1 U22438 ( .A1(n20434), .A2(n20458), .ZN(n20435) );
  NOR2_X1 U22439 ( .A1(n20436), .A2(n20435), .ZN(n20444) );
  AOI211_X1 U22440 ( .C1(n20436), .C2(n20435), .A(n20444), .B(n21205), .ZN(
        n20437) );
  AOI211_X1 U22441 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n20442), .A(n20438), 
        .B(n20437), .ZN(n20440) );
  NAND2_X1 U22442 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n20448) );
  OAI211_X1 U22443 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n20460), .B(n20448), .ZN(n20439) );
  NAND3_X1 U22444 ( .A1(n20441), .A2(n20440), .A3(n20439), .ZN(P3_U2643) );
  NOR2_X1 U22445 ( .A1(n20457), .A2(n20448), .ZN(n20461) );
  INV_X1 U22446 ( .A(n20461), .ZN(n20443) );
  AOI21_X1 U22447 ( .B1(n20443), .B2(n20488), .A(n20442), .ZN(n20479) );
  NOR2_X1 U22448 ( .A1(n20444), .A2(n20458), .ZN(n20445) );
  NOR2_X1 U22449 ( .A1(n20446), .A2(n20445), .ZN(n20459) );
  AOI211_X1 U22450 ( .C1(n20446), .C2(n20445), .A(n20459), .B(n21205), .ZN(
        n20450) );
  NAND2_X1 U22451 ( .A1(n20460), .A2(n20457), .ZN(n20447) );
  OAI22_X1 U22452 ( .A1(n11314), .A2(n20484), .B1(n20448), .B2(n20447), .ZN(
        n20449) );
  AOI211_X1 U22453 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n20472), .A(n20450), .B(
        n20449), .ZN(n20456) );
  NAND2_X1 U22454 ( .A1(n20454), .A2(n20453), .ZN(n20465) );
  NAND2_X1 U22455 ( .A1(n20451), .A2(n20465), .ZN(n20468) );
  INV_X1 U22456 ( .A(n20468), .ZN(n20452) );
  OAI21_X1 U22457 ( .B1(n20454), .B2(n20453), .A(n20452), .ZN(n20455) );
  OAI211_X1 U22458 ( .C1(n20479), .C2(n20457), .A(n20456), .B(n20455), .ZN(
        P3_U2642) );
  XOR2_X1 U22459 ( .A(n20475), .B(n20474), .Z(n20464) );
  NAND2_X1 U22460 ( .A1(n20461), .A2(n20460), .ZN(n20469) );
  NOR2_X1 U22461 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20469), .ZN(n20476) );
  OAI22_X1 U22462 ( .A1(n20479), .A2(n20470), .B1(n11315), .B2(n20484), .ZN(
        n20462) );
  AOI211_X1 U22463 ( .C1(n20464), .C2(n20463), .A(n20476), .B(n20462), .ZN(
        n20467) );
  NOR2_X1 U22464 ( .A1(n20486), .A2(n20465), .ZN(n20482) );
  OAI21_X1 U22465 ( .B1(n20472), .B2(n20482), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20466) );
  OAI211_X1 U22466 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n20468), .A(n20467), .B(
        n20466), .ZN(P3_U2641) );
  NOR3_X1 U22467 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20470), .A3(n20469), 
        .ZN(n20471) );
  AOI21_X1 U22468 ( .B1(n20472), .B2(P3_EBX_REG_31__SCAN_IN), .A(n20471), .ZN(
        n20483) );
  INV_X1 U22469 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20481) );
  INV_X1 U22470 ( .A(n20476), .ZN(n20478) );
  AOI21_X1 U22471 ( .B1(n20479), .B2(n20478), .A(n20477), .ZN(n20480) );
  NAND2_X1 U22472 ( .A1(n20487), .A2(n20486), .ZN(n20489) );
  AOI22_X1 U22473 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n20489), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n20488), .ZN(n20492) );
  NAND3_X1 U22474 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20490), .A3(
        n20703), .ZN(n20491) );
  OAI211_X1 U22475 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20493), .A(
        n20492), .B(n20491), .ZN(P3_U2671) );
  NAND2_X1 U22476 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n20504) );
  NOR4_X1 U22477 ( .A1(n20502), .A2(n20501), .A3(n20546), .A4(n20527), .ZN(
        n20503) );
  NOR2_X1 U22478 ( .A1(n20592), .A2(n20657), .ZN(n20656) );
  NAND3_X1 U22479 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n20656), .ZN(n20524) );
  NAND2_X1 U22480 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n20518), .ZN(n20513) );
  NOR2_X1 U22481 ( .A1(n20504), .A2(n20513), .ZN(n20645) );
  INV_X1 U22482 ( .A(n20513), .ZN(n20516) );
  AOI22_X1 U22483 ( .A1(n20516), .A2(P3_EAX_REG_12__SCAN_IN), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n20658), .ZN(n20508) );
  OAI222_X1 U22484 ( .A1(n20676), .A2(n20509), .B1(n20645), .B2(n20508), .C1(
        n20673), .C2(n20507), .ZN(P3_U2722) );
  NAND2_X1 U22485 ( .A1(n20513), .A2(P3_EAX_REG_12__SCAN_IN), .ZN(n20512) );
  AOI22_X1 U22486 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20667), .B1(n20631), .B2(
        n20510), .ZN(n20511) );
  OAI221_X1 U22487 ( .B1(n20513), .B2(P3_EAX_REG_12__SCAN_IN), .C1(n20512), 
        .C2(n20663), .A(n20511), .ZN(P3_U2723) );
  AOI21_X1 U22488 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20658), .A(n20518), .ZN(
        n20515) );
  OAI222_X1 U22489 ( .A1(n20676), .A2(n20517), .B1(n20516), .B2(n20515), .C1(
        n20673), .C2(n20514), .ZN(P3_U2724) );
  AOI211_X1 U22490 ( .C1(n20554), .C2(n20524), .A(n20663), .B(n20518), .ZN(
        n20519) );
  AOI21_X1 U22491 ( .B1(n20631), .B2(n20520), .A(n20519), .ZN(n20521) );
  OAI21_X1 U22492 ( .B1(n20522), .B2(n20676), .A(n20521), .ZN(P3_U2725) );
  AOI22_X1 U22493 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20667), .B1(n20631), .B2(
        n20523), .ZN(n20526) );
  OAI211_X1 U22494 ( .C1(n20556), .C2(P3_EAX_REG_9__SCAN_IN), .A(n20658), .B(
        n20524), .ZN(n20525) );
  NAND2_X1 U22495 ( .A1(n20526), .A2(n20525), .ZN(P3_U2726) );
  NAND3_X1 U22496 ( .A1(n20671), .A2(n20662), .A3(P3_EAX_REG_2__SCAN_IN), .ZN(
        n20547) );
  NAND3_X1 U22497 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(n20539), .ZN(n20530) );
  NOR2_X1 U22498 ( .A1(n20527), .A2(n20530), .ZN(n20533) );
  AOI21_X1 U22499 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20658), .A(n20533), .ZN(
        n20528) );
  OAI222_X1 U22500 ( .A1(n20676), .A2(n20529), .B1(n20656), .B2(n20528), .C1(
        n20673), .C2(n21021), .ZN(P3_U2728) );
  INV_X1 U22501 ( .A(n20530), .ZN(n20537) );
  AOI21_X1 U22502 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20658), .A(n20537), .ZN(
        n20532) );
  OAI222_X1 U22503 ( .A1(n20534), .A2(n20676), .B1(n20533), .B2(n20532), .C1(
        n20673), .C2(n20531), .ZN(P3_U2729) );
  AOI22_X1 U22504 ( .A1(n20539), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n20658), .ZN(n20536) );
  OAI222_X1 U22505 ( .A1(n20538), .A2(n20676), .B1(n20537), .B2(n20536), .C1(
        n20673), .C2(n20535), .ZN(P3_U2730) );
  AND2_X1 U22506 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20539), .ZN(n20542) );
  AOI21_X1 U22507 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20658), .A(n20539), .ZN(
        n20541) );
  OAI222_X1 U22508 ( .A1(n20543), .A2(n20676), .B1(n20542), .B2(n20541), .C1(
        n20673), .C2(n20540), .ZN(P3_U2731) );
  NAND2_X1 U22509 ( .A1(n20658), .A2(n20547), .ZN(n20549) );
  AOI22_X1 U22510 ( .A1(n20667), .A2(BUF2_REG_3__SCAN_IN), .B1(n20631), .B2(
        n20544), .ZN(n20545) );
  OAI221_X1 U22511 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20547), .C1(n20546), 
        .C2(n20549), .A(n20545), .ZN(P3_U2732) );
  NOR2_X1 U22512 ( .A1(n20662), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n20548) );
  OAI222_X1 U22513 ( .A1(n20676), .A2(n20551), .B1(n20673), .B2(n20550), .C1(
        n20549), .C2(n20548), .ZN(P3_U2733) );
  NOR4_X1 U22514 ( .A1(n20554), .A2(n20644), .A3(n20553), .A4(n20552), .ZN(
        n20555) );
  NAND2_X1 U22515 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20586), .ZN(n20582) );
  NAND2_X1 U22516 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20576), .ZN(n20564) );
  NAND2_X1 U22517 ( .A1(n20564), .A2(P3_EAX_REG_21__SCAN_IN), .ZN(n20563) );
  NOR2_X2 U22518 ( .A1(n20557), .A2(n20658), .ZN(n20639) );
  NAND2_X1 U22519 ( .A1(n20558), .A2(n20663), .ZN(n20637) );
  OAI22_X1 U22520 ( .A1(n20560), .A2(n20673), .B1(n20559), .B2(n20637), .ZN(
        n20561) );
  AOI21_X1 U22521 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n20639), .A(n20561), .ZN(
        n20562) );
  OAI221_X1 U22522 ( .B1(n20564), .B2(P3_EAX_REG_21__SCAN_IN), .C1(n20563), 
        .C2(n20663), .A(n20562), .ZN(P3_U2714) );
  AOI22_X1 U22523 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20638), .ZN(n20566) );
  OAI211_X1 U22524 ( .C1(n20576), .C2(P3_EAX_REG_20__SCAN_IN), .A(n20658), .B(
        n20564), .ZN(n20565) );
  OAI211_X1 U22525 ( .C1(n20567), .C2(n20673), .A(n20566), .B(n20565), .ZN(
        P3_U2715) );
  INV_X1 U22526 ( .A(n20633), .ZN(n20572) );
  OAI22_X1 U22527 ( .A1(n20663), .A2(n20570), .B1(n20592), .B2(n20569), .ZN(
        n20571) );
  AOI22_X1 U22528 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20638), .B1(n20572), .B2(
        n20571), .ZN(n20575) );
  AOI22_X1 U22529 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20639), .B1(n20631), .B2(
        n20573), .ZN(n20574) );
  NAND2_X1 U22530 ( .A1(n20575), .A2(n20574), .ZN(P3_U2713) );
  AOI22_X1 U22531 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20638), .ZN(n20580) );
  AOI211_X1 U22532 ( .C1(n20577), .C2(n20582), .A(n20576), .B(n20663), .ZN(
        n20578) );
  INV_X1 U22533 ( .A(n20578), .ZN(n20579) );
  OAI211_X1 U22534 ( .C1(n20581), .C2(n20673), .A(n20580), .B(n20579), .ZN(
        P3_U2716) );
  AOI22_X1 U22535 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20638), .ZN(n20584) );
  OAI211_X1 U22536 ( .C1(n20586), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20658), .B(
        n20582), .ZN(n20583) );
  OAI211_X1 U22537 ( .C1(n20585), .C2(n20673), .A(n20584), .B(n20583), .ZN(
        P3_U2717) );
  AOI22_X1 U22538 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20638), .ZN(n20589) );
  INV_X1 U22539 ( .A(n20586), .ZN(n20587) );
  OAI211_X1 U22540 ( .C1(n11281), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20658), .B(
        n20587), .ZN(n20588) );
  OAI211_X1 U22541 ( .C1(n20590), .C2(n20673), .A(n20589), .B(n20588), .ZN(
        P3_U2718) );
  AOI22_X1 U22542 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20639), .B1(n20631), .B2(
        n20591), .ZN(n20595) );
  NAND2_X1 U22543 ( .A1(n20633), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20632) );
  OAI211_X1 U22544 ( .C1(n20593), .C2(P3_EAX_REG_25__SCAN_IN), .A(n20658), .B(
        n11022), .ZN(n20594) );
  OAI211_X1 U22545 ( .C1(n20637), .C2(n20596), .A(n20595), .B(n20594), .ZN(
        P3_U2710) );
  AOI22_X1 U22546 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20638), .ZN(n20600) );
  NOR2_X2 U22547 ( .A1(n11022), .A2(n20597), .ZN(n20621) );
  AOI211_X1 U22548 ( .C1(n20597), .C2(n11022), .A(n20621), .B(n20663), .ZN(
        n20598) );
  INV_X1 U22549 ( .A(n20598), .ZN(n20599) );
  OAI211_X1 U22550 ( .C1(n20601), .C2(n20673), .A(n20600), .B(n20599), .ZN(
        P3_U2709) );
  NAND2_X1 U22551 ( .A1(n20605), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20604) );
  NAND2_X1 U22552 ( .A1(n20604), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n20603) );
  NAND2_X1 U22553 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n20638), .ZN(n20602) );
  OAI221_X1 U22554 ( .B1(n20604), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n20603), 
        .C2(n20663), .A(n20602), .ZN(P3_U2704) );
  AOI22_X1 U22555 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20638), .ZN(n20607) );
  OAI211_X1 U22556 ( .C1(n20605), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20658), .B(
        n20604), .ZN(n20606) );
  OAI211_X1 U22557 ( .C1(n20608), .C2(n20673), .A(n20607), .B(n20606), .ZN(
        P3_U2705) );
  AOI22_X1 U22558 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20639), .B1(n20631), .B2(
        n20609), .ZN(n20612) );
  OAI211_X1 U22559 ( .C1(n11037), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20658), .B(
        n20610), .ZN(n20611) );
  OAI211_X1 U22560 ( .C1(n20637), .C2(n20613), .A(n20612), .B(n20611), .ZN(
        P3_U2706) );
  AOI22_X1 U22561 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20638), .ZN(n20617) );
  AOI211_X1 U22562 ( .C1(n20614), .C2(n20620), .A(n11037), .B(n20663), .ZN(
        n20615) );
  INV_X1 U22563 ( .A(n20615), .ZN(n20616) );
  OAI211_X1 U22564 ( .C1(n20618), .C2(n20673), .A(n20617), .B(n20616), .ZN(
        P3_U2707) );
  INV_X1 U22565 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n20624) );
  AOI22_X1 U22566 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20639), .B1(n20631), .B2(
        n20619), .ZN(n20623) );
  OAI211_X1 U22567 ( .C1(n20621), .C2(P3_EAX_REG_27__SCAN_IN), .A(n20658), .B(
        n20620), .ZN(n20622) );
  OAI211_X1 U22568 ( .C1(n20637), .C2(n20624), .A(n20623), .B(n20622), .ZN(
        P3_U2708) );
  AOI22_X1 U22569 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20638), .ZN(n20628) );
  OAI211_X1 U22570 ( .C1(n20626), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20658), .B(
        n20625), .ZN(n20627) );
  OAI211_X1 U22571 ( .C1(n20629), .C2(n20673), .A(n20628), .B(n20627), .ZN(
        P3_U2711) );
  AOI22_X1 U22572 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20639), .B1(n20631), .B2(
        n20630), .ZN(n20635) );
  OAI211_X1 U22573 ( .C1(n20633), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20658), .B(
        n20632), .ZN(n20634) );
  OAI211_X1 U22574 ( .C1(n20637), .C2(n20636), .A(n20635), .B(n20634), .ZN(
        P3_U2712) );
  AOI22_X1 U22575 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20639), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20638), .ZN(n20642) );
  OAI211_X1 U22576 ( .C1(n20649), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20658), .B(
        n20640), .ZN(n20641) );
  OAI211_X1 U22577 ( .C1(n20643), .C2(n20673), .A(n20642), .B(n20641), .ZN(
        P3_U2719) );
  AOI22_X1 U22578 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20667), .B1(n20645), .B2(
        n20644), .ZN(n20647) );
  NAND3_X1 U22579 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n20658), .A3(n20651), 
        .ZN(n20646) );
  OAI211_X1 U22580 ( .C1(n20648), .C2(n20673), .A(n20647), .B(n20646), .ZN(
        P3_U2721) );
  AOI211_X1 U22581 ( .C1(n20651), .C2(n20650), .A(n20663), .B(n20649), .ZN(
        n20652) );
  AOI21_X1 U22582 ( .B1(n20667), .B2(BUF2_REG_15__SCAN_IN), .A(n20652), .ZN(
        n20653) );
  OAI21_X1 U22583 ( .B1(n20654), .B2(n20673), .A(n20653), .ZN(P3_U2720) );
  AOI22_X1 U22584 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20667), .B1(n20656), .B2(
        n20655), .ZN(n20660) );
  NAND3_X1 U22585 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n20658), .A3(n20657), .ZN(
        n20659) );
  OAI211_X1 U22586 ( .C1(n20661), .C2(n20673), .A(n20660), .B(n20659), .ZN(
        P3_U2727) );
  AOI211_X1 U22587 ( .C1(n20665), .C2(n20664), .A(n20663), .B(n20662), .ZN(
        n20666) );
  AOI21_X1 U22588 ( .B1(n20667), .B2(BUF2_REG_1__SCAN_IN), .A(n20666), .ZN(
        n20668) );
  OAI21_X1 U22589 ( .B1(n20669), .B2(n20673), .A(n20668), .ZN(P3_U2734) );
  AOI21_X1 U22590 ( .B1(n20671), .B2(n20670), .A(P3_EAX_REG_0__SCAN_IN), .ZN(
        n20674) );
  OAI222_X1 U22591 ( .A1(n20677), .A2(n20676), .B1(n20675), .B2(n20674), .C1(
        n20673), .C2(n20672), .ZN(P3_U2735) );
  NOR2_X1 U22592 ( .A1(n20678), .A2(n21068), .ZN(n20682) );
  AOI22_X1 U22593 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21138), .B1(
        n20682), .B2(n20680), .ZN(n21170) );
  INV_X1 U22594 ( .A(n20710), .ZN(n21209) );
  AOI222_X1 U22595 ( .A1(n20862), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21170), 
        .B2(n20728), .C1(n20680), .C2(n21209), .ZN(n20679) );
  AOI22_X1 U22596 ( .A1(n20733), .A2(n20680), .B1(n20679), .B2(n20730), .ZN(
        P3_U3290) );
  NOR3_X1 U22597 ( .A1(n20692), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        n20681), .ZN(n20711) );
  OAI22_X1 U22598 ( .A1(n20682), .A2(n20683), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20711), .ZN(n21168) );
  INV_X1 U22599 ( .A(n20683), .ZN(n20686) );
  AOI22_X1 U22600 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20684), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n20783), .ZN(n20701) );
  NOR2_X1 U22601 ( .A1(n20685), .A2(n20862), .ZN(n20700) );
  AOI222_X1 U22602 ( .A1(n21168), .A2(n20728), .B1(n20686), .B2(n21209), .C1(
        n20701), .C2(n20700), .ZN(n20687) );
  AOI22_X1 U22603 ( .A1(n20733), .A2(n20712), .B1(n20687), .B2(n20730), .ZN(
        P3_U3289) );
  NAND2_X1 U22604 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20713), .ZN(
        n20709) );
  NAND2_X1 U22605 ( .A1(n20712), .A2(n21165), .ZN(n20698) );
  NOR2_X1 U22606 ( .A1(n20712), .A2(n21165), .ZN(n20695) );
  OAI22_X1 U22607 ( .A1(n20691), .A2(n20690), .B1(n20689), .B2(n20688), .ZN(
        n20722) );
  AOI211_X1 U22608 ( .C1(n20712), .C2(n20692), .A(n20717), .B(n20722), .ZN(
        n20694) );
  AOI21_X1 U22609 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21068), .A(
        n20692), .ZN(n20693) );
  OAI222_X1 U22610 ( .A1(n20696), .A2(n20695), .B1(n20709), .B2(n20694), .C1(
        n20693), .C2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U22611 ( .A1(n21184), .A2(n20699), .B1(n20698), .B2(n20697), .ZN(
        n21164) );
  INV_X1 U22612 ( .A(n20700), .ZN(n20702) );
  OAI22_X1 U22613 ( .A1(n21164), .A2(n20703), .B1(n20702), .B2(n20701), .ZN(
        n20707) );
  NAND2_X1 U22614 ( .A1(n20704), .A2(n21209), .ZN(n20705) );
  OAI21_X1 U22615 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20705), .A(
        n20730), .ZN(n20706) );
  OAI22_X1 U22616 ( .A1(n20707), .A2(n20706), .B1(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20730), .ZN(n20708) );
  OAI21_X1 U22617 ( .B1(n20710), .B2(n20709), .A(n20708), .ZN(P3_U3288) );
  OR2_X1 U22618 ( .A1(n20712), .A2(n20711), .ZN(n20726) );
  NOR2_X1 U22619 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20732), .ZN(
        n20718) );
  NAND2_X1 U22620 ( .A1(n21165), .A2(n20713), .ZN(n20715) );
  AOI22_X1 U22621 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20713), .ZN(n20716) );
  AOI22_X1 U22622 ( .A1(n20718), .A2(n20717), .B1(n21184), .B2(n20716), .ZN(
        n20725) );
  AOI22_X1 U22623 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n20720), .B2(n20719), .ZN(
        n20723) );
  OAI211_X1 U22624 ( .C1(n20723), .C2(n20722), .A(n20721), .B(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20724) );
  OAI211_X1 U22625 ( .C1(n20727), .C2(n20726), .A(n20725), .B(n20724), .ZN(
        n21189) );
  AOI22_X1 U22626 ( .A1(n21209), .A2(n20729), .B1(n20728), .B2(n21189), .ZN(
        n20731) );
  AOI22_X1 U22627 ( .A1(n20733), .A2(n20732), .B1(n20731), .B2(n20730), .ZN(
        P3_U3285) );
  NAND2_X1 U22628 ( .A1(n21180), .A2(n20738), .ZN(n20735) );
  OAI22_X1 U22629 ( .A1(n20736), .A2(n20735), .B1(n21183), .B2(n20734), .ZN(
        n20745) );
  INV_X1 U22630 ( .A(n20737), .ZN(n20742) );
  XNOR2_X1 U22631 ( .A(n20738), .B(n20746), .ZN(n20740) );
  OAI21_X1 U22632 ( .B1(n20740), .B2(n20739), .A(n21198), .ZN(n21160) );
  NOR3_X1 U22633 ( .A1(n20742), .A2(n20741), .A3(n21160), .ZN(n20744) );
  AOI211_X1 U22634 ( .C1(n20746), .C2(n20745), .A(n20744), .B(n20743), .ZN(
        n20747) );
  AOI221_X4 U22635 ( .B1(n20748), .B2(n20747), .C1(n21183), .C2(n20747), .A(
        n21218), .ZN(n21136) );
  AOI22_X1 U22636 ( .A1(n21065), .A2(n20750), .B1(n21182), .B2(n20859), .ZN(
        n20874) );
  NAND2_X1 U22637 ( .A1(n21083), .A2(n20752), .ZN(n20753) );
  NOR3_X1 U22638 ( .A1(n20814), .A2(n20795), .A3(n20823), .ZN(n20826) );
  INV_X1 U22639 ( .A(n20826), .ZN(n20751) );
  NAND2_X1 U22640 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20800) );
  NOR2_X1 U22641 ( .A1(n20751), .A2(n20800), .ZN(n20815) );
  NAND2_X1 U22642 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20815), .ZN(
        n20841) );
  NOR2_X1 U22643 ( .A1(n20840), .A2(n20841), .ZN(n21137) );
  NAND2_X1 U22644 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21137), .ZN(
        n20861) );
  NOR2_X1 U22645 ( .A1(n20753), .A2(n20861), .ZN(n20976) );
  AOI21_X1 U22646 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20801) );
  INV_X1 U22647 ( .A(n20801), .ZN(n20786) );
  NAND2_X1 U22648 ( .A1(n20826), .A2(n20786), .ZN(n20816) );
  NOR2_X1 U22649 ( .A1(n20839), .A2(n20816), .ZN(n20843) );
  NAND3_X1 U22650 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n20843), .ZN(n20858) );
  NOR2_X1 U22651 ( .A1(n20755), .A2(n20858), .ZN(n21088) );
  AND2_X1 U22652 ( .A1(n20752), .A2(n21088), .ZN(n20757) );
  NAND2_X1 U22653 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20976), .ZN(
        n21067) );
  INV_X1 U22654 ( .A(n21067), .ZN(n20761) );
  AOI222_X1 U22655 ( .A1(n20893), .A2(n20976), .B1(n20757), .B2(n21184), .C1(
        n21068), .C2(n20761), .ZN(n20988) );
  OAI21_X1 U22656 ( .B1(n20874), .B2(n20753), .A(n20988), .ZN(n20926) );
  NAND2_X1 U22657 ( .A1(n21136), .A2(n20926), .ZN(n21081) );
  INV_X1 U22658 ( .A(n20754), .ZN(n20767) );
  NOR2_X1 U22659 ( .A1(n20755), .A2(n20861), .ZN(n20929) );
  AND2_X1 U22660 ( .A1(n20929), .A2(n20756), .ZN(n20758) );
  OAI22_X1 U22661 ( .A1(n21138), .A2(n20758), .B1(n20757), .B2(n21090), .ZN(
        n21066) );
  NOR2_X1 U22662 ( .A1(n21184), .A2(n20893), .ZN(n21128) );
  OAI22_X1 U22663 ( .A1(n20762), .A2(n21128), .B1(n20759), .B2(n21026), .ZN(
        n20760) );
  AOI211_X1 U22664 ( .C1(n21065), .C2(n21040), .A(n21066), .B(n20760), .ZN(
        n20931) );
  NAND2_X1 U22665 ( .A1(n20762), .A2(n20761), .ZN(n20763) );
  AOI21_X1 U22666 ( .B1(n21068), .B2(n20763), .A(n21092), .ZN(n20765) );
  AOI211_X1 U22667 ( .C1(n20931), .C2(n20765), .A(n21156), .B(n20764), .ZN(
        n20766) );
  AOI21_X1 U22668 ( .B1(n21152), .B2(n20767), .A(n20766), .ZN(n20769) );
  OAI211_X1 U22669 ( .C1(n20770), .C2(n21081), .A(n20769), .B(n20768), .ZN(
        P3_U2841) );
  INV_X1 U22670 ( .A(n20955), .ZN(n21016) );
  AND2_X1 U22671 ( .A1(n21156), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n20772) );
  NOR2_X1 U22672 ( .A1(n21184), .A2(n21068), .ZN(n21076) );
  AOI221_X1 U22673 ( .B1(n21076), .B2(n20862), .C1(n21138), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21092), .ZN(n20771) );
  AOI211_X1 U22674 ( .C1(n21049), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n20772), .B(n20771), .ZN(n20773) );
  OAI221_X1 U22675 ( .B1(n20775), .B2(n21016), .C1(n20774), .C2(n20846), .A(
        n20773), .ZN(P3_U2862) );
  AOI22_X1 U22676 ( .A1(n21156), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n20955), 
        .B2(n20776), .ZN(n20782) );
  AOI211_X1 U22677 ( .C1(n21138), .C2(n20862), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n21111), .ZN(n20780) );
  OR2_X1 U22678 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21076), .ZN(
        n20777) );
  OAI22_X1 U22679 ( .A1(n21179), .A2(n20778), .B1(n20783), .B2(n20777), .ZN(
        n20779) );
  OAI21_X1 U22680 ( .B1(n20780), .B2(n20779), .A(n21136), .ZN(n20781) );
  OAI211_X1 U22681 ( .C1(n21118), .C2(n20783), .A(n20782), .B(n20781), .ZN(
        P3_U2861) );
  AOI21_X1 U22682 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21068), .A(
        n20893), .ZN(n20799) );
  NOR2_X1 U22683 ( .A1(n20783), .A2(n20799), .ZN(n20790) );
  INV_X1 U22684 ( .A(n21085), .ZN(n21141) );
  NAND3_X1 U22685 ( .A1(n21184), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20784) );
  NAND2_X1 U22686 ( .A1(n21068), .A2(n20862), .ZN(n20928) );
  OAI211_X1 U22687 ( .C1(n21141), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20784), .B(n20928), .ZN(n20788) );
  OAI22_X1 U22688 ( .A1(n21090), .A2(n20786), .B1(n21179), .B2(n20785), .ZN(
        n20787) );
  AOI221_X1 U22689 ( .B1(n20790), .B2(n20789), .C1(n20788), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n20787), .ZN(n20794) );
  AOI22_X1 U22690 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21049), .B1(
        n20955), .B2(n20791), .ZN(n20793) );
  OAI211_X1 U22691 ( .C1(n20794), .C2(n21092), .A(n20793), .B(n20792), .ZN(
        P3_U2860) );
  OAI22_X1 U22692 ( .A1(n21129), .A2(n20796), .B1(n20795), .B2(n21118), .ZN(
        n20797) );
  AOI21_X1 U22693 ( .B1(n20955), .B2(n20798), .A(n20797), .ZN(n20804) );
  OAI22_X1 U22694 ( .A1(n20801), .A2(n21090), .B1(n20800), .B2(n20799), .ZN(
        n20825) );
  AOI22_X1 U22695 ( .A1(n21184), .A2(n20801), .B1(n21085), .B2(n20800), .ZN(
        n20802) );
  NAND3_X1 U22696 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20802), .A3(
        n20928), .ZN(n20806) );
  OAI211_X1 U22697 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20825), .A(
        n21136), .B(n20806), .ZN(n20803) );
  OAI211_X1 U22698 ( .C1(n20805), .C2(n20846), .A(n20804), .B(n20803), .ZN(
        P3_U2859) );
  NAND3_X1 U22699 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21059), .A3(
        n20806), .ZN(n20808) );
  NAND3_X1 U22700 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20814), .A3(
        n20825), .ZN(n20807) );
  OAI211_X1 U22701 ( .C1(n20809), .C2(n21179), .A(n20808), .B(n20807), .ZN(
        n20811) );
  AOI22_X1 U22702 ( .A1(n21136), .A2(n20811), .B1(n20955), .B2(n20810), .ZN(
        n20813) );
  OAI211_X1 U22703 ( .C1(n21118), .C2(n20814), .A(n20813), .B(n20812), .ZN(
        P3_U2858) );
  NAND4_X1 U22704 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21136), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A4(n20825), .ZN(n20824) );
  OAI211_X1 U22705 ( .C1(n21141), .C2(n20815), .A(n21136), .B(n20928), .ZN(
        n20817) );
  OAI221_X1 U22706 ( .B1(n20817), .B2(n21184), .C1(n20817), .C2(n20816), .A(
        n21129), .ZN(n20827) );
  NOR2_X1 U22707 ( .A1(n20846), .A2(n20818), .ZN(n20819) );
  AOI211_X1 U22708 ( .C1(n20955), .C2(n20821), .A(n20820), .B(n20819), .ZN(
        n20822) );
  OAI221_X1 U22709 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n20824), .C1(
        n20823), .C2(n20827), .A(n20822), .ZN(P3_U2857) );
  NAND2_X1 U22710 ( .A1(n20826), .A2(n20825), .ZN(n20838) );
  NOR2_X1 U22711 ( .A1(n21092), .A2(n20838), .ZN(n20829) );
  INV_X1 U22712 ( .A(n20827), .ZN(n20828) );
  MUX2_X1 U22713 ( .A(n20829), .B(n20828), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n20830) );
  AOI21_X1 U22714 ( .B1(n20955), .B2(n20831), .A(n20830), .ZN(n20833) );
  NAND2_X1 U22715 ( .A1(n21156), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n20832) );
  OAI211_X1 U22716 ( .C1(n20846), .C2(n20834), .A(n20833), .B(n20832), .ZN(
        P3_U2856) );
  OAI22_X1 U22717 ( .A1(n21129), .A2(n20835), .B1(n20840), .B2(n21118), .ZN(
        n20836) );
  AOI21_X1 U22718 ( .B1(n20955), .B2(n20837), .A(n20836), .ZN(n20845) );
  NOR2_X1 U22719 ( .A1(n20839), .A2(n20838), .ZN(n20867) );
  AOI21_X1 U22720 ( .B1(n21085), .B2(n20841), .A(n20840), .ZN(n20842) );
  OAI211_X1 U22721 ( .C1(n20843), .C2(n21090), .A(n20842), .B(n20928), .ZN(
        n20849) );
  OAI211_X1 U22722 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n20867), .A(
        n21136), .B(n20849), .ZN(n20844) );
  OAI211_X1 U22723 ( .C1(n20847), .C2(n20846), .A(n20845), .B(n20844), .ZN(
        P3_U2855) );
  AOI22_X1 U22724 ( .A1(n21065), .A2(n20857), .B1(n21182), .B2(n20848), .ZN(
        n20853) );
  NAND3_X1 U22725 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21059), .A3(
        n20849), .ZN(n20852) );
  NAND3_X1 U22726 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20867), .A3(
        n20850), .ZN(n20851) );
  NAND3_X1 U22727 ( .A1(n20853), .A2(n20852), .A3(n20851), .ZN(n20854) );
  AOI22_X1 U22728 ( .A1(n21136), .A2(n20854), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21049), .ZN(n20856) );
  OAI211_X1 U22729 ( .C1(n21133), .C2(n20857), .A(n20856), .B(n20855), .ZN(
        P3_U2854) );
  NAND2_X1 U22730 ( .A1(n21184), .A2(n20858), .ZN(n20906) );
  OAI21_X1 U22731 ( .B1(n20859), .B2(n21026), .A(n20906), .ZN(n21144) );
  NAND2_X1 U22732 ( .A1(n20893), .A2(n20861), .ZN(n21126) );
  OAI21_X1 U22733 ( .B1(n20860), .B2(n21090), .A(n21126), .ZN(n20891) );
  AOI211_X1 U22734 ( .C1(n20893), .C2(n20865), .A(n21144), .B(n20891), .ZN(
        n20880) );
  INV_X1 U22735 ( .A(n21065), .ZN(n21044) );
  NAND2_X1 U22736 ( .A1(n21044), .A2(n21026), .ZN(n21094) );
  NOR2_X1 U22737 ( .A1(n20862), .A2(n20861), .ZN(n21140) );
  NAND2_X1 U22738 ( .A1(n21065), .A2(n20863), .ZN(n21135) );
  OAI221_X1 U22739 ( .B1(n21142), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n21142), .C2(n21140), .A(n21135), .ZN(n20864) );
  AOI211_X1 U22740 ( .C1(n20865), .C2(n21094), .A(n21092), .B(n20864), .ZN(
        n21127) );
  OAI211_X1 U22741 ( .C1(n21142), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n20880), .B(n21127), .ZN(n20866) );
  NAND2_X1 U22742 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n20866), .ZN(
        n20872) );
  NAND3_X1 U22743 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n20867), .ZN(n20912) );
  AOI22_X1 U22744 ( .A1(n21152), .A2(n20869), .B1(n21150), .B2(n20868), .ZN(
        n20870) );
  OAI221_X1 U22745 ( .B1(n21156), .B2(n20872), .C1(n21129), .C2(n20871), .A(
        n20870), .ZN(P3_U2851) );
  AOI21_X1 U22746 ( .B1(n20874), .B2(n20912), .A(n20873), .ZN(n20875) );
  INV_X1 U22747 ( .A(n20875), .ZN(n20882) );
  AOI21_X1 U22748 ( .B1(n20876), .B2(n21140), .A(n21142), .ZN(n20888) );
  NAND2_X1 U22749 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20878) );
  AOI22_X1 U22750 ( .A1(n20893), .A2(n20878), .B1(n20877), .B2(n21094), .ZN(
        n20879) );
  NAND3_X1 U22751 ( .A1(n20880), .A2(n20879), .A3(n21135), .ZN(n21121) );
  NOR2_X1 U22752 ( .A1(n20888), .A2(n21121), .ZN(n20881) );
  MUX2_X1 U22753 ( .A(n20882), .B(n20881), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n20886) );
  AOI22_X1 U22754 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21049), .B1(
        n21152), .B2(n20883), .ZN(n20885) );
  OAI211_X1 U22755 ( .C1(n21092), .C2(n20886), .A(n20885), .B(n20884), .ZN(
        P3_U2850) );
  AOI22_X1 U22756 ( .A1(n21156), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n21152), 
        .B2(n20887), .ZN(n20902) );
  NOR2_X1 U22757 ( .A1(n20892), .A2(n20912), .ZN(n20896) );
  AOI21_X1 U22758 ( .B1(n21184), .B2(n20889), .A(n20888), .ZN(n21119) );
  OAI211_X1 U22759 ( .C1(n21076), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n20906), .B(n21119), .ZN(n20890) );
  AOI211_X1 U22760 ( .C1(n20893), .C2(n20892), .A(n20891), .B(n20890), .ZN(
        n20894) );
  INV_X1 U22761 ( .A(n20894), .ZN(n20895) );
  MUX2_X1 U22762 ( .A(n20896), .B(n20895), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n20900) );
  OAI22_X1 U22763 ( .A1(n21044), .A2(n20898), .B1(n21026), .B2(n20897), .ZN(
        n20899) );
  OAI21_X1 U22764 ( .B1(n20900), .B2(n20899), .A(n21136), .ZN(n20901) );
  OAI211_X1 U22765 ( .C1(n21118), .C2(n20903), .A(n20902), .B(n20901), .ZN(
        P3_U2848) );
  AOI21_X1 U22766 ( .B1(n20908), .B2(n21140), .A(n21142), .ZN(n20904) );
  INV_X1 U22767 ( .A(n20904), .ZN(n20905) );
  AND4_X1 U22768 ( .A1(n21126), .A2(n20906), .A3(n20905), .A4(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n20913) );
  NOR2_X1 U22769 ( .A1(n21084), .A2(n21026), .ZN(n20914) );
  OAI21_X1 U22770 ( .B1(n20915), .B2(n21044), .A(n21136), .ZN(n20907) );
  NOR2_X1 U22771 ( .A1(n20914), .A2(n20907), .ZN(n21110) );
  OAI211_X1 U22772 ( .C1(n20908), .C2(n21128), .A(n20913), .B(n21110), .ZN(
        n20909) );
  NAND2_X1 U22773 ( .A1(n21129), .A2(n20909), .ZN(n21108) );
  AOI22_X1 U22774 ( .A1(n21156), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n21152), 
        .B2(n20910), .ZN(n20923) );
  NOR3_X1 U22775 ( .A1(n20913), .A2(n20912), .A3(n20911), .ZN(n20921) );
  INV_X1 U22776 ( .A(n20914), .ZN(n20918) );
  OR2_X1 U22777 ( .A1(n21044), .A2(n20915), .ZN(n20916) );
  OAI22_X1 U22778 ( .A1(n20919), .A2(n20918), .B1(n20917), .B2(n20916), .ZN(
        n20920) );
  OAI21_X1 U22779 ( .B1(n20921), .B2(n20920), .A(n21136), .ZN(n20922) );
  OAI211_X1 U22780 ( .C1(n20924), .C2(n21108), .A(n20923), .B(n20922), .ZN(
        P3_U2847) );
  AOI22_X1 U22781 ( .A1(n21156), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n21152), 
        .B2(n20925), .ZN(n20935) );
  NAND2_X1 U22782 ( .A1(n20927), .A2(n20926), .ZN(n21055) );
  INV_X1 U22783 ( .A(n21055), .ZN(n20933) );
  NAND2_X1 U22784 ( .A1(n20929), .A2(n20928), .ZN(n21086) );
  NOR2_X1 U22785 ( .A1(n20938), .A2(n21086), .ZN(n20979) );
  INV_X1 U22786 ( .A(n20979), .ZN(n20965) );
  NAND2_X1 U22787 ( .A1(n21068), .A2(n20965), .ZN(n20930) );
  OAI211_X1 U22788 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n21128), .A(
        n20931), .B(n20930), .ZN(n20932) );
  OAI221_X1 U22789 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n20933), 
        .C1(n21048), .C2(n20932), .A(n21136), .ZN(n20934) );
  OAI211_X1 U22790 ( .C1(n21118), .C2(n21048), .A(n20935), .B(n20934), .ZN(
        P3_U2840) );
  NOR2_X1 U22791 ( .A1(n20988), .A2(n20987), .ZN(n20943) );
  AND2_X1 U22792 ( .A1(n20937), .A2(n20936), .ZN(n20942) );
  INV_X1 U22793 ( .A(n20938), .ZN(n20939) );
  AOI21_X1 U22794 ( .B1(n21088), .B2(n20939), .A(n21090), .ZN(n21046) );
  NAND2_X1 U22795 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20940) );
  NOR2_X1 U22796 ( .A1(n21141), .A2(n20979), .ZN(n21022) );
  NOR3_X1 U22797 ( .A1(n21046), .A2(n20940), .A3(n21022), .ZN(n20941) );
  NOR2_X1 U22798 ( .A1(n20941), .A2(n21111), .ZN(n20958) );
  AOI222_X1 U22799 ( .A1(n20944), .A2(n21065), .B1(n20943), .B2(n20942), .C1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n20958), .ZN(n20951) );
  INV_X1 U22800 ( .A(n20945), .ZN(n20946) );
  OAI22_X1 U22801 ( .A1(n20947), .A2(n21016), .B1(n21133), .B2(n20946), .ZN(
        n20948) );
  AOI211_X1 U22802 ( .C1(n21049), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n20949), .B(n20948), .ZN(n20950) );
  OAI21_X1 U22803 ( .B1(n20951), .B2(n21092), .A(n20950), .ZN(P3_U2837) );
  INV_X1 U22804 ( .A(n20952), .ZN(n20964) );
  NAND2_X1 U22805 ( .A1(n21156), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n20963) );
  NOR2_X1 U22806 ( .A1(n21055), .A2(n20953), .ZN(n20969) );
  NAND2_X1 U22807 ( .A1(n20955), .A2(n20954), .ZN(n20970) );
  NAND2_X1 U22808 ( .A1(n21065), .A2(n20956), .ZN(n20966) );
  OAI211_X1 U22809 ( .C1(n21111), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n20966), .ZN(n20957) );
  OAI21_X1 U22810 ( .B1(n20958), .B2(n20957), .A(n21136), .ZN(n20959) );
  OAI211_X1 U22811 ( .C1(n21118), .C2(n20960), .A(n20970), .B(n20959), .ZN(
        n20961) );
  OAI21_X1 U22812 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n20969), .A(
        n20961), .ZN(n20962) );
  OAI211_X1 U22813 ( .C1(n20964), .C2(n21133), .A(n20963), .B(n20962), .ZN(
        P3_U2836) );
  NAND4_X1 U22814 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20978) );
  AOI21_X1 U22815 ( .B1(n21184), .B2(n20978), .A(n21046), .ZN(n21023) );
  OAI21_X1 U22816 ( .B1(n20965), .B2(n20978), .A(n21085), .ZN(n20967) );
  NAND4_X1 U22817 ( .A1(n21023), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n20967), .A4(n20966), .ZN(n20968) );
  AOI22_X1 U22818 ( .A1(n21136), .A2(n20968), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21049), .ZN(n20971) );
  NAND2_X1 U22819 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n20969), .ZN(
        n21032) );
  AOI22_X1 U22820 ( .A1(n20971), .A2(n20970), .B1(n21032), .B2(n21031), .ZN(
        n20972) );
  AOI21_X1 U22821 ( .B1(n21152), .B2(n20973), .A(n20972), .ZN(n20975) );
  NAND2_X1 U22822 ( .A1(n20975), .A2(n20974), .ZN(P3_U2835) );
  NOR2_X1 U22823 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21090), .ZN(
        n21030) );
  INV_X1 U22824 ( .A(n20976), .ZN(n20977) );
  NOR3_X1 U22825 ( .A1(n20977), .A2(n20987), .A3(n20986), .ZN(n20982) );
  NOR2_X1 U22826 ( .A1(n21031), .A2(n20978), .ZN(n21024) );
  AOI21_X1 U22827 ( .B1(n20979), .B2(n21024), .A(n21142), .ZN(n20980) );
  INV_X1 U22828 ( .A(n20980), .ZN(n20981) );
  OAI211_X1 U22829 ( .C1(n21138), .C2(n20982), .A(n21023), .B(n20981), .ZN(
        n20994) );
  AOI22_X1 U22830 ( .A1(n21156), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n20985), 
        .B2(n21129), .ZN(n20992) );
  INV_X1 U22831 ( .A(n21027), .ZN(n20990) );
  NOR3_X1 U22832 ( .A1(n20988), .A2(n20987), .A3(n20986), .ZN(n21006) );
  AOI21_X1 U22833 ( .B1(n21025), .B2(n21065), .A(n21006), .ZN(n20989) );
  OAI21_X1 U22834 ( .B1(n21026), .B2(n20990), .A(n20989), .ZN(n20996) );
  NAND3_X1 U22835 ( .A1(n21136), .A2(n21004), .A3(n20996), .ZN(n20991) );
  OAI211_X1 U22836 ( .C1(n20993), .C2(n21133), .A(n20992), .B(n20991), .ZN(
        P3_U2833) );
  AOI211_X1 U22837 ( .C1(n21059), .C2(n20995), .A(n21005), .B(n20994), .ZN(
        n21011) );
  AOI21_X1 U22838 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n20996), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n20997) );
  AOI21_X1 U22839 ( .B1(n20998), .B2(n21011), .A(n20997), .ZN(n20999) );
  AOI22_X1 U22840 ( .A1(n21136), .A2(n20999), .B1(n21049), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21001) );
  OAI211_X1 U22841 ( .C1(n21002), .C2(n21133), .A(n21001), .B(n21000), .ZN(
        P3_U2832) );
  AOI21_X1 U22842 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21049), .A(
        n21003), .ZN(n21015) );
  NAND2_X1 U22843 ( .A1(n21059), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n21010) );
  NOR3_X1 U22844 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21005), .A3(
        n21004), .ZN(n21007) );
  AOI22_X1 U22845 ( .A1(n21065), .A2(n21008), .B1(n21007), .B2(n21006), .ZN(
        n21009) );
  OAI21_X1 U22846 ( .B1(n21011), .B2(n21010), .A(n21009), .ZN(n21013) );
  AOI22_X1 U22847 ( .A1(n21136), .A2(n21013), .B1(n21152), .B2(n21012), .ZN(
        n21014) );
  OAI211_X1 U22848 ( .C1(n21017), .C2(n21016), .A(n21015), .B(n21014), .ZN(
        P3_U2831) );
  NOR2_X1 U22849 ( .A1(n21049), .A2(n21022), .ZN(n21043) );
  OAI211_X1 U22850 ( .C1(n21141), .C2(n21024), .A(n21043), .B(n21023), .ZN(
        n21029) );
  OAI22_X1 U22851 ( .A1(n21027), .A2(n21026), .B1(n21025), .B2(n21044), .ZN(
        n21028) );
  OAI22_X1 U22852 ( .A1(n21034), .A2(n21033), .B1(n21032), .B2(n21031), .ZN(
        n21035) );
  OAI221_X1 U22853 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21136), 
        .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21035), .A(n21129), .ZN(
        n21039) );
  NOR2_X1 U22854 ( .A1(n21054), .A2(n21040), .ZN(n21045) );
  OAI21_X1 U22855 ( .B1(n21054), .B2(n21041), .A(n21182), .ZN(n21042) );
  OAI211_X1 U22856 ( .C1(n21045), .C2(n21044), .A(n21043), .B(n21042), .ZN(
        n21058) );
  NOR2_X1 U22857 ( .A1(n21058), .A2(n21046), .ZN(n21047) );
  AOI21_X1 U22858 ( .B1(n21047), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n21156), .ZN(n21057) );
  NOR3_X1 U22859 ( .A1(n21049), .A2(n21048), .A3(n21055), .ZN(n21051) );
  AOI221_X1 U22860 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21057), 
        .C1(n21051), .C2(n21057), .A(n21050), .ZN(n21052) );
  OAI21_X1 U22861 ( .B1(n21133), .B2(n21053), .A(n21052), .ZN(P3_U2839) );
  NOR4_X1 U22862 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21055), .A3(
        n21092), .A4(n21054), .ZN(n21056) );
  AOI21_X1 U22863 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21156), .A(n21056), 
        .ZN(n21061) );
  OAI211_X1 U22864 ( .C1(n21059), .C2(n21058), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21057), .ZN(n21060) );
  OAI211_X1 U22865 ( .C1(n21062), .C2(n21133), .A(n21061), .B(n21060), .ZN(
        P3_U2838) );
  AOI22_X1 U22866 ( .A1(n21065), .A2(n21064), .B1(n21182), .B2(n21063), .ZN(
        n21070) );
  AOI211_X1 U22867 ( .C1(n21068), .C2(n21067), .A(n21092), .B(n21066), .ZN(
        n21069) );
  AOI21_X1 U22868 ( .B1(n21070), .B2(n21069), .A(n21156), .ZN(n21078) );
  AOI22_X1 U22869 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21078), .B1(
        n21152), .B2(n21071), .ZN(n21073) );
  OAI211_X1 U22870 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21081), .A(
        n21073), .B(n21072), .ZN(P3_U2843) );
  AOI22_X1 U22871 ( .A1(n21156), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n21152), 
        .B2(n21074), .ZN(n21080) );
  NOR3_X1 U22872 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21076), .A3(
        n21075), .ZN(n21077) );
  OAI21_X1 U22873 ( .B1(n21078), .B2(n21077), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21079) );
  OAI211_X1 U22874 ( .C1(n21082), .C2(n21081), .A(n21080), .B(n21079), .ZN(
        P3_U2842) );
  NAND2_X1 U22875 ( .A1(n21083), .A2(n21150), .ZN(n21116) );
  NAND3_X1 U22876 ( .A1(n21084), .A2(n21089), .A3(n21135), .ZN(n21093) );
  OAI21_X1 U22877 ( .B1(n21109), .B2(n21086), .A(n21085), .ZN(n21087) );
  OAI221_X1 U22878 ( .B1(n21090), .B2(n21089), .C1(n21090), .C2(n21088), .A(
        n21087), .ZN(n21091) );
  AOI211_X1 U22879 ( .C1(n21094), .C2(n21093), .A(n21092), .B(n21091), .ZN(
        n21102) );
  AOI221_X1 U22880 ( .B1(n21141), .B2(n21102), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n21102), .A(n21095), .ZN(
        n21096) );
  AOI22_X1 U22881 ( .A1(n21097), .A2(n21152), .B1(n21096), .B2(n21129), .ZN(
        n21099) );
  OAI211_X1 U22882 ( .C1(n21116), .C2(n21100), .A(n21099), .B(n21098), .ZN(
        P3_U2844) );
  NOR3_X1 U22883 ( .A1(n21156), .A2(n21102), .A3(n21101), .ZN(n21104) );
  NOR3_X1 U22884 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21109), .A3(
        n21116), .ZN(n21103) );
  AOI211_X1 U22885 ( .C1(n21152), .C2(n21105), .A(n21104), .B(n21103), .ZN(
        n21106) );
  OAI21_X1 U22886 ( .B1(n21129), .B2(n21107), .A(n21106), .ZN(P3_U2845) );
  AOI211_X1 U22887 ( .C1(n21111), .C2(n21110), .A(n21109), .B(n21108), .ZN(
        n21112) );
  AOI211_X1 U22888 ( .C1(n21152), .C2(n21114), .A(n21113), .B(n21112), .ZN(
        n21115) );
  OAI21_X1 U22889 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21116), .A(
        n21115), .ZN(P3_U2846) );
  AOI22_X1 U22890 ( .A1(n21156), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21150), 
        .B2(n21117), .ZN(n21123) );
  NAND2_X1 U22891 ( .A1(n21119), .A2(n21118), .ZN(n21120) );
  OAI211_X1 U22892 ( .C1(n21121), .C2(n21120), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21129), .ZN(n21122) );
  OAI211_X1 U22893 ( .C1(n21124), .C2(n21133), .A(n21123), .B(n21122), .ZN(
        P3_U2849) );
  NOR2_X1 U22894 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21149), .ZN(
        n21125) );
  AOI22_X1 U22895 ( .A1(n21156), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21150), 
        .B2(n21125), .ZN(n21132) );
  OAI211_X1 U22896 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21128), .A(
        n21127), .B(n21126), .ZN(n21130) );
  OAI211_X1 U22897 ( .C1(n21144), .C2(n21130), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21129), .ZN(n21131) );
  OAI211_X1 U22898 ( .C1(n21134), .C2(n21133), .A(n21132), .B(n21131), .ZN(
        P3_U2852) );
  OAI211_X1 U22899 ( .C1(n21138), .C2(n21137), .A(n21136), .B(n21135), .ZN(
        n21139) );
  INV_X1 U22900 ( .A(n21139), .ZN(n21147) );
  AOI211_X1 U22901 ( .C1(n21142), .C2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n21141), .B(n21140), .ZN(n21143) );
  INV_X1 U22902 ( .A(n21143), .ZN(n21146) );
  INV_X1 U22903 ( .A(n21144), .ZN(n21145) );
  NAND3_X1 U22904 ( .A1(n21147), .A2(n21146), .A3(n21145), .ZN(n21148) );
  NAND2_X1 U22905 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21148), .ZN(
        n21155) );
  AOI22_X1 U22906 ( .A1(n21152), .A2(n21151), .B1(n21150), .B2(n21149), .ZN(
        n21153) );
  OAI221_X1 U22907 ( .B1(n21156), .B2(n21155), .C1(n21129), .C2(n21154), .A(
        n21153), .ZN(P3_U2853) );
  NAND2_X1 U22908 ( .A1(n21628), .A2(n18302), .ZN(n21204) );
  INV_X1 U22909 ( .A(n21157), .ZN(n21203) );
  NOR2_X1 U22910 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .ZN(
        n21163) );
  INV_X1 U22911 ( .A(n21158), .ZN(n21159) );
  NAND3_X1 U22912 ( .A1(n21178), .A2(n21160), .A3(n21159), .ZN(n21220) );
  OAI211_X1 U22913 ( .C1(n21163), .C2(n21220), .A(n21162), .B(n21161), .ZN(
        n21194) );
  INV_X1 U22914 ( .A(n21195), .ZN(n21188) );
  AOI22_X1 U22915 ( .A1(n21195), .A2(n21165), .B1(n21164), .B2(n21188), .ZN(
        n21185) );
  OR3_X1 U22916 ( .A1(n21170), .A2(n21169), .A3(n21166), .ZN(n21167) );
  AOI22_X1 U22917 ( .A1(n21170), .A2(n21169), .B1(n21168), .B2(n21167), .ZN(
        n21172) );
  OAI21_X1 U22918 ( .B1(n21195), .B2(n21172), .A(n21171), .ZN(n21173) );
  AOI222_X1 U22919 ( .A1(n21185), .A2(n21174), .B1(n21185), .B2(n21173), .C1(
        n21174), .C2(n21173), .ZN(n21192) );
  NAND2_X1 U22920 ( .A1(n21176), .A2(n21175), .ZN(n21191) );
  OAI22_X1 U22921 ( .A1(n21180), .A2(n21179), .B1(n21178), .B2(n21177), .ZN(
        n21181) );
  AOI221_X1 U22922 ( .B1(n21184), .B2(n21183), .C1(n21182), .C2(n21183), .A(
        n21181), .ZN(n21223) );
  INV_X1 U22923 ( .A(n21185), .ZN(n21186) );
  OAI221_X1 U22924 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n21192), .A(n21186), .ZN(
        n21187) );
  OAI221_X1 U22925 ( .B1(n21195), .B2(n21189), .C1(n21188), .C2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n21187), .ZN(n21190) );
  OAI211_X1 U22926 ( .C1(n21192), .C2(n21191), .A(n21223), .B(n21190), .ZN(
        n21193) );
  AOI211_X1 U22927 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21195), .A(
        n21194), .B(n21193), .ZN(n21219) );
  OAI211_X1 U22928 ( .C1(n21197), .C2(n21196), .A(n21221), .B(n21219), .ZN(
        n21207) );
  OAI21_X1 U22929 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n21198), .A(n21207), 
        .ZN(n21212) );
  INV_X1 U22930 ( .A(n21212), .ZN(n21200) );
  NAND3_X1 U22931 ( .A1(n21201), .A2(n21200), .A3(n21199), .ZN(n21202) );
  NAND4_X1 U22932 ( .A1(n21205), .A2(n21204), .A3(n21203), .A4(n21202), .ZN(
        P3_U2997) );
  OAI221_X1 U22933 ( .B1(n21208), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21208), 
        .C2(n21207), .A(n21206), .ZN(P3_U3282) );
  AOI22_X1 U22934 ( .A1(n21210), .A2(n21209), .B1(n21628), .B2(n18302), .ZN(
        n21211) );
  INV_X1 U22935 ( .A(n21211), .ZN(n21215) );
  NOR2_X1 U22936 ( .A1(n21213), .A2(n21212), .ZN(n21214) );
  MUX2_X1 U22937 ( .A(n21215), .B(n21214), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21217) );
  OAI211_X1 U22938 ( .C1(n21219), .C2(n21218), .A(n21217), .B(n21216), .ZN(
        P3_U2996) );
  NAND2_X1 U22939 ( .A1(n21221), .A2(n21220), .ZN(n21225) );
  NAND2_X1 U22940 ( .A1(n21225), .A2(P3_MORE_REG_SCAN_IN), .ZN(n21222) );
  OAI21_X1 U22941 ( .B1(n21225), .B2(n21223), .A(n21222), .ZN(P3_U3295) );
  AOI21_X1 U22942 ( .B1(n21225), .B2(P3_FLUSH_REG_SCAN_IN), .A(n21224), .ZN(
        n21226) );
  INV_X1 U22943 ( .A(n21226), .ZN(P3_U2637) );
  AOI211_X1 U22944 ( .C1(n21230), .C2(n21229), .A(n21228), .B(n21227), .ZN(
        n21236) );
  OAI211_X1 U22945 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21232), .A(n21231), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21233) );
  AOI21_X1 U22946 ( .B1(n21233), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21556), 
        .ZN(n21235) );
  NAND2_X1 U22947 ( .A1(n21236), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21234) );
  OAI21_X1 U22948 ( .B1(n21236), .B2(n21235), .A(n21234), .ZN(P1_U3485) );
  NAND2_X1 U22949 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21240), .ZN(
        n21243) );
  INV_X1 U22950 ( .A(n21245), .ZN(n21237) );
  OAI22_X1 U22951 ( .A1(n21238), .A2(n21243), .B1(n21367), .B2(n21237), .ZN(
        n21330) );
  OAI221_X1 U22952 ( .B1(n21330), .B2(n21415), .C1(n21330), .C2(n21240), .A(
        n21254), .ZN(n21251) );
  INV_X1 U22953 ( .A(n21238), .ZN(n21413) );
  AOI21_X1 U22954 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21240), .A(
        n21239), .ZN(n21241) );
  AOI211_X1 U22955 ( .C1(n21413), .C2(n21243), .A(n21242), .B(n21241), .ZN(
        n21244) );
  OAI21_X1 U22956 ( .B1(n21245), .B2(n21367), .A(n21244), .ZN(n21252) );
  AOI22_X1 U22957 ( .A1(n21246), .A2(n21411), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21252), .ZN(n21250) );
  NAND2_X1 U22958 ( .A1(n21390), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n21249) );
  NAND2_X1 U22959 ( .A1(n21409), .A2(n21247), .ZN(n21248) );
  NAND4_X1 U22960 ( .A1(n21251), .A2(n21250), .A3(n21249), .A4(n21248), .ZN(
        P1_U3018) );
  AOI21_X1 U22961 ( .B1(n21254), .B2(n21330), .A(n21252), .ZN(n21262) );
  AOI22_X1 U22962 ( .A1(n21308), .A2(n21310), .B1(n21325), .B2(n21253), .ZN(
        n21319) );
  NOR4_X1 U22963 ( .A1(n21319), .A2(n21255), .A3(n21254), .A4(n21309), .ZN(
        n21258) );
  OAI22_X1 U22964 ( .A1(n21256), .A2(n21335), .B1(n21389), .B2(n21464), .ZN(
        n21257) );
  AOI21_X1 U22965 ( .B1(n21258), .B2(n21261), .A(n21257), .ZN(n21260) );
  NAND2_X1 U22966 ( .A1(n21390), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21259) );
  OAI211_X1 U22967 ( .C1(n21262), .C2(n21261), .A(n21260), .B(n21259), .ZN(
        P1_U3017) );
  NOR2_X1 U22968 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21263), .ZN(
        n21269) );
  INV_X1 U22969 ( .A(n21264), .ZN(n21267) );
  OAI22_X1 U22970 ( .A1(n21267), .A2(n21335), .B1(n21266), .B2(n21265), .ZN(
        n21268) );
  AOI21_X1 U22971 ( .B1(n21269), .B2(n21282), .A(n21268), .ZN(n21271) );
  OAI211_X1 U22972 ( .C1(n21389), .C2(n21272), .A(n21271), .B(n21270), .ZN(
        P1_U3026) );
  INV_X1 U22973 ( .A(n21273), .ZN(n21433) );
  INV_X1 U22974 ( .A(n21274), .ZN(n21281) );
  INV_X1 U22975 ( .A(n21275), .ZN(n21279) );
  OAI211_X1 U22976 ( .C1(n21277), .C2(n21328), .A(n21283), .B(n21276), .ZN(
        n21278) );
  AOI21_X1 U22977 ( .B1(n21278), .B2(n21337), .A(n21414), .ZN(n21289) );
  OAI22_X1 U22978 ( .A1(n21279), .A2(n21335), .B1(n13546), .B2(n21289), .ZN(
        n21280) );
  AOI211_X1 U22979 ( .C1(n21409), .C2(n21433), .A(n21281), .B(n21280), .ZN(
        n21284) );
  NAND3_X1 U22980 ( .A1(n21283), .A2(n13546), .A3(n21282), .ZN(n21288) );
  NAND2_X1 U22981 ( .A1(n21284), .A2(n21288), .ZN(P1_U3024) );
  INV_X1 U22982 ( .A(n21285), .ZN(n21292) );
  NOR3_X1 U22983 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21287), .A3(
        n21286), .ZN(n21291) );
  AOI21_X1 U22984 ( .B1(n21289), .B2(n21288), .A(n14484), .ZN(n21290) );
  AOI211_X1 U22985 ( .C1(n21292), .C2(n21411), .A(n21291), .B(n21290), .ZN(
        n21294) );
  NAND2_X1 U22986 ( .A1(n21390), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21293) );
  OAI211_X1 U22987 ( .C1(n21389), .C2(n21295), .A(n21294), .B(n21293), .ZN(
        P1_U3023) );
  OAI22_X1 U22988 ( .A1(n21401), .A2(n21297), .B1(n21389), .B2(n21296), .ZN(
        n21298) );
  AOI21_X1 U22989 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n21299), .A(
        n21298), .ZN(n21303) );
  OAI211_X1 U22990 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n21301), .B(n21300), .ZN(
        n21302) );
  OAI211_X1 U22991 ( .C1(n21304), .C2(n21335), .A(n21303), .B(n21302), .ZN(
        P1_U3021) );
  NOR2_X1 U22992 ( .A1(n21401), .A2(n21305), .ZN(n21315) );
  NOR2_X1 U22993 ( .A1(n21319), .A2(n21309), .ZN(n21313) );
  NAND2_X1 U22994 ( .A1(n21325), .A2(n21306), .ZN(n21307) );
  OAI211_X1 U22995 ( .C1(n21308), .C2(n21328), .A(n21327), .B(n21307), .ZN(
        n21321) );
  AOI21_X1 U22996 ( .B1(n21310), .B2(n21309), .A(n21321), .ZN(n21311) );
  INV_X1 U22997 ( .A(n21311), .ZN(n21312) );
  MUX2_X1 U22998 ( .A(n21313), .B(n21312), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n21314) );
  AOI211_X1 U22999 ( .C1(n21409), .C2(n21452), .A(n21315), .B(n21314), .ZN(
        n21316) );
  OAI21_X1 U23000 ( .B1(n21317), .B2(n21335), .A(n21316), .ZN(P1_U3019) );
  OAI22_X1 U23001 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21319), .B1(
        n21318), .B2(n21335), .ZN(n21320) );
  AOI21_X1 U23002 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21321), .A(
        n21320), .ZN(n21323) );
  OAI211_X1 U23003 ( .C1(n21389), .C2(n21445), .A(n21323), .B(n21322), .ZN(
        P1_U3020) );
  NAND2_X1 U23004 ( .A1(n21325), .A2(n21324), .ZN(n21326) );
  OAI211_X1 U23005 ( .C1(n21329), .C2(n21328), .A(n21327), .B(n21326), .ZN(
        n21353) );
  AOI22_X1 U23006 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21353), .B1(
        n21390), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n21334) );
  NAND2_X1 U23007 ( .A1(n21331), .A2(n21330), .ZN(n21358) );
  NAND2_X1 U23008 ( .A1(n21332), .A2(n21358), .ZN(n21351) );
  AOI22_X1 U23009 ( .A1(n21479), .A2(n21409), .B1(n13569), .B2(n21351), .ZN(
        n21333) );
  OAI211_X1 U23010 ( .C1(n21336), .C2(n21335), .A(n21334), .B(n21333), .ZN(
        P1_U3016) );
  NAND2_X1 U23011 ( .A1(n15558), .A2(n21351), .ZN(n21342) );
  AOI21_X1 U23012 ( .B1(n21343), .B2(n21337), .A(n21353), .ZN(n21349) );
  OAI22_X1 U23013 ( .A1(n21349), .A2(n15558), .B1(n21389), .B2(n21504), .ZN(
        n21338) );
  AOI21_X1 U23014 ( .B1(n21339), .B2(n21411), .A(n21338), .ZN(n21341) );
  NAND2_X1 U23015 ( .A1(n21390), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n21340) );
  OAI211_X1 U23016 ( .C1(n21343), .C2(n21342), .A(n21341), .B(n21340), .ZN(
        P1_U3013) );
  NOR2_X1 U23017 ( .A1(n13569), .A2(n15552), .ZN(n21350) );
  AOI21_X1 U23018 ( .B1(n21350), .B2(n21351), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21348) );
  AOI22_X1 U23019 ( .A1(n21409), .A2(n21345), .B1(n21411), .B2(n21344), .ZN(
        n21347) );
  NAND2_X1 U23020 ( .A1(n21390), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n21346) );
  OAI211_X1 U23021 ( .C1(n21349), .C2(n21348), .A(n21347), .B(n21346), .ZN(
        P1_U3014) );
  AOI21_X1 U23022 ( .B1(n13569), .B2(n15552), .A(n21350), .ZN(n21352) );
  AOI22_X1 U23023 ( .A1(n21390), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n21352), 
        .B2(n21351), .ZN(n21356) );
  AOI22_X1 U23024 ( .A1(n21354), .A2(n21411), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21353), .ZN(n21355) );
  OAI211_X1 U23025 ( .C1(n21389), .C2(n21357), .A(n21356), .B(n21355), .ZN(
        P1_U3015) );
  NOR2_X1 U23026 ( .A1(n21359), .A2(n21358), .ZN(n21363) );
  NOR2_X1 U23027 ( .A1(n21360), .A2(n21363), .ZN(n21382) );
  NOR3_X1 U23028 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21382), .A3(
        n21361), .ZN(n21362) );
  AOI21_X1 U23029 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n21390), .A(n21362), 
        .ZN(n21372) );
  NOR2_X1 U23030 ( .A1(n21415), .A2(n21363), .ZN(n21368) );
  INV_X1 U23031 ( .A(n21364), .ZN(n21365) );
  OAI21_X1 U23032 ( .B1(n21367), .B2(n21366), .A(n21365), .ZN(n21373) );
  INV_X1 U23033 ( .A(n21373), .ZN(n21384) );
  OAI21_X1 U23034 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21368), .A(
        n21384), .ZN(n21370) );
  AOI22_X1 U23035 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21370), .B1(
        n21411), .B2(n21369), .ZN(n21371) );
  OAI211_X1 U23036 ( .C1(n21389), .C2(n21516), .A(n21372), .B(n21371), .ZN(
        P1_U3011) );
  AOI22_X1 U23037 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21373), .B1(
        n21390), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n21377) );
  AOI22_X1 U23038 ( .A1(n21409), .A2(n21375), .B1(n21411), .B2(n21374), .ZN(
        n21376) );
  OAI211_X1 U23039 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21382), .A(
        n21377), .B(n21376), .ZN(P1_U3012) );
  NOR2_X1 U23040 ( .A1(n21401), .A2(n21523), .ZN(n21380) );
  NOR3_X1 U23041 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21382), .A3(
        n21378), .ZN(n21379) );
  AOI211_X1 U23042 ( .C1(n21381), .C2(n21411), .A(n21380), .B(n21379), .ZN(
        n21388) );
  NAND2_X1 U23043 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21383) );
  NOR3_X1 U23044 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21382), .A3(
        n21383), .ZN(n21391) );
  INV_X1 U23045 ( .A(n21383), .ZN(n21386) );
  OAI21_X1 U23046 ( .B1(n21386), .B2(n21385), .A(n21384), .ZN(n21396) );
  OAI21_X1 U23047 ( .B1(n21391), .B2(n21396), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21387) );
  OAI211_X1 U23048 ( .C1(n21389), .C2(n21528), .A(n21388), .B(n21387), .ZN(
        P1_U3009) );
  AND2_X1 U23049 ( .A1(n21390), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n21392) );
  AOI211_X1 U23050 ( .C1(n21411), .C2(n21393), .A(n21392), .B(n21391), .ZN(
        n21398) );
  INV_X1 U23051 ( .A(n21394), .ZN(n21395) );
  AOI22_X1 U23052 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21396), .B1(
        n21409), .B2(n21395), .ZN(n21397) );
  NAND2_X1 U23053 ( .A1(n21398), .A2(n21397), .ZN(P1_U3010) );
  AOI22_X1 U23054 ( .A1(n21400), .A2(n21411), .B1(n21409), .B2(n21399), .ZN(
        n21407) );
  NOR2_X1 U23055 ( .A1(n21401), .A2(n21534), .ZN(n21402) );
  AOI221_X1 U23056 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21405), 
        .C1(n21404), .C2(n21403), .A(n21402), .ZN(n21406) );
  NAND2_X1 U23057 ( .A1(n21407), .A2(n21406), .ZN(P1_U3008) );
  AOI22_X1 U23058 ( .A1(n21411), .A2(n21410), .B1(n21409), .B2(n21408), .ZN(
        n21419) );
  INV_X1 U23059 ( .A(n21412), .ZN(n21418) );
  OAI22_X1 U23060 ( .A1(n21415), .A2(n21414), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21413), .ZN(n21416) );
  NAND4_X1 U23061 ( .A1(n21419), .A2(n21418), .A3(n21417), .A4(n21416), .ZN(
        P1_U3031) );
  OAI22_X1 U23062 ( .A1(n21421), .A2(n21505), .B1(n21535), .B2(n21420), .ZN(
        n21422) );
  AOI211_X1 U23063 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21495), .B(n21422), .ZN(n21431) );
  INV_X1 U23064 ( .A(n21423), .ZN(n21429) );
  NAND4_X1 U23065 ( .A1(n21509), .A2(n21424), .A3(P1_REIP_REG_6__SCAN_IN), 
        .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n21443) );
  NAND2_X1 U23066 ( .A1(n21443), .A2(n21485), .ZN(n21438) );
  INV_X1 U23067 ( .A(n21438), .ZN(n21428) );
  NAND3_X1 U23068 ( .A1(n21509), .A2(n21424), .A3(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n21425) );
  NAND2_X1 U23069 ( .A1(n21426), .A2(n21425), .ZN(n21427) );
  AOI22_X1 U23070 ( .A1(n21429), .A2(n21525), .B1(n21428), .B2(n21427), .ZN(
        n21430) );
  OAI211_X1 U23071 ( .C1(n21432), .C2(n21519), .A(n21431), .B(n21430), .ZN(
        P1_U2834) );
  AOI22_X1 U23072 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n21529), .B1(n21490), .B2(
        n21433), .ZN(n21434) );
  OAI21_X1 U23073 ( .B1(n21435), .B2(n21519), .A(n21434), .ZN(n21436) );
  AOI211_X1 U23074 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21495), .B(n21436), .ZN(n21442) );
  INV_X1 U23075 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21437) );
  NOR2_X1 U23076 ( .A1(n21438), .A2(n21437), .ZN(n21439) );
  AOI21_X1 U23077 ( .B1(n21440), .B2(n21525), .A(n21439), .ZN(n21441) );
  OAI211_X1 U23078 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n21443), .A(n21442), .B(
        n21441), .ZN(P1_U2833) );
  NOR2_X1 U23079 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21453), .ZN(n21459) );
  AOI22_X1 U23080 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n21529), .B1(n21444), 
        .B2(n21459), .ZN(n21451) );
  OAI22_X1 U23081 ( .A1(n21446), .A2(n21519), .B1(n21535), .B2(n21445), .ZN(
        n21447) );
  AOI211_X1 U23082 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21495), .B(n21447), .ZN(n21450) );
  AOI22_X1 U23083 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21458), .B1(n21525), 
        .B2(n21448), .ZN(n21449) );
  NAND3_X1 U23084 ( .A1(n21451), .A2(n21450), .A3(n21449), .ZN(P1_U2829) );
  AOI22_X1 U23085 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(n21529), .B1(n21490), 
        .B2(n21452), .ZN(n21463) );
  NOR3_X1 U23086 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n21454), .A3(n21453), 
        .ZN(n21455) );
  AOI211_X1 U23087 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21495), .B(n21455), .ZN(n21462) );
  AOI22_X1 U23088 ( .A1(n21457), .A2(n21530), .B1(n21525), .B2(n21456), .ZN(
        n21461) );
  OAI21_X1 U23089 ( .B1(n21459), .B2(n21458), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n21460) );
  NAND4_X1 U23090 ( .A1(n21463), .A2(n21462), .A3(n21461), .A4(n21460), .ZN(
        P1_U2828) );
  OAI22_X1 U23091 ( .A1(n21465), .A2(n21505), .B1(n21535), .B2(n21464), .ZN(
        n21466) );
  AOI211_X1 U23092 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21495), .B(n21466), .ZN(n21472) );
  AOI22_X1 U23093 ( .A1(n21468), .A2(n21525), .B1(n21530), .B2(n21467), .ZN(
        n21471) );
  OAI221_X1 U23094 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n21475), .C1(n21469), 
        .C2(n21473), .A(n21485), .ZN(n21470) );
  NAND3_X1 U23095 ( .A1(n21472), .A2(n21471), .A3(n21470), .ZN(P1_U2826) );
  NAND2_X1 U23096 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n21474) );
  NOR2_X1 U23097 ( .A1(n21474), .A2(n21473), .ZN(n21484) );
  AOI22_X1 U23098 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n21475), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n21485), .ZN(n21483) );
  AOI22_X1 U23099 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n21517), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(n21529), .ZN(n21476) );
  INV_X1 U23100 ( .A(n21476), .ZN(n21477) );
  AOI211_X1 U23101 ( .C1(n21530), .C2(n21478), .A(n21495), .B(n21477), .ZN(
        n21482) );
  AOI22_X1 U23102 ( .A1(n21480), .A2(n21525), .B1(n21490), .B2(n21479), .ZN(
        n21481) );
  OAI211_X1 U23103 ( .C1(n21484), .C2(n21483), .A(n21482), .B(n21481), .ZN(
        P1_U2825) );
  AOI21_X1 U23104 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n21485), .A(n21484), 
        .ZN(n21493) );
  OAI22_X1 U23105 ( .A1(n21487), .A2(n21519), .B1(n21486), .B2(n21505), .ZN(
        n21488) );
  AOI211_X1 U23106 ( .C1(n21517), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21495), .B(n21488), .ZN(n21492) );
  AOI22_X1 U23107 ( .A1(n21638), .A2(n21525), .B1(n21490), .B2(n21489), .ZN(
        n21491) );
  OAI211_X1 U23108 ( .C1(n21494), .C2(n21493), .A(n21492), .B(n21491), .ZN(
        P1_U2824) );
  AOI21_X1 U23109 ( .B1(n21517), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21495), .ZN(n21496) );
  INV_X1 U23110 ( .A(n21496), .ZN(n21500) );
  OAI22_X1 U23111 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n21498), .B1(n21497), 
        .B2(n21519), .ZN(n21499) );
  AOI211_X1 U23112 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n21529), .A(n21500), .B(
        n21499), .ZN(n21503) );
  AOI22_X1 U23113 ( .A1(n21642), .A2(n21525), .B1(n21501), .B2(
        P1_REIP_REG_18__SCAN_IN), .ZN(n21502) );
  OAI211_X1 U23114 ( .C1(n21535), .C2(n21504), .A(n21503), .B(n21502), .ZN(
        P1_U2822) );
  OAI22_X1 U23115 ( .A1(n21507), .A2(n21519), .B1(n21506), .B2(n21505), .ZN(
        n21514) );
  AOI21_X1 U23116 ( .B1(n21509), .B2(n21508), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n21511) );
  OAI22_X1 U23117 ( .A1(n21512), .A2(n21537), .B1(n21511), .B2(n21510), .ZN(
        n21513) );
  AOI211_X1 U23118 ( .C1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n21517), .A(
        n21514), .B(n21513), .ZN(n21515) );
  OAI21_X1 U23119 ( .B1(n21535), .B2(n21516), .A(n21515), .ZN(P1_U2820) );
  AOI22_X1 U23120 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21517), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(n21529), .ZN(n21518) );
  OAI21_X1 U23121 ( .B1(n21520), .B2(n21519), .A(n21518), .ZN(n21521) );
  AOI221_X1 U23122 ( .B1(n21524), .B2(n21523), .C1(n21522), .C2(
        P1_REIP_REG_22__SCAN_IN), .A(n21521), .ZN(n21527) );
  NAND2_X1 U23123 ( .A1(n21654), .A2(n21525), .ZN(n21526) );
  OAI211_X1 U23124 ( .C1(n21528), .C2(n21535), .A(n21527), .B(n21526), .ZN(
        P1_U2818) );
  AOI22_X1 U23125 ( .A1(n21531), .A2(n21530), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n21529), .ZN(n21543) );
  INV_X1 U23126 ( .A(n21532), .ZN(n21541) );
  NAND2_X1 U23127 ( .A1(n21534), .A2(n21533), .ZN(n21540) );
  OAI22_X1 U23128 ( .A1(n21538), .A2(n21537), .B1(n21536), .B2(n21535), .ZN(
        n21539) );
  AOI21_X1 U23129 ( .B1(n21541), .B2(n21540), .A(n21539), .ZN(n21542) );
  OAI211_X1 U23130 ( .C1(n21545), .C2(n21544), .A(n21543), .B(n21542), .ZN(
        P1_U2817) );
  OAI21_X1 U23131 ( .B1(n21548), .B2(n21547), .A(n21546), .ZN(P1_U2806) );
  NOR2_X1 U23132 ( .A1(n11213), .A2(n21549), .ZN(n21551) );
  OAI21_X1 U23133 ( .B1(n21551), .B2(n11847), .A(n21550), .ZN(P1_U3163) );
  OAI221_X1 U23134 ( .B1(n21805), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n21805), 
        .C2(n21553), .A(n21552), .ZN(P1_U3466) );
  INV_X1 U23135 ( .A(n21553), .ZN(n21554) );
  AOI21_X1 U23136 ( .B1(n21556), .B2(n21555), .A(n21554), .ZN(n21557) );
  OAI22_X1 U23137 ( .A1(n21559), .A2(n21558), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21557), .ZN(n21560) );
  OAI21_X1 U23138 ( .B1(n21562), .B2(n21561), .A(n21560), .ZN(P1_U3161) );
  OAI21_X1 U23139 ( .B1(n21564), .B2(n21829), .A(n21563), .ZN(P1_U2805) );
  AOI21_X1 U23140 ( .B1(n21566), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21565), 
        .ZN(n21567) );
  INV_X1 U23141 ( .A(n21567), .ZN(P1_U3465) );
  INV_X1 U23142 ( .A(n21568), .ZN(n21570) );
  OAI21_X1 U23143 ( .B1(n21572), .B2(n21569), .A(n21570), .ZN(P2_U2818) );
  OAI21_X1 U23144 ( .B1(n21572), .B2(n21571), .A(n21570), .ZN(P2_U3592) );
  INV_X1 U23145 ( .A(n21573), .ZN(n21575) );
  OAI21_X1 U23146 ( .B1(n21577), .B2(n21574), .A(n21575), .ZN(P3_U2636) );
  OAI21_X1 U23147 ( .B1(n21577), .B2(n21576), .A(n21575), .ZN(P3_U3281) );
  INV_X1 U23148 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21617) );
  AOI21_X1 U23149 ( .B1(HOLD), .B2(n21578), .A(n21617), .ZN(n21579) );
  AOI21_X1 U23150 ( .B1(n21628), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21614), 
        .ZN(n21635) );
  AOI21_X1 U23151 ( .B1(n21625), .B2(NA), .A(n21622), .ZN(n21627) );
  OAI22_X1 U23152 ( .A1(n21621), .A2(n21579), .B1(n21635), .B2(n21627), .ZN(
        P3_U3029) );
  AOI21_X1 U23153 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n21585), .A(n21618), .ZN(n21581) );
  AOI21_X1 U23154 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .A(n21581), .ZN(n21584) );
  AOI22_X1 U23155 ( .A1(n21586), .A2(n21607), .B1(n21581), .B2(n21580), .ZN(
        n21583) );
  NOR2_X1 U23156 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21607), .ZN(n21582) );
  AOI21_X1 U23157 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21586), .A(n21591), 
        .ZN(n21593) );
  OAI33_X1 U23158 ( .A1(n21591), .A2(n21584), .A3(n21583), .B1(n21585), .B2(
        n21582), .B3(n21593), .ZN(P1_U3196) );
  OAI21_X1 U23159 ( .B1(n21585), .B2(n21618), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21589) );
  OAI221_X1 U23160 ( .B1(n21586), .B2(HOLD), .C1(n21586), .C2(n21585), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n21588) );
  OAI211_X1 U23161 ( .C1(n21591), .C2(n21589), .A(n21588), .B(n21587), .ZN(
        P1_U3195) );
  NOR2_X1 U23162 ( .A1(n11627), .A2(n21618), .ZN(n21590) );
  AOI211_X1 U23163 ( .C1(NA), .C2(n21591), .A(n21590), .B(n21589), .ZN(n21592)
         );
  OAI22_X1 U23164 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21593), .B1(n22246), 
        .B2(n21592), .ZN(P1_U3194) );
  NAND2_X1 U23165 ( .A1(n21594), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21608) );
  OAI221_X1 U23166 ( .B1(n21608), .B2(P2_STATE_REG_2__SCAN_IN), .C1(
        P2_STATE_REG_0__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21595) );
  INV_X1 U23167 ( .A(n21595), .ZN(n21599) );
  INV_X1 U23168 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21606) );
  AOI22_X1 U23169 ( .A1(HOLD), .A2(n21596), .B1(NA), .B2(n21606), .ZN(n21597)
         );
  OAI22_X1 U23170 ( .A1(n21600), .A2(n21599), .B1(n21598), .B2(n21597), .ZN(
        P2_U3209) );
  NAND2_X1 U23171 ( .A1(n21601), .A2(HOLD), .ZN(n21603) );
  OAI211_X1 U23172 ( .C1(n21612), .C2(n21618), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21602) );
  NAND4_X1 U23173 ( .A1(n21604), .A2(n21603), .A3(n21608), .A4(n21602), .ZN(
        P2_U3210) );
  INV_X1 U23174 ( .A(n21608), .ZN(n21605) );
  AOI221_X1 U23175 ( .B1(HOLD), .B2(P2_STATE_REG_0__SCAN_IN), .C1(n21607), 
        .C2(n21606), .A(n21605), .ZN(n21613) );
  OAI22_X1 U23176 ( .A1(NA), .A2(n21608), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21609) );
  OAI211_X1 U23177 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21609), .ZN(n21610) );
  OAI211_X1 U23178 ( .C1(n21613), .C2(n21612), .A(n21611), .B(n21610), .ZN(
        P2_U3211) );
  NAND2_X1 U23179 ( .A1(HOLD), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n21620) );
  INV_X1 U23180 ( .A(n21620), .ZN(n21632) );
  NOR2_X1 U23181 ( .A1(n21632), .A2(n21614), .ZN(n21616) );
  AOI21_X1 U23182 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(n21616), .A(n21615), .ZN(n21626) );
  NAND2_X1 U23183 ( .A1(n21618), .A2(n21617), .ZN(n21630) );
  OAI221_X1 U23184 ( .B1(n21628), .B2(n21620), .C1(n21628), .C2(n21630), .A(
        n21619), .ZN(n21624) );
  OAI21_X1 U23185 ( .B1(n21628), .B2(n21622), .A(n21621), .ZN(n21623) );
  OAI221_X1 U23186 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21626), .C1(n21625), 
        .C2(n21624), .A(n21623), .ZN(P3_U3030) );
  INV_X1 U23187 ( .A(n21627), .ZN(n21634) );
  NAND2_X1 U23188 ( .A1(n21628), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n21629) );
  OAI22_X1 U23189 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n21629), .ZN(n21631) );
  OAI211_X1 U23190 ( .C1(n21632), .C2(n21631), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(n21630), .ZN(n21633) );
  OAI21_X1 U23191 ( .B1(n21635), .B2(n21634), .A(n21633), .ZN(P3_U3031) );
  INV_X1 U23192 ( .A(n21636), .ZN(n21651) );
  AOI22_X1 U23193 ( .A1(n21651), .A2(n21637), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n21649), .ZN(n21640) );
  AOI22_X1 U23194 ( .A1(n21638), .A2(n21653), .B1(n21652), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n21639) );
  OAI211_X1 U23195 ( .C1(n21657), .C2(n21676), .A(n21640), .B(n21639), .ZN(
        P1_U2888) );
  AOI22_X1 U23196 ( .A1(n21651), .A2(n21641), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n21649), .ZN(n21644) );
  AOI22_X1 U23197 ( .A1(n21642), .A2(n21653), .B1(n21652), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n21643) );
  OAI211_X1 U23198 ( .C1(n21657), .C2(n21904), .A(n21644), .B(n21643), .ZN(
        P1_U2886) );
  AOI22_X1 U23199 ( .A1(n21651), .A2(n21645), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n21649), .ZN(n21648) );
  AOI22_X1 U23200 ( .A1(n21646), .A2(n21653), .B1(n21652), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n21647) );
  OAI211_X1 U23201 ( .C1(n21657), .C2(n21993), .A(n21648), .B(n21647), .ZN(
        P1_U2884) );
  AOI22_X1 U23202 ( .A1(n21651), .A2(n21650), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n21649), .ZN(n21656) );
  AOI22_X1 U23203 ( .A1(n21654), .A2(n21653), .B1(n21652), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n21655) );
  OAI211_X1 U23204 ( .C1(n21657), .C2(n22086), .A(n21656), .B(n21655), .ZN(
        P1_U2882) );
  INV_X1 U23205 ( .A(n21752), .ZN(n21658) );
  INV_X1 U23206 ( .A(n22143), .ZN(n21659) );
  NAND2_X1 U23207 ( .A1(n21659), .A2(n21852), .ZN(n21660) );
  NAND2_X1 U23208 ( .A1(n21852), .A2(n21829), .ZN(n21795) );
  OAI21_X1 U23209 ( .B1(n21660), .B2(n22238), .A(n21795), .ZN(n21673) );
  OR2_X1 U23210 ( .A1(n21753), .A2(n11214), .ZN(n21690) );
  INV_X1 U23211 ( .A(n13964), .ZN(n21832) );
  NOR2_X1 U23212 ( .A1(n21690), .A2(n21832), .ZN(n21670) );
  NOR2_X1 U23213 ( .A1(n21668), .A2(n11847), .ZN(n21775) );
  INV_X1 U23214 ( .A(n21773), .ZN(n21755) );
  NOR2_X1 U23215 ( .A1(n21754), .A2(n21755), .ZN(n21714) );
  INV_X1 U23216 ( .A(n21845), .ZN(n21808) );
  NAND2_X2 U23217 ( .A1(n21664), .A2(n21662), .ZN(n22136) );
  NAND2_X2 U23218 ( .A1(n21664), .A2(n21663), .ZN(n22134) );
  OAI22_X2 U23219 ( .A1(n21665), .A2(n22136), .B1(n16343), .B2(n22134), .ZN(
        n21837) );
  NOR2_X2 U23220 ( .A1(n22132), .A2(n21667), .ZN(n21844) );
  NOR3_X1 U23221 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21683) );
  INV_X1 U23222 ( .A(n21683), .ZN(n21680) );
  NOR2_X1 U23223 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21680), .ZN(
        n22133) );
  AOI22_X1 U23224 ( .A1(n22238), .A2(n21837), .B1(n21844), .B2(n22133), .ZN(
        n21678) );
  INV_X1 U23225 ( .A(n21668), .ZN(n21669) );
  NOR2_X1 U23226 ( .A1(n21669), .A2(n11847), .ZN(n21799) );
  INV_X1 U23227 ( .A(n21670), .ZN(n21672) );
  INV_X1 U23228 ( .A(n22133), .ZN(n21671) );
  AOI22_X1 U23229 ( .A1(n21673), .A2(n21672), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21671), .ZN(n21674) );
  OAI211_X1 U23230 ( .C1(n21714), .C2(n11847), .A(n21780), .B(n21674), .ZN(
        n22137) );
  OAI22_X2 U23231 ( .A1(n21676), .A2(n22136), .B1(n21675), .B2(n22134), .ZN(
        n21853) );
  AOI22_X1 U23232 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n21853), .ZN(n21677) );
  OAI211_X1 U23233 ( .C1(n22140), .C2(n21808), .A(n21678), .B(n21677), .ZN(
        P1_U3033) );
  INV_X1 U23234 ( .A(n21853), .ZN(n21840) );
  INV_X1 U23235 ( .A(n21690), .ZN(n21700) );
  INV_X1 U23236 ( .A(n21679), .ZN(n21811) );
  NOR2_X1 U23237 ( .A1(n21810), .A2(n21680), .ZN(n22141) );
  AOI21_X1 U23238 ( .B1(n21700), .B2(n21811), .A(n22141), .ZN(n21681) );
  OAI22_X1 U23239 ( .A1(n21681), .A2(n21850), .B1(n21680), .B2(n11847), .ZN(
        n22142) );
  AOI22_X1 U23240 ( .A1(n22142), .A2(n21845), .B1(n21844), .B2(n22141), .ZN(
        n21685) );
  OAI21_X1 U23241 ( .B1(n21711), .B2(n21829), .A(n21681), .ZN(n21682) );
  OAI221_X1 U23242 ( .B1(n21852), .B2(n21683), .C1(n21850), .C2(n21682), .A(
        n21848), .ZN(n22144) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n21837), .ZN(n21684) );
  OAI211_X1 U23244 ( .C1(n21840), .C2(n22149), .A(n21685), .B(n21684), .ZN(
        P1_U3041) );
  INV_X1 U23245 ( .A(n21821), .ZN(n21688) );
  NAND2_X1 U23246 ( .A1(n22149), .A2(n21852), .ZN(n21689) );
  OAI21_X1 U23247 ( .B1(n22156), .B2(n21689), .A(n21795), .ZN(n21693) );
  NOR2_X1 U23248 ( .A1(n21690), .A2(n13964), .ZN(n21695) );
  INV_X1 U23249 ( .A(n21837), .ZN(n21856) );
  INV_X1 U23250 ( .A(n21844), .ZN(n21691) );
  NOR3_X1 U23251 ( .A1(n21823), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21706) );
  NAND2_X1 U23252 ( .A1(n21810), .A2(n21706), .ZN(n22147) );
  OAI22_X1 U23253 ( .A1(n22149), .A2(n21856), .B1(n21691), .B2(n22147), .ZN(
        n21692) );
  INV_X1 U23254 ( .A(n21692), .ZN(n21698) );
  INV_X1 U23255 ( .A(n21693), .ZN(n21696) );
  NOR2_X1 U23256 ( .A1(n11525), .A2(n11847), .ZN(n21735) );
  AOI21_X1 U23257 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22147), .A(n21735), 
        .ZN(n21694) );
  OAI211_X1 U23258 ( .C1(n21696), .C2(n21695), .A(n21694), .B(n21780), .ZN(
        n22151) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22151), .B1(
        n22156), .B2(n21853), .ZN(n21697) );
  OAI211_X1 U23260 ( .C1(n22154), .C2(n21808), .A(n21698), .B(n21697), .ZN(
        P1_U3049) );
  INV_X1 U23261 ( .A(n21706), .ZN(n21704) );
  NOR2_X1 U23262 ( .A1(n21810), .A2(n21704), .ZN(n22155) );
  AOI21_X1 U23263 ( .B1(n21700), .B2(n11087), .A(n22155), .ZN(n21708) );
  AOI21_X1 U23264 ( .B1(n21702), .B2(n21701), .A(n21850), .ZN(n21709) );
  INV_X1 U23265 ( .A(n21709), .ZN(n21703) );
  OAI22_X1 U23266 ( .A1(n11847), .A2(n21704), .B1(n21708), .B2(n21703), .ZN(
        n21705) );
  AOI22_X1 U23267 ( .A1(n22156), .A2(n21837), .B1(n21844), .B2(n22155), .ZN(
        n21713) );
  OAI21_X1 U23268 ( .B1(n21852), .B2(n21706), .A(n21848), .ZN(n21707) );
  AOI21_X1 U23269 ( .B1(n21709), .B2(n21708), .A(n21707), .ZN(n21710) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22157), .B1(
        n22163), .B2(n21853), .ZN(n21712) );
  OAI211_X1 U23271 ( .C1(n22160), .C2(n21808), .A(n21713), .B(n21712), .ZN(
        P1_U3057) );
  NOR3_X1 U23272 ( .A1(n21824), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21728) );
  INV_X1 U23273 ( .A(n21728), .ZN(n21724) );
  NOR2_X1 U23274 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21724), .ZN(
        n22162) );
  INV_X1 U23275 ( .A(n21714), .ZN(n21717) );
  INV_X1 U23276 ( .A(n21799), .ZN(n21827) );
  OR2_X1 U23277 ( .A1(n13802), .A2(n21715), .ZN(n21733) );
  INV_X1 U23278 ( .A(n21733), .ZN(n21744) );
  NAND3_X1 U23279 ( .A1(n21744), .A2(n21852), .A3(n13964), .ZN(n21716) );
  OAI21_X1 U23280 ( .B1(n21717), .B2(n21827), .A(n21716), .ZN(n22161) );
  AOI22_X1 U23281 ( .A1(n21844), .A2(n22162), .B1(n21845), .B2(n22161), .ZN(
        n21723) );
  INV_X1 U23282 ( .A(n22163), .ZN(n21718) );
  AOI21_X1 U23283 ( .B1(n21718), .B2(n22172), .A(n21829), .ZN(n21719) );
  AOI21_X1 U23284 ( .B1(n21744), .B2(n13964), .A(n21719), .ZN(n21720) );
  NOR2_X1 U23285 ( .A1(n21720), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21721) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n21837), .ZN(n21722) );
  OAI211_X1 U23287 ( .C1(n21840), .C2(n22172), .A(n21723), .B(n21722), .ZN(
        P1_U3065) );
  NOR2_X1 U23288 ( .A1(n21810), .A2(n21724), .ZN(n22167) );
  AOI21_X1 U23289 ( .B1(n21744), .B2(n21811), .A(n22167), .ZN(n21725) );
  OAI22_X1 U23290 ( .A1(n21725), .A2(n21850), .B1(n21724), .B2(n11847), .ZN(
        n22168) );
  AOI22_X1 U23291 ( .A1(n21845), .A2(n22168), .B1(n21844), .B2(n22167), .ZN(
        n21730) );
  INV_X1 U23292 ( .A(n21742), .ZN(n21726) );
  OAI21_X1 U23293 ( .B1(n21726), .B2(n21829), .A(n21725), .ZN(n21727) );
  OAI221_X1 U23294 ( .B1(n21852), .B2(n21728), .C1(n21850), .C2(n21727), .A(
        n21848), .ZN(n22169) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n21853), .ZN(n21729) );
  OAI211_X1 U23296 ( .C1(n21856), .C2(n22172), .A(n21730), .B(n21729), .ZN(
        P1_U3073) );
  INV_X1 U23297 ( .A(n22174), .ZN(n21731) );
  NAND2_X1 U23298 ( .A1(n21731), .A2(n21852), .ZN(n21732) );
  OAI21_X1 U23299 ( .B1(n21732), .B2(n22181), .A(n21795), .ZN(n21737) );
  NOR2_X1 U23300 ( .A1(n21733), .A2(n13964), .ZN(n21734) );
  NOR3_X1 U23301 ( .A1(n21824), .A2(n21823), .A3(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21749) );
  INV_X1 U23302 ( .A(n21749), .ZN(n21745) );
  NOR2_X1 U23303 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21745), .ZN(
        n22173) );
  AOI22_X1 U23304 ( .A1(n22174), .A2(n21837), .B1(n22173), .B2(n21844), .ZN(
        n21740) );
  INV_X1 U23305 ( .A(n21734), .ZN(n21736) );
  AOI21_X1 U23306 ( .B1(n21737), .B2(n21736), .A(n21735), .ZN(n21738) );
  OAI211_X1 U23307 ( .C1(n22173), .C2(n21805), .A(n21835), .B(n21738), .ZN(
        n22175) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n21853), .ZN(n21739) );
  OAI211_X1 U23309 ( .C1(n22178), .C2(n21808), .A(n21740), .B(n21739), .ZN(
        P1_U3081) );
  NOR2_X1 U23310 ( .A1(n21743), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22179) );
  AOI21_X1 U23311 ( .B1(n21744), .B2(n11087), .A(n22179), .ZN(n21747) );
  OAI22_X1 U23312 ( .A1(n21747), .A2(n21850), .B1(n21745), .B2(n11847), .ZN(
        n22180) );
  AOI22_X1 U23313 ( .A1(n22180), .A2(n21845), .B1(n21844), .B2(n22179), .ZN(
        n21751) );
  NAND2_X1 U23314 ( .A1(n21747), .A2(n21746), .ZN(n21748) );
  OAI221_X1 U23315 ( .B1(n21852), .B2(n21749), .C1(n21850), .C2(n21748), .A(
        n21848), .ZN(n22182) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n21837), .ZN(n21750) );
  OAI211_X1 U23317 ( .C1(n21840), .C2(n22185), .A(n21751), .B(n21750), .ZN(
        P1_U3089) );
  AND2_X1 U23318 ( .A1(n21753), .A2(n13802), .ZN(n21783) );
  NOR3_X1 U23319 ( .A1(n21825), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21767) );
  INV_X1 U23320 ( .A(n21767), .ZN(n21764) );
  NOR2_X1 U23321 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21764), .ZN(
        n22186) );
  AOI21_X1 U23322 ( .B1(n21783), .B2(n13964), .A(n22186), .ZN(n21759) );
  INV_X1 U23323 ( .A(n21754), .ZN(n21756) );
  NOR2_X1 U23324 ( .A1(n21756), .A2(n21755), .ZN(n21798) );
  INV_X1 U23325 ( .A(n21798), .ZN(n21801) );
  INV_X1 U23326 ( .A(n21775), .ZN(n21757) );
  OAI22_X1 U23327 ( .A1(n21759), .A2(n21850), .B1(n21801), .B2(n21757), .ZN(
        n22187) );
  AOI22_X1 U23328 ( .A1(n22187), .A2(n21845), .B1(n21844), .B2(n22186), .ZN(
        n21763) );
  INV_X1 U23329 ( .A(n22197), .ZN(n21758) );
  OAI21_X1 U23330 ( .B1(n21758), .B2(n22188), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21760) );
  NAND2_X1 U23331 ( .A1(n21760), .A2(n21759), .ZN(n21761) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n21837), .ZN(n21762) );
  OAI211_X1 U23333 ( .C1(n21840), .C2(n22197), .A(n21763), .B(n21762), .ZN(
        P1_U3097) );
  NOR2_X1 U23334 ( .A1(n21810), .A2(n21764), .ZN(n22192) );
  AOI21_X1 U23335 ( .B1(n21783), .B2(n21811), .A(n22192), .ZN(n21765) );
  OAI22_X1 U23336 ( .A1(n21765), .A2(n21850), .B1(n21764), .B2(n11847), .ZN(
        n22193) );
  AOI22_X1 U23337 ( .A1(n22193), .A2(n21845), .B1(n21844), .B2(n22192), .ZN(
        n21769) );
  INV_X1 U23338 ( .A(n21770), .ZN(n21790) );
  OAI21_X1 U23339 ( .B1(n21790), .B2(n21829), .A(n21765), .ZN(n21766) );
  OAI221_X1 U23340 ( .B1(n21852), .B2(n21767), .C1(n21850), .C2(n21766), .A(
        n21848), .ZN(n22194) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n21853), .ZN(n21768) );
  OAI211_X1 U23342 ( .C1(n21856), .C2(n22197), .A(n21769), .B(n21768), .ZN(
        P1_U3105) );
  INV_X1 U23343 ( .A(n22199), .ZN(n21771) );
  NAND3_X1 U23344 ( .A1(n21771), .A2(n21852), .A3(n22210), .ZN(n21772) );
  NAND2_X1 U23345 ( .A1(n21772), .A2(n21795), .ZN(n21778) );
  OR2_X1 U23346 ( .A1(n21773), .A2(n21825), .ZN(n21828) );
  INV_X1 U23347 ( .A(n21828), .ZN(n21774) );
  NOR3_X1 U23348 ( .A1(n21825), .A2(n21823), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21787) );
  NAND2_X1 U23349 ( .A1(n21810), .A2(n21787), .ZN(n22061) );
  INV_X1 U23350 ( .A(n22061), .ZN(n22198) );
  AOI22_X1 U23351 ( .A1(n22199), .A2(n21837), .B1(n21844), .B2(n22198), .ZN(
        n21782) );
  INV_X1 U23352 ( .A(n21776), .ZN(n21777) );
  AOI22_X1 U23353 ( .A1(n21778), .A2(n21777), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22061), .ZN(n21779) );
  NAND2_X1 U23354 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21828), .ZN(n21834) );
  NAND3_X1 U23355 ( .A1(n21780), .A2(n21779), .A3(n21834), .ZN(n22201) );
  INV_X1 U23356 ( .A(n22210), .ZN(n22200) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22201), .B1(
        n22200), .B2(n21853), .ZN(n21781) );
  OAI211_X1 U23358 ( .C1(n22204), .C2(n21808), .A(n21782), .B(n21781), .ZN(
        P1_U3113) );
  INV_X1 U23359 ( .A(n21787), .ZN(n21784) );
  NOR2_X1 U23360 ( .A1(n21810), .A2(n21784), .ZN(n22205) );
  AOI21_X1 U23361 ( .B1(n21783), .B2(n11087), .A(n22205), .ZN(n21785) );
  OAI22_X1 U23362 ( .A1(n21785), .A2(n21850), .B1(n21784), .B2(n11847), .ZN(
        n22206) );
  AOI22_X1 U23363 ( .A1(n21845), .A2(n22206), .B1(n21844), .B2(n22205), .ZN(
        n21792) );
  NOR3_X1 U23364 ( .A1(n21790), .A2(n21850), .A3(n21786), .ZN(n21788) );
  AOI22_X1 U23365 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n22213), .B2(n21853), .ZN(n21791) );
  OAI211_X1 U23366 ( .C1(n21856), .C2(n22210), .A(n21792), .B(n21791), .ZN(
        P1_U3121) );
  INV_X1 U23367 ( .A(n22213), .ZN(n21794) );
  NAND3_X1 U23368 ( .A1(n21794), .A2(n21852), .A3(n22224), .ZN(n21796) );
  NAND2_X1 U23369 ( .A1(n21796), .A2(n21795), .ZN(n21803) );
  OR2_X1 U23370 ( .A1(n13802), .A2(n21797), .ZN(n21809) );
  NOR2_X1 U23371 ( .A1(n21809), .A2(n21832), .ZN(n21800) );
  INV_X1 U23372 ( .A(n22224), .ZN(n22212) );
  NOR3_X1 U23373 ( .A1(n21824), .A2(n21825), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21815) );
  INV_X1 U23374 ( .A(n21815), .ZN(n21812) );
  NOR2_X1 U23375 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21812), .ZN(
        n22211) );
  AOI22_X1 U23376 ( .A1(n22212), .A2(n21853), .B1(n21844), .B2(n22211), .ZN(
        n21807) );
  INV_X1 U23377 ( .A(n21800), .ZN(n21802) );
  AOI22_X1 U23378 ( .A1(n21803), .A2(n21802), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21801), .ZN(n21804) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n21837), .ZN(n21806) );
  OAI211_X1 U23380 ( .C1(n22218), .C2(n21808), .A(n21807), .B(n21806), .ZN(
        P1_U3129) );
  INV_X1 U23381 ( .A(n21809), .ZN(n21842) );
  NOR2_X1 U23382 ( .A1(n21810), .A2(n21812), .ZN(n22219) );
  AOI21_X1 U23383 ( .B1(n21842), .B2(n21811), .A(n22219), .ZN(n21813) );
  OAI22_X1 U23384 ( .A1(n21813), .A2(n21850), .B1(n21812), .B2(n11847), .ZN(
        n22220) );
  AOI22_X1 U23385 ( .A1(n21845), .A2(n22220), .B1(n21844), .B2(n22219), .ZN(
        n21820) );
  INV_X1 U23386 ( .A(n21822), .ZN(n21818) );
  OAI21_X1 U23387 ( .B1(n21818), .B2(n21829), .A(n21813), .ZN(n21814) );
  OAI221_X1 U23388 ( .B1(n21852), .B2(n21815), .C1(n21850), .C2(n21814), .A(
        n21848), .ZN(n22221) );
  INV_X1 U23389 ( .A(n21816), .ZN(n21817) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n21853), .ZN(n21819) );
  OAI211_X1 U23391 ( .C1(n21856), .C2(n22224), .A(n21820), .B(n21819), .ZN(
        P1_U3137) );
  NOR3_X1 U23392 ( .A1(n21825), .A2(n21824), .A3(n21823), .ZN(n21851) );
  INV_X1 U23393 ( .A(n21851), .ZN(n21843) );
  NOR2_X1 U23394 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21843), .ZN(
        n22226) );
  NAND3_X1 U23395 ( .A1(n21842), .A2(n21832), .A3(n21852), .ZN(n21826) );
  OAI21_X1 U23396 ( .B1(n21828), .B2(n21827), .A(n21826), .ZN(n22225) );
  AOI22_X1 U23397 ( .A1(n21844), .A2(n22226), .B1(n21845), .B2(n22225), .ZN(
        n21839) );
  INV_X1 U23398 ( .A(n22228), .ZN(n21830) );
  AOI21_X1 U23399 ( .B1(n21830), .B2(n22242), .A(n21829), .ZN(n21831) );
  AOI21_X1 U23400 ( .B1(n21842), .B2(n21832), .A(n21831), .ZN(n21833) );
  NOR2_X1 U23401 ( .A1(n21833), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21836) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n21837), .ZN(n21838) );
  OAI211_X1 U23403 ( .C1(n21840), .C2(n22242), .A(n21839), .B(n21838), .ZN(
        P1_U3145) );
  INV_X1 U23404 ( .A(n21841), .ZN(n22233) );
  AOI21_X1 U23405 ( .B1(n21842), .B2(n11087), .A(n22233), .ZN(n21847) );
  OAI22_X1 U23406 ( .A1(n21847), .A2(n21850), .B1(n21843), .B2(n11847), .ZN(
        n22236) );
  AOI22_X1 U23407 ( .A1(n22236), .A2(n21845), .B1(n21844), .B2(n22233), .ZN(
        n21855) );
  NAND2_X1 U23408 ( .A1(n21847), .A2(n21846), .ZN(n21849) );
  OAI221_X1 U23409 ( .B1(n21852), .B2(n21851), .C1(n21850), .C2(n21849), .A(
        n21848), .ZN(n22239) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n21853), .ZN(n21854) );
  OAI211_X1 U23411 ( .C1(n21856), .C2(n22242), .A(n21855), .B(n21854), .ZN(
        P1_U3153) );
  OAI22_X2 U23412 ( .A1(n21858), .A2(n22134), .B1(n15835), .B2(n22136), .ZN(
        n21890) );
  NOR2_X2 U23413 ( .A1(n22132), .A2(n21859), .ZN(n21894) );
  AOI22_X1 U23414 ( .A1(n22238), .A2(n21890), .B1(n21894), .B2(n22133), .ZN(
        n21862) );
  OAI22_X2 U23415 ( .A1(n15861), .A2(n22136), .B1(n21860), .B2(n22134), .ZN(
        n21896) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n21896), .ZN(n21861) );
  OAI211_X1 U23417 ( .C1(n22140), .C2(n21887), .A(n21862), .B(n21861), .ZN(
        P1_U3034) );
  INV_X1 U23418 ( .A(n21896), .ZN(n21893) );
  AOI22_X1 U23419 ( .A1(n22142), .A2(n21895), .B1(n21894), .B2(n22141), .ZN(
        n21864) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n21890), .ZN(n21863) );
  OAI211_X1 U23421 ( .C1(n21893), .C2(n22149), .A(n21864), .B(n21863), .ZN(
        P1_U3042) );
  INV_X1 U23422 ( .A(n22147), .ZN(n22091) );
  AOI22_X1 U23423 ( .A1(n22156), .A2(n21896), .B1(n21894), .B2(n22091), .ZN(
        n21866) );
  INV_X1 U23424 ( .A(n22149), .ZN(n22092) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22151), .B1(
        n22092), .B2(n21890), .ZN(n21865) );
  OAI211_X1 U23426 ( .C1(n22154), .C2(n21887), .A(n21866), .B(n21865), .ZN(
        P1_U3050) );
  AOI22_X1 U23427 ( .A1(n22163), .A2(n21896), .B1(n21894), .B2(n22155), .ZN(
        n21868) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22157), .B1(
        n22156), .B2(n21890), .ZN(n21867) );
  OAI211_X1 U23429 ( .C1(n22160), .C2(n21887), .A(n21868), .B(n21867), .ZN(
        P1_U3058) );
  AOI22_X1 U23430 ( .A1(n21894), .A2(n22162), .B1(n21895), .B2(n22161), .ZN(
        n21870) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n21890), .ZN(n21869) );
  OAI211_X1 U23432 ( .C1(n21893), .C2(n22172), .A(n21870), .B(n21869), .ZN(
        P1_U3066) );
  INV_X1 U23433 ( .A(n21890), .ZN(n21899) );
  AOI22_X1 U23434 ( .A1(n21895), .A2(n22168), .B1(n21894), .B2(n22167), .ZN(
        n21872) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n21896), .ZN(n21871) );
  OAI211_X1 U23436 ( .C1(n21899), .C2(n22172), .A(n21872), .B(n21871), .ZN(
        P1_U3074) );
  AOI22_X1 U23437 ( .A1(n22181), .A2(n21896), .B1(n21894), .B2(n22173), .ZN(
        n21874) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22175), .B1(
        n22174), .B2(n21890), .ZN(n21873) );
  OAI211_X1 U23439 ( .C1(n22178), .C2(n21887), .A(n21874), .B(n21873), .ZN(
        P1_U3082) );
  AOI22_X1 U23440 ( .A1(n22180), .A2(n21895), .B1(n21894), .B2(n22179), .ZN(
        n21876) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n21890), .ZN(n21875) );
  OAI211_X1 U23442 ( .C1(n21893), .C2(n22185), .A(n21876), .B(n21875), .ZN(
        P1_U3090) );
  AOI22_X1 U23443 ( .A1(n22187), .A2(n21895), .B1(n21894), .B2(n22186), .ZN(
        n21878) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n21890), .ZN(n21877) );
  OAI211_X1 U23445 ( .C1(n21893), .C2(n22197), .A(n21878), .B(n21877), .ZN(
        P1_U3098) );
  AOI22_X1 U23446 ( .A1(n22193), .A2(n21895), .B1(n21894), .B2(n22192), .ZN(
        n21880) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n21896), .ZN(n21879) );
  OAI211_X1 U23448 ( .C1(n21899), .C2(n22197), .A(n21880), .B(n21879), .ZN(
        P1_U3106) );
  AOI22_X1 U23449 ( .A1(n22199), .A2(n21890), .B1(n21894), .B2(n22198), .ZN(
        n21882) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22201), .B1(
        n22200), .B2(n21896), .ZN(n21881) );
  OAI211_X1 U23451 ( .C1(n22204), .C2(n21887), .A(n21882), .B(n21881), .ZN(
        P1_U3114) );
  AOI22_X1 U23452 ( .A1(n21895), .A2(n22206), .B1(n21894), .B2(n22205), .ZN(
        n21884) );
  AOI22_X1 U23453 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n22213), .B2(n21896), .ZN(n21883) );
  OAI211_X1 U23454 ( .C1(n21899), .C2(n22210), .A(n21884), .B(n21883), .ZN(
        P1_U3122) );
  AOI22_X1 U23455 ( .A1(n22212), .A2(n21896), .B1(n21894), .B2(n22211), .ZN(
        n21886) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n21890), .ZN(n21885) );
  OAI211_X1 U23457 ( .C1(n22218), .C2(n21887), .A(n21886), .B(n21885), .ZN(
        P1_U3130) );
  AOI22_X1 U23458 ( .A1(n21895), .A2(n22220), .B1(n21894), .B2(n22219), .ZN(
        n21889) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n21896), .ZN(n21888) );
  OAI211_X1 U23460 ( .C1(n21899), .C2(n22224), .A(n21889), .B(n21888), .ZN(
        P1_U3138) );
  AOI22_X1 U23461 ( .A1(n21894), .A2(n22226), .B1(n21895), .B2(n22225), .ZN(
        n21892) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n21890), .ZN(n21891) );
  OAI211_X1 U23463 ( .C1(n21893), .C2(n22242), .A(n21892), .B(n21891), .ZN(
        P1_U3146) );
  AOI22_X1 U23464 ( .A1(n22236), .A2(n21895), .B1(n21894), .B2(n22233), .ZN(
        n21898) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n21896), .ZN(n21897) );
  OAI211_X1 U23466 ( .C1(n21899), .C2(n22242), .A(n21898), .B(n21897), .ZN(
        P1_U3154) );
  INV_X1 U23467 ( .A(n21939), .ZN(n21931) );
  OAI22_X2 U23468 ( .A1(n21901), .A2(n22134), .B1(n15830), .B2(n22136), .ZN(
        n21934) );
  NOR2_X2 U23469 ( .A1(n22132), .A2(n21902), .ZN(n21938) );
  AOI22_X1 U23470 ( .A1(n22238), .A2(n21934), .B1(n21938), .B2(n22133), .ZN(
        n21906) );
  OAI22_X2 U23471 ( .A1(n21904), .A2(n22136), .B1(n21903), .B2(n22134), .ZN(
        n21940) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n21940), .ZN(n21905) );
  OAI211_X1 U23473 ( .C1(n22140), .C2(n21931), .A(n21906), .B(n21905), .ZN(
        P1_U3035) );
  INV_X1 U23474 ( .A(n21940), .ZN(n21937) );
  AOI22_X1 U23475 ( .A1(n22142), .A2(n21939), .B1(n21938), .B2(n22141), .ZN(
        n21908) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n21934), .ZN(n21907) );
  OAI211_X1 U23477 ( .C1(n21937), .C2(n22149), .A(n21908), .B(n21907), .ZN(
        P1_U3043) );
  AOI22_X1 U23478 ( .A1(n22156), .A2(n21940), .B1(n21938), .B2(n22091), .ZN(
        n21910) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22151), .B1(
        n22092), .B2(n21934), .ZN(n21909) );
  OAI211_X1 U23480 ( .C1(n22154), .C2(n21931), .A(n21910), .B(n21909), .ZN(
        P1_U3051) );
  AOI22_X1 U23481 ( .A1(n22163), .A2(n21940), .B1(n21938), .B2(n22155), .ZN(
        n21912) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22157), .B1(
        n22156), .B2(n21934), .ZN(n21911) );
  OAI211_X1 U23483 ( .C1(n22160), .C2(n21931), .A(n21912), .B(n21911), .ZN(
        P1_U3059) );
  AOI22_X1 U23484 ( .A1(n21938), .A2(n22162), .B1(n21939), .B2(n22161), .ZN(
        n21914) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n21934), .ZN(n21913) );
  OAI211_X1 U23486 ( .C1(n21937), .C2(n22172), .A(n21914), .B(n21913), .ZN(
        P1_U3067) );
  INV_X1 U23487 ( .A(n21934), .ZN(n21943) );
  AOI22_X1 U23488 ( .A1(n21939), .A2(n22168), .B1(n21938), .B2(n22167), .ZN(
        n21916) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n21940), .ZN(n21915) );
  OAI211_X1 U23490 ( .C1(n21943), .C2(n22172), .A(n21916), .B(n21915), .ZN(
        P1_U3075) );
  AOI22_X1 U23491 ( .A1(n22174), .A2(n21934), .B1(n22173), .B2(n21938), .ZN(
        n21918) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n21940), .ZN(n21917) );
  OAI211_X1 U23493 ( .C1(n22178), .C2(n21931), .A(n21918), .B(n21917), .ZN(
        P1_U3083) );
  AOI22_X1 U23494 ( .A1(n22180), .A2(n21939), .B1(n21938), .B2(n22179), .ZN(
        n21920) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n21934), .ZN(n21919) );
  OAI211_X1 U23496 ( .C1(n21937), .C2(n22185), .A(n21920), .B(n21919), .ZN(
        P1_U3091) );
  AOI22_X1 U23497 ( .A1(n22187), .A2(n21939), .B1(n21938), .B2(n22186), .ZN(
        n21922) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n21934), .ZN(n21921) );
  OAI211_X1 U23499 ( .C1(n21937), .C2(n22197), .A(n21922), .B(n21921), .ZN(
        P1_U3099) );
  AOI22_X1 U23500 ( .A1(n22193), .A2(n21939), .B1(n21938), .B2(n22192), .ZN(
        n21924) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n21940), .ZN(n21923) );
  OAI211_X1 U23502 ( .C1(n21943), .C2(n22197), .A(n21924), .B(n21923), .ZN(
        P1_U3107) );
  AOI22_X1 U23503 ( .A1(n22199), .A2(n21934), .B1(n21938), .B2(n22198), .ZN(
        n21926) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22201), .B1(
        n22200), .B2(n21940), .ZN(n21925) );
  OAI211_X1 U23505 ( .C1(n22204), .C2(n21931), .A(n21926), .B(n21925), .ZN(
        P1_U3115) );
  AOI22_X1 U23506 ( .A1(n21939), .A2(n22206), .B1(n21938), .B2(n22205), .ZN(
        n21928) );
  AOI22_X1 U23507 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n22213), .B2(n21940), .ZN(n21927) );
  OAI211_X1 U23508 ( .C1(n21943), .C2(n22210), .A(n21928), .B(n21927), .ZN(
        P1_U3123) );
  AOI22_X1 U23509 ( .A1(n22212), .A2(n21940), .B1(n21938), .B2(n22211), .ZN(
        n21930) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n21934), .ZN(n21929) );
  OAI211_X1 U23511 ( .C1(n22218), .C2(n21931), .A(n21930), .B(n21929), .ZN(
        P1_U3131) );
  AOI22_X1 U23512 ( .A1(n21939), .A2(n22220), .B1(n21938), .B2(n22219), .ZN(
        n21933) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n21940), .ZN(n21932) );
  OAI211_X1 U23514 ( .C1(n21943), .C2(n22224), .A(n21933), .B(n21932), .ZN(
        P1_U3139) );
  AOI22_X1 U23515 ( .A1(n21938), .A2(n22226), .B1(n21939), .B2(n22225), .ZN(
        n21936) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n21934), .ZN(n21935) );
  OAI211_X1 U23517 ( .C1(n21937), .C2(n22242), .A(n21936), .B(n21935), .ZN(
        P1_U3147) );
  AOI22_X1 U23518 ( .A1(n22236), .A2(n21939), .B1(n21938), .B2(n22233), .ZN(
        n21942) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n21940), .ZN(n21941) );
  OAI211_X1 U23520 ( .C1(n21943), .C2(n22242), .A(n21942), .B(n21941), .ZN(
        P1_U3155) );
  INV_X1 U23521 ( .A(n21983), .ZN(n21976) );
  OAI22_X2 U23522 ( .A1(n21945), .A2(n22134), .B1(n15824), .B2(n22136), .ZN(
        n21979) );
  INV_X1 U23523 ( .A(n22132), .ZN(n22038) );
  NAND2_X1 U23524 ( .A1(n22038), .A2(n21946), .ZN(n21968) );
  AOI22_X1 U23525 ( .A1(n22238), .A2(n21979), .B1(n21984), .B2(n22133), .ZN(
        n21949) );
  OAI22_X2 U23526 ( .A1(n15856), .A2(n22136), .B1(n21947), .B2(n22134), .ZN(
        n21985) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n21985), .ZN(n21948) );
  OAI211_X1 U23528 ( .C1(n22140), .C2(n21976), .A(n21949), .B(n21948), .ZN(
        P1_U3036) );
  INV_X1 U23529 ( .A(n21985), .ZN(n21982) );
  AOI22_X1 U23530 ( .A1(n22142), .A2(n21983), .B1(n21984), .B2(n22141), .ZN(
        n21951) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n21979), .ZN(n21950) );
  OAI211_X1 U23532 ( .C1(n21982), .C2(n22149), .A(n21951), .B(n21950), .ZN(
        P1_U3044) );
  AOI22_X1 U23533 ( .A1(n22156), .A2(n21985), .B1(n21984), .B2(n22091), .ZN(
        n21953) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22151), .B1(
        n22092), .B2(n21979), .ZN(n21952) );
  OAI211_X1 U23535 ( .C1(n22154), .C2(n21976), .A(n21953), .B(n21952), .ZN(
        P1_U3052) );
  AOI22_X1 U23536 ( .A1(n22163), .A2(n21985), .B1(n21984), .B2(n22155), .ZN(
        n21955) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22157), .B1(
        n22156), .B2(n21979), .ZN(n21954) );
  OAI211_X1 U23538 ( .C1(n22160), .C2(n21976), .A(n21955), .B(n21954), .ZN(
        P1_U3060) );
  AOI22_X1 U23539 ( .A1(n21984), .A2(n22162), .B1(n21983), .B2(n22161), .ZN(
        n21957) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n21979), .ZN(n21956) );
  OAI211_X1 U23541 ( .C1(n21982), .C2(n22172), .A(n21957), .B(n21956), .ZN(
        P1_U3068) );
  INV_X1 U23542 ( .A(n21979), .ZN(n21988) );
  AOI22_X1 U23543 ( .A1(n21984), .A2(n22167), .B1(n22168), .B2(n21983), .ZN(
        n21959) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n21985), .ZN(n21958) );
  OAI211_X1 U23545 ( .C1(n21988), .C2(n22172), .A(n21959), .B(n21958), .ZN(
        P1_U3076) );
  AOI22_X1 U23546 ( .A1(n22174), .A2(n21979), .B1(n21984), .B2(n22173), .ZN(
        n21961) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n21985), .ZN(n21960) );
  OAI211_X1 U23548 ( .C1(n22178), .C2(n21976), .A(n21961), .B(n21960), .ZN(
        P1_U3084) );
  AOI22_X1 U23549 ( .A1(n21984), .A2(n22179), .B1(n22180), .B2(n21983), .ZN(
        n21963) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n21979), .ZN(n21962) );
  OAI211_X1 U23551 ( .C1(n21982), .C2(n22185), .A(n21963), .B(n21962), .ZN(
        P1_U3092) );
  AOI22_X1 U23552 ( .A1(n21983), .A2(n22187), .B1(n21984), .B2(n22186), .ZN(
        n21965) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n21979), .ZN(n21964) );
  OAI211_X1 U23554 ( .C1(n21982), .C2(n22197), .A(n21965), .B(n21964), .ZN(
        P1_U3100) );
  AOI22_X1 U23555 ( .A1(n21983), .A2(n22193), .B1(n21984), .B2(n22192), .ZN(
        n21967) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n21985), .ZN(n21966) );
  OAI211_X1 U23557 ( .C1(n21988), .C2(n22197), .A(n21967), .B(n21966), .ZN(
        P1_U3108) );
  OAI22_X1 U23558 ( .A1(n22210), .A2(n21982), .B1(n21968), .B2(n22061), .ZN(
        n21969) );
  INV_X1 U23559 ( .A(n21969), .ZN(n21971) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22201), .B1(
        n22199), .B2(n21979), .ZN(n21970) );
  OAI211_X1 U23561 ( .C1(n22204), .C2(n21976), .A(n21971), .B(n21970), .ZN(
        P1_U3116) );
  AOI22_X1 U23562 ( .A1(n21984), .A2(n22205), .B1(n22206), .B2(n21983), .ZN(
        n21973) );
  AOI22_X1 U23563 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n22213), .B2(n21985), .ZN(n21972) );
  OAI211_X1 U23564 ( .C1(n21988), .C2(n22210), .A(n21973), .B(n21972), .ZN(
        P1_U3124) );
  AOI22_X1 U23565 ( .A1(n22212), .A2(n21985), .B1(n21984), .B2(n22211), .ZN(
        n21975) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n21979), .ZN(n21974) );
  OAI211_X1 U23567 ( .C1(n22218), .C2(n21976), .A(n21975), .B(n21974), .ZN(
        P1_U3132) );
  AOI22_X1 U23568 ( .A1(n21984), .A2(n22219), .B1(n22220), .B2(n21983), .ZN(
        n21978) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n21985), .ZN(n21977) );
  OAI211_X1 U23570 ( .C1(n21988), .C2(n22224), .A(n21978), .B(n21977), .ZN(
        P1_U3140) );
  AOI22_X1 U23571 ( .A1(n21984), .A2(n22226), .B1(n21983), .B2(n22225), .ZN(
        n21981) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n21979), .ZN(n21980) );
  OAI211_X1 U23573 ( .C1(n21982), .C2(n22242), .A(n21981), .B(n21980), .ZN(
        P1_U3148) );
  AOI22_X1 U23574 ( .A1(n21984), .A2(n22233), .B1(n22236), .B2(n21983), .ZN(
        n21987) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n21985), .ZN(n21986) );
  OAI211_X1 U23576 ( .C1(n21988), .C2(n22242), .A(n21987), .B(n21986), .ZN(
        P1_U3156) );
  INV_X1 U23577 ( .A(n22029), .ZN(n22022) );
  OAI22_X2 U23578 ( .A1(n21990), .A2(n22134), .B1(n15817), .B2(n22136), .ZN(
        n22025) );
  NAND2_X1 U23579 ( .A1(n22038), .A2(n21991), .ZN(n22014) );
  AOI22_X1 U23580 ( .A1(n22238), .A2(n22025), .B1(n22030), .B2(n22133), .ZN(
        n21995) );
  OAI22_X2 U23581 ( .A1(n21993), .A2(n22136), .B1(n21992), .B2(n22134), .ZN(
        n22031) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n22031), .ZN(n21994) );
  OAI211_X1 U23583 ( .C1(n22140), .C2(n22022), .A(n21995), .B(n21994), .ZN(
        P1_U3037) );
  INV_X1 U23584 ( .A(n22031), .ZN(n22028) );
  AOI22_X1 U23585 ( .A1(n22142), .A2(n22029), .B1(n22030), .B2(n22141), .ZN(
        n21997) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n22025), .ZN(n21996) );
  OAI211_X1 U23587 ( .C1(n22028), .C2(n22149), .A(n21997), .B(n21996), .ZN(
        P1_U3045) );
  AOI22_X1 U23588 ( .A1(n22156), .A2(n22031), .B1(n22030), .B2(n22091), .ZN(
        n21999) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22151), .B1(
        n22092), .B2(n22025), .ZN(n21998) );
  OAI211_X1 U23590 ( .C1(n22154), .C2(n22022), .A(n21999), .B(n21998), .ZN(
        P1_U3053) );
  AOI22_X1 U23591 ( .A1(n22163), .A2(n22031), .B1(n22030), .B2(n22155), .ZN(
        n22001) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22157), .B1(
        n22156), .B2(n22025), .ZN(n22000) );
  OAI211_X1 U23593 ( .C1(n22160), .C2(n22022), .A(n22001), .B(n22000), .ZN(
        P1_U3061) );
  AOI22_X1 U23594 ( .A1(n22030), .A2(n22162), .B1(n22029), .B2(n22161), .ZN(
        n22003) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n22025), .ZN(n22002) );
  OAI211_X1 U23596 ( .C1(n22028), .C2(n22172), .A(n22003), .B(n22002), .ZN(
        P1_U3069) );
  INV_X1 U23597 ( .A(n22025), .ZN(n22034) );
  AOI22_X1 U23598 ( .A1(n22030), .A2(n22167), .B1(n22168), .B2(n22029), .ZN(
        n22005) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n22031), .ZN(n22004) );
  OAI211_X1 U23600 ( .C1(n22034), .C2(n22172), .A(n22005), .B(n22004), .ZN(
        P1_U3077) );
  AOI22_X1 U23601 ( .A1(n22174), .A2(n22025), .B1(n22030), .B2(n22173), .ZN(
        n22007) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22031), .ZN(n22006) );
  OAI211_X1 U23603 ( .C1(n22178), .C2(n22022), .A(n22007), .B(n22006), .ZN(
        P1_U3085) );
  AOI22_X1 U23604 ( .A1(n22030), .A2(n22179), .B1(n22180), .B2(n22029), .ZN(
        n22009) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n22025), .ZN(n22008) );
  OAI211_X1 U23606 ( .C1(n22028), .C2(n22185), .A(n22009), .B(n22008), .ZN(
        P1_U3093) );
  AOI22_X1 U23607 ( .A1(n22029), .A2(n22187), .B1(n22030), .B2(n22186), .ZN(
        n22011) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n22025), .ZN(n22010) );
  OAI211_X1 U23609 ( .C1(n22028), .C2(n22197), .A(n22011), .B(n22010), .ZN(
        P1_U3101) );
  AOI22_X1 U23610 ( .A1(n22029), .A2(n22193), .B1(n22030), .B2(n22192), .ZN(
        n22013) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n22031), .ZN(n22012) );
  OAI211_X1 U23612 ( .C1(n22034), .C2(n22197), .A(n22013), .B(n22012), .ZN(
        P1_U3109) );
  OAI22_X1 U23613 ( .A1(n22210), .A2(n22028), .B1(n22014), .B2(n22061), .ZN(
        n22015) );
  INV_X1 U23614 ( .A(n22015), .ZN(n22017) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22201), .B1(
        n22199), .B2(n22025), .ZN(n22016) );
  OAI211_X1 U23616 ( .C1(n22204), .C2(n22022), .A(n22017), .B(n22016), .ZN(
        P1_U3117) );
  AOI22_X1 U23617 ( .A1(n22030), .A2(n22205), .B1(n22206), .B2(n22029), .ZN(
        n22019) );
  AOI22_X1 U23618 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n22213), .B2(n22031), .ZN(n22018) );
  OAI211_X1 U23619 ( .C1(n22034), .C2(n22210), .A(n22019), .B(n22018), .ZN(
        P1_U3125) );
  AOI22_X1 U23620 ( .A1(n22212), .A2(n22031), .B1(n22030), .B2(n22211), .ZN(
        n22021) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n22025), .ZN(n22020) );
  OAI211_X1 U23622 ( .C1(n22218), .C2(n22022), .A(n22021), .B(n22020), .ZN(
        P1_U3133) );
  AOI22_X1 U23623 ( .A1(n22030), .A2(n22219), .B1(n22220), .B2(n22029), .ZN(
        n22024) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n22031), .ZN(n22023) );
  OAI211_X1 U23625 ( .C1(n22034), .C2(n22224), .A(n22024), .B(n22023), .ZN(
        P1_U3141) );
  AOI22_X1 U23626 ( .A1(n22030), .A2(n22226), .B1(n22029), .B2(n22225), .ZN(
        n22027) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n22025), .ZN(n22026) );
  OAI211_X1 U23628 ( .C1(n22028), .C2(n22242), .A(n22027), .B(n22026), .ZN(
        P1_U3149) );
  AOI22_X1 U23629 ( .A1(n22030), .A2(n22233), .B1(n22236), .B2(n22029), .ZN(
        n22033) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n22031), .ZN(n22032) );
  OAI211_X1 U23631 ( .C1(n22034), .C2(n22242), .A(n22033), .B(n22032), .ZN(
        P1_U3157) );
  INV_X1 U23632 ( .A(n22077), .ZN(n22070) );
  OAI22_X2 U23633 ( .A1(n22036), .A2(n22134), .B1(n15810), .B2(n22136), .ZN(
        n22073) );
  NAND2_X1 U23634 ( .A1(n22038), .A2(n22037), .ZN(n22062) );
  AOI22_X1 U23635 ( .A1(n22238), .A2(n22073), .B1(n22078), .B2(n22133), .ZN(
        n22041) );
  OAI22_X2 U23636 ( .A1(n15850), .A2(n22136), .B1(n22039), .B2(n22134), .ZN(
        n22079) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n22079), .ZN(n22040) );
  OAI211_X1 U23638 ( .C1(n22140), .C2(n22070), .A(n22041), .B(n22040), .ZN(
        P1_U3038) );
  INV_X1 U23639 ( .A(n22079), .ZN(n22076) );
  AOI22_X1 U23640 ( .A1(n22142), .A2(n22077), .B1(n22078), .B2(n22141), .ZN(
        n22043) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n22073), .ZN(n22042) );
  OAI211_X1 U23642 ( .C1(n22076), .C2(n22149), .A(n22043), .B(n22042), .ZN(
        P1_U3046) );
  INV_X1 U23643 ( .A(n22073), .ZN(n22082) );
  OAI22_X1 U23644 ( .A1(n22149), .A2(n22082), .B1(n22062), .B2(n22147), .ZN(
        n22044) );
  INV_X1 U23645 ( .A(n22044), .ZN(n22046) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22151), .B1(
        n22156), .B2(n22079), .ZN(n22045) );
  OAI211_X1 U23647 ( .C1(n22154), .C2(n22070), .A(n22046), .B(n22045), .ZN(
        P1_U3054) );
  AOI22_X1 U23648 ( .A1(n22156), .A2(n22073), .B1(n22078), .B2(n22155), .ZN(
        n22048) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22157), .B1(
        n22163), .B2(n22079), .ZN(n22047) );
  OAI211_X1 U23650 ( .C1(n22160), .C2(n22070), .A(n22048), .B(n22047), .ZN(
        P1_U3062) );
  AOI22_X1 U23651 ( .A1(n22078), .A2(n22162), .B1(n22077), .B2(n22161), .ZN(
        n22050) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n22073), .ZN(n22049) );
  OAI211_X1 U23653 ( .C1(n22076), .C2(n22172), .A(n22050), .B(n22049), .ZN(
        P1_U3070) );
  AOI22_X1 U23654 ( .A1(n22078), .A2(n22167), .B1(n22168), .B2(n22077), .ZN(
        n22052) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n22079), .ZN(n22051) );
  OAI211_X1 U23656 ( .C1(n22082), .C2(n22172), .A(n22052), .B(n22051), .ZN(
        P1_U3078) );
  AOI22_X1 U23657 ( .A1(n22181), .A2(n22079), .B1(n22078), .B2(n22173), .ZN(
        n22054) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22175), .B1(
        n22174), .B2(n22073), .ZN(n22053) );
  OAI211_X1 U23659 ( .C1(n22178), .C2(n22070), .A(n22054), .B(n22053), .ZN(
        P1_U3086) );
  AOI22_X1 U23660 ( .A1(n22078), .A2(n22179), .B1(n22180), .B2(n22077), .ZN(
        n22056) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n22073), .ZN(n22055) );
  OAI211_X1 U23662 ( .C1(n22076), .C2(n22185), .A(n22056), .B(n22055), .ZN(
        P1_U3094) );
  AOI22_X1 U23663 ( .A1(n22077), .A2(n22187), .B1(n22078), .B2(n22186), .ZN(
        n22058) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n22073), .ZN(n22057) );
  OAI211_X1 U23665 ( .C1(n22076), .C2(n22197), .A(n22058), .B(n22057), .ZN(
        P1_U3102) );
  AOI22_X1 U23666 ( .A1(n22077), .A2(n22193), .B1(n22078), .B2(n22192), .ZN(
        n22060) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n22079), .ZN(n22059) );
  OAI211_X1 U23668 ( .C1(n22082), .C2(n22197), .A(n22060), .B(n22059), .ZN(
        P1_U3110) );
  OAI22_X1 U23669 ( .A1(n22210), .A2(n22076), .B1(n22062), .B2(n22061), .ZN(
        n22063) );
  INV_X1 U23670 ( .A(n22063), .ZN(n22065) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22201), .B1(
        n22199), .B2(n22073), .ZN(n22064) );
  OAI211_X1 U23672 ( .C1(n22204), .C2(n22070), .A(n22065), .B(n22064), .ZN(
        P1_U3118) );
  AOI22_X1 U23673 ( .A1(n22078), .A2(n22205), .B1(n22206), .B2(n22077), .ZN(
        n22067) );
  AOI22_X1 U23674 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n22213), .B2(n22079), .ZN(n22066) );
  OAI211_X1 U23675 ( .C1(n22082), .C2(n22210), .A(n22067), .B(n22066), .ZN(
        P1_U3126) );
  AOI22_X1 U23676 ( .A1(n22212), .A2(n22079), .B1(n22078), .B2(n22211), .ZN(
        n22069) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n22073), .ZN(n22068) );
  OAI211_X1 U23678 ( .C1(n22218), .C2(n22070), .A(n22069), .B(n22068), .ZN(
        P1_U3134) );
  AOI22_X1 U23679 ( .A1(n22078), .A2(n22219), .B1(n22220), .B2(n22077), .ZN(
        n22072) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n22079), .ZN(n22071) );
  OAI211_X1 U23681 ( .C1(n22082), .C2(n22224), .A(n22072), .B(n22071), .ZN(
        P1_U3142) );
  AOI22_X1 U23682 ( .A1(n22078), .A2(n22226), .B1(n22077), .B2(n22225), .ZN(
        n22075) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n22073), .ZN(n22074) );
  OAI211_X1 U23684 ( .C1(n22076), .C2(n22242), .A(n22075), .B(n22074), .ZN(
        P1_U3150) );
  AOI22_X1 U23685 ( .A1(n22078), .A2(n22233), .B1(n22236), .B2(n22077), .ZN(
        n22081) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n22079), .ZN(n22080) );
  OAI211_X1 U23687 ( .C1(n22082), .C2(n22242), .A(n22081), .B(n22080), .ZN(
        P1_U3158) );
  OAI22_X2 U23688 ( .A1(n22084), .A2(n22134), .B1(n15804), .B2(n22136), .ZN(
        n22118) );
  NOR2_X2 U23689 ( .A1(n22132), .A2(n11656), .ZN(n22122) );
  AOI22_X1 U23690 ( .A1(n22238), .A2(n22118), .B1(n22122), .B2(n22133), .ZN(
        n22088) );
  OAI22_X2 U23691 ( .A1(n22086), .A2(n22136), .B1(n22085), .B2(n22134), .ZN(
        n22124) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n22124), .ZN(n22087) );
  OAI211_X1 U23693 ( .C1(n22140), .C2(n22115), .A(n22088), .B(n22087), .ZN(
        P1_U3039) );
  INV_X1 U23694 ( .A(n22124), .ZN(n22121) );
  AOI22_X1 U23695 ( .A1(n22142), .A2(n22123), .B1(n22122), .B2(n22141), .ZN(
        n22090) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n22118), .ZN(n22089) );
  OAI211_X1 U23697 ( .C1(n22121), .C2(n22149), .A(n22090), .B(n22089), .ZN(
        P1_U3047) );
  AOI22_X1 U23698 ( .A1(n22156), .A2(n22124), .B1(n22122), .B2(n22091), .ZN(
        n22094) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22151), .B1(
        n22092), .B2(n22118), .ZN(n22093) );
  OAI211_X1 U23700 ( .C1(n22154), .C2(n22115), .A(n22094), .B(n22093), .ZN(
        P1_U3055) );
  AOI22_X1 U23701 ( .A1(n22163), .A2(n22124), .B1(n22122), .B2(n22155), .ZN(
        n22096) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22157), .B1(
        n22156), .B2(n22118), .ZN(n22095) );
  OAI211_X1 U23703 ( .C1(n22160), .C2(n22115), .A(n22096), .B(n22095), .ZN(
        P1_U3063) );
  AOI22_X1 U23704 ( .A1(n22122), .A2(n22162), .B1(n22123), .B2(n22161), .ZN(
        n22098) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n22118), .ZN(n22097) );
  OAI211_X1 U23706 ( .C1(n22121), .C2(n22172), .A(n22098), .B(n22097), .ZN(
        P1_U3071) );
  INV_X1 U23707 ( .A(n22118), .ZN(n22127) );
  AOI22_X1 U23708 ( .A1(n22123), .A2(n22168), .B1(n22122), .B2(n22167), .ZN(
        n22100) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n22124), .ZN(n22099) );
  OAI211_X1 U23710 ( .C1(n22127), .C2(n22172), .A(n22100), .B(n22099), .ZN(
        P1_U3079) );
  AOI22_X1 U23711 ( .A1(n22174), .A2(n22118), .B1(n22173), .B2(n22122), .ZN(
        n22102) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22175), .B1(
        n22181), .B2(n22124), .ZN(n22101) );
  OAI211_X1 U23713 ( .C1(n22178), .C2(n22115), .A(n22102), .B(n22101), .ZN(
        P1_U3087) );
  AOI22_X1 U23714 ( .A1(n22180), .A2(n22123), .B1(n22122), .B2(n22179), .ZN(
        n22104) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n22118), .ZN(n22103) );
  OAI211_X1 U23716 ( .C1(n22121), .C2(n22185), .A(n22104), .B(n22103), .ZN(
        P1_U3095) );
  AOI22_X1 U23717 ( .A1(n22187), .A2(n22123), .B1(n22122), .B2(n22186), .ZN(
        n22106) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n22118), .ZN(n22105) );
  OAI211_X1 U23719 ( .C1(n22121), .C2(n22197), .A(n22106), .B(n22105), .ZN(
        P1_U3103) );
  AOI22_X1 U23720 ( .A1(n22193), .A2(n22123), .B1(n22122), .B2(n22192), .ZN(
        n22108) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n22124), .ZN(n22107) );
  OAI211_X1 U23722 ( .C1(n22127), .C2(n22197), .A(n22108), .B(n22107), .ZN(
        P1_U3111) );
  AOI22_X1 U23723 ( .A1(n22199), .A2(n22118), .B1(n22122), .B2(n22198), .ZN(
        n22110) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22201), .B1(
        n22200), .B2(n22124), .ZN(n22109) );
  OAI211_X1 U23725 ( .C1(n22204), .C2(n22115), .A(n22110), .B(n22109), .ZN(
        P1_U3119) );
  AOI22_X1 U23726 ( .A1(n22123), .A2(n22206), .B1(n22122), .B2(n22205), .ZN(
        n22112) );
  AOI22_X1 U23727 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n22213), .B2(n22124), .ZN(n22111) );
  OAI211_X1 U23728 ( .C1(n22127), .C2(n22210), .A(n22112), .B(n22111), .ZN(
        P1_U3127) );
  AOI22_X1 U23729 ( .A1(n22212), .A2(n22124), .B1(n22122), .B2(n22211), .ZN(
        n22114) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n22118), .ZN(n22113) );
  OAI211_X1 U23731 ( .C1(n22218), .C2(n22115), .A(n22114), .B(n22113), .ZN(
        P1_U3135) );
  AOI22_X1 U23732 ( .A1(n22123), .A2(n22220), .B1(n22122), .B2(n22219), .ZN(
        n22117) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n22124), .ZN(n22116) );
  OAI211_X1 U23734 ( .C1(n22127), .C2(n22224), .A(n22117), .B(n22116), .ZN(
        P1_U3143) );
  AOI22_X1 U23735 ( .A1(n22122), .A2(n22226), .B1(n22123), .B2(n22225), .ZN(
        n22120) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n22118), .ZN(n22119) );
  OAI211_X1 U23737 ( .C1(n22121), .C2(n22242), .A(n22120), .B(n22119), .ZN(
        P1_U3151) );
  AOI22_X1 U23738 ( .A1(n22236), .A2(n22123), .B1(n22122), .B2(n22233), .ZN(
        n22126) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n22124), .ZN(n22125) );
  OAI211_X1 U23740 ( .C1(n22127), .C2(n22242), .A(n22126), .B(n22125), .ZN(
        P1_U3159) );
  INV_X1 U23741 ( .A(n22235), .ZN(n22217) );
  OAI22_X2 U23742 ( .A1(n12410), .A2(n22136), .B1(n22130), .B2(n22134), .ZN(
        n22227) );
  NOR2_X2 U23743 ( .A1(n22132), .A2(n22131), .ZN(n22234) );
  AOI22_X1 U23744 ( .A1(n22238), .A2(n22227), .B1(n22234), .B2(n22133), .ZN(
        n22139) );
  OAI22_X2 U23745 ( .A1(n15845), .A2(n22136), .B1(n22135), .B2(n22134), .ZN(
        n22237) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22137), .B1(
        n22143), .B2(n22237), .ZN(n22138) );
  OAI211_X1 U23747 ( .C1(n22140), .C2(n22217), .A(n22139), .B(n22138), .ZN(
        P1_U3040) );
  INV_X1 U23748 ( .A(n22237), .ZN(n22232) );
  AOI22_X1 U23749 ( .A1(n22142), .A2(n22235), .B1(n22234), .B2(n22141), .ZN(
        n22146) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22144), .B1(
        n22143), .B2(n22227), .ZN(n22145) );
  OAI211_X1 U23751 ( .C1(n22232), .C2(n22149), .A(n22146), .B(n22145), .ZN(
        P1_U3048) );
  INV_X1 U23752 ( .A(n22227), .ZN(n22243) );
  INV_X1 U23753 ( .A(n22234), .ZN(n22148) );
  OAI22_X1 U23754 ( .A1(n22149), .A2(n22243), .B1(n22148), .B2(n22147), .ZN(
        n22150) );
  INV_X1 U23755 ( .A(n22150), .ZN(n22153) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22151), .B1(
        n22156), .B2(n22237), .ZN(n22152) );
  OAI211_X1 U23757 ( .C1(n22154), .C2(n22217), .A(n22153), .B(n22152), .ZN(
        P1_U3056) );
  AOI22_X1 U23758 ( .A1(n22163), .A2(n22237), .B1(n22234), .B2(n22155), .ZN(
        n22159) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22157), .B1(
        n22156), .B2(n22227), .ZN(n22158) );
  OAI211_X1 U23760 ( .C1(n22160), .C2(n22217), .A(n22159), .B(n22158), .ZN(
        P1_U3064) );
  AOI22_X1 U23761 ( .A1(n22234), .A2(n22162), .B1(n22235), .B2(n22161), .ZN(
        n22166) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22164), .B1(
        n22163), .B2(n22227), .ZN(n22165) );
  OAI211_X1 U23763 ( .C1(n22232), .C2(n22172), .A(n22166), .B(n22165), .ZN(
        P1_U3072) );
  AOI22_X1 U23764 ( .A1(n22235), .A2(n22168), .B1(n22234), .B2(n22167), .ZN(
        n22171) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22169), .B1(
        n22174), .B2(n22237), .ZN(n22170) );
  OAI211_X1 U23766 ( .C1(n22243), .C2(n22172), .A(n22171), .B(n22170), .ZN(
        P1_U3080) );
  AOI22_X1 U23767 ( .A1(n22181), .A2(n22237), .B1(n22173), .B2(n22234), .ZN(
        n22177) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22175), .B1(
        n22174), .B2(n22227), .ZN(n22176) );
  OAI211_X1 U23769 ( .C1(n22178), .C2(n22217), .A(n22177), .B(n22176), .ZN(
        P1_U3088) );
  AOI22_X1 U23770 ( .A1(n22180), .A2(n22235), .B1(n22234), .B2(n22179), .ZN(
        n22184) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22182), .B1(
        n22181), .B2(n22227), .ZN(n22183) );
  OAI211_X1 U23772 ( .C1(n22232), .C2(n22185), .A(n22184), .B(n22183), .ZN(
        P1_U3096) );
  AOI22_X1 U23773 ( .A1(n22187), .A2(n22235), .B1(n22234), .B2(n22186), .ZN(
        n22191) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22189), .B1(
        n22188), .B2(n22227), .ZN(n22190) );
  OAI211_X1 U23775 ( .C1(n22232), .C2(n22197), .A(n22191), .B(n22190), .ZN(
        P1_U3104) );
  AOI22_X1 U23776 ( .A1(n22193), .A2(n22235), .B1(n22234), .B2(n22192), .ZN(
        n22196) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22194), .B1(
        n22199), .B2(n22237), .ZN(n22195) );
  OAI211_X1 U23778 ( .C1(n22243), .C2(n22197), .A(n22196), .B(n22195), .ZN(
        P1_U3112) );
  AOI22_X1 U23779 ( .A1(n22199), .A2(n22227), .B1(n22234), .B2(n22198), .ZN(
        n22203) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22201), .B1(
        n22200), .B2(n22237), .ZN(n22202) );
  OAI211_X1 U23781 ( .C1(n22204), .C2(n22217), .A(n22203), .B(n22202), .ZN(
        P1_U3120) );
  AOI22_X1 U23782 ( .A1(n22235), .A2(n22206), .B1(n22234), .B2(n22205), .ZN(
        n22209) );
  AOI22_X1 U23783 ( .A1(n22207), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n22213), .B2(n22237), .ZN(n22208) );
  OAI211_X1 U23784 ( .C1(n22243), .C2(n22210), .A(n22209), .B(n22208), .ZN(
        P1_U3128) );
  AOI22_X1 U23785 ( .A1(n22212), .A2(n22237), .B1(n22234), .B2(n22211), .ZN(
        n22216) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22214), .B1(
        n22213), .B2(n22227), .ZN(n22215) );
  OAI211_X1 U23787 ( .C1(n22218), .C2(n22217), .A(n22216), .B(n22215), .ZN(
        P1_U3136) );
  AOI22_X1 U23788 ( .A1(n22235), .A2(n22220), .B1(n22234), .B2(n22219), .ZN(
        n22223) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22221), .B1(
        n22228), .B2(n22237), .ZN(n22222) );
  OAI211_X1 U23790 ( .C1(n22243), .C2(n22224), .A(n22223), .B(n22222), .ZN(
        P1_U3144) );
  AOI22_X1 U23791 ( .A1(n22234), .A2(n22226), .B1(n22235), .B2(n22225), .ZN(
        n22231) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22229), .B1(
        n22228), .B2(n22227), .ZN(n22230) );
  OAI211_X1 U23793 ( .C1(n22232), .C2(n22242), .A(n22231), .B(n22230), .ZN(
        P1_U3152) );
  AOI22_X1 U23794 ( .A1(n22236), .A2(n22235), .B1(n22234), .B2(n22233), .ZN(
        n22241) );
  AOI22_X1 U23795 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22239), .B1(
        n22238), .B2(n22237), .ZN(n22240) );
  OAI211_X1 U23796 ( .C1(n22243), .C2(n22242), .A(n22241), .B(n22240), .ZN(
        P1_U3160) );
  AOI22_X1 U23797 ( .A1(n22246), .A2(n22245), .B1(n22244), .B2(n19831), .ZN(
        P1_U3486) );
  BUF_X1 U11354 ( .A(n15076), .Z(n17722) );
  CLKBUF_X3 U11193 ( .A(n15208), .Z(n10977) );
  CLKBUF_X1 U11083 ( .A(n12967), .Z(n10974) );
  NOR2_X2 U11386 ( .A1(n20713), .A2(n15040), .ZN(n15079) );
  BUF_X2 U11085 ( .A(n15065), .Z(n17723) );
  MUX2_X1 U11102 ( .A(n12335), .B(n11634), .S(n11633), .Z(n11635) );
  NAND2_X1 U11108 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20680), .ZN(
        n15041) );
  CLKBUF_X1 U11120 ( .A(n12967), .Z(n10975) );
  NAND2_X2 U11127 ( .A1(n21138), .A2(n21142), .ZN(n21085) );
  CLKBUF_X1 U11153 ( .A(n12967), .Z(n10973) );
  CLKBUF_X1 U11155 ( .A(n18557), .Z(n10997) );
  CLKBUF_X1 U11163 ( .A(n15065), .Z(n17741) );
  XNOR2_X1 U11171 ( .A(n17806), .B(n17807), .ZN(n18176) );
  CLKBUF_X1 U11351 ( .A(n17358), .Z(n17369) );
  CLKBUF_X1 U12255 ( .A(n12516), .Z(n15436) );
endmodule

