

module b14_C_AntiSAT_k_256_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047;

  INV_X2 U2486 ( .A(n4290), .ZN(n5040) );
  INV_X2 U2487 ( .A(n3687), .ZN(n3676) );
  INV_X1 U2488 ( .A(n2993), .ZN(n3144) );
  NAND2_X2 U2489 ( .A1(n2495), .A2(n2494), .ZN(n2725) );
  INV_X1 U2490 ( .A(n3689), .ZN(n3058) );
  INV_X1 U2491 ( .A(n3671), .ZN(n3686) );
  NAND2_X1 U2492 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  XNOR2_X2 U2493 ( .A(n4034), .B(n4048), .ZN(n4531) );
  NAND2_X2 U2494 ( .A1(n4522), .A2(n4033), .ZN(n4034) );
  OAI22_X2 U2495 ( .A1(n3622), .A2(n3621), .B1(n3620), .B2(n3619), .ZN(n3754)
         );
  XNOR2_X2 U2496 ( .A(n2492), .B(IR_REG_30__SCAN_IN), .ZN(n2493) );
  INV_X1 U2497 ( .A(n3997), .ZN(n3161) );
  OAI21_X1 U2499 ( .B1(n4135), .B2(n2270), .A(n2753), .ZN(n4115) );
  NOR2_X1 U2500 ( .A1(n4532), .A2(n4035), .ZN(n4544) );
  AND2_X1 U2501 ( .A1(n2386), .A2(n2385), .ZN(n4139) );
  NAND2_X1 U2502 ( .A1(n3835), .A2(n3483), .ZN(n3511) );
  NAND2_X1 U2503 ( .A1(n2384), .A2(n3946), .ZN(n3835) );
  NAND2_X1 U2504 ( .A1(n4551), .A2(n3943), .ZN(n2384) );
  NAND2_X1 U2505 ( .A1(n2429), .A2(n3924), .ZN(n3303) );
  NAND2_X1 U2506 ( .A1(n4468), .A2(n3321), .ZN(n4481) );
  NAND2_X1 U2507 ( .A1(n4469), .A2(REG1_REG_8__SCAN_IN), .ZN(n4468) );
  XNOR2_X1 U2508 ( .A(n3320), .B(n4472), .ZN(n4469) );
  NAND2_X1 U2509 ( .A1(n3118), .A2(n2520), .ZN(n3169) );
  OAI21_X1 U2510 ( .B1(n2383), .B2(n4452), .A(REG1_REG_7__SCAN_IN), .ZN(n2382)
         );
  NOR2_X1 U2511 ( .A1(n3886), .A2(n2530), .ZN(n2544) );
  NAND2_X1 U2512 ( .A1(n3919), .A2(n3916), .ZN(n3886) );
  NOR2_X1 U2513 ( .A1(n2944), .A2(n2959), .ZN(n3319) );
  AND4_X1 U2514 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n3068)
         );
  NAND4_X1 U2515 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .ZN(n3141)
         );
  AND4_X1 U2516 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .ZN(n3709)
         );
  NAND4_X1 U2517 ( .A1(n2537), .A2(n2536), .A3(n2535), .A4(n2534), .ZN(n3997)
         );
  INV_X1 U2518 ( .A(n2966), .ZN(n2309) );
  NAND2_X2 U2519 ( .A1(n2966), .A2(n2988), .ZN(n3687) );
  NAND2_X1 U2520 ( .A1(n3022), .A2(n2257), .ZN(n4019) );
  XNOR2_X1 U2521 ( .A(n2834), .B(IR_REG_24__SCAN_IN), .ZN(n2840) );
  OAI21_X1 U2522 ( .B1(n2352), .B2(n2529), .A(n2351), .ZN(n3140) );
  NAND2_X1 U2523 ( .A1(n2843), .A2(IR_REG_31__SCAN_IN), .ZN(n2834) );
  XNOR2_X1 U2524 ( .A(n2836), .B(IR_REG_26__SCAN_IN), .ZN(n2901) );
  AOI21_X1 U2525 ( .B1(n2684), .B2(IR_REG_31__SCAN_IN), .A(n2316), .ZN(n2315)
         );
  OR2_X1 U2526 ( .A1(n2829), .A2(n2490), .ZN(n2836) );
  AND2_X1 U2527 ( .A1(n2635), .A2(n2637), .ZN(n2682) );
  NAND2_X1 U2528 ( .A1(n2317), .A2(n4772), .ZN(n2316) );
  NAND2_X1 U2529 ( .A1(n2318), .A2(IR_REG_31__SCAN_IN), .ZN(n2317) );
  INV_X1 U2530 ( .A(IR_REG_3__SCAN_IN), .ZN(n2538) );
  NOR2_X1 U2531 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2356)
         );
  NOR2_X1 U2532 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2355)
         );
  AND3_X1 U2533 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2557) );
  XNOR2_X2 U2534 ( .A(n2778), .B(n4838), .ZN(n2782) );
  AND2_X4 U2535 ( .A1(n2493), .A2(n2494), .ZN(n2522) );
  NAND2_X1 U2536 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2505) );
  NOR2_X1 U2537 ( .A1(n2338), .A2(n2959), .ZN(n2337) );
  AND3_X1 U2538 ( .A1(n2680), .A2(n4889), .A3(n2679), .ZN(n2681) );
  INV_X1 U2539 ( .A(IR_REG_16__SCAN_IN), .ZN(n2679) );
  AND2_X1 U2540 ( .A1(n2463), .A2(n3288), .ZN(n2303) );
  OR2_X1 U2541 ( .A1(n3689), .A2(n4638), .ZN(n3671) );
  AND2_X1 U2542 ( .A1(n3692), .A2(n4092), .ZN(n3844) );
  INV_X1 U2543 ( .A(n2293), .ZN(n2292) );
  OAI21_X1 U2544 ( .B1(n2253), .B2(n2294), .A(n2707), .ZN(n2293) );
  OAI22_X1 U2545 ( .A1(n2404), .A2(n2403), .B1(n3404), .B2(n3413), .ZN(n2396)
         );
  OAI21_X1 U2546 ( .B1(n3210), .B2(n3209), .A(n3934), .ZN(n3275) );
  AND2_X1 U2547 ( .A1(n2244), .A2(n2296), .ZN(n2295) );
  INV_X1 U2548 ( .A(IR_REG_25__SCAN_IN), .ZN(n2296) );
  AND2_X1 U2549 ( .A1(n2485), .A2(n2486), .ZN(n2473) );
  INV_X1 U2550 ( .A(IR_REG_21__SCAN_IN), .ZN(n2486) );
  AOI21_X1 U2551 ( .B1(n2463), .B2(n2466), .A(n2307), .ZN(n2306) );
  INV_X1 U2552 ( .A(n3243), .ZN(n2307) );
  NOR2_X1 U2553 ( .A1(n2459), .A2(n2474), .ZN(n2458) );
  INV_X1 U2554 ( .A(n3797), .ZN(n2459) );
  NOR2_X1 U2555 ( .A1(n4428), .A2(n2334), .ZN(n2331) );
  NAND2_X1 U2556 ( .A1(n4474), .A2(n4475), .ZN(n4473) );
  NAND2_X1 U2557 ( .A1(n2344), .A2(n2343), .ZN(n2346) );
  OR2_X1 U2558 ( .A1(n3471), .A2(n4427), .ZN(n2344) );
  AND2_X1 U2559 ( .A1(n2347), .A2(n4426), .ZN(n2343) );
  NAND2_X1 U2560 ( .A1(n2285), .A2(n2282), .ZN(n4135) );
  AOI21_X1 U2561 ( .B1(n2283), .B2(n2287), .A(n2269), .ZN(n2282) );
  NAND2_X1 U2562 ( .A1(n4172), .A2(n2286), .ZN(n2285) );
  NOR2_X1 U2563 ( .A1(n2745), .A2(n2284), .ZN(n2283) );
  NAND2_X1 U2564 ( .A1(n3369), .A2(n3298), .ZN(n2584) );
  AND2_X1 U2565 ( .A1(n2408), .A2(n2407), .ZN(n3229) );
  NOR2_X1 U2566 ( .A1(n3996), .A2(n3215), .ZN(n2410) );
  NAND2_X1 U2567 ( .A1(n2301), .A2(n2299), .ZN(n2494) );
  NOR2_X1 U2568 ( .A1(n2491), .A2(n2300), .ZN(n2299) );
  OAI21_X1 U2569 ( .B1(n2823), .B2(IR_REG_28__SCAN_IN), .A(n2271), .ZN(n2301)
         );
  NOR2_X1 U2570 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2300)
         );
  NOR2_X1 U2571 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2358)
         );
  NOR2_X1 U2572 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2357)
         );
  AND2_X1 U2573 ( .A1(n2333), .A2(n2336), .ZN(n2332) );
  NAND2_X1 U2574 ( .A1(n2959), .A2(n2338), .ZN(n2336) );
  INV_X1 U2575 ( .A(n2337), .ZN(n2335) );
  INV_X1 U2576 ( .A(n3608), .ZN(n2325) );
  INV_X1 U2577 ( .A(n2699), .ZN(n2294) );
  INV_X1 U2578 ( .A(IR_REG_6__SCAN_IN), .ZN(n2594) );
  INV_X1 U2579 ( .A(n3778), .ZN(n2312) );
  OR2_X1 U2580 ( .A1(n3606), .A2(n2325), .ZN(n2322) );
  NAND2_X1 U2581 ( .A1(n2325), .A2(n3606), .ZN(n2324) );
  NAND2_X1 U2582 ( .A1(n2941), .A2(n2940), .ZN(n2942) );
  AND2_X1 U2583 ( .A1(n4018), .A2(n2379), .ZN(n2944) );
  NAND2_X1 U2584 ( .A1(n4429), .A2(REG1_REG_5__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U2585 ( .A1(n3341), .A2(n4458), .ZN(n3342) );
  NAND2_X1 U2586 ( .A1(n4139), .A2(n2814), .ZN(n4117) );
  AND2_X1 U2587 ( .A1(n4141), .A2(n4160), .ZN(n2745) );
  AND2_X1 U2588 ( .A1(n3899), .A2(n4155), .ZN(n3958) );
  NAND2_X1 U2589 ( .A1(n2813), .A2(n2812), .ZN(n4156) );
  NAND2_X1 U2590 ( .A1(n2292), .A2(n2294), .ZN(n2291) );
  OR2_X1 U2591 ( .A1(n2564), .A2(n2410), .ZN(n2406) );
  AOI21_X1 U2592 ( .B1(n2873), .B2(n2872), .A(n3844), .ZN(n2438) );
  AND2_X1 U2593 ( .A1(n4197), .A2(n2250), .ZN(n2371) );
  NAND2_X1 U2594 ( .A1(n4354), .A2(n3609), .ZN(n2369) );
  NAND2_X1 U2595 ( .A1(n3582), .A2(n3384), .ZN(n2361) );
  OR2_X1 U2596 ( .A1(n3312), .A2(n3371), .ZN(n3311) );
  INV_X1 U2597 ( .A(IR_REG_23__SCAN_IN), .ZN(n2833) );
  NAND2_X1 U2598 ( .A1(n2832), .A2(IR_REG_31__SCAN_IN), .ZN(n2841) );
  NOR2_X1 U2599 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2481)
         );
  INV_X1 U2600 ( .A(IR_REG_15__SCAN_IN), .ZN(n4889) );
  INV_X1 U2601 ( .A(IR_REG_2__SCAN_IN), .ZN(n2302) );
  NAND2_X1 U2602 ( .A1(n2260), .A2(n3238), .ZN(n2463) );
  INV_X1 U2603 ( .A(n3190), .ZN(n2467) );
  INV_X1 U2604 ( .A(n3185), .ZN(n2466) );
  INV_X1 U2605 ( .A(n2267), .ZN(n2443) );
  AND2_X1 U2606 ( .A1(n3625), .A2(n3624), .ZN(n3755) );
  NAND2_X1 U2607 ( .A1(n2470), .A2(n2468), .ZN(n3400) );
  NOR2_X1 U2608 ( .A1(n3368), .A2(n2469), .ZN(n2468) );
  INV_X1 U2609 ( .A(n2471), .ZN(n2469) );
  NOR2_X1 U2610 ( .A1(n2455), .A2(n2456), .ZN(n2453) );
  NOR2_X1 U2611 ( .A1(n3728), .A2(n2457), .ZN(n2456) );
  NOR2_X1 U2612 ( .A1(n3754), .A2(n2264), .ZN(n2461) );
  NAND2_X1 U2613 ( .A1(n3186), .A2(n3185), .ZN(n2465) );
  AND2_X1 U2614 ( .A1(n3982), .A2(n4423), .ZN(n2979) );
  AND2_X1 U2615 ( .A1(n2901), .A2(n4422), .ZN(n2449) );
  NAND2_X1 U2616 ( .A1(n4019), .A2(n4020), .ZN(n4018) );
  NOR2_X1 U2617 ( .A1(n2946), .A2(n2947), .ZN(n3318) );
  XNOR2_X1 U2618 ( .A(n3342), .B(n4472), .ZN(n4464) );
  NAND2_X1 U2619 ( .A1(n4473), .A2(n3344), .ZN(n3345) );
  NAND2_X1 U2620 ( .A1(n4480), .A2(n3322), .ZN(n3323) );
  NAND2_X1 U2621 ( .A1(n4486), .A2(REG1_REG_10__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U2622 ( .A1(n4501), .A2(n2275), .ZN(n3325) );
  NAND2_X1 U2623 ( .A1(n3334), .A2(REG1_REG_11__SCAN_IN), .ZN(n2275) );
  XNOR2_X1 U2624 ( .A(n2377), .B(n4029), .ZN(n3475) );
  NAND2_X1 U2625 ( .A1(n3474), .A2(n2378), .ZN(n2377) );
  NAND2_X1 U2626 ( .A1(n4427), .A2(REG1_REG_13__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U2627 ( .A1(n3475), .A2(REG1_REG_14__SCAN_IN), .ZN(n4031) );
  NOR2_X1 U2628 ( .A1(n4517), .A2(n2354), .ZN(n4049) );
  AND2_X1 U2629 ( .A1(n4047), .A2(REG2_REG_15__SCAN_IN), .ZN(n2354) );
  OAI22_X1 U2630 ( .A1(n4104), .A2(n2768), .B1(n4125), .B2(n4305), .ZN(n2865)
         );
  AOI21_X1 U2631 ( .B1(n4117), .B2(n3856), .A(n3967), .ZN(n4101) );
  OAI21_X1 U2632 ( .B1(n4115), .B2(n3902), .A(n3903), .ZN(n4104) );
  NAND2_X1 U2633 ( .A1(n2416), .A2(n2415), .ZN(n4172) );
  OR2_X1 U2634 ( .A1(n2419), .A2(n2730), .ZN(n2415) );
  NOR2_X1 U2635 ( .A1(n2730), .A2(n2418), .ZN(n2417) );
  INV_X1 U2636 ( .A(n4141), .ZN(n4183) );
  NAND2_X1 U2637 ( .A1(n4217), .A2(n2719), .ZN(n2420) );
  NOR2_X1 U2638 ( .A1(n4284), .A2(n4256), .ZN(n4241) );
  NAND2_X1 U2639 ( .A1(n3600), .A2(n2688), .ZN(n2414) );
  NAND2_X1 U2640 ( .A1(n2414), .A2(n2253), .ZN(n4270) );
  NOR2_X1 U2641 ( .A1(n2265), .A2(n2428), .ZN(n2427) );
  NAND2_X1 U2642 ( .A1(n2391), .A2(n2395), .ZN(n4549) );
  INV_X1 U2643 ( .A(n2392), .ZN(n2391) );
  OAI21_X1 U2644 ( .B1(n2396), .B2(n2393), .A(n2259), .ZN(n2392) );
  NAND2_X1 U2645 ( .A1(n2795), .A2(n3941), .ZN(n4551) );
  OAI21_X1 U2646 ( .B1(n3303), .B2(n3932), .A(n3926), .ZN(n3377) );
  NOR2_X1 U2647 ( .A1(n2585), .A2(n2405), .ZN(n2404) );
  INV_X1 U2648 ( .A(n2575), .ZN(n2405) );
  INV_X1 U2649 ( .A(IR_REG_20__SCAN_IN), .ZN(n4838) );
  NOR2_X1 U2650 ( .A1(n2544), .A2(n3154), .ZN(n2542) );
  NAND2_X1 U2651 ( .A1(n2547), .A2(n2546), .ZN(n2412) );
  NAND2_X1 U2652 ( .A1(n3155), .A2(n2545), .ZN(n2546) );
  NAND2_X1 U2653 ( .A1(n2685), .A2(n2319), .ZN(n2318) );
  INV_X1 U2654 ( .A(IR_REG_18__SCAN_IN), .ZN(n2319) );
  INV_X1 U2655 ( .A(IR_REG_19__SCAN_IN), .ZN(n4772) );
  INV_X1 U2656 ( .A(n4552), .ZN(n4298) );
  NAND2_X1 U2657 ( .A1(n4164), .A2(n2364), .ZN(n4126) );
  AND2_X1 U2658 ( .A1(n4184), .A2(n4166), .ZN(n4164) );
  AND2_X1 U2659 ( .A1(n2782), .A2(n4599), .ZN(n4638) );
  AND2_X1 U2660 ( .A1(n2431), .A2(n2488), .ZN(n2430) );
  NOR2_X1 U2661 ( .A1(IR_REG_27__SCAN_IN), .A2(n2489), .ZN(n2431) );
  OR2_X1 U2662 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2489)
         );
  NAND2_X1 U2663 ( .A1(n2841), .A2(n2833), .ZN(n2843) );
  NAND2_X1 U2664 ( .A1(n2473), .A2(n2635), .ZN(n2831) );
  AND4_X1 U2665 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n2485)
         );
  NOR2_X1 U2666 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2484)
         );
  NOR2_X1 U2667 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2483)
         );
  NOR2_X1 U2668 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2482)
         );
  INV_X1 U2669 ( .A(IR_REG_13__SCAN_IN), .ZN(n2637) );
  NOR2_X1 U2670 ( .A1(n2553), .A2(IR_REG_5__SCAN_IN), .ZN(n2596) );
  NOR2_X1 U2671 ( .A1(n2256), .A2(n2298), .ZN(n3369) );
  AND4_X1 U2672 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(n3451)
         );
  AND2_X1 U2673 ( .A1(n2697), .A2(n2696), .ZN(n3758) );
  INV_X1 U2674 ( .A(n3292), .ZN(n3298) );
  NAND2_X1 U2675 ( .A1(n2513), .A2(REG1_REG_1__SCAN_IN), .ZN(n2498) );
  OR2_X1 U2676 ( .A1(n2725), .A2(n2496), .ZN(n2497) );
  INV_X1 U2677 ( .A(n4438), .ZN(n3802) );
  AND4_X1 U2678 ( .A1(n2647), .A2(n2646), .A3(n2645), .A4(n2644), .ZN(n3824)
         );
  OAI21_X1 U2679 ( .B1(n3721), .B2(n2693), .A(n2736), .ZN(n4194) );
  NAND2_X1 U2680 ( .A1(n2718), .A2(n2717), .ZN(n4236) );
  AOI22_X1 U2681 ( .A1(n2702), .A2(REG0_REG_19__SCAN_IN), .B1(n2817), .B2(
        REG1_REG_19__SCAN_IN), .ZN(n2704) );
  INV_X1 U2682 ( .A(n4436), .ZN(n4281) );
  NAND2_X1 U2683 ( .A1(n2817), .A2(REG1_REG_5__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U2684 ( .A1(n2920), .A2(n2919), .ZN(n3016) );
  NAND2_X1 U2685 ( .A1(n2332), .A2(n2335), .ZN(n2330) );
  NOR2_X1 U2686 ( .A1(n2329), .A2(n2331), .ZN(n2328) );
  NAND2_X1 U2687 ( .A1(n4481), .A2(n4482), .ZN(n4480) );
  NAND2_X1 U2688 ( .A1(n2346), .A2(n2345), .ZN(n3472) );
  NAND2_X1 U2689 ( .A1(n2342), .A2(n2341), .ZN(n2345) );
  AOI21_X1 U2690 ( .B1(n2347), .B2(n4427), .A(n4426), .ZN(n2341) );
  NOR2_X1 U2691 ( .A1(n3473), .A2(n3472), .ZN(n4044) );
  XNOR2_X1 U2692 ( .A(n4049), .B(n4048), .ZN(n4528) );
  NAND2_X1 U2693 ( .A1(n4528), .A2(n3531), .ZN(n4527) );
  XNOR2_X1 U2694 ( .A(n2339), .B(n4066), .ZN(n4071) );
  NOR2_X1 U2695 ( .A1(n4063), .A2(n2274), .ZN(n2339) );
  AND2_X1 U2696 ( .A1(n4001), .A2(n2924), .ZN(n4507) );
  INV_X1 U2697 ( .A(n4346), .ZN(n4657) );
  NAND2_X1 U2698 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2380)
         );
  INV_X1 U2699 ( .A(IR_REG_24__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U2700 ( .A1(n3807), .A2(n2446), .ZN(n2445) );
  INV_X1 U2701 ( .A(n3746), .ZN(n2446) );
  NAND2_X1 U2702 ( .A1(n2445), .A2(n3745), .ZN(n2444) );
  INV_X1 U2703 ( .A(n2458), .ZN(n2457) );
  OAI21_X1 U2704 ( .B1(n3728), .B2(n2462), .A(n3637), .ZN(n2455) );
  OR2_X1 U2705 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  NAND2_X1 U2706 ( .A1(n4495), .A2(n3347), .ZN(n3348) );
  INV_X1 U2707 ( .A(n2737), .ZN(n2284) );
  NOR2_X1 U2708 ( .A1(n2288), .A2(n2745), .ZN(n2286) );
  INV_X1 U2709 ( .A(n2719), .ZN(n2418) );
  INV_X1 U2710 ( .A(n2424), .ZN(n2422) );
  AOI21_X1 U2711 ( .B1(n3889), .B2(n2426), .A(n2425), .ZN(n2424) );
  INV_X1 U2712 ( .A(n3833), .ZN(n2426) );
  INV_X1 U2713 ( .A(n2649), .ZN(n2428) );
  NAND2_X1 U2714 ( .A1(n2403), .A2(n2394), .ZN(n2393) );
  INV_X1 U2715 ( .A(n2607), .ZN(n2394) );
  INV_X1 U2716 ( .A(IR_REG_14__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U2717 ( .A1(n4102), .A2(n4282), .ZN(n2435) );
  AND2_X1 U2718 ( .A1(n4164), .A2(n2273), .ZN(n2876) );
  NOR2_X1 U2719 ( .A1(n4121), .A2(n4147), .ZN(n2364) );
  AND2_X1 U2720 ( .A1(n4200), .A2(n2248), .ZN(n2419) );
  NOR2_X1 U2721 ( .A1(n2376), .A2(n3281), .ZN(n2374) );
  NAND2_X1 U2722 ( .A1(n3252), .A2(n3078), .ZN(n2376) );
  INV_X1 U2723 ( .A(n3178), .ZN(n2375) );
  NAND2_X1 U2724 ( .A1(n2388), .A2(n3909), .ZN(n3120) );
  NAND2_X1 U2725 ( .A1(n2390), .A2(n2389), .ZN(n2388) );
  INV_X1 U2726 ( .A(n2786), .ZN(n2390) );
  INV_X1 U2727 ( .A(IR_REG_26__SCAN_IN), .ZN(n2488) );
  INV_X1 U2728 ( .A(IR_REG_28__SCAN_IN), .ZN(n2824) );
  NAND2_X1 U2729 ( .A1(n2502), .A2(n2501), .ZN(n2823) );
  INV_X1 U2730 ( .A(n2503), .ZN(n2502) );
  OR2_X1 U2731 ( .A1(n2615), .A2(IR_REG_10__SCAN_IN), .ZN(n2616) );
  AND2_X1 U2732 ( .A1(n2596), .A2(n2595), .ZN(n2605) );
  AND3_X1 U2733 ( .A1(n2594), .A2(n4904), .A3(n2593), .ZN(n2595) );
  INV_X1 U2734 ( .A(IR_REG_7__SCAN_IN), .ZN(n4904) );
  INV_X1 U2735 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U2736 ( .A1(n2662), .A2(REG3_REG_16__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U2737 ( .A1(n3363), .A2(n3364), .ZN(n2471) );
  OAI211_X1 U2738 ( .C1(n2306), .C2(n2305), .A(n2304), .B(n2472), .ZN(n2470)
         );
  OR2_X1 U2739 ( .A1(n3363), .A2(n3364), .ZN(n2472) );
  INV_X1 U2740 ( .A(n3992), .ZN(n4555) );
  NAND2_X1 U2741 ( .A1(n3777), .A2(n3778), .ZN(n3776) );
  INV_X1 U2742 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2628) );
  OR3_X1 U2743 ( .A1(n2721), .A2(n3738), .A3(n2720), .ZN(n2731) );
  OAI21_X1 U2744 ( .B1(n3777), .B2(n2313), .A(n2310), .ZN(n2314) );
  NAND2_X1 U2745 ( .A1(n2266), .A2(n3780), .ZN(n2313) );
  AND2_X1 U2746 ( .A1(n2311), .A2(n2268), .ZN(n2310) );
  NAND2_X1 U2747 ( .A1(n3041), .A2(n3042), .ZN(n3063) );
  NOR2_X2 U2748 ( .A1(n2642), .A2(n2641), .ZN(n2650) );
  NAND2_X1 U2749 ( .A1(n2817), .A2(REG1_REG_14__SCAN_IN), .ZN(n2645) );
  INV_X1 U2750 ( .A(n2324), .ZN(n2323) );
  AND2_X1 U2751 ( .A1(n3613), .A2(n2322), .ZN(n2321) );
  NAND2_X1 U2752 ( .A1(n2320), .A2(n2324), .ZN(n3614) );
  NAND2_X1 U2753 ( .A1(n3607), .A2(n2322), .ZN(n2320) );
  AND2_X1 U2754 ( .A1(n2775), .A2(n2774), .ZN(n3692) );
  NAND2_X1 U2755 ( .A1(n4008), .A2(n4007), .ZN(n4006) );
  XNOR2_X1 U2756 ( .A(n2942), .B(n3026), .ZN(n3023) );
  NAND2_X1 U2757 ( .A1(n3023), .A2(REG1_REG_4__SCAN_IN), .ZN(n3022) );
  INV_X1 U2758 ( .A(n4023), .ZN(n2334) );
  INV_X1 U2759 ( .A(n2958), .ZN(n2338) );
  INV_X1 U2760 ( .A(n2332), .ZN(n2329) );
  NAND2_X1 U2761 ( .A1(n4463), .A2(n3343), .ZN(n4474) );
  NAND2_X1 U2762 ( .A1(n4487), .A2(n3346), .ZN(n4496) );
  NAND2_X1 U2763 ( .A1(n4496), .A2(n4497), .ZN(n4495) );
  XNOR2_X1 U2764 ( .A(n3348), .B(n4516), .ZN(n4508) );
  OR2_X1 U2765 ( .A1(n3470), .A2(REG2_REG_13__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U2766 ( .A1(n2876), .A2(n3848), .ZN(n4297) );
  NAND2_X1 U2767 ( .A1(n4100), .A2(n2816), .ZN(n2873) );
  AND2_X1 U2768 ( .A1(n2529), .A2(DATAI_28_), .ZN(n4092) );
  OR2_X1 U2769 ( .A1(n4163), .A2(n4313), .ZN(n2753) );
  NAND2_X1 U2770 ( .A1(n4156), .A2(n3958), .ZN(n2386) );
  INV_X1 U2771 ( .A(n4242), .ZN(n3782) );
  NAND2_X1 U2772 ( .A1(n2709), .A2(REG3_REG_20__SCAN_IN), .ZN(n2721) );
  AOI21_X1 U2773 ( .B1(n2414), .B2(n2292), .A(n2290), .ZN(n2289) );
  NAND2_X1 U2774 ( .A1(n2291), .A2(n2708), .ZN(n2290) );
  AND2_X1 U2775 ( .A1(n2529), .A2(DATAI_20_), .ZN(n4242) );
  NAND2_X1 U2776 ( .A1(n2423), .A2(n2424), .ZN(n4230) );
  NAND2_X1 U2777 ( .A1(n2805), .A2(n3833), .ZN(n3526) );
  OAI21_X1 U2778 ( .B1(n4549), .B2(n2279), .A(n2276), .ZN(n3428) );
  AOI21_X1 U2779 ( .B1(n2278), .B2(n2277), .A(n2281), .ZN(n2276) );
  INV_X1 U2780 ( .A(n4550), .ZN(n2277) );
  OR2_X1 U2781 ( .A1(n2598), .A2(n3403), .ZN(n2609) );
  INV_X1 U2782 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U2783 ( .A1(n2398), .A2(n2402), .ZN(n3376) );
  NAND2_X1 U2784 ( .A1(n2400), .A2(n2399), .ZN(n2398) );
  NAND2_X1 U2785 ( .A1(n3260), .A2(n3927), .ZN(n2429) );
  NAND2_X1 U2786 ( .A1(n2577), .A2(REG3_REG_8__SCAN_IN), .ZN(n2587) );
  NOR2_X1 U2787 ( .A1(n3178), .A2(n2372), .ZN(n3267) );
  NAND2_X1 U2788 ( .A1(n2374), .A2(n3239), .ZN(n2372) );
  INV_X1 U2789 ( .A(IR_REG_11__SCAN_IN), .ZN(n4868) );
  AND2_X1 U2790 ( .A1(n3003), .A2(n2979), .ZN(n4558) );
  AND2_X1 U2791 ( .A1(n2992), .A2(n2979), .ZN(n4282) );
  NAND2_X1 U2792 ( .A1(n2790), .A2(n3915), .ZN(n3158) );
  NAND2_X1 U2793 ( .A1(n2387), .A2(n3910), .ZN(n3170) );
  NAND2_X1 U2794 ( .A1(n3120), .A2(n3119), .ZN(n2387) );
  AND2_X1 U2795 ( .A1(n3915), .A2(n3912), .ZN(n3888) );
  INV_X1 U2796 ( .A(n3140), .ZN(n3136) );
  AND2_X1 U2797 ( .A1(n3136), .A2(n4601), .ZN(n3134) );
  INV_X1 U2798 ( .A(n4558), .ZN(n4274) );
  NOR2_X1 U2799 ( .A1(n4297), .A2(n4299), .ZN(n4296) );
  AOI21_X1 U2800 ( .B1(n2436), .B2(n4254), .A(n2433), .ZN(n4082) );
  NAND2_X1 U2801 ( .A1(n2435), .A2(n2434), .ZN(n2433) );
  XNOR2_X1 U2802 ( .A(n2438), .B(n2437), .ZN(n2436) );
  NAND2_X1 U2803 ( .A1(n3845), .A2(n4075), .ZN(n2434) );
  NAND2_X1 U2804 ( .A1(n4164), .A2(n4313), .ZN(n4145) );
  AND2_X1 U2805 ( .A1(n4241), .A2(n2251), .ZN(n4184) );
  AND2_X1 U2806 ( .A1(n2420), .A2(n2419), .ZN(n4328) );
  NAND2_X1 U2807 ( .A1(n4241), .A2(n2250), .ZN(n4218) );
  INV_X1 U2808 ( .A(n2369), .ZN(n2368) );
  NOR3_X1 U2809 ( .A1(n4367), .A2(n4439), .A3(n3826), .ZN(n4360) );
  NOR2_X1 U2810 ( .A1(n4367), .A2(n3826), .ZN(n3533) );
  NAND2_X1 U2811 ( .A1(n2360), .A2(n3576), .ZN(n2359) );
  INV_X1 U2812 ( .A(n2361), .ZN(n2360) );
  NOR3_X1 U2813 ( .A1(n3311), .A2(n4567), .A3(n2361), .ZN(n3439) );
  NOR3_X1 U2814 ( .A1(n3311), .A2(n4567), .A3(n3406), .ZN(n4565) );
  NAND2_X1 U2815 ( .A1(n2375), .A2(n2374), .ZN(n3278) );
  NOR2_X1 U2816 ( .A1(n3178), .A2(n3159), .ZN(n3212) );
  NAND2_X1 U2817 ( .A1(n2375), .A2(n2373), .ZN(n3280) );
  INV_X1 U2818 ( .A(n2376), .ZN(n2373) );
  INV_X1 U2819 ( .A(n3215), .ZN(n3252) );
  NAND2_X1 U2820 ( .A1(n3128), .A2(n3134), .ZN(n3176) );
  OR2_X1 U2821 ( .A1(n3176), .A2(n3175), .ZN(n3178) );
  NAND2_X1 U2822 ( .A1(n2503), .A2(IR_REG_31__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U2823 ( .A1(n2830), .A2(n2439), .ZN(n2839) );
  INV_X1 U2824 ( .A(n2841), .ZN(n2842) );
  NAND2_X1 U2825 ( .A1(n2777), .A2(IR_REG_31__SCAN_IN), .ZN(n2778) );
  AND2_X1 U2826 ( .A1(n2669), .A2(n2659), .ZN(n4047) );
  NAND2_X1 U2827 ( .A1(n2308), .A2(n2306), .ZN(n3289) );
  NAND2_X1 U2828 ( .A1(n2464), .A2(n2463), .ZN(n2308) );
  INV_X1 U2829 ( .A(n3993), .ZN(n3404) );
  AOI21_X1 U2830 ( .B1(n2460), .B2(n2458), .A(n3796), .ZN(n3729) );
  INV_X1 U2831 ( .A(n2461), .ZN(n2460) );
  OAI22_X1 U2832 ( .A1(n3710), .A2(n3711), .B1(n3685), .B2(n3684), .ZN(n3696)
         );
  NAND2_X1 U2833 ( .A1(n3289), .A2(n3288), .ZN(n3365) );
  INV_X1 U2834 ( .A(n3461), .ZN(n3582) );
  AND2_X1 U2835 ( .A1(n2755), .A2(n2747), .ZN(n4146) );
  AND4_X1 U2836 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .ZN(n4436)
         );
  OAI21_X1 U2837 ( .B1(n2529), .B2(n2452), .A(n2363), .ZN(n3705) );
  NAND2_X1 U2838 ( .A1(n2529), .A2(DATAI_0_), .ZN(n2363) );
  INV_X1 U2839 ( .A(n3541), .ZN(n3576) );
  NAND2_X1 U2840 ( .A1(n2441), .A2(n3037), .ZN(n3047) );
  NAND2_X1 U2841 ( .A1(n2440), .A2(n3063), .ZN(n3046) );
  NOR2_X1 U2842 ( .A1(n2461), .A2(n2474), .ZN(n3799) );
  INV_X1 U2843 ( .A(n4448), .ZN(n3804) );
  AND4_X1 U2844 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n3262)
         );
  NAND2_X1 U2845 ( .A1(n2465), .A2(n3190), .ZN(n3237) );
  OR2_X1 U2846 ( .A1(n2756), .A2(n2762), .ZN(n4129) );
  OAI21_X1 U2847 ( .B1(n3744), .B2(n3745), .A(n3746), .ZN(n3809) );
  AND4_X1 U2848 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n3823)
         );
  INV_X1 U2849 ( .A(n3816), .ZN(n4443) );
  NAND2_X1 U2850 ( .A1(n2987), .A2(n4264), .ZN(n4438) );
  NAND2_X1 U2851 ( .A1(n2817), .A2(REG1_REG_31__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U2852 ( .A1(n2822), .A2(n2821), .ZN(n3987) );
  INV_X1 U2853 ( .A(n4163), .ZN(n4122) );
  NAND2_X1 U2854 ( .A1(n2744), .A2(n2743), .ZN(n4141) );
  INV_X1 U2855 ( .A(n3823), .ZN(n3989) );
  NAND4_X1 U2856 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n3612)
         );
  INV_X1 U2857 ( .A(n3451), .ZN(n3991) );
  INV_X1 U2858 ( .A(n3369), .ZN(n3305) );
  INV_X1 U2859 ( .A(n3262), .ZN(n3994) );
  NAND2_X1 U2860 ( .A1(n2817), .A2(REG1_REG_6__SCAN_IN), .ZN(n2559) );
  OR2_X1 U2861 ( .A1(n2725), .A2(n2533), .ZN(n2536) );
  OR2_X1 U2862 ( .A1(n2725), .A2(n2506), .ZN(n2509) );
  OAI21_X1 U2863 ( .B1(n2353), .B2(n2917), .A(n2350), .ZN(n4011) );
  NAND2_X1 U2864 ( .A1(n4011), .A2(n2918), .ZN(n4010) );
  XNOR2_X1 U2865 ( .A(n2951), .B(n2929), .ZN(n2950) );
  INV_X1 U2866 ( .A(n4430), .ZN(n3026) );
  NAND2_X1 U2867 ( .A1(n4022), .A2(n2331), .ZN(n2327) );
  NAND2_X1 U2868 ( .A1(n4021), .A2(n2958), .ZN(n3338) );
  XNOR2_X1 U2869 ( .A(n3345), .B(n4491), .ZN(n4488) );
  NAND2_X1 U2870 ( .A1(n4485), .A2(n3324), .ZN(n4502) );
  NAND2_X1 U2871 ( .A1(n4502), .A2(n4503), .ZN(n4501) );
  INV_X1 U2872 ( .A(n2377), .ZN(n4030) );
  INV_X1 U2873 ( .A(n2346), .ZN(n4045) );
  NAND2_X1 U2874 ( .A1(n4527), .A2(n4050), .ZN(n4536) );
  NOR2_X1 U2875 ( .A1(n4052), .A2(n4053), .ZN(n4063) );
  NAND2_X1 U2876 ( .A1(n4537), .A2(n2340), .ZN(n4052) );
  NAND2_X1 U2877 ( .A1(n4584), .A2(n4846), .ZN(n2340) );
  OAI21_X1 U2878 ( .B1(n4172), .B2(n2737), .A(n2287), .ZN(n4154) );
  AND2_X1 U2879 ( .A1(n2420), .A2(n2248), .ZN(n4201) );
  NAND2_X1 U2880 ( .A1(n4241), .A2(n3782), .ZN(n4341) );
  NAND2_X1 U2881 ( .A1(n4270), .A2(n2699), .ZN(n4248) );
  NAND2_X1 U2882 ( .A1(n2414), .A2(n2689), .ZN(n4272) );
  NAND2_X1 U2883 ( .A1(n3481), .A2(n2649), .ZN(n3510) );
  OR2_X1 U2884 ( .A1(n2247), .A2(n3555), .ZN(n4367) );
  NAND2_X1 U2885 ( .A1(n4549), .A2(n4550), .ZN(n2280) );
  NAND2_X1 U2886 ( .A1(n2401), .A2(n2584), .ZN(n3308) );
  NAND2_X1 U2887 ( .A1(n2576), .A2(n2404), .ZN(n2401) );
  NAND2_X1 U2888 ( .A1(n2411), .A2(n2409), .ZN(n3274) );
  INV_X1 U2889 ( .A(n2410), .ZN(n2409) );
  NAND2_X1 U2890 ( .A1(n2413), .A2(n2412), .ZN(n3220) );
  OR2_X1 U2891 ( .A1(n2986), .A2(n2985), .ZN(n4264) );
  NAND2_X1 U2892 ( .A1(n2777), .A2(n2706), .ZN(n4069) );
  OAI21_X1 U2893 ( .B1(n2684), .B2(n2318), .A(IR_REG_31__SCAN_IN), .ZN(n2705)
         );
  INV_X1 U2894 ( .A(n4263), .ZN(n5032) );
  INV_X1 U2895 ( .A(n4264), .ZN(n5034) );
  INV_X1 U2896 ( .A(n3705), .ZN(n4601) );
  AND2_X1 U2897 ( .A1(n2784), .A2(n3877), .ZN(n4599) );
  AND2_X1 U2898 ( .A1(n4290), .A2(n4298), .ZN(n4148) );
  OAI21_X1 U2899 ( .B1(n4107), .B2(n4305), .A(n2365), .ZN(n4381) );
  NAND2_X1 U2900 ( .A1(n2900), .A2(n2983), .ZN(n4582) );
  INV_X1 U2901 ( .A(n3003), .ZN(n2992) );
  AND2_X1 U2902 ( .A1(n3052), .A2(STATE_REG_SCAN_IN), .ZN(n4583) );
  XNOR2_X1 U2903 ( .A(n2780), .B(IR_REG_22__SCAN_IN), .ZN(n3982) );
  XNOR2_X1 U2904 ( .A(n2779), .B(IR_REG_21__SCAN_IN), .ZN(n4423) );
  AND2_X1 U2905 ( .A1(n2556), .A2(n2555), .ZN(n4429) );
  AND2_X1 U2906 ( .A1(n2541), .A2(n2540), .ZN(n4431) );
  XNOR2_X1 U2907 ( .A(n2518), .B(IR_REG_2__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U2908 ( .A1(n2452), .A2(n2451), .ZN(n2450) );
  CLKBUF_X2 U2909 ( .A(n2909), .Z(U4043) );
  OAI211_X1 U2910 ( .C1(n4022), .C2(n2335), .A(n2332), .B(n2327), .ZN(n2960)
         );
  OR2_X1 U2911 ( .A1(n4091), .A2(n4358), .ZN(n2858) );
  OR2_X1 U2912 ( .A1(n4091), .A2(n4417), .ZN(n2863) );
  NAND2_X1 U2913 ( .A1(n2349), .A2(n2348), .ZN(U3351) );
  NAND2_X1 U2914 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2348) );
  MUX2_X2 U2915 ( .A(n2505), .B(n2504), .S(n2870), .Z(n2529) );
  OAI21_X1 U2916 ( .B1(n3607), .B2(n2323), .A(n2321), .ZN(n3819) );
  AND2_X1 U2917 ( .A1(n2448), .A2(n2447), .ZN(n3744) );
  AND3_X1 U2918 ( .A1(n4771), .A2(n2487), .A3(n2833), .ZN(n2244) );
  NAND2_X1 U2919 ( .A1(n3996), .A2(n3215), .ZN(n2245) );
  OR2_X1 U2920 ( .A1(n2455), .A2(n2264), .ZN(n2246) );
  OR3_X1 U2921 ( .A1(n3311), .A2(n2359), .A3(n4567), .ZN(n2247) );
  OR2_X1 U2922 ( .A1(n4236), .A2(n3650), .ZN(n2248) );
  OR2_X1 U2923 ( .A1(n2684), .A2(IR_REG_17__SCAN_IN), .ZN(n2249) );
  INV_X1 U2924 ( .A(n4452), .ZN(n4598) );
  AND2_X1 U2925 ( .A1(n3782), .A2(n4335), .ZN(n2250) );
  INV_X1 U2926 ( .A(n3334), .ZN(n4591) );
  AND2_X1 U2927 ( .A1(n2618), .A2(n2626), .ZN(n3334) );
  INV_X1 U2928 ( .A(n2857), .ZN(n4285) );
  AND2_X1 U2929 ( .A1(n2371), .A2(n4186), .ZN(n2251) );
  AND2_X1 U2930 ( .A1(n2364), .A2(n4305), .ZN(n2252) );
  AND3_X1 U2931 ( .A1(n2473), .A2(n2295), .A3(n2635), .ZN(n2829) );
  AND2_X1 U2932 ( .A1(n4276), .A2(n2689), .ZN(n2253) );
  XNOR2_X1 U2933 ( .A(n2380), .B(IR_REG_1__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U2934 ( .A1(n3776), .A2(n3780), .ZN(n3734) );
  OR2_X1 U2935 ( .A1(n4557), .A2(n3461), .ZN(n2254) );
  AOI21_X1 U2936 ( .B1(n3717), .B2(n3669), .A(n3668), .ZN(n3765) );
  OR2_X1 U2937 ( .A1(n3993), .A2(n3371), .ZN(n2255) );
  AND2_X1 U2938 ( .A1(n2817), .A2(REG1_REG_8__SCAN_IN), .ZN(n2256) );
  OR2_X1 U2939 ( .A1(n2943), .A2(n3026), .ZN(n2257) );
  INV_X1 U2940 ( .A(IR_REG_27__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U2941 ( .A1(n2635), .A2(n2485), .ZN(n2258) );
  NAND2_X1 U2942 ( .A1(n4555), .A2(n3384), .ZN(n2259) );
  INV_X1 U2943 ( .A(n2279), .ZN(n2278) );
  NAND2_X1 U2944 ( .A1(n2619), .A2(n2254), .ZN(n2279) );
  NOR2_X1 U2945 ( .A1(n2798), .A2(n3582), .ZN(n2281) );
  INV_X1 U2946 ( .A(n2403), .ZN(n2399) );
  NAND2_X1 U2947 ( .A1(n2255), .A2(n2584), .ZN(n2403) );
  OR2_X1 U2948 ( .A1(n3236), .A2(n2467), .ZN(n2260) );
  AND2_X1 U2949 ( .A1(n3921), .A2(n2793), .ZN(n2261) );
  INV_X1 U2950 ( .A(n3288), .ZN(n2305) );
  NOR2_X1 U2951 ( .A1(n3953), .A2(n2422), .ZN(n2262) );
  AND2_X1 U2952 ( .A1(n2444), .A2(n2443), .ZN(n2263) );
  INV_X1 U2953 ( .A(IR_REG_31__SCAN_IN), .ZN(n2490) );
  INV_X1 U2954 ( .A(IR_REG_1__SCAN_IN), .ZN(n2451) );
  AND2_X1 U2955 ( .A1(n3756), .A2(n3755), .ZN(n2264) );
  INV_X1 U2956 ( .A(n3875), .ZN(n2437) );
  NOR2_X1 U2957 ( .A1(n3612), .A2(n3826), .ZN(n2265) );
  NAND2_X1 U2958 ( .A1(n4164), .A2(n2252), .ZN(n2365) );
  INV_X1 U2959 ( .A(n3906), .ZN(n2389) );
  NAND2_X1 U2960 ( .A1(n3736), .A2(n3735), .ZN(n2266) );
  MUX2_X1 U2961 ( .A(n4430), .B(DATAI_4_), .S(n2529), .Z(n3159) );
  AND2_X1 U2962 ( .A1(n3680), .A2(n3679), .ZN(n2267) );
  NAND2_X1 U2963 ( .A1(n3653), .A2(n3652), .ZN(n2268) );
  INV_X1 U2964 ( .A(n2288), .ZN(n2287) );
  INV_X1 U2965 ( .A(n3898), .ZN(n2385) );
  AND2_X1 U2966 ( .A1(n4183), .A2(n4166), .ZN(n2269) );
  NOR2_X1 U2967 ( .A1(n3614), .A2(n3613), .ZN(n3818) );
  NOR2_X1 U2968 ( .A1(n4122), .A2(n4147), .ZN(n2270) );
  AND2_X1 U2969 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2271)
         );
  INV_X1 U2970 ( .A(n2788), .ZN(n3119) );
  NOR2_X1 U2971 ( .A1(n3311), .A2(n3406), .ZN(n2362) );
  AND2_X1 U2972 ( .A1(n4241), .A2(n2371), .ZN(n2272) );
  INV_X1 U2973 ( .A(n3836), .ZN(n2425) );
  NAND2_X1 U2974 ( .A1(n2280), .A2(n2619), .ZN(n3438) );
  NAND2_X1 U2975 ( .A1(n2576), .A2(n2575), .ZN(n3259) );
  NAND2_X1 U2976 ( .A1(n2470), .A2(n2471), .ZN(n3366) );
  NOR2_X1 U2977 ( .A1(n4367), .A2(n2367), .ZN(n2370) );
  INV_X1 U2978 ( .A(n2366), .ZN(n4283) );
  NOR3_X1 U2979 ( .A1(n4367), .A2(n4439), .A3(n2369), .ZN(n2366) );
  INV_X1 U2980 ( .A(n3796), .ZN(n2462) );
  INV_X1 U2981 ( .A(IR_REG_17__SCAN_IN), .ZN(n2685) );
  INV_X1 U2982 ( .A(n4439), .ZN(n3617) );
  NAND2_X1 U2983 ( .A1(n2517), .A2(n2477), .ZN(n2993) );
  INV_X1 U2984 ( .A(n3068), .ZN(n2915) );
  AND2_X1 U2985 ( .A1(n2529), .A2(DATAI_27_), .ZN(n4108) );
  INV_X1 U2986 ( .A(n4108), .ZN(n4305) );
  INV_X1 U2987 ( .A(n4186), .ZN(n4180) );
  NAND2_X1 U2988 ( .A1(n2529), .A2(DATAI_23_), .ZN(n4186) );
  AND2_X1 U2989 ( .A1(n2529), .A2(DATAI_21_), .ZN(n3650) );
  INV_X1 U2990 ( .A(n4147), .ZN(n4313) );
  AND2_X1 U2991 ( .A1(n2529), .A2(DATAI_25_), .ZN(n4147) );
  INV_X1 U2992 ( .A(n4092), .ZN(n3690) );
  AND2_X1 U2993 ( .A1(n2252), .A2(n3690), .ZN(n2273) );
  AND2_X1 U2994 ( .A1(n4064), .A2(REG2_REG_18__SCAN_IN), .ZN(n2274) );
  AND2_X1 U2995 ( .A1(n2686), .A2(n2249), .ZN(n4051) );
  INV_X1 U2996 ( .A(n4051), .ZN(n4584) );
  INV_X1 U2997 ( .A(IR_REG_0__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U2998 ( .A1(n2930), .A2(REG1_REG_3__SCAN_IN), .ZN(n2941) );
  NAND2_X1 U2999 ( .A1(n3330), .A2(n3329), .ZN(n3474) );
  NOR2_X2 U3000 ( .A1(n4531), .A2(REG1_REG_16__SCAN_IN), .ZN(n4532) );
  NAND2_X1 U3001 ( .A1(n4523), .A2(n4524), .ZN(n4522) );
  NOR2_X1 U3002 ( .A1(n3771), .A2(n4186), .ZN(n2288) );
  INV_X1 U3003 ( .A(n2289), .ZN(n4226) );
  AOI22_X1 U3004 ( .A1(n2702), .A2(REG0_REG_18__SCAN_IN), .B1(n2817), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n2697) );
  NAND4_X1 U3005 ( .A1(n2473), .A2(n2295), .A3(n2635), .A4(n2488), .ZN(n2503)
         );
  NAND3_X1 U3006 ( .A1(n2473), .A2(n2635), .A3(n2244), .ZN(n2297) );
  NAND3_X1 U3007 ( .A1(n2580), .A2(n2581), .A3(n2579), .ZN(n2298) );
  NAND3_X1 U3008 ( .A1(n2452), .A2(n2451), .A3(n2302), .ZN(n2527) );
  INV_X1 U3009 ( .A(n2527), .ZN(n2479) );
  NAND2_X1 U3010 ( .A1(n2464), .A2(n2303), .ZN(n2304) );
  OAI21_X1 U3011 ( .B1(n2464), .B2(n2466), .A(n2463), .ZN(n3244) );
  NAND2_X4 U3012 ( .A1(n2309), .A2(n3054), .ZN(n3691) );
  NAND2_X2 U3013 ( .A1(n2782), .A2(n4423), .ZN(n2966) );
  NAND3_X1 U3014 ( .A1(n2266), .A2(n3780), .A3(n2312), .ZN(n2311) );
  INV_X1 U3015 ( .A(n2314), .ZN(n3789) );
  INV_X1 U3016 ( .A(n2315), .ZN(n2777) );
  NOR2_X1 U3017 ( .A1(n3553), .A2(n2476), .ZN(n3607) );
  NAND2_X1 U3018 ( .A1(n4022), .A2(n2328), .ZN(n2326) );
  OAI211_X1 U3019 ( .C1(n4022), .C2(n2330), .A(REG2_REG_6__SCAN_IN), .B(n2326), 
        .ZN(n3339) );
  NAND2_X1 U3020 ( .A1(n4022), .A2(n4023), .ZN(n4021) );
  NAND2_X1 U3021 ( .A1(n2337), .A2(n2334), .ZN(n2333) );
  NAND2_X1 U3022 ( .A1(n3471), .A2(n2347), .ZN(n2342) );
  NAND2_X1 U3023 ( .A1(n2353), .A2(n2917), .ZN(n2350) );
  NAND2_X1 U3024 ( .A1(n2353), .A2(REG2_REG_1__SCAN_IN), .ZN(n3013) );
  NAND2_X1 U3025 ( .A1(n2353), .A2(REG1_REG_1__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U3026 ( .A1(n2353), .A2(STATE_REG_SCAN_IN), .ZN(n2349) );
  XNOR2_X1 U3027 ( .A(n2353), .B(n2926), .ZN(n4008) );
  NAND2_X1 U3028 ( .A1(n2529), .A2(DATAI_1_), .ZN(n2351) );
  INV_X1 U3029 ( .A(n2353), .ZN(n2352) );
  NAND2_X1 U3030 ( .A1(n4017), .A2(n2353), .ZN(n4016) );
  NAND2_X1 U3031 ( .A1(n4538), .A2(n4536), .ZN(n4537) );
  AOI21_X1 U3032 ( .B1(n4071), .B2(n4507), .A(n4070), .ZN(n4072) );
  NAND2_X1 U3033 ( .A1(n3349), .A2(n4506), .ZN(n3470) );
  NAND4_X1 U3034 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), .ZN(n2480)
         );
  INV_X1 U3035 ( .A(n2362), .ZN(n4566) );
  INV_X1 U3036 ( .A(n2365), .ZN(n4106) );
  NAND3_X1 U3037 ( .A1(n3617), .A2(n2368), .A3(n4285), .ZN(n2367) );
  INV_X1 U3038 ( .A(n2370), .ZN(n4284) );
  INV_X1 U3039 ( .A(n2383), .ZN(n4455) );
  NAND2_X1 U3040 ( .A1(n2382), .A2(n2381), .ZN(n3320) );
  NAND2_X1 U3041 ( .A1(n2383), .A2(n4452), .ZN(n2381) );
  OR2_X1 U3042 ( .A1(n3318), .A2(n3319), .ZN(n2383) );
  NAND2_X1 U3043 ( .A1(n2576), .A2(n2397), .ZN(n2395) );
  NOR2_X1 U3044 ( .A1(n2396), .A2(n2607), .ZN(n2397) );
  INV_X1 U3045 ( .A(n2576), .ZN(n2400) );
  INV_X1 U3046 ( .A(n2396), .ZN(n2402) );
  NAND2_X1 U3047 ( .A1(n2406), .A2(n2563), .ZN(n2408) );
  NAND3_X1 U3048 ( .A1(n2245), .A2(n2413), .A3(n2412), .ZN(n2411) );
  NAND4_X1 U3049 ( .A1(n2413), .A2(n2245), .A3(n2412), .A4(n2563), .ZN(n2407)
         );
  NAND2_X1 U3050 ( .A1(n2543), .A2(n2542), .ZN(n2413) );
  NAND2_X1 U3051 ( .A1(n4217), .A2(n2417), .ZN(n2416) );
  NAND2_X1 U3052 ( .A1(n2792), .A2(n2261), .ZN(n2794) );
  NAND2_X1 U3053 ( .A1(n2792), .A2(n3921), .ZN(n2421) );
  XNOR2_X1 U3054 ( .A(n2421), .B(n3922), .ZN(n3228) );
  NAND2_X1 U3055 ( .A1(n2423), .A2(n2262), .ZN(n4174) );
  OR2_X2 U3056 ( .A1(n2805), .A2(n3525), .ZN(n2423) );
  NAND2_X1 U3057 ( .A1(n3481), .A2(n2427), .ZN(n2661) );
  NAND2_X1 U3058 ( .A1(n3482), .A2(n3892), .ZN(n3481) );
  OAI21_X2 U3059 ( .B1(n3158), .B2(n2791), .A(n3919), .ZN(n3210) );
  NAND2_X1 U3060 ( .A1(n2829), .A2(n2430), .ZN(n2432) );
  INV_X1 U3061 ( .A(n2432), .ZN(n2491) );
  INV_X1 U3062 ( .A(n2829), .ZN(n2439) );
  NAND4_X1 U3063 ( .A1(n2441), .A2(n3037), .A3(n2440), .A4(n3063), .ZN(n3064)
         );
  NAND2_X1 U3064 ( .A1(n3044), .A2(n3043), .ZN(n2440) );
  NAND2_X1 U3065 ( .A1(n3033), .A2(n3034), .ZN(n2441) );
  NAND2_X1 U3066 ( .A1(n2442), .A2(n2263), .ZN(n3710) );
  NAND3_X1 U3067 ( .A1(n2448), .A2(n2447), .A3(n2445), .ZN(n2442) );
  NAND2_X1 U3068 ( .A1(n3766), .A2(n3768), .ZN(n2447) );
  INV_X1 U3069 ( .A(n3765), .ZN(n2448) );
  INV_X1 U3070 ( .A(n3054), .ZN(n2972) );
  INV_X4 U3071 ( .A(n3691), .ZN(n3681) );
  NAND2_X2 U3072 ( .A1(n2840), .A2(n2449), .ZN(n3054) );
  NAND2_X1 U3073 ( .A1(IR_REG_31__SCAN_IN), .A2(n2450), .ZN(n2518) );
  NOR2_X2 U3074 ( .A1(n2454), .A2(n2453), .ZN(n3777) );
  NOR2_X1 U3075 ( .A1(n3754), .A2(n2246), .ZN(n2454) );
  NAND2_X1 U3076 ( .A1(n3186), .A2(n3238), .ZN(n2464) );
  OR2_X1 U3077 ( .A1(n2831), .A2(IR_REG_22__SCAN_IN), .ZN(n2832) );
  INV_X1 U3078 ( .A(n2493), .ZN(n2495) );
  NAND2_X1 U3079 ( .A1(n2837), .A2(n2901), .ZN(n2900) );
  AND2_X1 U3080 ( .A1(n3627), .A2(n3626), .ZN(n2474) );
  AND2_X1 U3081 ( .A1(n2538), .A2(n2478), .ZN(n2475) );
  INV_X1 U3082 ( .A(n4358), .ZN(n2879) );
  INV_X1 U3083 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3084 ( .A1(n4645), .A2(n4638), .ZN(n4417) );
  INV_X1 U3085 ( .A(n4417), .ZN(n2884) );
  NAND2_X1 U3086 ( .A1(n3552), .A2(n3565), .ZN(n2476) );
  OR2_X1 U3087 ( .A1(n3844), .A2(n3850), .ZN(n3864) );
  INV_X1 U3088 ( .A(n3864), .ZN(n2776) );
  AND3_X1 U3089 ( .A1(n2516), .A2(n2515), .A3(n2514), .ZN(n2477) );
  INV_X1 U3090 ( .A(n4200), .ZN(n2729) );
  NAND2_X1 U3091 ( .A1(n2728), .A2(n2727), .ZN(n4214) );
  INV_X1 U3092 ( .A(IR_REG_4__SCAN_IN), .ZN(n2478) );
  INV_X1 U3093 ( .A(IR_REG_22__SCAN_IN), .ZN(n2487) );
  INV_X1 U3094 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U3095 ( .A1(n3709), .A2(n3140), .ZN(n3909) );
  INV_X1 U3096 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2565) );
  INV_X1 U3097 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2690) );
  OR2_X1 U3098 ( .A1(n2787), .A2(n3671), .ZN(n2974) );
  NOR2_X1 U3099 ( .A1(n2731), .A2(n3722), .ZN(n2738) );
  AND2_X1 U3100 ( .A1(n4083), .A2(n2770), .ZN(n3697) );
  NOR2_X1 U3101 ( .A1(n2755), .A2(n2754), .ZN(n2762) );
  INV_X1 U3102 ( .A(n4135), .ZN(n4136) );
  NOR2_X1 U3103 ( .A1(n3739), .A2(n4197), .ZN(n2730) );
  INV_X1 U3104 ( .A(n4557), .ZN(n2798) );
  OR2_X1 U3105 ( .A1(n2587), .A2(n2586), .ZN(n2598) );
  INV_X1 U3106 ( .A(n3121), .ZN(n3128) );
  INV_X1 U3107 ( .A(n2983), .ZN(n2986) );
  AND2_X1 U3108 ( .A1(n3719), .A2(n3720), .ZN(n3662) );
  NOR2_X1 U3109 ( .A1(n2691), .A2(n2690), .ZN(n2700) );
  INV_X1 U3110 ( .A(n4214), .ZN(n3739) );
  OR2_X1 U3111 ( .A1(n2746), .A2(n3749), .ZN(n2755) );
  OR2_X1 U3112 ( .A1(n2673), .A2(n2672), .ZN(n2691) );
  OR2_X1 U3113 ( .A1(n2629), .A2(n2628), .ZN(n2642) );
  OR2_X1 U3114 ( .A1(n2991), .A2(n3981), .ZN(n2994) );
  INV_X1 U3115 ( .A(n3810), .ZN(n4434) );
  AND2_X1 U3116 ( .A1(n2762), .A2(REG3_REG_27__SCAN_IN), .ZN(n2769) );
  INV_X1 U3117 ( .A(n4431), .ZN(n2929) );
  INV_X1 U3118 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3403) );
  AND2_X1 U3119 ( .A1(n2752), .A2(n2751), .ZN(n4163) );
  AND2_X1 U3120 ( .A1(n3900), .A2(n4175), .ZN(n4212) );
  INV_X1 U3121 ( .A(n4282), .ZN(n4554) );
  INV_X1 U3122 ( .A(n4127), .ZN(n4121) );
  NAND2_X1 U3123 ( .A1(n3267), .A2(n3298), .ZN(n3312) );
  NAND2_X1 U3124 ( .A1(n4424), .A2(n4599), .ZN(n4552) );
  AND2_X1 U3125 ( .A1(n3053), .A2(n2983), .ZN(n3093) );
  OR2_X1 U3126 ( .A1(n2605), .A2(n2490), .ZN(n2597) );
  AND2_X1 U3127 ( .A1(n2700), .A2(REG3_REG_19__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U3128 ( .A1(n3107), .A2(n3106), .ZN(n3186) );
  INV_X1 U3129 ( .A(n4197), .ZN(n4203) );
  NAND2_X1 U3130 ( .A1(n2557), .A2(REG3_REG_6__SCAN_IN), .ZN(n2566) );
  AND2_X1 U3131 ( .A1(n2650), .A2(REG3_REG_15__SCAN_IN), .ZN(n2662) );
  OR2_X1 U3132 ( .A1(n2769), .A2(n2763), .ZN(n4110) );
  XNOR2_X1 U3133 ( .A(n2825), .B(n2824), .ZN(n3003) );
  AND2_X1 U3134 ( .A1(n4001), .A2(n3998), .ZN(n4542) );
  OAI21_X1 U3135 ( .B1(n4129), .B2(n2693), .A(n2760), .ZN(n4142) );
  OAI211_X1 U3136 ( .C1(n4244), .C2(n2693), .A(n2712), .B(n2711), .ZN(n4213)
         );
  NAND4_X1 U3137 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(n3557)
         );
  INV_X1 U3138 ( .A(n4293), .ZN(n5045) );
  NAND2_X1 U3139 ( .A1(n3095), .A2(n4264), .ZN(n4290) );
  OAI22_X1 U3140 ( .A1(n2900), .A2(D_REG_0__SCAN_IN), .B1(n2901), .B2(n2840), 
        .ZN(n3092) );
  INV_X1 U3141 ( .A(n4084), .ZN(n2885) );
  NAND2_X1 U3142 ( .A1(n3382), .A2(n4606), .ZN(n4619) );
  AND2_X1 U3143 ( .A1(n2782), .A2(n2783), .ZN(n4639) );
  AND2_X1 U3144 ( .A1(n3054), .A2(n4583), .ZN(n2983) );
  AND2_X1 U3145 ( .A1(n2582), .A2(n2574), .ZN(n4452) );
  AND2_X1 U3146 ( .A1(n2908), .A2(n2923), .ZN(n4541) );
  INV_X1 U3147 ( .A(n3814), .ZN(n4435) );
  OR2_X1 U31480 ( .A1(n2991), .A2(n2982), .ZN(n3816) );
  NAND2_X1 U31490 ( .A1(n3057), .A2(STATE_REG_SCAN_IN), .ZN(n4448) );
  INV_X1 U3150 ( .A(n3692), .ZN(n4102) );
  OAI211_X1 U3151 ( .C1(n4265), .C2(n2693), .A(n2704), .B(n2703), .ZN(n4235)
         );
  NAND4_X1 U3152 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n4557)
         );
  NAND2_X1 U3153 ( .A1(n4001), .A2(n3003), .ZN(n4548) );
  OR2_X1 U3154 ( .A1(n4288), .A2(n4631), .ZN(n4263) );
  NOR2_X1 U3155 ( .A1(n2860), .A2(n3092), .ZN(n4346) );
  NAND2_X1 U3156 ( .A1(n4659), .A2(n4638), .ZN(n4358) );
  INV_X2 U3157 ( .A(n4657), .ZN(n4659) );
  AND3_X1 U3158 ( .A1(n4623), .A2(n4622), .A3(n4621), .ZN(n4654) );
  OR2_X1 U3159 ( .A1(n2860), .A2(n2977), .ZN(n4643) );
  INV_X1 U3160 ( .A(n4582), .ZN(n4581) );
  INV_X1 U3161 ( .A(n2494), .ZN(n4421) );
  INV_X1 U3162 ( .A(n3354), .ZN(n4427) );
  INV_X1 U3163 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2856) );
  NAND2_X1 U3164 ( .A1(n2479), .A2(n2475), .ZN(n2553) );
  NOR2_X2 U3165 ( .A1(n2553), .A2(n2480), .ZN(n2635) );
  AND2_X2 U3166 ( .A1(n4421), .A2(n2493), .ZN(n2531) );
  NAND2_X1 U3167 ( .A1(n2531), .A2(REG3_REG_1__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3168 ( .A1(n2522), .A2(REG2_REG_1__SCAN_IN), .ZN(n2499) );
  NOR2_X1 U3169 ( .A1(n2494), .A2(n2493), .ZN(n2513) );
  INV_X1 U3170 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2496) );
  INV_X1 U3171 ( .A(n3709), .ZN(n2511) );
  NAND2_X1 U3172 ( .A1(n2501), .A2(n2824), .ZN(n2504) );
  NAND2_X1 U3173 ( .A1(n2511), .A2(n3136), .ZN(n3907) );
  NAND2_X1 U3174 ( .A1(n3907), .A2(n3909), .ZN(n2786) );
  NAND2_X1 U3175 ( .A1(n2531), .A2(REG3_REG_0__SCAN_IN), .ZN(n2510) );
  INV_X1 U3176 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3177 ( .A1(n2513), .A2(REG1_REG_0__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3178 ( .A1(n2522), .A2(REG2_REG_0__SCAN_IN), .ZN(n2507) );
  AND2_X1 U3179 ( .A1(n3141), .A2(n3705), .ZN(n3137) );
  NAND2_X1 U3180 ( .A1(n2786), .A2(n3137), .ZN(n3139) );
  NAND2_X1 U3181 ( .A1(n2511), .A2(n3140), .ZN(n2512) );
  NAND2_X1 U3182 ( .A1(n3139), .A2(n2512), .ZN(n3116) );
  INV_X1 U3183 ( .A(n3116), .ZN(n2519) );
  CLKBUF_X3 U3184 ( .A(n2513), .Z(n2817) );
  NAND2_X1 U3185 ( .A1(n2817), .A2(REG1_REG_2__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3186 ( .A1(n2531), .A2(REG3_REG_2__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U3187 ( .A1(n2522), .A2(REG2_REG_2__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U3188 ( .A1(n2702), .A2(REG0_REG_2__SCAN_IN), .ZN(n2514) );
  MUX2_X1 U3189 ( .A(n4432), .B(DATAI_2_), .S(n2529), .Z(n3121) );
  NAND2_X1 U3190 ( .A1(n2993), .A2(n3128), .ZN(n3913) );
  NAND2_X1 U3191 ( .A1(n3144), .A2(n3121), .ZN(n3910) );
  NAND2_X1 U3192 ( .A1(n3913), .A2(n3910), .ZN(n2788) );
  NAND2_X1 U3193 ( .A1(n2519), .A2(n2788), .ZN(n3118) );
  NAND2_X1 U3194 ( .A1(n3144), .A2(n3128), .ZN(n2520) );
  INV_X1 U3195 ( .A(n3169), .ZN(n2543) );
  INV_X1 U3196 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2521) );
  XNOR2_X1 U3197 ( .A(n2521), .B(REG3_REG_3__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U3198 ( .A1(n2531), .A2(n3074), .ZN(n2526) );
  NAND2_X1 U3199 ( .A1(n2702), .A2(REG0_REG_4__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U3200 ( .A1(n2817), .A2(REG1_REG_4__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3201 ( .A1(n2522), .A2(REG2_REG_4__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3202 ( .A1(n2527), .A2(IR_REG_31__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U3203 ( .A1(n2539), .A2(n2538), .ZN(n2541) );
  NAND2_X1 U3204 ( .A1(n2541), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  XNOR2_X1 U3205 ( .A(n2528), .B(IR_REG_4__SCAN_IN), .ZN(n4430) );
  INV_X1 U3206 ( .A(n3159), .ZN(n3078) );
  NAND2_X1 U3207 ( .A1(n2915), .A2(n3078), .ZN(n3919) );
  NAND2_X1 U3208 ( .A1(n3068), .A2(n3159), .ZN(n3916) );
  NAND2_X1 U3209 ( .A1(n2915), .A2(n3159), .ZN(n2545) );
  INV_X1 U32100 ( .A(n2545), .ZN(n2530) );
  INV_X1 U32110 ( .A(n2531), .ZN(n2693) );
  INV_X1 U32120 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32130 ( .A1(n2531), .A2(n2532), .ZN(n2537) );
  INV_X1 U32140 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32150 ( .A1(n2817), .A2(REG1_REG_3__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32160 ( .A1(n2522), .A2(REG2_REG_3__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32170 ( .A1(n2539), .A2(n2538), .ZN(n2540) );
  MUX2_X1 U32180 ( .A(n4431), .B(DATAI_3_), .S(n2529), .Z(n3175) );
  NOR2_X1 U32190 ( .A1(n3997), .A2(n3175), .ZN(n3154) );
  INV_X1 U32200 ( .A(n2544), .ZN(n2547) );
  NAND2_X1 U32210 ( .A1(n3997), .A2(n3175), .ZN(n3155) );
  AOI21_X1 U32220 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2548) );
  NOR2_X1 U32230 ( .A1(n2548), .A2(n2557), .ZN(n3216) );
  NAND2_X1 U32240 ( .A1(n2531), .A2(n3216), .ZN(n2552) );
  NAND2_X1 U32250 ( .A1(n2702), .A2(REG0_REG_5__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32260 ( .A1(n2522), .A2(REG2_REG_5__SCAN_IN), .ZN(n2549) );
  NAND4_X1 U32270 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n3996)
         );
  NAND2_X1 U32280 ( .A1(n2553), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  MUX2_X1 U32290 ( .A(IR_REG_31__SCAN_IN), .B(n2554), .S(IR_REG_5__SCAN_IN), 
        .Z(n2556) );
  INV_X1 U32300 ( .A(n2596), .ZN(n2555) );
  MUX2_X1 U32310 ( .A(n4429), .B(DATAI_5_), .S(n2529), .Z(n3215) );
  OAI21_X1 U32320 ( .B1(n2557), .B2(REG3_REG_6__SCAN_IN), .A(n2566), .ZN(n3208) );
  INV_X1 U32330 ( .A(n3208), .ZN(n5035) );
  NAND2_X1 U32340 ( .A1(n2531), .A2(n5035), .ZN(n2561) );
  NAND2_X1 U32350 ( .A1(n2702), .A2(REG0_REG_6__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32360 ( .A1(n2522), .A2(REG2_REG_6__SCAN_IN), .ZN(n2558) );
  NAND4_X1 U32370 ( .A1(n2561), .A2(n2560), .A3(n2559), .A4(n2558), .ZN(n3995)
         );
  OR2_X1 U32380 ( .A1(n2596), .A2(n2490), .ZN(n2562) );
  XNOR2_X1 U32390 ( .A(n2562), .B(IR_REG_6__SCAN_IN), .ZN(n4428) );
  MUX2_X1 U32400 ( .A(n4428), .B(DATAI_6_), .S(n2529), .Z(n3281) );
  NOR2_X1 U32410 ( .A1(n3995), .A2(n3281), .ZN(n2564) );
  NAND2_X1 U32420 ( .A1(n3995), .A2(n3281), .ZN(n2563) );
  NOR2_X2 U32430 ( .A1(n2566), .A2(n2565), .ZN(n2577) );
  AND2_X1 U32440 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  NOR2_X1 U32450 ( .A1(n2577), .A2(n2567), .ZN(n3232) );
  NAND2_X1 U32460 ( .A1(n2531), .A2(n3232), .ZN(n2571) );
  NAND2_X1 U32470 ( .A1(n2702), .A2(REG0_REG_7__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U32480 ( .A1(n2817), .A2(REG1_REG_7__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U32490 ( .A1(n2522), .A2(REG2_REG_7__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32500 ( .A1(n2596), .A2(n2594), .ZN(n2572) );
  NAND2_X1 U32510 ( .A1(n2572), .A2(IR_REG_31__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32520 ( .A1(n2573), .A2(n4904), .ZN(n2582) );
  OR2_X1 U32530 ( .A1(n2573), .A2(n4904), .ZN(n2574) );
  MUX2_X1 U32540 ( .A(n4452), .B(DATAI_7_), .S(n2529), .Z(n3247) );
  NAND2_X1 U32550 ( .A1(n3262), .A2(n3247), .ZN(n2793) );
  INV_X1 U32560 ( .A(n3247), .ZN(n3239) );
  NAND2_X1 U32570 ( .A1(n3994), .A2(n3239), .ZN(n3925) );
  NAND2_X1 U32580 ( .A1(n2793), .A2(n3925), .ZN(n3885) );
  NAND2_X1 U32590 ( .A1(n3229), .A2(n3885), .ZN(n2576) );
  NAND2_X1 U32600 ( .A1(n3994), .A2(n3247), .ZN(n2575) );
  OR2_X1 U32610 ( .A1(n2577), .A2(REG3_REG_8__SCAN_IN), .ZN(n2578) );
  AND2_X1 U32620 ( .A1(n2587), .A2(n2578), .ZN(n3300) );
  NAND2_X1 U32630 ( .A1(n2531), .A2(n3300), .ZN(n2581) );
  NAND2_X1 U32640 ( .A1(n2702), .A2(REG0_REG_8__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U32650 ( .A1(n2522), .A2(REG2_REG_8__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32660 ( .A1(n2582), .A2(IR_REG_31__SCAN_IN), .ZN(n2583) );
  XNOR2_X1 U32670 ( .A(n2583), .B(IR_REG_8__SCAN_IN), .ZN(n4596) );
  MUX2_X1 U32680 ( .A(n4596), .B(DATAI_8_), .S(n2529), .Z(n3292) );
  AND2_X1 U32690 ( .A1(n3305), .A2(n3292), .ZN(n2585) );
  NAND2_X1 U32700 ( .A1(n2587), .A2(n2586), .ZN(n2588) );
  NAND2_X1 U32710 ( .A1(n2598), .A2(n2588), .ZN(n3310) );
  INV_X1 U32720 ( .A(n3310), .ZN(n3372) );
  NAND2_X1 U32730 ( .A1(n2531), .A2(n3372), .ZN(n2592) );
  NAND2_X1 U32740 ( .A1(n2702), .A2(REG0_REG_9__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U32750 ( .A1(n2817), .A2(REG1_REG_9__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U32760 ( .A1(n2522), .A2(REG2_REG_9__SCAN_IN), .ZN(n2589) );
  NAND4_X1 U32770 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n3993)
         );
  INV_X1 U32780 ( .A(IR_REG_8__SCAN_IN), .ZN(n2593) );
  XNOR2_X1 U32790 ( .A(n2597), .B(IR_REG_9__SCAN_IN), .ZN(n3336) );
  MUX2_X1 U32800 ( .A(n3336), .B(DATAI_9_), .S(n2529), .Z(n3371) );
  INV_X1 U32810 ( .A(n3371), .ZN(n3413) );
  NAND2_X1 U32820 ( .A1(n2598), .A2(n3403), .ZN(n2599) );
  AND2_X1 U32830 ( .A1(n2609), .A2(n2599), .ZN(n3386) );
  NAND2_X1 U32840 ( .A1(n2531), .A2(n3386), .ZN(n2603) );
  NAND2_X1 U32850 ( .A1(n2702), .A2(REG0_REG_10__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U32860 ( .A1(n2817), .A2(REG1_REG_10__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U32870 ( .A1(n2522), .A2(REG2_REG_10__SCAN_IN), .ZN(n2600) );
  NAND4_X1 U32880 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n3992)
         );
  INV_X1 U32890 ( .A(IR_REG_9__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U32900 ( .A1(n2605), .A2(n2604), .ZN(n2615) );
  NAND2_X1 U32910 ( .A1(n2615), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  XNOR2_X1 U32920 ( .A(n2606), .B(IR_REG_10__SCAN_IN), .ZN(n4592) );
  MUX2_X1 U32930 ( .A(n4592), .B(DATAI_10_), .S(n2529), .Z(n3406) );
  AND2_X1 U32940 ( .A1(n3992), .A2(n3406), .ZN(n2607) );
  INV_X1 U32950 ( .A(n3406), .ZN(n3384) );
  NOR2_X2 U32960 ( .A1(n2609), .A2(n2608), .ZN(n2620) );
  AND2_X1 U32970 ( .A1(n2609), .A2(n2608), .ZN(n2610) );
  NOR2_X1 U32980 ( .A1(n2620), .A2(n2610), .ZN(n4564) );
  NAND2_X1 U32990 ( .A1(n2531), .A2(n4564), .ZN(n2614) );
  NAND2_X1 U33000 ( .A1(n2702), .A2(REG0_REG_11__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33010 ( .A1(n2817), .A2(REG1_REG_11__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U33020 ( .A1(n2522), .A2(REG2_REG_11__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33030 ( .A1(n2616), .A2(IR_REG_31__SCAN_IN), .ZN(n2617) );
  OR2_X1 U33040 ( .A1(n2617), .A2(n4868), .ZN(n2618) );
  NAND2_X1 U33050 ( .A1(n2617), .A2(n4868), .ZN(n2626) );
  MUX2_X1 U33060 ( .A(n3334), .B(DATAI_11_), .S(n2529), .Z(n4567) );
  NAND2_X1 U33070 ( .A1(n3451), .A2(n4567), .ZN(n3420) );
  INV_X1 U33080 ( .A(n4567), .ZN(n4553) );
  NAND2_X1 U33090 ( .A1(n3991), .A2(n4553), .ZN(n3422) );
  NAND2_X1 U33100 ( .A1(n3420), .A2(n3422), .ZN(n4550) );
  NAND2_X1 U33110 ( .A1(n3451), .A2(n4553), .ZN(n2619) );
  OR2_X1 U33120 ( .A1(n2620), .A2(REG3_REG_12__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U33130 ( .A1(n2620), .A2(REG3_REG_12__SCAN_IN), .ZN(n2629) );
  AND2_X1 U33140 ( .A1(n2621), .A2(n2629), .ZN(n3467) );
  NAND2_X1 U33150 ( .A1(n2531), .A2(n3467), .ZN(n2625) );
  NAND2_X1 U33160 ( .A1(n2702), .A2(REG0_REG_12__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33170 ( .A1(n2817), .A2(REG1_REG_12__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U33180 ( .A1(n2522), .A2(REG2_REG_12__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U33190 ( .A1(n2626), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  XNOR2_X1 U33200 ( .A(n2627), .B(IR_REG_12__SCAN_IN), .ZN(n4588) );
  MUX2_X1 U33210 ( .A(n4588), .B(DATAI_12_), .S(n2529), .Z(n3461) );
  NAND2_X1 U33220 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
  AND2_X1 U33230 ( .A1(n2642), .A2(n2630), .ZN(n3578) );
  NAND2_X1 U33240 ( .A1(n2531), .A2(n3578), .ZN(n2634) );
  NAND2_X1 U33250 ( .A1(n2702), .A2(REG0_REG_13__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U33260 ( .A1(n2817), .A2(REG1_REG_13__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U33270 ( .A1(n2522), .A2(REG2_REG_13__SCAN_IN), .ZN(n2631) );
  NOR2_X1 U33280 ( .A1(n2635), .A2(n2490), .ZN(n2636) );
  MUX2_X1 U33290 ( .A(n2490), .B(n2636), .S(IR_REG_13__SCAN_IN), .Z(n2638) );
  OR2_X1 U33300 ( .A1(n2638), .A2(n2682), .ZN(n3354) );
  MUX2_X1 U33310 ( .A(n4427), .B(DATAI_13_), .S(n2529), .Z(n3541) );
  AND2_X1 U33320 ( .A1(n3557), .A2(n3541), .ZN(n2640) );
  INV_X1 U33330 ( .A(n3557), .ZN(n3487) );
  NAND2_X1 U33340 ( .A1(n3487), .A2(n3576), .ZN(n2639) );
  OAI21_X1 U33350 ( .B1(n3428), .B2(n2640), .A(n2639), .ZN(n3482) );
  AND2_X1 U33360 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  NOR2_X1 U33370 ( .A1(n2650), .A2(n2643), .ZN(n3562) );
  NAND2_X1 U33380 ( .A1(n2531), .A2(n3562), .ZN(n2647) );
  NAND2_X1 U33390 ( .A1(n2702), .A2(REG0_REG_14__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U33400 ( .A1(n2522), .A2(REG2_REG_14__SCAN_IN), .ZN(n2644) );
  OR2_X1 U33410 ( .A1(n2682), .A2(n2490), .ZN(n2648) );
  XNOR2_X1 U33420 ( .A(n2648), .B(IR_REG_14__SCAN_IN), .ZN(n4426) );
  MUX2_X1 U33430 ( .A(n4426), .B(DATAI_14_), .S(n2529), .Z(n3555) );
  NAND2_X1 U33440 ( .A1(n3824), .A2(n3555), .ZN(n3831) );
  INV_X1 U33450 ( .A(n3824), .ZN(n3990) );
  INV_X1 U33460 ( .A(n3555), .ZN(n3560) );
  NAND2_X1 U33470 ( .A1(n3990), .A2(n3560), .ZN(n3832) );
  NAND2_X1 U33480 ( .A1(n3831), .A2(n3832), .ZN(n3892) );
  NAND2_X1 U33490 ( .A1(n3824), .A2(n3560), .ZN(n2649) );
  NOR2_X1 U33500 ( .A1(n2650), .A2(REG3_REG_15__SCAN_IN), .ZN(n2651) );
  OR2_X1 U33510 ( .A1(n2662), .A2(n2651), .ZN(n3829) );
  INV_X1 U33520 ( .A(n3829), .ZN(n2652) );
  NAND2_X1 U3353 ( .A1(n2531), .A2(n2652), .ZN(n2656) );
  NAND2_X1 U33540 ( .A1(n2702), .A2(REG0_REG_15__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3355 ( .A1(n2817), .A2(REG1_REG_15__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3356 ( .A1(n2522), .A2(REG2_REG_15__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3357 ( .A1(n2682), .A2(n2680), .ZN(n2657) );
  NAND2_X1 U3358 ( .A1(n2657), .A2(IR_REG_31__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3359 ( .A1(n2658), .A2(n4889), .ZN(n2669) );
  OR2_X1 U3360 ( .A1(n2658), .A2(n4889), .ZN(n2659) );
  MUX2_X1 U3361 ( .A(n4047), .B(DATAI_15_), .S(n2529), .Z(n3826) );
  NAND2_X1 U3362 ( .A1(n3612), .A2(n3826), .ZN(n2660) );
  NAND2_X1 U3363 ( .A1(n2661), .A2(n2660), .ZN(n3524) );
  OR2_X1 U3364 ( .A1(n2662), .A2(REG3_REG_16__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3365 ( .A1(n2673), .A2(n2663), .ZN(n4447) );
  INV_X1 U3366 ( .A(n4447), .ZN(n2664) );
  NAND2_X1 U3367 ( .A1(n2531), .A2(n2664), .ZN(n2668) );
  NAND2_X1 U3368 ( .A1(n2702), .A2(REG0_REG_16__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3369 ( .A1(n2817), .A2(REG1_REG_16__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3370 ( .A1(n2522), .A2(REG2_REG_16__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3371 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  XNOR2_X1 U3372 ( .A(n2670), .B(IR_REG_16__SCAN_IN), .ZN(n4048) );
  MUX2_X1 U3373 ( .A(n4048), .B(DATAI_16_), .S(n2529), .Z(n4439) );
  NAND2_X1 U3374 ( .A1(n3823), .A2(n4439), .ZN(n3952) );
  NAND2_X1 U3375 ( .A1(n3989), .A2(n3617), .ZN(n3836) );
  NAND2_X1 U3376 ( .A1(n3952), .A2(n3836), .ZN(n3525) );
  NAND2_X1 U3377 ( .A1(n3524), .A2(n3525), .ZN(n3523) );
  NAND2_X1 U3378 ( .A1(n3989), .A2(n4439), .ZN(n2671) );
  NAND2_X1 U3379 ( .A1(n3523), .A2(n2671), .ZN(n3600) );
  NAND2_X1 U3380 ( .A1(n2673), .A2(n2672), .ZN(n2674) );
  AND2_X1 U3381 ( .A1(n2691), .A2(n2674), .ZN(n3761) );
  NAND2_X1 U3382 ( .A1(n2531), .A2(n3761), .ZN(n2678) );
  NAND2_X1 U3383 ( .A1(n2702), .A2(REG0_REG_17__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3384 ( .A1(n2817), .A2(REG1_REG_17__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3385 ( .A1(n2522), .A2(REG2_REG_17__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3386 ( .A1(n2682), .A2(n2681), .ZN(n2684) );
  NAND2_X1 U3387 ( .A1(n2684), .A2(IR_REG_31__SCAN_IN), .ZN(n2683) );
  MUX2_X1 U3388 ( .A(IR_REG_31__SCAN_IN), .B(n2683), .S(IR_REG_17__SCAN_IN), 
        .Z(n2686) );
  INV_X1 U3389 ( .A(DATAI_17_), .ZN(n2687) );
  MUX2_X1 U3390 ( .A(n4584), .B(n2687), .S(n2529), .Z(n4354) );
  NAND2_X1 U3391 ( .A1(n4436), .A2(n4354), .ZN(n2688) );
  INV_X1 U3392 ( .A(n4354), .ZN(n3760) );
  NAND2_X1 U3393 ( .A1(n4281), .A2(n3760), .ZN(n2689) );
  AND2_X1 U3394 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  OR2_X1 U3395 ( .A1(n2692), .A2(n2700), .ZN(n3800) );
  NAND2_X1 U3396 ( .A1(n2522), .A2(REG2_REG_18__SCAN_IN), .ZN(n2694) );
  OAI21_X1 U3397 ( .B1(n3800), .B2(n2693), .A(n2694), .ZN(n2695) );
  INV_X1 U3398 ( .A(n2695), .ZN(n2696) );
  NAND2_X1 U3399 ( .A1(n2249), .A2(IR_REG_31__SCAN_IN), .ZN(n2698) );
  XNOR2_X1 U3400 ( .A(n2698), .B(IR_REG_18__SCAN_IN), .ZN(n4064) );
  MUX2_X1 U3401 ( .A(n4064), .B(DATAI_18_), .S(n2529), .Z(n2857) );
  NAND2_X1 U3402 ( .A1(n3758), .A2(n2857), .ZN(n4249) );
  INV_X1 U3403 ( .A(n3758), .ZN(n4257) );
  NAND2_X1 U3404 ( .A1(n4257), .A2(n4285), .ZN(n4250) );
  NAND2_X1 U3405 ( .A1(n4249), .A2(n4250), .ZN(n4276) );
  INV_X1 U3406 ( .A(n4276), .ZN(n4273) );
  NAND2_X1 U3407 ( .A1(n3758), .A2(n4285), .ZN(n2699) );
  NOR2_X1 U3408 ( .A1(n2700), .A2(REG3_REG_19__SCAN_IN), .ZN(n2701) );
  OR2_X1 U3409 ( .A1(n2709), .A2(n2701), .ZN(n4265) );
  NAND2_X1 U3410 ( .A1(n2522), .A2(REG2_REG_19__SCAN_IN), .ZN(n2703) );
  OR2_X1 U3411 ( .A1(n2705), .A2(n4772), .ZN(n2706) );
  INV_X1 U3412 ( .A(n4069), .ZN(n4425) );
  MUX2_X1 U3413 ( .A(n4425), .B(DATAI_19_), .S(n2529), .Z(n4256) );
  NAND2_X1 U3414 ( .A1(n4235), .A2(n4256), .ZN(n2707) );
  OR2_X1 U3415 ( .A1(n4235), .A2(n4256), .ZN(n2708) );
  OR2_X1 U3416 ( .A1(n2709), .A2(REG3_REG_20__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U3417 ( .A1(n2721), .A2(n2710), .ZN(n4244) );
  AOI22_X1 U3418 ( .A1(n2702), .A2(REG0_REG_20__SCAN_IN), .B1(n2817), .B2(
        REG1_REG_20__SCAN_IN), .ZN(n2712) );
  NAND2_X1 U3419 ( .A1(n2522), .A2(REG2_REG_20__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3420 ( .A1(n4213), .A2(n4242), .ZN(n3868) );
  NAND2_X1 U3421 ( .A1(n4226), .A2(n3868), .ZN(n2713) );
  OR2_X1 U3422 ( .A1(n4213), .A2(n4242), .ZN(n3869) );
  NAND2_X1 U3423 ( .A1(n2713), .A2(n3869), .ZN(n4217) );
  XNOR2_X1 U3424 ( .A(n2721), .B(REG3_REG_21__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U3425 ( .A1(n4220), .A2(n2531), .ZN(n2718) );
  INV_X1 U3426 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U3427 ( .A1(n2817), .A2(REG1_REG_21__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3428 ( .A1(n2522), .A2(REG2_REG_21__SCAN_IN), .ZN(n2714) );
  OAI211_X1 U3429 ( .C1(n2725), .C2(n4405), .A(n2715), .B(n2714), .ZN(n2716)
         );
  INV_X1 U3430 ( .A(n2716), .ZN(n2717) );
  NAND2_X1 U3431 ( .A1(n4236), .A2(n3650), .ZN(n2719) );
  INV_X1 U3432 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3738) );
  INV_X1 U3433 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2720) );
  OAI21_X1 U3434 ( .B1(n2721), .B2(n3738), .A(n2720), .ZN(n2722) );
  AND2_X1 U3435 ( .A1(n2722), .A2(n2731), .ZN(n4204) );
  NAND2_X1 U3436 ( .A1(n4204), .A2(n2531), .ZN(n2728) );
  INV_X1 U3437 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U3438 ( .A1(n2817), .A2(REG1_REG_22__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3439 ( .A1(n2522), .A2(REG2_REG_22__SCAN_IN), .ZN(n2723) );
  OAI211_X1 U3440 ( .C1(n2725), .C2(n4401), .A(n2724), .B(n2723), .ZN(n2726)
         );
  INV_X1 U3441 ( .A(n2726), .ZN(n2727) );
  NAND2_X1 U3442 ( .A1(n2529), .A2(DATAI_22_), .ZN(n4197) );
  NAND2_X1 U3443 ( .A1(n3739), .A2(n4203), .ZN(n4176) );
  NAND2_X1 U3444 ( .A1(n4214), .A2(n4197), .ZN(n2811) );
  NAND2_X1 U3445 ( .A1(n4176), .A2(n2811), .ZN(n4200) );
  INV_X1 U3446 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3722) );
  AND2_X1 U3447 ( .A1(n2731), .A2(n3722), .ZN(n2732) );
  OR2_X1 U3448 ( .A1(n2732), .A2(n2738), .ZN(n3721) );
  INV_X1 U3449 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U3450 ( .A1(n2817), .A2(REG1_REG_23__SCAN_IN), .ZN(n2734) );
  NAND2_X1 U3451 ( .A1(n2522), .A2(REG2_REG_23__SCAN_IN), .ZN(n2733) );
  OAI211_X1 U3452 ( .C1(n2725), .C2(n4395), .A(n2734), .B(n2733), .ZN(n2735)
         );
  INV_X1 U3453 ( .A(n2735), .ZN(n2736) );
  NOR2_X1 U3454 ( .A1(n4194), .A2(n4180), .ZN(n2737) );
  INV_X1 U3455 ( .A(n4194), .ZN(n3771) );
  NAND2_X1 U3456 ( .A1(n2738), .A2(REG3_REG_24__SCAN_IN), .ZN(n2746) );
  OR2_X1 U3457 ( .A1(n2738), .A2(REG3_REG_24__SCAN_IN), .ZN(n2739) );
  AND2_X1 U34580 ( .A1(n2746), .A2(n2739), .ZN(n4167) );
  NAND2_X1 U34590 ( .A1(n4167), .A2(n2531), .ZN(n2744) );
  INV_X1 U3460 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U3461 ( .A1(n2817), .A2(REG1_REG_24__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U3462 ( .A1(n2522), .A2(REG2_REG_24__SCAN_IN), .ZN(n2740) );
  OAI211_X1 U3463 ( .C1(n2725), .C2(n4391), .A(n2741), .B(n2740), .ZN(n2742)
         );
  INV_X1 U3464 ( .A(n2742), .ZN(n2743) );
  NAND2_X1 U3465 ( .A1(n2529), .A2(DATAI_24_), .ZN(n4166) );
  INV_X1 U3466 ( .A(n4166), .ZN(n4160) );
  INV_X1 U34670 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3749) );
  NAND2_X1 U3468 ( .A1(n2746), .A2(n3749), .ZN(n2747) );
  NAND2_X1 U34690 ( .A1(n4146), .A2(n2531), .ZN(n2752) );
  INV_X1 U3470 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U34710 ( .A1(n2817), .A2(REG1_REG_25__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U3472 ( .A1(n2522), .A2(REG2_REG_25__SCAN_IN), .ZN(n2748) );
  OAI211_X1 U34730 ( .C1(n2725), .C2(n4387), .A(n2749), .B(n2748), .ZN(n2750)
         );
  INV_X1 U3474 ( .A(n2750), .ZN(n2751) );
  INV_X1 U34750 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2754) );
  AND2_X1 U3476 ( .A1(n2755), .A2(n2754), .ZN(n2756) );
  INV_X1 U34770 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U3478 ( .A1(n2817), .A2(REG1_REG_26__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U34790 ( .A1(n2522), .A2(REG2_REG_26__SCAN_IN), .ZN(n2757) );
  OAI211_X1 U3480 ( .C1(n2725), .C2(n4383), .A(n2758), .B(n2757), .ZN(n2759)
         );
  INV_X1 U34810 ( .A(n2759), .ZN(n2760) );
  NAND2_X1 U3482 ( .A1(n2529), .A2(DATAI_26_), .ZN(n4127) );
  AND2_X1 U34830 ( .A1(n4142), .A2(n4121), .ZN(n3902) );
  INV_X1 U3484 ( .A(n4142), .ZN(n2761) );
  NAND2_X1 U34850 ( .A1(n2761), .A2(n4127), .ZN(n3903) );
  NOR2_X1 U3486 ( .A1(n2762), .A2(REG3_REG_27__SCAN_IN), .ZN(n2763) );
  INV_X1 U34870 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U3488 ( .A1(n2817), .A2(REG1_REG_27__SCAN_IN), .ZN(n2765) );
  NAND2_X1 U34890 ( .A1(n2522), .A2(REG2_REG_27__SCAN_IN), .ZN(n2764) );
  OAI211_X1 U3490 ( .C1(n2725), .C2(n4379), .A(n2765), .B(n2764), .ZN(n2766)
         );
  INV_X1 U34910 ( .A(n2766), .ZN(n2767) );
  OAI21_X2 U3492 ( .B1(n4110), .B2(n2693), .A(n2767), .ZN(n3988) );
  NOR2_X1 U34930 ( .A1(n3988), .A2(n4108), .ZN(n2768) );
  INV_X1 U3494 ( .A(n3988), .ZN(n4125) );
  NAND2_X1 U34950 ( .A1(n2769), .A2(REG3_REG_28__SCAN_IN), .ZN(n4083) );
  OR2_X1 U3496 ( .A1(n2769), .A2(REG3_REG_28__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U34970 ( .A1(n3697), .A2(n2531), .ZN(n2775) );
  INV_X1 U3498 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2862) );
  NAND2_X1 U34990 ( .A1(n2817), .A2(REG1_REG_28__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U3500 ( .A1(n2522), .A2(REG2_REG_28__SCAN_IN), .ZN(n2771) );
  OAI211_X1 U35010 ( .C1(n2725), .C2(n2862), .A(n2772), .B(n2771), .ZN(n2773)
         );
  INV_X1 U3502 ( .A(n2773), .ZN(n2774) );
  NOR2_X1 U35030 ( .A1(n3692), .A2(n4092), .ZN(n3850) );
  XNOR2_X1 U3504 ( .A(n2865), .B(n2776), .ZN(n4090) );
  NAND2_X1 U35050 ( .A1(n2258), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U35060 ( .A1(n2831), .A2(IR_REG_31__SCAN_IN), .ZN(n2780) );
  XNOR2_X1 U35070 ( .A(n2966), .B(n3982), .ZN(n2781) );
  NAND2_X1 U35080 ( .A1(n2781), .A2(n4069), .ZN(n3382) );
  NOR2_X1 U35090 ( .A1(n4069), .A2(n3982), .ZN(n2783) );
  INV_X1 U35100 ( .A(n4639), .ZN(n4606) );
  INV_X1 U35110 ( .A(n2782), .ZN(n4424) );
  INV_X1 U35120 ( .A(n3982), .ZN(n2784) );
  INV_X1 U35130 ( .A(n4423), .ZN(n3877) );
  NAND2_X1 U35140 ( .A1(n4424), .A2(n4423), .ZN(n3861) );
  OR2_X1 U35150 ( .A1(n4069), .A2(n2784), .ZN(n2785) );
  NAND2_X2 U35160 ( .A1(n3861), .A2(n2785), .ZN(n4254) );
  INV_X1 U35170 ( .A(n3141), .ZN(n2787) );
  NAND2_X1 U35180 ( .A1(n2787), .A2(n3705), .ZN(n3906) );
  NAND2_X1 U35190 ( .A1(n3161), .A2(n3175), .ZN(n3915) );
  INV_X1 U35200 ( .A(n3175), .ZN(n2789) );
  NAND2_X1 U35210 ( .A1(n3997), .A2(n2789), .ZN(n3912) );
  NAND2_X1 U35220 ( .A1(n3170), .A2(n3888), .ZN(n2790) );
  INV_X1 U35230 ( .A(n3916), .ZN(n2791) );
  AND2_X1 U35240 ( .A1(n3996), .A2(n3252), .ZN(n3209) );
  INV_X1 U35250 ( .A(n3996), .ZN(n3203) );
  NAND2_X1 U35260 ( .A1(n3203), .A2(n3215), .ZN(n3934) );
  INV_X1 U35270 ( .A(n3281), .ZN(n5038) );
  NAND2_X1 U35280 ( .A1(n3995), .A2(n5038), .ZN(n3935) );
  NAND2_X1 U35290 ( .A1(n3275), .A2(n3935), .ZN(n2792) );
  INV_X1 U35300 ( .A(n3995), .ZN(n3245) );
  NAND2_X1 U35310 ( .A1(n3245), .A2(n3281), .ZN(n3921) );
  NAND2_X1 U35320 ( .A1(n2794), .A2(n3925), .ZN(n3260) );
  NAND2_X1 U35330 ( .A1(n3369), .A2(n3292), .ZN(n3927) );
  NAND2_X1 U35340 ( .A1(n3305), .A2(n3298), .ZN(n3924) );
  AND2_X1 U35350 ( .A1(n3993), .A2(n3413), .ZN(n3932) );
  NAND2_X1 U35360 ( .A1(n3404), .A2(n3371), .ZN(n3926) );
  NAND2_X1 U35370 ( .A1(n3992), .A2(n3384), .ZN(n3942) );
  NAND2_X1 U35380 ( .A1(n3377), .A2(n3942), .ZN(n2795) );
  NAND2_X1 U35390 ( .A1(n4555), .A2(n3406), .ZN(n3941) );
  NAND2_X1 U35400 ( .A1(n4557), .A2(n3582), .ZN(n3434) );
  NAND2_X1 U35410 ( .A1(n3557), .A2(n3576), .ZN(n2796) );
  NAND2_X1 U35420 ( .A1(n3434), .A2(n2796), .ZN(n2799) );
  INV_X1 U35430 ( .A(n3422), .ZN(n2797) );
  NOR2_X1 U35440 ( .A1(n2799), .A2(n2797), .ZN(n3943) );
  NAND2_X1 U35450 ( .A1(n2798), .A2(n3461), .ZN(n3435) );
  NAND2_X1 U35460 ( .A1(n3420), .A2(n3435), .ZN(n2802) );
  INV_X1 U35470 ( .A(n2799), .ZN(n2801) );
  NOR2_X1 U35480 ( .A1(n3557), .A2(n3576), .ZN(n2800) );
  AOI21_X1 U35490 ( .B1(n2802), .B2(n2801), .A(n2800), .ZN(n3946) );
  INV_X1 U35500 ( .A(n3892), .ZN(n3483) );
  INV_X1 U35510 ( .A(n3612), .ZN(n4433) );
  NAND2_X1 U35520 ( .A1(n4433), .A2(n3826), .ZN(n3834) );
  INV_X1 U35530 ( .A(n3826), .ZN(n3609) );
  NAND2_X1 U35540 ( .A1(n3612), .A2(n3609), .ZN(n3833) );
  NAND2_X1 U35550 ( .A1(n3834), .A2(n3833), .ZN(n3891) );
  INV_X1 U35560 ( .A(n3831), .ZN(n2803) );
  NOR2_X1 U35570 ( .A1(n3891), .A2(n2803), .ZN(n2804) );
  NAND2_X1 U35580 ( .A1(n3511), .A2(n2804), .ZN(n2805) );
  INV_X1 U35590 ( .A(n3525), .ZN(n3889) );
  INV_X1 U35600 ( .A(n4256), .ZN(n4262) );
  NAND2_X1 U35610 ( .A1(n4235), .A2(n4262), .ZN(n2806) );
  AND2_X1 U35620 ( .A1(n2806), .A2(n4250), .ZN(n4232) );
  NAND2_X1 U35630 ( .A1(n4213), .A2(n3782), .ZN(n2809) );
  NAND2_X1 U35640 ( .A1(n4281), .A2(n4354), .ZN(n4227) );
  NAND3_X1 U35650 ( .A1(n4232), .A2(n2809), .A3(n4227), .ZN(n3953) );
  INV_X1 U35660 ( .A(n4232), .ZN(n2807) );
  OAI22_X1 U35670 ( .A1(n2807), .A2(n4249), .B1(n4235), .B2(n4262), .ZN(n4231)
         );
  NAND2_X1 U35680 ( .A1(n4436), .A2(n3760), .ZN(n4228) );
  OAI22_X1 U35690 ( .A1(n2807), .A2(n4228), .B1(n4213), .B2(n3782), .ZN(n2808)
         );
  OR2_X1 U35700 ( .A1(n4231), .A2(n2808), .ZN(n2810) );
  NAND2_X1 U35710 ( .A1(n2810), .A2(n2809), .ZN(n4173) );
  INV_X1 U35720 ( .A(n3650), .ZN(n4335) );
  OR2_X1 U35730 ( .A1(n4236), .A2(n4335), .ZN(n4175) );
  AND2_X1 U35740 ( .A1(n4176), .A2(n4175), .ZN(n3959) );
  AND2_X1 U35750 ( .A1(n4173), .A2(n3959), .ZN(n3838) );
  NAND2_X1 U35760 ( .A1(n4174), .A2(n3838), .ZN(n2813) );
  NAND2_X1 U35770 ( .A1(n4194), .A2(n4186), .ZN(n3867) );
  NAND2_X1 U35780 ( .A1(n3867), .A2(n2811), .ZN(n3830) );
  AND2_X1 U35790 ( .A1(n4236), .A2(n4335), .ZN(n3960) );
  AND2_X1 U35800 ( .A1(n4176), .A2(n3960), .ZN(n3841) );
  NOR2_X1 U35810 ( .A1(n3830), .A2(n3841), .ZN(n2812) );
  NAND2_X1 U3582 ( .A1(n4183), .A2(n4160), .ZN(n3899) );
  OR2_X1 U3583 ( .A1(n4194), .A2(n4186), .ZN(n4155) );
  AND2_X1 U3584 ( .A1(n4141), .A2(n4166), .ZN(n3898) );
  NOR2_X1 U3585 ( .A1(n4163), .A2(n4147), .ZN(n3866) );
  INV_X1 U3586 ( .A(n3866), .ZN(n2814) );
  OR2_X1 U3587 ( .A1(n4142), .A2(n4127), .ZN(n2815) );
  NAND2_X1 U3588 ( .A1(n4163), .A2(n4147), .ZN(n4116) );
  NAND2_X1 U3589 ( .A1(n2815), .A2(n4116), .ZN(n3962) );
  INV_X1 U3590 ( .A(n3962), .ZN(n3856) );
  NAND2_X1 U3591 ( .A1(n4142), .A2(n4127), .ZN(n3851) );
  INV_X1 U3592 ( .A(n3851), .ZN(n3967) );
  XNOR2_X1 U3593 ( .A(n3988), .B(n4108), .ZN(n4105) );
  NAND2_X1 U3594 ( .A1(n4101), .A2(n4105), .ZN(n4100) );
  NOR2_X1 U3595 ( .A1(n3988), .A2(n4305), .ZN(n3843) );
  INV_X1 U3596 ( .A(n3843), .ZN(n2816) );
  XOR2_X1 U3597 ( .A(n3864), .B(n2873), .Z(n2826) );
  OR2_X1 U3598 ( .A1(n4083), .A2(n2693), .ZN(n2822) );
  INV_X1 U3599 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2883) );
  NAND2_X1 U3600 ( .A1(n2817), .A2(REG1_REG_29__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U3601 ( .A1(n2522), .A2(REG2_REG_29__SCAN_IN), .ZN(n2818) );
  OAI211_X1 U3602 ( .C1(n2725), .C2(n2883), .A(n2819), .B(n2818), .ZN(n2820)
         );
  INV_X1 U3603 ( .A(n2820), .ZN(n2821) );
  NAND2_X1 U3604 ( .A1(n2823), .A2(IR_REG_31__SCAN_IN), .ZN(n2825) );
  AOI222_X1 U3605 ( .A1(n4254), .A2(n2826), .B1(n3987), .B2(n4558), .C1(n3988), 
        .C2(n4282), .ZN(n4099) );
  OAI21_X1 U3606 ( .B1(n3690), .B2(n4552), .A(n4099), .ZN(n2827) );
  AOI21_X1 U3607 ( .B1(n4090), .B2(n4619), .A(n2827), .ZN(n2861) );
  NAND2_X1 U3608 ( .A1(n2297), .A2(IR_REG_31__SCAN_IN), .ZN(n2828) );
  MUX2_X1 U3609 ( .A(IR_REG_31__SCAN_IN), .B(n2828), .S(IR_REG_25__SCAN_IN), 
        .Z(n2830) );
  NAND2_X1 U3610 ( .A1(n2839), .A2(B_REG_SCAN_IN), .ZN(n2835) );
  MUX2_X1 U3611 ( .A(n2835), .B(B_REG_SCAN_IN), .S(n2840), .Z(n2837) );
  INV_X1 U3612 ( .A(n2901), .ZN(n2904) );
  NAND2_X1 U3613 ( .A1(n2904), .A2(n2839), .ZN(n2838) );
  OAI21_X1 U3614 ( .B1(n2900), .B2(D_REG_1__SCAN_IN), .A(n2838), .ZN(n2976) );
  NAND2_X1 U3615 ( .A1(n2782), .A2(n4069), .ZN(n2978) );
  NAND2_X1 U3616 ( .A1(n2978), .A2(n2979), .ZN(n3053) );
  INV_X1 U3617 ( .A(n2839), .ZN(n4422) );
  NAND2_X1 U3618 ( .A1(n2842), .A2(IR_REG_23__SCAN_IN), .ZN(n2844) );
  NAND2_X1 U3619 ( .A1(n2844), .A2(n2843), .ZN(n3052) );
  INV_X1 U3620 ( .A(n2900), .ZN(n2855) );
  NOR4_X1 U3621 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2853) );
  NOR4_X1 U3622 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2852) );
  INV_X1 U3623 ( .A(D_REG_27__SCAN_IN), .ZN(n4769) );
  INV_X1 U3624 ( .A(D_REG_26__SCAN_IN), .ZN(n4579) );
  INV_X1 U3625 ( .A(D_REG_17__SCAN_IN), .ZN(n4580) );
  INV_X1 U3626 ( .A(D_REG_13__SCAN_IN), .ZN(n4773) );
  NAND4_X1 U3627 ( .A1(n4769), .A2(n4579), .A3(n4580), .A4(n4773), .ZN(n2850)
         );
  NOR4_X1 U3628 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2848) );
  NOR4_X1 U3629 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2847) );
  NOR4_X1 U3630 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2846) );
  NOR4_X1 U3631 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2845) );
  NAND4_X1 U3632 ( .A1(n2848), .A2(n2847), .A3(n2846), .A4(n2845), .ZN(n2849)
         );
  NOR4_X1 U3633 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2850), 
        .A4(n2849), .ZN(n2851) );
  NAND3_X1 U3634 ( .A1(n2853), .A2(n2852), .A3(n2851), .ZN(n2854) );
  NAND2_X1 U3635 ( .A1(n2855), .A2(n2854), .ZN(n3091) );
  NAND2_X1 U3636 ( .A1(n4639), .A2(n3877), .ZN(n2985) );
  NAND4_X1 U3637 ( .A1(n2976), .A2(n3093), .A3(n3091), .A4(n2985), .ZN(n2860)
         );
  MUX2_X1 U3638 ( .A(n2856), .B(n2861), .S(n4659), .Z(n2859) );
  INV_X1 U3639 ( .A(n2876), .ZN(n2877) );
  OAI21_X1 U3640 ( .B1(n4106), .B2(n3690), .A(n2877), .ZN(n4091) );
  NAND2_X1 U3641 ( .A1(n2859), .A2(n2858), .ZN(U3546) );
  INV_X1 U3642 ( .A(n3092), .ZN(n2977) );
  INV_X2 U3643 ( .A(n4643), .ZN(n4645) );
  MUX2_X1 U3644 ( .A(n2862), .B(n2861), .S(n4645), .Z(n2864) );
  NAND2_X1 U3645 ( .A1(n2864), .A2(n2863), .ZN(U3514) );
  INV_X1 U3646 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2875) );
  AOI22_X1 U3647 ( .A1(n2865), .A2(n3864), .B1(n4092), .B2(n4102), .ZN(n2866)
         );
  NAND2_X1 U3648 ( .A1(n2529), .A2(DATAI_29_), .ZN(n3848) );
  XOR2_X1 U3649 ( .A(n3848), .B(n3987), .Z(n3875) );
  XNOR2_X1 U3650 ( .A(n2866), .B(n2437), .ZN(n4080) );
  INV_X1 U3651 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2869) );
  NAND2_X1 U3652 ( .A1(n2817), .A2(REG1_REG_30__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U3653 ( .A1(n2522), .A2(REG2_REG_30__SCAN_IN), .ZN(n2867) );
  OAI211_X1 U3654 ( .C1(n2725), .C2(n2869), .A(n2868), .B(n2867), .ZN(n3845)
         );
  XNOR2_X1 U3655 ( .A(n2870), .B(IR_REG_27__SCAN_IN), .ZN(n3004) );
  NAND2_X1 U3656 ( .A1(n3004), .A2(B_REG_SCAN_IN), .ZN(n2871) );
  AND2_X1 U3657 ( .A1(n4558), .A2(n2871), .ZN(n4075) );
  INV_X1 U3658 ( .A(n3850), .ZN(n2872) );
  OAI21_X1 U3659 ( .B1(n3848), .B2(n4552), .A(n4082), .ZN(n2874) );
  AOI21_X1 U3660 ( .B1(n4080), .B2(n4619), .A(n2874), .ZN(n2882) );
  MUX2_X1 U3661 ( .A(n2875), .B(n2882), .S(n4659), .Z(n2881) );
  INV_X1 U3662 ( .A(n3848), .ZN(n4081) );
  NAND2_X1 U3663 ( .A1(n2877), .A2(n4081), .ZN(n2878) );
  NAND2_X1 U3664 ( .A1(n4297), .A2(n2878), .ZN(n4084) );
  NAND2_X1 U3665 ( .A1(n2885), .A2(n2879), .ZN(n2880) );
  NAND2_X1 U3666 ( .A1(n2881), .A2(n2880), .ZN(U3547) );
  MUX2_X1 U3667 ( .A(n2883), .B(n2882), .S(n4645), .Z(n2887) );
  NAND2_X1 U3668 ( .A1(n2885), .A2(n2884), .ZN(n2886) );
  NAND2_X1 U3669 ( .A1(n2887), .A2(n2886), .ZN(U3515) );
  INV_X1 U3670 ( .A(n4583), .ZN(n2989) );
  NOR2_X1 U3671 ( .A1(n3054), .A2(n2989), .ZN(n2909) );
  INV_X2 U3672 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3673 ( .A(DATAI_22_), .ZN(n4902) );
  NAND2_X1 U3674 ( .A1(n3982), .A2(STATE_REG_SCAN_IN), .ZN(n2888) );
  OAI21_X1 U3675 ( .B1(STATE_REG_SCAN_IN), .B2(n4902), .A(n2888), .ZN(U3330)
         );
  INV_X1 U3676 ( .A(DATAI_18_), .ZN(n2890) );
  NAND2_X1 U3677 ( .A1(n4064), .A2(STATE_REG_SCAN_IN), .ZN(n2889) );
  OAI21_X1 U3678 ( .B1(STATE_REG_SCAN_IN), .B2(n2890), .A(n2889), .ZN(U3334)
         );
  INV_X1 U3679 ( .A(DATAI_26_), .ZN(n2892) );
  NAND2_X1 U3680 ( .A1(n2901), .A2(STATE_REG_SCAN_IN), .ZN(n2891) );
  OAI21_X1 U3681 ( .B1(STATE_REG_SCAN_IN), .B2(n2892), .A(n2891), .ZN(U3326)
         );
  INV_X1 U3682 ( .A(DATAI_24_), .ZN(n4739) );
  NAND2_X1 U3683 ( .A1(n2840), .A2(STATE_REG_SCAN_IN), .ZN(n2893) );
  OAI21_X1 U3684 ( .B1(STATE_REG_SCAN_IN), .B2(n4739), .A(n2893), .ZN(U3328)
         );
  INV_X1 U3685 ( .A(DATAI_27_), .ZN(n4735) );
  NAND2_X1 U3686 ( .A1(n3004), .A2(STATE_REG_SCAN_IN), .ZN(n2894) );
  OAI21_X1 U3687 ( .B1(STATE_REG_SCAN_IN), .B2(n4735), .A(n2894), .ZN(U3325)
         );
  INV_X1 U3688 ( .A(DATAI_31_), .ZN(n2897) );
  INV_X1 U3689 ( .A(IR_REG_30__SCAN_IN), .ZN(n2895) );
  NAND4_X1 U3690 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .A4(n2895), .ZN(n2896) );
  OAI21_X1 U3691 ( .B1(STATE_REG_SCAN_IN), .B2(n2897), .A(n2896), .ZN(U3321)
         );
  INV_X1 U3692 ( .A(DATAI_30_), .ZN(n4733) );
  NAND2_X1 U3693 ( .A1(n2493), .A2(STATE_REG_SCAN_IN), .ZN(n2898) );
  OAI21_X1 U3694 ( .B1(STATE_REG_SCAN_IN), .B2(n4733), .A(n2898), .ZN(U3322)
         );
  INV_X1 U3695 ( .A(DATAI_28_), .ZN(n4736) );
  NAND2_X1 U3696 ( .A1(n2992), .A2(STATE_REG_SCAN_IN), .ZN(n2899) );
  OAI21_X1 U3697 ( .B1(STATE_REG_SCAN_IN), .B2(n4736), .A(n2899), .ZN(U3324)
         );
  INV_X1 U3698 ( .A(D_REG_1__SCAN_IN), .ZN(n2903) );
  NOR3_X1 U3699 ( .A1(n2989), .A2(n2901), .A3(n4422), .ZN(n2902) );
  AOI21_X1 U3700 ( .B1(n4582), .B2(n2903), .A(n2902), .ZN(U3459) );
  NAND2_X1 U3701 ( .A1(n2904), .A2(n4583), .ZN(n2905) );
  OAI22_X1 U3702 ( .A1(n4581), .A2(D_REG_0__SCAN_IN), .B1(n2840), .B2(n2905), 
        .ZN(n2906) );
  INV_X1 U3703 ( .A(n2906), .ZN(U3458) );
  NAND2_X1 U3704 ( .A1(n2979), .A2(n3052), .ZN(n2907) );
  AND2_X1 U3705 ( .A1(n2529), .A2(n2907), .ZN(n2922) );
  INV_X1 U3706 ( .A(n2922), .ZN(n2908) );
  OR2_X1 U3707 ( .A1(n3052), .A2(U3149), .ZN(n3985) );
  NAND2_X1 U3708 ( .A1(n2986), .A2(n3985), .ZN(n2923) );
  NOR2_X1 U3709 ( .A1(n4541), .A2(U4043), .ZN(U3148) );
  INV_X1 U3710 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4899) );
  INV_X1 U3711 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4371) );
  NAND2_X1 U3712 ( .A1(n2522), .A2(REG2_REG_31__SCAN_IN), .ZN(n2910) );
  OAI211_X1 U3713 ( .C1(n2725), .C2(n4371), .A(n2911), .B(n2910), .ZN(n4076)
         );
  NAND2_X1 U3714 ( .A1(n4076), .A2(U4043), .ZN(n2913) );
  OAI21_X1 U3715 ( .B1(n2909), .B2(n4899), .A(n2913), .ZN(U3581) );
  INV_X1 U3716 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4811) );
  NAND2_X1 U3717 ( .A1(n3141), .A2(U4043), .ZN(n2914) );
  OAI21_X1 U3718 ( .B1(n2909), .B2(n4811), .A(n2914), .ZN(U3550) );
  INV_X1 U3719 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U3720 ( .A1(n2915), .A2(U4043), .ZN(n2916) );
  OAI21_X1 U3721 ( .B1(n2909), .B2(n4858), .A(n2916), .ZN(U3554) );
  INV_X1 U3722 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3012) );
  MUX2_X1 U3723 ( .A(REG2_REG_2__SCAN_IN), .B(n3012), .S(n4432), .Z(n2920) );
  INV_X1 U3724 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2917) );
  AND2_X1 U3725 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2918)
         );
  NAND2_X1 U3726 ( .A1(n4010), .A2(n3013), .ZN(n2919) );
  NAND2_X1 U3727 ( .A1(n4432), .A2(REG2_REG_2__SCAN_IN), .ZN(n2921) );
  NAND2_X1 U3728 ( .A1(n3016), .A2(n2921), .ZN(n2951) );
  XNOR2_X1 U3729 ( .A(n2950), .B(REG2_REG_3__SCAN_IN), .ZN(n2933) );
  AND2_X1 U3730 ( .A1(n2923), .A2(n2922), .ZN(n4001) );
  INV_X1 U3731 ( .A(n3004), .ZN(n3998) );
  OR2_X1 U3732 ( .A1(n3998), .A2(n3003), .ZN(n3980) );
  INV_X1 U3733 ( .A(n3980), .ZN(n2924) );
  INV_X1 U3734 ( .A(n4507), .ZN(n4535) );
  NOR2_X1 U3735 ( .A1(STATE_REG_SCAN_IN), .A2(n2532), .ZN(n3070) );
  NOR2_X1 U3736 ( .A1(n4548), .A2(n2929), .ZN(n2925) );
  AOI211_X1 U3737 ( .C1(n4541), .C2(ADDR_REG_3__SCAN_IN), .A(n3070), .B(n2925), 
        .ZN(n2932) );
  INV_X1 U3738 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4649) );
  MUX2_X1 U3739 ( .A(REG1_REG_2__SCAN_IN), .B(n4649), .S(n4432), .Z(n3011) );
  INV_X1 U3740 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2926) );
  AND2_X1 U3741 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4007)
         );
  NAND2_X1 U3742 ( .A1(n4006), .A2(n2927), .ZN(n3010) );
  NAND2_X1 U3743 ( .A1(n3011), .A2(n3010), .ZN(n3009) );
  NAND2_X1 U3744 ( .A1(n4432), .A2(REG1_REG_2__SCAN_IN), .ZN(n2928) );
  NAND2_X1 U3745 ( .A1(n3009), .A2(n2928), .ZN(n2939) );
  XNOR2_X1 U3746 ( .A(n2939), .B(n2929), .ZN(n2930) );
  OAI211_X1 U3747 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2930), .A(n4542), .B(n2941), 
        .ZN(n2931) );
  OAI211_X1 U3748 ( .C1(n2933), .C2(n4535), .A(n2932), .B(n2931), .ZN(U3243)
         );
  INV_X1 U3749 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4925) );
  NAND2_X1 U3750 ( .A1(n3845), .A2(U4043), .ZN(n2934) );
  OAI21_X1 U3751 ( .B1(n2909), .B2(n4925), .A(n2934), .ZN(U3580) );
  INV_X1 U3752 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4818) );
  NAND2_X1 U3753 ( .A1(n3305), .A2(U4043), .ZN(n2935) );
  OAI21_X1 U3754 ( .B1(n2909), .B2(n4818), .A(n2935), .ZN(U3558) );
  INV_X1 U3755 ( .A(n4548), .ZN(n4017) );
  INV_X1 U3756 ( .A(n4541), .ZN(n4477) );
  INV_X1 U3757 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n2938) );
  INV_X1 U3758 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2936) );
  NOR2_X1 U3759 ( .A1(STATE_REG_SCAN_IN), .A2(n2936), .ZN(n3205) );
  INV_X1 U3760 ( .A(n3205), .ZN(n2937) );
  OAI21_X1 U3761 ( .B1(n4477), .B2(n2938), .A(n2937), .ZN(n2949) );
  INV_X1 U3762 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2947) );
  NAND2_X1 U3763 ( .A1(n2939), .A2(n4431), .ZN(n2940) );
  INV_X1 U3764 ( .A(n2942), .ZN(n2943) );
  XOR2_X1 U3765 ( .A(n4429), .B(REG1_REG_5__SCAN_IN), .Z(n4020) );
  INV_X1 U3766 ( .A(n4428), .ZN(n2959) );
  AOI21_X1 U3767 ( .B1(n2944), .B2(n2959), .A(n3319), .ZN(n2945) );
  INV_X1 U3768 ( .A(n2945), .ZN(n2946) );
  INV_X1 U3769 ( .A(n4542), .ZN(n4074) );
  AOI211_X1 U3770 ( .C1(n2947), .C2(n2946), .A(n3318), .B(n4074), .ZN(n2948)
         );
  AOI211_X1 U3771 ( .C1(n4017), .C2(n4428), .A(n2949), .B(n2948), .ZN(n2962)
         );
  NAND2_X1 U3772 ( .A1(n2950), .A2(REG2_REG_3__SCAN_IN), .ZN(n2953) );
  NAND2_X1 U3773 ( .A1(n2951), .A2(n4431), .ZN(n2952) );
  NAND2_X1 U3774 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  XNOR2_X1 U3775 ( .A(n2954), .B(n3026), .ZN(n3021) );
  NAND2_X1 U3776 ( .A1(n3021), .A2(REG2_REG_4__SCAN_IN), .ZN(n2956) );
  NAND2_X1 U3777 ( .A1(n2954), .A2(n4430), .ZN(n2955) );
  NAND2_X1 U3778 ( .A1(n2956), .A2(n2955), .ZN(n4022) );
  INV_X1 U3779 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2957) );
  MUX2_X1 U3780 ( .A(REG2_REG_5__SCAN_IN), .B(n2957), .S(n4429), .Z(n4023) );
  NAND2_X1 U3781 ( .A1(n4429), .A2(REG2_REG_5__SCAN_IN), .ZN(n2958) );
  OAI211_X1 U3782 ( .C1(n2960), .C2(REG2_REG_6__SCAN_IN), .A(n4507), .B(n3339), 
        .ZN(n2961) );
  NAND2_X1 U3783 ( .A1(n2962), .A2(n2961), .ZN(U3246) );
  INV_X1 U3784 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U3785 ( .A1(n3612), .A2(U4043), .ZN(n2963) );
  OAI21_X1 U3786 ( .B1(n2909), .B2(n4845), .A(n2963), .ZN(U3565) );
  INV_X1 U3787 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U3788 ( .A1(n3557), .A2(U4043), .ZN(n2964) );
  OAI21_X1 U3789 ( .B1(n2909), .B2(n4821), .A(n2964), .ZN(U3563) );
  INV_X1 U3790 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U3791 ( .A1(n4213), .A2(U4043), .ZN(n2965) );
  OAI21_X1 U3792 ( .B1(n2909), .B2(n4820), .A(n2965), .ZN(U3570) );
  NAND2_X4 U3793 ( .A1(n2966), .A2(n3054), .ZN(n3689) );
  OAI22_X1 U3794 ( .A1(n3709), .A2(n3691), .B1(n3136), .B2(n3689), .ZN(n2967)
         );
  NAND2_X1 U3795 ( .A1(n4069), .A2(n3982), .ZN(n2988) );
  XNOR2_X1 U3796 ( .A(n2967), .B(n3687), .ZN(n3036) );
  OR2_X1 U3797 ( .A1(n3709), .A2(n3671), .ZN(n2969) );
  NAND2_X1 U3798 ( .A1(n3140), .A2(n3681), .ZN(n2968) );
  NAND2_X1 U3799 ( .A1(n2969), .A2(n2968), .ZN(n3035) );
  XNOR2_X1 U3800 ( .A(n3036), .B(n3035), .ZN(n3031) );
  AND2_X1 U3801 ( .A1(n3705), .A2(n3058), .ZN(n2970) );
  AOI21_X1 U3802 ( .B1(n3141), .B2(n3681), .A(n2970), .ZN(n2975) );
  NAND2_X1 U3803 ( .A1(n2972), .A2(REG1_REG_0__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3804 ( .A1(n2975), .A2(n2971), .ZN(n3001) );
  AOI22_X1 U3805 ( .A1(n3705), .A2(n3681), .B1(IR_REG_0__SCAN_IN), .B2(n2972), 
        .ZN(n2973) );
  NAND2_X1 U3806 ( .A1(n2974), .A2(n2973), .ZN(n3002) );
  AOI22_X1 U3807 ( .A1(n3001), .A2(n3002), .B1(n3676), .B2(n2975), .ZN(n3032)
         );
  XNOR2_X1 U3808 ( .A(n3031), .B(n3032), .ZN(n2997) );
  INV_X1 U3809 ( .A(n2976), .ZN(n3094) );
  NAND3_X1 U3810 ( .A1(n2977), .A2(n3094), .A3(n3091), .ZN(n2991) );
  NAND2_X1 U3811 ( .A1(n2978), .A2(n4599), .ZN(n2981) );
  INV_X1 U3812 ( .A(n2979), .ZN(n2980) );
  NAND3_X1 U3813 ( .A1(n2981), .A2(n2983), .A3(n2980), .ZN(n2982) );
  NAND2_X1 U3814 ( .A1(n2991), .A2(n2985), .ZN(n3056) );
  NAND2_X1 U3815 ( .A1(n3056), .A2(n3093), .ZN(n3706) );
  NAND2_X1 U3816 ( .A1(n4298), .A2(n2983), .ZN(n2984) );
  OR2_X1 U3817 ( .A1(n2991), .A2(n2984), .ZN(n2987) );
  AOI22_X1 U3818 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3706), .B1(n4438), .B2(n3140), .ZN(n2996) );
  NOR2_X1 U3819 ( .A1(n2989), .A2(n2988), .ZN(n2990) );
  NAND2_X1 U3820 ( .A1(n3681), .A2(n2990), .ZN(n3981) );
  NOR2_X2 U3821 ( .A1(n2994), .A2(n2992), .ZN(n3814) );
  NOR2_X2 U3822 ( .A1(n2994), .A2(n3003), .ZN(n3810) );
  AOI22_X1 U3823 ( .A1(n3814), .A2(n2993), .B1(n3810), .B2(n3141), .ZN(n2995)
         );
  OAI211_X1 U3824 ( .C1(n2997), .C2(n3816), .A(n2996), .B(n2995), .ZN(U3219)
         );
  INV_X1 U3825 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4823) );
  NAND2_X1 U3826 ( .A1(n4194), .A2(U4043), .ZN(n2998) );
  OAI21_X1 U3827 ( .B1(n2909), .B2(n4823), .A(n2998), .ZN(U3573) );
  INV_X1 U3828 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2999) );
  AND2_X1 U3829 ( .A1(n3004), .A2(n2999), .ZN(n3000) );
  OR2_X1 U3830 ( .A1(n3000), .A2(n3003), .ZN(n3999) );
  NAND2_X1 U3831 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4009) );
  OAI21_X1 U3832 ( .B1(n3980), .B2(n4009), .A(n2909), .ZN(n3006) );
  XOR2_X1 U3833 ( .A(n3002), .B(n3001), .Z(n3704) );
  NOR3_X1 U3834 ( .A1(n3704), .A2(n3004), .A3(n3003), .ZN(n3005) );
  AOI211_X1 U3835 ( .C1(n2452), .C2(n3999), .A(n3006), .B(n3005), .ZN(n3027)
         );
  INV_X1 U3836 ( .A(n4432), .ZN(n3008) );
  AOI22_X1 U3837 ( .A1(n4541), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3007) );
  OAI21_X1 U3838 ( .B1(n3008), .B2(n4548), .A(n3007), .ZN(n3020) );
  OAI211_X1 U3839 ( .C1(n3011), .C2(n3010), .A(n4542), .B(n3009), .ZN(n3018)
         );
  MUX2_X1 U3840 ( .A(n3012), .B(REG2_REG_2__SCAN_IN), .S(n4432), .Z(n3014) );
  NAND3_X1 U3841 ( .A1(n3014), .A2(n4010), .A3(n3013), .ZN(n3015) );
  NAND3_X1 U3842 ( .A1(n4507), .A2(n3016), .A3(n3015), .ZN(n3017) );
  NAND2_X1 U3843 ( .A1(n3018), .A2(n3017), .ZN(n3019) );
  OR3_X1 U3844 ( .A1(n3027), .A2(n3020), .A3(n3019), .ZN(U3242) );
  XOR2_X1 U3845 ( .A(REG2_REG_4__SCAN_IN), .B(n3021), .Z(n3029) );
  OAI211_X1 U3846 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3023), .A(n4542), .B(n3022), 
        .ZN(n3025) );
  AND2_X1 U3847 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3088) );
  AOI21_X1 U3848 ( .B1(n4541), .B2(ADDR_REG_4__SCAN_IN), .A(n3088), .ZN(n3024)
         );
  OAI211_X1 U3849 ( .C1(n4548), .C2(n3026), .A(n3025), .B(n3024), .ZN(n3028)
         );
  AOI211_X1 U3850 ( .C1(n4507), .C2(n3029), .A(n3028), .B(n3027), .ZN(n3030)
         );
  INV_X1 U3851 ( .A(n3030), .ZN(U3244) );
  INV_X1 U3852 ( .A(n3031), .ZN(n3034) );
  INV_X1 U3853 ( .A(n3032), .ZN(n3033) );
  NAND2_X1 U3854 ( .A1(n3036), .A2(n3035), .ZN(n3037) );
  OAI22_X1 U3855 ( .A1(n3144), .A2(n3691), .B1(n3128), .B2(n3689), .ZN(n3038)
         );
  XNOR2_X1 U3856 ( .A(n3038), .B(n3676), .ZN(n3041) );
  OR2_X1 U3857 ( .A1(n3144), .A2(n3671), .ZN(n3040) );
  NAND2_X1 U3858 ( .A1(n3121), .A2(n3681), .ZN(n3039) );
  AND2_X1 U3859 ( .A1(n3040), .A2(n3039), .ZN(n3042) );
  INV_X1 U3860 ( .A(n3041), .ZN(n3044) );
  INV_X1 U3861 ( .A(n3042), .ZN(n3043) );
  INV_X1 U3862 ( .A(n3064), .ZN(n3045) );
  AOI21_X1 U3863 ( .B1(n3047), .B2(n3046), .A(n3045), .ZN(n3050) );
  AOI22_X1 U3864 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3706), .B1(n4438), .B2(n3121), .ZN(n3049) );
  AOI22_X1 U3865 ( .A1(n3810), .A2(n2511), .B1(n3814), .B2(n3997), .ZN(n3048)
         );
  OAI211_X1 U3866 ( .C1(n3050), .C2(n3816), .A(n3049), .B(n3048), .ZN(U3234)
         );
  INV_X1 U3867 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U3868 ( .A1(n4122), .A2(U4043), .ZN(n3051) );
  OAI21_X1 U3869 ( .B1(n2909), .B2(n4842), .A(n3051), .ZN(U3575) );
  AND3_X1 U3870 ( .A1(n3054), .A2(n3053), .A3(n3052), .ZN(n3055) );
  NAND2_X1 U3871 ( .A1(n3056), .A2(n3055), .ZN(n3057) );
  NAND2_X1 U3872 ( .A1(n3997), .A2(n3681), .ZN(n3060) );
  NAND2_X1 U3873 ( .A1(n3175), .A2(n3058), .ZN(n3059) );
  NAND2_X1 U3874 ( .A1(n3060), .A2(n3059), .ZN(n3061) );
  XNOR2_X1 U3875 ( .A(n3061), .B(n3687), .ZN(n3075) );
  AND2_X1 U3876 ( .A1(n3175), .A2(n3681), .ZN(n3062) );
  AOI21_X1 U3877 ( .B1(n3997), .B2(n3686), .A(n3062), .ZN(n3076) );
  XNOR2_X1 U3878 ( .A(n3075), .B(n3076), .ZN(n3066) );
  NAND2_X1 U3879 ( .A1(n3064), .A2(n3063), .ZN(n3065) );
  NAND2_X1 U3880 ( .A1(n3065), .A2(n3066), .ZN(n3084) );
  OAI21_X1 U3881 ( .B1(n3066), .B2(n3065), .A(n3084), .ZN(n3067) );
  NAND2_X1 U3882 ( .A1(n3067), .A2(n4443), .ZN(n3072) );
  OAI22_X1 U3883 ( .A1(n3068), .A2(n4435), .B1(n4434), .B2(n3144), .ZN(n3069)
         );
  AOI211_X1 U3884 ( .C1(n3175), .C2(n4438), .A(n3070), .B(n3069), .ZN(n3071)
         );
  OAI211_X1 U3885 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4448), .A(n3072), .B(n3071), 
        .ZN(U3215) );
  INV_X1 U3886 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U3887 ( .A1(n4142), .A2(U4043), .ZN(n3073) );
  OAI21_X1 U3888 ( .B1(U4043), .B2(n4900), .A(n3073), .ZN(U3576) );
  INV_X1 U3889 ( .A(n3074), .ZN(n3153) );
  INV_X1 U3890 ( .A(n3075), .ZN(n3077) );
  NAND2_X1 U3891 ( .A1(n3077), .A2(n3076), .ZN(n3082) );
  AND2_X1 U3892 ( .A1(n3084), .A2(n3082), .ZN(n3086) );
  OAI22_X1 U3893 ( .A1(n3068), .A2(n3691), .B1(n3078), .B2(n3689), .ZN(n3079)
         );
  XNOR2_X1 U3894 ( .A(n3079), .B(n3676), .ZN(n3103) );
  OR2_X1 U3895 ( .A1(n3068), .A2(n3671), .ZN(n3081) );
  NAND2_X1 U3896 ( .A1(n3159), .A2(n3681), .ZN(n3080) );
  NAND2_X1 U3897 ( .A1(n3081), .A2(n3080), .ZN(n3104) );
  XNOR2_X1 U3898 ( .A(n3103), .B(n3104), .ZN(n3085) );
  AND2_X1 U3899 ( .A1(n3082), .A2(n3085), .ZN(n3083) );
  NAND2_X1 U3900 ( .A1(n3084), .A2(n3083), .ZN(n3107) );
  OAI211_X1 U3901 ( .C1(n3086), .C2(n3085), .A(n4443), .B(n3107), .ZN(n3090)
         );
  OAI22_X1 U3902 ( .A1(n3161), .A2(n4434), .B1(n4435), .B2(n3203), .ZN(n3087)
         );
  AOI211_X1 U3903 ( .C1(n3159), .C2(n4438), .A(n3088), .B(n3087), .ZN(n3089)
         );
  OAI211_X1 U3904 ( .C1(n4448), .C2(n3153), .A(n3090), .B(n3089), .ZN(U3227)
         );
  NAND4_X1 U3905 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3095)
         );
  NAND2_X1 U3906 ( .A1(n4290), .A2(n4069), .ZN(n4288) );
  INV_X1 U3907 ( .A(n4288), .ZN(n3096) );
  AOI21_X1 U3908 ( .B1(n3096), .B2(n4599), .A(n4148), .ZN(n3102) );
  INV_X1 U3909 ( .A(n3382), .ZN(n4563) );
  NAND2_X1 U3910 ( .A1(n3141), .A2(n4601), .ZN(n3908) );
  NAND2_X1 U3911 ( .A1(n3906), .A2(n3908), .ZN(n4604) );
  OAI21_X1 U3912 ( .B1(n4563), .B2(n4254), .A(n4604), .ZN(n3097) );
  OAI21_X1 U3913 ( .B1(n3709), .B2(n4274), .A(n3097), .ZN(n4602) );
  INV_X1 U3914 ( .A(n4604), .ZN(n3099) );
  OR2_X1 U3915 ( .A1(n2966), .A2(n4069), .ZN(n3221) );
  NOR2_X1 U3916 ( .A1(n5040), .A2(n3221), .ZN(n4573) );
  INV_X1 U3917 ( .A(n4573), .ZN(n3132) );
  AOI22_X1 U3918 ( .A1(n5040), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n5034), .ZN(n3098) );
  OAI21_X1 U3919 ( .B1(n3099), .B2(n3132), .A(n3098), .ZN(n3100) );
  AOI21_X1 U3920 ( .B1(n4290), .B2(n4602), .A(n3100), .ZN(n3101) );
  OAI21_X1 U3921 ( .B1(n3102), .B2(n4601), .A(n3101), .ZN(U3290) );
  INV_X1 U3922 ( .A(n3103), .ZN(n3105) );
  NAND2_X1 U3923 ( .A1(n3105), .A2(n3104), .ZN(n3106) );
  NAND2_X1 U3924 ( .A1(n3996), .A2(n3681), .ZN(n3109) );
  NAND2_X1 U3925 ( .A1(n3215), .A2(n3058), .ZN(n3108) );
  NAND2_X1 U3926 ( .A1(n3109), .A2(n3108), .ZN(n3110) );
  XNOR2_X1 U3927 ( .A(n3110), .B(n3687), .ZN(n3189) );
  AND2_X1 U3928 ( .A1(n3215), .A2(n3681), .ZN(n3111) );
  AOI21_X1 U3929 ( .B1(n3996), .B2(n3686), .A(n3111), .ZN(n3187) );
  XNOR2_X1 U3930 ( .A(n3189), .B(n3187), .ZN(n3185) );
  XNOR2_X1 U3931 ( .A(n3186), .B(n3185), .ZN(n3115) );
  AND2_X1 U3932 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4024) );
  OAI22_X1 U3933 ( .A1(n3068), .A2(n4434), .B1(n4435), .B2(n3245), .ZN(n3112)
         );
  AOI211_X1 U3934 ( .C1(n3215), .C2(n4438), .A(n4024), .B(n3112), .ZN(n3114)
         );
  NAND2_X1 U3935 ( .A1(n3804), .A2(n3216), .ZN(n3113) );
  OAI211_X1 U3936 ( .C1(n3115), .C2(n3816), .A(n3114), .B(n3113), .ZN(U3224)
         );
  NAND2_X1 U3937 ( .A1(n3116), .A2(n3119), .ZN(n3117) );
  NAND2_X1 U3938 ( .A1(n3118), .A2(n3117), .ZN(n4614) );
  INV_X1 U3939 ( .A(n4614), .ZN(n3133) );
  XNOR2_X1 U3940 ( .A(n3120), .B(n2788), .ZN(n3126) );
  INV_X1 U3941 ( .A(n4254), .ZN(n4560) );
  NAND2_X1 U3942 ( .A1(n4614), .A2(n4563), .ZN(n3125) );
  AOI22_X1 U3943 ( .A1(n3997), .A2(n4558), .B1(n4298), .B2(n3121), .ZN(n3122)
         );
  OAI21_X1 U3944 ( .B1(n3709), .B2(n4554), .A(n3122), .ZN(n3123) );
  INV_X1 U3945 ( .A(n3123), .ZN(n3124) );
  OAI211_X1 U3946 ( .C1(n3126), .C2(n4560), .A(n3125), .B(n3124), .ZN(n4612)
         );
  MUX2_X1 U3947 ( .A(n4612), .B(REG2_REG_2__SCAN_IN), .S(n5040), .Z(n3127) );
  INV_X1 U3948 ( .A(n3127), .ZN(n3131) );
  INV_X1 U3949 ( .A(n4638), .ZN(n4631) );
  INV_X1 U3950 ( .A(n3176), .ZN(n4610) );
  NOR2_X1 U3951 ( .A1(n3134), .A2(n3128), .ZN(n4611) );
  NOR3_X1 U3952 ( .A1(n4263), .A2(n4610), .A3(n4611), .ZN(n3129) );
  AOI21_X1 U3953 ( .B1(n5034), .B2(REG3_REG_2__SCAN_IN), .A(n3129), .ZN(n3130)
         );
  OAI211_X1 U3954 ( .C1(n3133), .C2(n3132), .A(n3131), .B(n3130), .ZN(U3288)
         );
  INV_X1 U3955 ( .A(n3134), .ZN(n3135) );
  OAI21_X1 U3956 ( .B1(n4601), .B2(n3136), .A(n3135), .ZN(n4605) );
  OR2_X1 U3957 ( .A1(n2786), .A2(n3137), .ZN(n3138) );
  NAND2_X1 U3958 ( .A1(n3139), .A2(n3138), .ZN(n4607) );
  NAND2_X1 U3959 ( .A1(n3140), .A2(n4298), .ZN(n3143) );
  NAND2_X1 U3960 ( .A1(n3141), .A2(n4282), .ZN(n3142) );
  OAI211_X1 U3961 ( .C1(n3144), .C2(n4274), .A(n3143), .B(n3142), .ZN(n3145)
         );
  INV_X1 U3962 ( .A(n3145), .ZN(n3148) );
  XNOR2_X1 U3963 ( .A(n2786), .B(n3906), .ZN(n3146) );
  NAND2_X1 U3964 ( .A1(n3146), .A2(n4254), .ZN(n3147) );
  OAI211_X1 U3965 ( .C1(n4607), .C2(n3382), .A(n3148), .B(n3147), .ZN(n4609)
         );
  MUX2_X1 U3966 ( .A(n4609), .B(REG2_REG_1__SCAN_IN), .S(n5040), .Z(n3149) );
  INV_X1 U3967 ( .A(n3149), .ZN(n3152) );
  INV_X1 U3968 ( .A(n4607), .ZN(n3150) );
  AOI22_X1 U3969 ( .A1(n3150), .A2(n4573), .B1(REG3_REG_1__SCAN_IN), .B2(n5034), .ZN(n3151) );
  OAI211_X1 U3970 ( .C1(n4263), .C2(n4605), .A(n3152), .B(n3151), .ZN(U3289)
         );
  AOI211_X1 U3971 ( .C1(n3159), .C2(n3178), .A(n4631), .B(n3212), .ZN(n4616)
         );
  NOR2_X1 U3972 ( .A1(n4264), .A2(n3153), .ZN(n3165) );
  OR2_X1 U3973 ( .A1(n3169), .A2(n3154), .ZN(n3156) );
  NAND2_X1 U3974 ( .A1(n3156), .A2(n3155), .ZN(n3157) );
  XNOR2_X1 U3975 ( .A(n3157), .B(n3886), .ZN(n3166) );
  XOR2_X1 U3976 ( .A(n3886), .B(n3158), .Z(n3163) );
  AOI22_X1 U3977 ( .A1(n3996), .A2(n4558), .B1(n4298), .B2(n3159), .ZN(n3160)
         );
  OAI21_X1 U3978 ( .B1(n3161), .B2(n4554), .A(n3160), .ZN(n3162) );
  AOI21_X1 U3979 ( .B1(n3163), .B2(n4254), .A(n3162), .ZN(n3164) );
  OAI21_X1 U3980 ( .B1(n3382), .B2(n3166), .A(n3164), .ZN(n4615) );
  AOI211_X1 U3981 ( .C1(n4616), .C2(n4069), .A(n3165), .B(n4615), .ZN(n3168)
         );
  INV_X1 U3982 ( .A(n3166), .ZN(n4617) );
  AOI22_X1 U3983 ( .A1(n4617), .A2(n4573), .B1(REG2_REG_4__SCAN_IN), .B2(n5040), .ZN(n3167) );
  OAI21_X1 U3984 ( .B1(n3168), .B2(n5040), .A(n3167), .ZN(U3286) );
  XNOR2_X1 U3985 ( .A(n3169), .B(n3888), .ZN(n4570) );
  XNOR2_X1 U3986 ( .A(n3170), .B(n3888), .ZN(n3174) );
  AOI22_X1 U3987 ( .A1(n2993), .A2(n4282), .B1(n3175), .B2(n4298), .ZN(n3171)
         );
  OAI21_X1 U3988 ( .B1(n3068), .B2(n4274), .A(n3171), .ZN(n3173) );
  NOR2_X1 U3989 ( .A1(n4570), .A2(n3382), .ZN(n3172) );
  AOI211_X1 U3990 ( .C1(n3174), .C2(n4254), .A(n3173), .B(n3172), .ZN(n4577)
         );
  OAI21_X1 U3991 ( .B1(n4570), .B2(n4606), .A(n4577), .ZN(n3183) );
  NAND2_X1 U3992 ( .A1(n3176), .A2(n3175), .ZN(n3177) );
  NAND2_X1 U3993 ( .A1(n3178), .A2(n3177), .ZN(n4571) );
  OAI22_X1 U3994 ( .A1(n4417), .A2(n4571), .B1(n4645), .B2(n2533), .ZN(n3179)
         );
  AOI21_X1 U3995 ( .B1(n3183), .B2(n4645), .A(n3179), .ZN(n3180) );
  INV_X1 U3996 ( .A(n3180), .ZN(U3473) );
  INV_X1 U3997 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3181) );
  OAI22_X1 U3998 ( .A1(n4358), .A2(n4571), .B1(n4659), .B2(n3181), .ZN(n3182)
         );
  AOI21_X1 U3999 ( .B1(n3183), .B2(n4659), .A(n3182), .ZN(n3184) );
  INV_X1 U4000 ( .A(n3184), .ZN(U3521) );
  INV_X1 U4001 ( .A(n3187), .ZN(n3188) );
  NAND2_X1 U4002 ( .A1(n3189), .A2(n3188), .ZN(n3190) );
  NAND2_X1 U4003 ( .A1(n3995), .A2(n3681), .ZN(n3192) );
  NAND2_X1 U4004 ( .A1(n3281), .A2(n3058), .ZN(n3191) );
  NAND2_X1 U4005 ( .A1(n3192), .A2(n3191), .ZN(n3193) );
  XNOR2_X1 U4006 ( .A(n3193), .B(n3687), .ZN(n3196) );
  NAND2_X1 U4007 ( .A1(n3995), .A2(n3686), .ZN(n3195) );
  NAND2_X1 U4008 ( .A1(n3281), .A2(n3681), .ZN(n3194) );
  NAND2_X1 U4009 ( .A1(n3195), .A2(n3194), .ZN(n3197) );
  AND2_X1 U4010 ( .A1(n3196), .A2(n3197), .ZN(n3236) );
  INV_X1 U4011 ( .A(n3236), .ZN(n3200) );
  INV_X1 U4012 ( .A(n3196), .ZN(n3199) );
  INV_X1 U4013 ( .A(n3197), .ZN(n3198) );
  NAND2_X1 U4014 ( .A1(n3199), .A2(n3198), .ZN(n3238) );
  NAND2_X1 U4015 ( .A1(n3200), .A2(n3238), .ZN(n3201) );
  XNOR2_X1 U4016 ( .A(n3237), .B(n3201), .ZN(n3202) );
  NAND2_X1 U4017 ( .A1(n3202), .A2(n4443), .ZN(n3207) );
  OAI22_X1 U4018 ( .A1(n3203), .A2(n4434), .B1(n4435), .B2(n3262), .ZN(n3204)
         );
  AOI211_X1 U4019 ( .C1(n3281), .C2(n4438), .A(n3205), .B(n3204), .ZN(n3206)
         );
  OAI211_X1 U4020 ( .C1(n4448), .C2(n3208), .A(n3207), .B(n3206), .ZN(U3236)
         );
  INV_X1 U4021 ( .A(n3209), .ZN(n3918) );
  NAND2_X1 U4022 ( .A1(n3918), .A2(n3934), .ZN(n3884) );
  XNOR2_X1 U4023 ( .A(n3210), .B(n3884), .ZN(n3211) );
  AOI222_X1 U4024 ( .A1(n4254), .A2(n3211), .B1(n3995), .B2(n4558), .C1(n2915), 
        .C2(n4282), .ZN(n3251) );
  INV_X1 U4025 ( .A(n3212), .ZN(n3214) );
  INV_X1 U4026 ( .A(n3280), .ZN(n3213) );
  AOI21_X1 U4027 ( .B1(n3215), .B2(n3214), .A(n3213), .ZN(n3256) );
  INV_X1 U4028 ( .A(n4148), .ZN(n5039) );
  NOR2_X1 U4029 ( .A1(n5039), .A2(n3252), .ZN(n3219) );
  INV_X1 U4030 ( .A(n3216), .ZN(n3217) );
  OAI22_X1 U4031 ( .A1(n4290), .A2(n2957), .B1(n3217), .B2(n4264), .ZN(n3218)
         );
  AOI211_X1 U4032 ( .C1(n3256), .C2(n5032), .A(n3219), .B(n3218), .ZN(n3224)
         );
  XOR2_X1 U4033 ( .A(n3884), .B(n3220), .Z(n3254) );
  NAND2_X1 U4034 ( .A1(n3382), .A2(n3221), .ZN(n3222) );
  NAND2_X1 U4035 ( .A1(n4290), .A2(n3222), .ZN(n4293) );
  NAND2_X1 U4036 ( .A1(n3254), .A2(n5045), .ZN(n3223) );
  OAI211_X1 U4037 ( .C1(n3251), .C2(n5040), .A(n3224), .B(n3223), .ZN(U3285)
         );
  INV_X1 U4038 ( .A(n3885), .ZN(n3922) );
  NAND2_X1 U4039 ( .A1(n3995), .A2(n4282), .ZN(n3226) );
  NAND2_X1 U4040 ( .A1(n3305), .A2(n4558), .ZN(n3225) );
  OAI211_X1 U4041 ( .C1(n4552), .C2(n3239), .A(n3226), .B(n3225), .ZN(n3227)
         );
  AOI21_X1 U4042 ( .B1(n3228), .B2(n4254), .A(n3227), .ZN(n4623) );
  XNOR2_X1 U40430 ( .A(n3229), .B(n3922), .ZN(n4620) );
  NAND2_X1 U4044 ( .A1(n3278), .A2(n3247), .ZN(n3230) );
  NAND2_X1 U4045 ( .A1(n3230), .A2(n4638), .ZN(n3231) );
  OR2_X1 U4046 ( .A1(n3267), .A2(n3231), .ZN(n4622) );
  NOR2_X1 U4047 ( .A1(n4622), .A2(n4288), .ZN(n3234) );
  INV_X1 U4048 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3337) );
  INV_X1 U4049 ( .A(n3232), .ZN(n3250) );
  OAI22_X1 U4050 ( .A1(n4290), .A2(n3337), .B1(n3250), .B2(n4264), .ZN(n3233)
         );
  AOI211_X1 U4051 ( .C1(n4620), .C2(n5045), .A(n3234), .B(n3233), .ZN(n3235)
         );
  OAI21_X1 U4052 ( .B1(n5040), .B2(n4623), .A(n3235), .ZN(U3283) );
  OAI22_X1 U4053 ( .A1(n3262), .A2(n3691), .B1(n3689), .B2(n3239), .ZN(n3240)
         );
  XNOR2_X1 U4054 ( .A(n3240), .B(n3676), .ZN(n3285) );
  OR2_X1 U4055 ( .A1(n3262), .A2(n3671), .ZN(n3242) );
  NAND2_X1 U4056 ( .A1(n3247), .A2(n3681), .ZN(n3241) );
  NAND2_X1 U4057 ( .A1(n3242), .A2(n3241), .ZN(n3286) );
  XNOR2_X1 U4058 ( .A(n3285), .B(n3286), .ZN(n3243) );
  OAI211_X1 U4059 ( .C1(n3244), .C2(n3243), .A(n3289), .B(n4443), .ZN(n3249)
         );
  AND2_X1 U4060 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4457) );
  OAI22_X1 U4061 ( .A1(n3245), .A2(n4434), .B1(n4435), .B2(n3369), .ZN(n3246)
         );
  AOI211_X1 U4062 ( .C1(n3247), .C2(n4438), .A(n4457), .B(n3246), .ZN(n3248)
         );
  OAI211_X1 U4063 ( .C1(n4448), .C2(n3250), .A(n3249), .B(n3248), .ZN(U3210)
         );
  OAI21_X1 U4064 ( .B1(n3252), .B2(n4552), .A(n3251), .ZN(n3253) );
  AOI21_X1 U4065 ( .B1(n3254), .B2(n4619), .A(n3253), .ZN(n3258) );
  AOI22_X1 U4066 ( .A1(n3256), .A2(n2879), .B1(REG1_REG_5__SCAN_IN), .B2(n4657), .ZN(n3255) );
  OAI21_X1 U4067 ( .B1(n3258), .B2(n4657), .A(n3255), .ZN(U3523) );
  AOI22_X1 U4068 ( .A1(n3256), .A2(n2884), .B1(REG0_REG_5__SCAN_IN), .B2(n4643), .ZN(n3257) );
  OAI21_X1 U4069 ( .B1(n3258), .B2(n4643), .A(n3257), .ZN(U3477) );
  NAND2_X1 U4070 ( .A1(n3927), .A2(n3924), .ZN(n3882) );
  XNOR2_X1 U4071 ( .A(n3259), .B(n3882), .ZN(n3266) );
  XNOR2_X1 U4072 ( .A(n3260), .B(n3882), .ZN(n3264) );
  AOI22_X1 U4073 ( .A1(n3993), .A2(n4558), .B1(n4298), .B2(n3292), .ZN(n3261)
         );
  OAI21_X1 U4074 ( .B1(n3262), .B2(n4554), .A(n3261), .ZN(n3263) );
  AOI21_X1 U4075 ( .B1(n3264), .B2(n4254), .A(n3263), .ZN(n3265) );
  OAI21_X1 U4076 ( .B1(n3266), .B2(n3382), .A(n3265), .ZN(n4627) );
  INV_X1 U4077 ( .A(n4627), .ZN(n3273) );
  INV_X1 U4078 ( .A(n3266), .ZN(n4629) );
  NOR2_X1 U4079 ( .A1(n3267), .A2(n3298), .ZN(n4626) );
  INV_X1 U4080 ( .A(n3312), .ZN(n4625) );
  NOR3_X1 U4081 ( .A1(n4626), .A2(n4625), .A3(n4263), .ZN(n3271) );
  INV_X1 U4082 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3269) );
  INV_X1 U4083 ( .A(n3300), .ZN(n3268) );
  OAI22_X1 U4084 ( .A1(n4290), .A2(n3269), .B1(n3268), .B2(n4264), .ZN(n3270)
         );
  AOI211_X1 U4085 ( .C1(n4629), .C2(n4573), .A(n3271), .B(n3270), .ZN(n3272)
         );
  OAI21_X1 U4086 ( .B1(n3273), .B2(n5040), .A(n3272), .ZN(U3282) );
  AND2_X1 U4087 ( .A1(n3921), .A2(n3935), .ZN(n3887) );
  XOR2_X1 U4088 ( .A(n3887), .B(n3274), .Z(n5044) );
  XNOR2_X1 U4089 ( .A(n3275), .B(n3887), .ZN(n3276) );
  AOI222_X1 U4090 ( .A1(n4254), .A2(n3276), .B1(n3994), .B2(n4558), .C1(n3996), 
        .C2(n4282), .ZN(n5041) );
  OAI21_X1 U4091 ( .B1(n5038), .B2(n4552), .A(n5041), .ZN(n3277) );
  AOI21_X1 U4092 ( .B1(n4619), .B2(n5044), .A(n3277), .ZN(n3284) );
  INV_X1 U4093 ( .A(n3278), .ZN(n3279) );
  AOI21_X1 U4094 ( .B1(n3281), .B2(n3280), .A(n3279), .ZN(n5033) );
  AOI22_X1 U4095 ( .A1(n5033), .A2(n2884), .B1(n4643), .B2(REG0_REG_6__SCAN_IN), .ZN(n3282) );
  OAI21_X1 U4096 ( .B1(n3284), .B2(n4643), .A(n3282), .ZN(U3479) );
  AOI22_X1 U4097 ( .A1(n5033), .A2(n2879), .B1(n4657), .B2(REG1_REG_6__SCAN_IN), .ZN(n3283) );
  OAI21_X1 U4098 ( .B1(n3284), .B2(n4657), .A(n3283), .ZN(U3524) );
  INV_X1 U4099 ( .A(n3285), .ZN(n3287) );
  NAND2_X1 U4100 ( .A1(n3287), .A2(n3286), .ZN(n3288) );
  NAND2_X1 U4101 ( .A1(n3305), .A2(n3686), .ZN(n3291) );
  NAND2_X1 U4102 ( .A1(n3292), .A2(n3681), .ZN(n3290) );
  NAND2_X1 U4103 ( .A1(n3291), .A2(n3290), .ZN(n3364) );
  NAND2_X1 U4104 ( .A1(n3305), .A2(n3681), .ZN(n3294) );
  NAND2_X1 U4105 ( .A1(n3292), .A2(n3058), .ZN(n3293) );
  NAND2_X1 U4106 ( .A1(n3294), .A2(n3293), .ZN(n3295) );
  XNOR2_X1 U4107 ( .A(n3295), .B(n3687), .ZN(n3363) );
  XOR2_X1 U4108 ( .A(n3364), .B(n3363), .Z(n3296) );
  XNOR2_X1 U4109 ( .A(n3365), .B(n3296), .ZN(n3302) );
  AOI22_X1 U4110 ( .A1(n3810), .A2(n3994), .B1(n3814), .B2(n3993), .ZN(n3297)
         );
  NAND2_X1 U4111 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4465) );
  OAI211_X1 U4112 ( .C1(n3802), .C2(n3298), .A(n3297), .B(n4465), .ZN(n3299)
         );
  AOI21_X1 U4113 ( .B1(n3300), .B2(n3804), .A(n3299), .ZN(n3301) );
  OAI21_X1 U4114 ( .B1(n3302), .B2(n3816), .A(n3301), .ZN(U3218) );
  INV_X1 U4115 ( .A(n3932), .ZN(n3936) );
  AND2_X1 U4116 ( .A1(n3936), .A2(n3926), .ZN(n3890) );
  INV_X1 U4117 ( .A(n3890), .ZN(n3309) );
  XNOR2_X1 U4118 ( .A(n3303), .B(n3309), .ZN(n3304) );
  NAND2_X1 U4119 ( .A1(n3304), .A2(n4254), .ZN(n3307) );
  AOI22_X1 U4120 ( .A1(n4282), .A2(n3305), .B1(n3992), .B2(n4558), .ZN(n3306)
         );
  AND2_X1 U4121 ( .A1(n3307), .A2(n3306), .ZN(n3412) );
  XNOR2_X1 U4122 ( .A(n3308), .B(n3309), .ZN(n3410) );
  INV_X1 U4123 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3335) );
  OAI22_X1 U4124 ( .A1(n3310), .A2(n4264), .B1(n3335), .B2(n4290), .ZN(n3315)
         );
  INV_X1 U4125 ( .A(n3311), .ZN(n3385) );
  AOI21_X1 U4126 ( .B1(n3371), .B2(n3312), .A(n3385), .ZN(n3418) );
  INV_X1 U4127 ( .A(n3418), .ZN(n3313) );
  OAI22_X1 U4128 ( .A1(n3313), .A2(n4263), .B1(n3413), .B2(n5039), .ZN(n3314)
         );
  AOI211_X1 U4129 ( .C1(n3410), .C2(n5045), .A(n3315), .B(n3314), .ZN(n3316)
         );
  OAI21_X1 U4130 ( .B1(n5040), .B2(n3412), .A(n3316), .ZN(U3281) );
  INV_X1 U4131 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U4132 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3334), .B1(n4591), .B2(
        n4797), .ZN(n4503) );
  NAND2_X1 U4133 ( .A1(n3336), .A2(REG1_REG_9__SCAN_IN), .ZN(n3322) );
  INV_X1 U4134 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3317) );
  INV_X1 U4135 ( .A(n3336), .ZN(n4595) );
  AOI22_X1 U4136 ( .A1(n3336), .A2(REG1_REG_9__SCAN_IN), .B1(n3317), .B2(n4595), .ZN(n4482) );
  INV_X1 U4137 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U4138 ( .A1(n4596), .A2(n3320), .ZN(n3321) );
  INV_X1 U4139 ( .A(n4596), .ZN(n4472) );
  NAND2_X1 U4140 ( .A1(n4592), .A2(n3323), .ZN(n3324) );
  INV_X1 U4141 ( .A(n4592), .ZN(n4491) );
  XNOR2_X1 U4142 ( .A(n3323), .B(n4491), .ZN(n4486) );
  NAND2_X1 U4143 ( .A1(n4588), .A2(n3325), .ZN(n3326) );
  INV_X1 U4144 ( .A(n4588), .ZN(n4516) );
  XNOR2_X1 U4145 ( .A(n3325), .B(n4516), .ZN(n4513) );
  NAND2_X1 U4146 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U4147 ( .A1(n3326), .A2(n4512), .ZN(n3330) );
  INV_X1 U4148 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3328) );
  NOR2_X1 U4149 ( .A1(n3354), .A2(n3328), .ZN(n3327) );
  AOI21_X1 U4150 ( .B1(n3328), .B2(n3354), .A(n3327), .ZN(n3329) );
  OAI211_X1 U4151 ( .C1(n3330), .C2(n3329), .A(n3474), .B(n4542), .ZN(n3358)
         );
  INV_X1 U4152 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3332) );
  NOR2_X1 U4153 ( .A1(n3354), .A2(n3332), .ZN(n3331) );
  AOI21_X1 U4154 ( .B1(n3332), .B2(n3354), .A(n3331), .ZN(n3351) );
  NAND2_X1 U4155 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3334), .ZN(n3347) );
  INV_X1 U4156 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4157 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3334), .B1(n4591), .B2(
        n3333), .ZN(n4497) );
  NAND2_X1 U4158 ( .A1(n3336), .A2(REG2_REG_9__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4159 ( .A1(n3336), .A2(REG2_REG_9__SCAN_IN), .B1(n3335), .B2(n4595), .ZN(n4475) );
  NAND2_X1 U4160 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4452), .ZN(n3341) );
  AOI22_X1 U4161 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4452), .B1(n4598), .B2(n3337), .ZN(n4460) );
  NAND2_X1 U4162 ( .A1(n3338), .A2(n4428), .ZN(n3340) );
  NAND2_X1 U4163 ( .A1(n3340), .A2(n3339), .ZN(n4459) );
  NAND2_X1 U4164 ( .A1(n4460), .A2(n4459), .ZN(n4458) );
  NAND2_X1 U4165 ( .A1(n4596), .A2(n3342), .ZN(n3343) );
  NAND2_X1 U4166 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4464), .ZN(n4463) );
  NAND2_X1 U4167 ( .A1(n4592), .A2(n3345), .ZN(n3346) );
  NAND2_X1 U4168 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U4169 ( .A1(n4588), .A2(n3348), .ZN(n3349) );
  NAND2_X1 U4170 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4508), .ZN(n4506) );
  OAI21_X1 U4171 ( .B1(n3351), .B2(n3470), .A(n4507), .ZN(n3350) );
  AOI21_X1 U4172 ( .B1(n3351), .B2(n3470), .A(n3350), .ZN(n3356) );
  NAND2_X1 U4173 ( .A1(REG3_REG_13__SCAN_IN), .A2(U3149), .ZN(n3574) );
  INV_X1 U4174 ( .A(n3574), .ZN(n3352) );
  AOI21_X1 U4175 ( .B1(n4541), .B2(ADDR_REG_13__SCAN_IN), .A(n3352), .ZN(n3353) );
  OAI21_X1 U4176 ( .B1(n4548), .B2(n3354), .A(n3353), .ZN(n3355) );
  NOR2_X1 U4177 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  NAND2_X1 U4178 ( .A1(n3358), .A2(n3357), .ZN(U3253) );
  NAND2_X1 U4179 ( .A1(n3993), .A2(n3681), .ZN(n3360) );
  NAND2_X1 U4180 ( .A1(n3371), .A2(n3058), .ZN(n3359) );
  NAND2_X1 U4181 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  XNOR2_X1 U4182 ( .A(n3361), .B(n3676), .ZN(n3393) );
  AND2_X1 U4183 ( .A1(n3371), .A2(n3681), .ZN(n3362) );
  AOI21_X1 U4184 ( .B1(n3993), .B2(n3686), .A(n3362), .ZN(n3392) );
  XNOR2_X1 U4185 ( .A(n3393), .B(n3392), .ZN(n3368) );
  INV_X1 U4186 ( .A(n3400), .ZN(n3367) );
  AOI21_X1 U4187 ( .B1(n3368), .B2(n3366), .A(n3367), .ZN(n3375) );
  NOR2_X1 U4188 ( .A1(STATE_REG_SCAN_IN), .A2(n2586), .ZN(n4479) );
  OAI22_X1 U4189 ( .A1(n3369), .A2(n4434), .B1(n4435), .B2(n4555), .ZN(n3370)
         );
  AOI211_X1 U4190 ( .C1(n3371), .C2(n4438), .A(n4479), .B(n3370), .ZN(n3374)
         );
  NAND2_X1 U4191 ( .A1(n3804), .A2(n3372), .ZN(n3373) );
  OAI211_X1 U4192 ( .C1(n3375), .C2(n3816), .A(n3374), .B(n3373), .ZN(U3228)
         );
  NAND2_X1 U4193 ( .A1(n3941), .A2(n3942), .ZN(n3883) );
  XNOR2_X1 U4194 ( .A(n3376), .B(n3883), .ZN(n3383) );
  XOR2_X1 U4195 ( .A(n3883), .B(n3377), .Z(n3380) );
  AOI22_X1 U4196 ( .A1(n3991), .A2(n4558), .B1(n4298), .B2(n3406), .ZN(n3378)
         );
  OAI21_X1 U4197 ( .B1(n3404), .B2(n4554), .A(n3378), .ZN(n3379) );
  AOI21_X1 U4198 ( .B1(n3380), .B2(n4254), .A(n3379), .ZN(n3381) );
  OAI21_X1 U4199 ( .B1(n3383), .B2(n3382), .A(n3381), .ZN(n4633) );
  INV_X1 U4200 ( .A(n4633), .ZN(n3391) );
  INV_X1 U4201 ( .A(n3383), .ZN(n4635) );
  NOR2_X1 U4202 ( .A1(n3385), .A2(n3384), .ZN(n4632) );
  NOR3_X1 U4203 ( .A1(n4632), .A2(n2362), .A3(n4263), .ZN(n3389) );
  INV_X1 U4204 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3387) );
  INV_X1 U4205 ( .A(n3386), .ZN(n3409) );
  OAI22_X1 U4206 ( .A1(n4290), .A2(n3387), .B1(n3409), .B2(n4264), .ZN(n3388)
         );
  AOI211_X1 U4207 ( .C1(n4635), .C2(n4573), .A(n3389), .B(n3388), .ZN(n3390)
         );
  OAI21_X1 U4208 ( .B1(n3391), .B2(n5040), .A(n3390), .ZN(U3280) );
  NAND2_X1 U4209 ( .A1(n3393), .A2(n3392), .ZN(n3398) );
  AND2_X1 U4210 ( .A1(n3400), .A2(n3398), .ZN(n3402) );
  NAND2_X1 U4211 ( .A1(n3992), .A2(n3681), .ZN(n3395) );
  NAND2_X1 U4212 ( .A1(n3406), .A2(n3058), .ZN(n3394) );
  NAND2_X1 U4213 ( .A1(n3395), .A2(n3394), .ZN(n3396) );
  XNOR2_X1 U4214 ( .A(n3396), .B(n3687), .ZN(n3447) );
  AND2_X1 U4215 ( .A1(n3406), .A2(n3681), .ZN(n3397) );
  AOI21_X1 U4216 ( .B1(n3992), .B2(n3686), .A(n3397), .ZN(n3445) );
  XNOR2_X1 U4217 ( .A(n3447), .B(n3445), .ZN(n3401) );
  AND2_X1 U4218 ( .A1(n3401), .A2(n3398), .ZN(n3399) );
  NAND2_X1 U4219 ( .A1(n3400), .A2(n3399), .ZN(n3449) );
  OAI211_X1 U4220 ( .C1(n3402), .C2(n3401), .A(n4443), .B(n3449), .ZN(n3408)
         );
  NOR2_X1 U4221 ( .A1(STATE_REG_SCAN_IN), .A2(n3403), .ZN(n4493) );
  OAI22_X1 U4222 ( .A1(n3404), .A2(n4434), .B1(n4435), .B2(n3451), .ZN(n3405)
         );
  AOI211_X1 U4223 ( .C1(n3406), .C2(n4438), .A(n4493), .B(n3405), .ZN(n3407)
         );
  OAI211_X1 U4224 ( .C1(n4448), .C2(n3409), .A(n3408), .B(n3407), .ZN(U3214)
         );
  NAND2_X1 U4225 ( .A1(n3410), .A2(n4619), .ZN(n3411) );
  OAI211_X1 U4226 ( .C1(n4552), .C2(n3413), .A(n3412), .B(n3411), .ZN(n3416)
         );
  MUX2_X1 U4227 ( .A(REG0_REG_9__SCAN_IN), .B(n3416), .S(n4645), .Z(n3414) );
  AOI21_X1 U4228 ( .B1(n3418), .B2(n2884), .A(n3414), .ZN(n3415) );
  INV_X1 U4229 ( .A(n3415), .ZN(U3485) );
  MUX2_X1 U4230 ( .A(REG1_REG_9__SCAN_IN), .B(n3416), .S(n4659), .Z(n3417) );
  AOI21_X1 U4231 ( .B1(n2879), .B2(n3418), .A(n3417), .ZN(n3419) );
  INV_X1 U4232 ( .A(n3419), .ZN(U3527) );
  INV_X1 U4233 ( .A(n3420), .ZN(n3421) );
  AOI21_X1 U4234 ( .B1(n4551), .B2(n3422), .A(n3421), .ZN(n3436) );
  INV_X1 U4235 ( .A(n3434), .ZN(n3423) );
  AOI21_X1 U4236 ( .B1(n3436), .B2(n3435), .A(n3423), .ZN(n3424) );
  XNOR2_X1 U4237 ( .A(n3557), .B(n3576), .ZN(n3881) );
  XNOR2_X1 U4238 ( .A(n3424), .B(n3881), .ZN(n3427) );
  OAI22_X1 U4239 ( .A1(n3824), .A2(n4274), .B1(n4552), .B2(n3576), .ZN(n3425)
         );
  AOI21_X1 U4240 ( .B1(n4282), .B2(n4557), .A(n3425), .ZN(n3426) );
  OAI21_X1 U4241 ( .B1(n3427), .B2(n4560), .A(n3426), .ZN(n3493) );
  INV_X1 U4242 ( .A(n3493), .ZN(n3433) );
  XOR2_X1 U4243 ( .A(n3881), .B(n3428), .Z(n3494) );
  OR2_X1 U4244 ( .A1(n3439), .A2(n3576), .ZN(n3429) );
  NAND2_X1 U4245 ( .A1(n2247), .A2(n3429), .ZN(n3499) );
  AOI22_X1 U4246 ( .A1(n5040), .A2(REG2_REG_13__SCAN_IN), .B1(n3578), .B2(
        n5034), .ZN(n3430) );
  OAI21_X1 U4247 ( .B1(n3499), .B2(n4263), .A(n3430), .ZN(n3431) );
  AOI21_X1 U4248 ( .B1(n3494), .B2(n5045), .A(n3431), .ZN(n3432) );
  OAI21_X1 U4249 ( .B1(n5040), .B2(n3433), .A(n3432), .ZN(U3277) );
  AND2_X1 U4250 ( .A1(n3435), .A2(n3434), .ZN(n3879) );
  XOR2_X1 U4251 ( .A(n3879), .B(n3436), .Z(n3437) );
  AOI222_X1 U4252 ( .A1(n4254), .A2(n3437), .B1(n3557), .B2(n4558), .C1(n3991), 
        .C2(n4282), .ZN(n3581) );
  XOR2_X1 U4253 ( .A(n3879), .B(n3438), .Z(n3584) );
  INV_X1 U4254 ( .A(n3439), .ZN(n3440) );
  OAI21_X1 U4255 ( .B1(n4565), .B2(n3582), .A(n3440), .ZN(n3589) );
  AOI22_X1 U4256 ( .A1(n5040), .A2(REG2_REG_12__SCAN_IN), .B1(n3467), .B2(
        n5034), .ZN(n3442) );
  NAND2_X1 U4257 ( .A1(n4148), .A2(n3461), .ZN(n3441) );
  OAI211_X1 U4258 ( .C1(n3589), .C2(n4263), .A(n3442), .B(n3441), .ZN(n3443)
         );
  AOI21_X1 U4259 ( .B1(n3584), .B2(n5045), .A(n3443), .ZN(n3444) );
  OAI21_X1 U4260 ( .B1(n3581), .B2(n5040), .A(n3444), .ZN(U3278) );
  INV_X1 U4261 ( .A(n3445), .ZN(n3446) );
  NAND2_X1 U4262 ( .A1(n3447), .A2(n3446), .ZN(n3448) );
  NAND2_X1 U4263 ( .A1(n3449), .A2(n3448), .ZN(n3502) );
  OAI22_X1 U4264 ( .A1(n3451), .A2(n3691), .B1(n3689), .B2(n4553), .ZN(n3450)
         );
  XNOR2_X1 U4265 ( .A(n3450), .B(n3676), .ZN(n3454) );
  OR2_X1 U4266 ( .A1(n3451), .A2(n3671), .ZN(n3453) );
  NAND2_X1 U4267 ( .A1(n4567), .A2(n3681), .ZN(n3452) );
  AND2_X1 U4268 ( .A1(n3453), .A2(n3452), .ZN(n3455) );
  NAND2_X1 U4269 ( .A1(n3454), .A2(n3455), .ZN(n3503) );
  NAND2_X1 U4270 ( .A1(n3502), .A2(n3503), .ZN(n3501) );
  INV_X1 U4271 ( .A(n3454), .ZN(n3457) );
  INV_X1 U4272 ( .A(n3455), .ZN(n3456) );
  NAND2_X1 U4273 ( .A1(n3457), .A2(n3456), .ZN(n3505) );
  NAND2_X1 U4274 ( .A1(n3501), .A2(n3505), .ZN(n3546) );
  NAND2_X1 U4275 ( .A1(n4557), .A2(n3681), .ZN(n3459) );
  NAND2_X1 U4276 ( .A1(n3461), .A2(n3058), .ZN(n3458) );
  NAND2_X1 U4277 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  XNOR2_X1 U4278 ( .A(n3460), .B(n3687), .ZN(n3568) );
  NAND2_X1 U4279 ( .A1(n4557), .A2(n3686), .ZN(n3463) );
  NAND2_X1 U4280 ( .A1(n3461), .A2(n3681), .ZN(n3462) );
  NAND2_X1 U4281 ( .A1(n3463), .A2(n3462), .ZN(n3567) );
  INV_X1 U4282 ( .A(n3567), .ZN(n3547) );
  XNOR2_X1 U4283 ( .A(n3568), .B(n3547), .ZN(n3464) );
  XNOR2_X1 U4284 ( .A(n3546), .B(n3464), .ZN(n3469) );
  AOI22_X1 U4285 ( .A1(n3810), .A2(n3991), .B1(n3814), .B2(n3557), .ZN(n3465)
         );
  NAND2_X1 U4286 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4509) );
  OAI211_X1 U4287 ( .C1(n3802), .C2(n3582), .A(n3465), .B(n4509), .ZN(n3466)
         );
  AOI21_X1 U4288 ( .B1(n3467), .B2(n3804), .A(n3466), .ZN(n3468) );
  OAI21_X1 U4289 ( .B1(n3469), .B2(n3816), .A(n3468), .ZN(U3221) );
  INV_X1 U4290 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3473) );
  INV_X1 U4291 ( .A(n4426), .ZN(n4029) );
  AND2_X1 U4292 ( .A1(n3470), .A2(REG2_REG_13__SCAN_IN), .ZN(n3471) );
  AOI211_X1 U4293 ( .C1(n3473), .C2(n3472), .A(n4044), .B(n4535), .ZN(n3480)
         );
  OAI211_X1 U4294 ( .C1(REG1_REG_14__SCAN_IN), .C2(n3475), .A(n4542), .B(n4031), .ZN(n3478) );
  NAND2_X1 U4295 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3558) );
  INV_X1 U4296 ( .A(n3558), .ZN(n3476) );
  AOI21_X1 U4297 ( .B1(n4541), .B2(ADDR_REG_14__SCAN_IN), .A(n3476), .ZN(n3477) );
  OAI211_X1 U4298 ( .C1(n4548), .C2(n4029), .A(n3478), .B(n3477), .ZN(n3479)
         );
  OR2_X1 U4299 ( .A1(n3480), .A2(n3479), .ZN(U3254) );
  OAI21_X1 U4300 ( .B1(n3482), .B2(n3892), .A(n3481), .ZN(n4365) );
  OAI21_X1 U4301 ( .B1(n3483), .B2(n3835), .A(n3511), .ZN(n3484) );
  NAND2_X1 U4302 ( .A1(n3484), .A2(n4254), .ZN(n3486) );
  AOI22_X1 U4303 ( .A1(n3612), .A2(n4558), .B1(n4298), .B2(n3555), .ZN(n3485)
         );
  OAI211_X1 U4304 ( .C1(n3487), .C2(n4554), .A(n3486), .B(n3485), .ZN(n3488)
         );
  AOI21_X1 U4305 ( .B1(n4365), .B2(n4563), .A(n3488), .ZN(n4369) );
  NAND2_X1 U4306 ( .A1(n2247), .A2(n3555), .ZN(n4366) );
  AND3_X1 U4307 ( .A1(n4367), .A2(n5032), .A3(n4366), .ZN(n3491) );
  INV_X1 U4308 ( .A(n3562), .ZN(n3489) );
  OAI22_X1 U4309 ( .A1(n4290), .A2(n3473), .B1(n3489), .B2(n4264), .ZN(n3490)
         );
  AOI211_X1 U4310 ( .C1(n4365), .C2(n4573), .A(n3491), .B(n3490), .ZN(n3492)
         );
  OAI21_X1 U4311 ( .B1(n4369), .B2(n5040), .A(n3492), .ZN(U3276) );
  INV_X1 U4312 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3495) );
  AOI21_X1 U4313 ( .B1(n3494), .B2(n4619), .A(n3493), .ZN(n3497) );
  MUX2_X1 U4314 ( .A(n3495), .B(n3497), .S(n4645), .Z(n3496) );
  OAI21_X1 U4315 ( .B1(n3499), .B2(n4417), .A(n3496), .ZN(U3493) );
  MUX2_X1 U4316 ( .A(n3328), .B(n3497), .S(n4659), .Z(n3498) );
  OAI21_X1 U4317 ( .B1(n4358), .B2(n3499), .A(n3498), .ZN(U3531) );
  AOI22_X1 U4318 ( .A1(n3810), .A2(n3992), .B1(n3814), .B2(n4557), .ZN(n3500)
         );
  NAND2_X1 U4319 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4499) );
  OAI211_X1 U4320 ( .C1(n3802), .C2(n4553), .A(n3500), .B(n4499), .ZN(n3508)
         );
  INV_X1 U4321 ( .A(n3501), .ZN(n3506) );
  AOI21_X1 U4322 ( .B1(n3505), .B2(n3503), .A(n3502), .ZN(n3504) );
  AOI211_X1 U4323 ( .C1(n3506), .C2(n3505), .A(n3816), .B(n3504), .ZN(n3507)
         );
  AOI211_X1 U4324 ( .C1(n3804), .C2(n4564), .A(n3508), .B(n3507), .ZN(n3509)
         );
  INV_X1 U4325 ( .A(n3509), .ZN(U3233) );
  XNOR2_X1 U4326 ( .A(n3510), .B(n3891), .ZN(n3592) );
  NAND2_X1 U4327 ( .A1(n3511), .A2(n3831), .ZN(n3513) );
  INV_X1 U4328 ( .A(n3891), .ZN(n3512) );
  XNOR2_X1 U4329 ( .A(n3513), .B(n3512), .ZN(n3515) );
  OAI22_X1 U4330 ( .A1(n3824), .A2(n4554), .B1(n3823), .B2(n4274), .ZN(n3514)
         );
  AOI21_X1 U4331 ( .B1(n3515), .B2(n4254), .A(n3514), .ZN(n3590) );
  NOR2_X1 U4332 ( .A1(n3590), .A2(n5040), .ZN(n3521) );
  AND2_X1 U4333 ( .A1(n4367), .A2(n3826), .ZN(n3516) );
  OR2_X1 U4334 ( .A1(n3516), .A2(n3533), .ZN(n3597) );
  INV_X1 U4335 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3517) );
  OAI22_X1 U4336 ( .A1(n4290), .A2(n3517), .B1(n3829), .B2(n4264), .ZN(n3518)
         );
  AOI21_X1 U4337 ( .B1(n3826), .B2(n4148), .A(n3518), .ZN(n3519) );
  OAI21_X1 U4338 ( .B1(n3597), .B2(n4263), .A(n3519), .ZN(n3520) );
  AOI211_X1 U4339 ( .C1(n3592), .C2(n5045), .A(n3521), .B(n3520), .ZN(n3522)
         );
  INV_X1 U4340 ( .A(n3522), .ZN(U3275) );
  OAI21_X1 U4341 ( .B1(n3524), .B2(n3525), .A(n3523), .ZN(n4364) );
  XNOR2_X1 U4342 ( .A(n3526), .B(n3525), .ZN(n3530) );
  NAND2_X1 U4343 ( .A1(n4439), .A2(n4298), .ZN(n3528) );
  NAND2_X1 U4344 ( .A1(n3612), .A2(n4282), .ZN(n3527) );
  OAI211_X1 U4345 ( .C1(n4436), .C2(n4274), .A(n3528), .B(n3527), .ZN(n3529)
         );
  AOI21_X1 U4346 ( .B1(n3530), .B2(n4254), .A(n3529), .ZN(n4362) );
  INV_X1 U4347 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3531) );
  OAI22_X1 U4348 ( .A1(n4290), .A2(n3531), .B1(n4447), .B2(n4264), .ZN(n3532)
         );
  INV_X1 U4349 ( .A(n3532), .ZN(n3535) );
  NOR2_X1 U4350 ( .A1(n3533), .A2(n3617), .ZN(n4359) );
  OR3_X1 U4351 ( .A1(n4360), .A2(n4359), .A3(n4263), .ZN(n3534) );
  OAI211_X1 U4352 ( .C1(n4362), .C2(n5040), .A(n3535), .B(n3534), .ZN(n3536)
         );
  INV_X1 U4353 ( .A(n3536), .ZN(n3537) );
  OAI21_X1 U4354 ( .B1(n4364), .B2(n4293), .A(n3537), .ZN(U3274) );
  NAND2_X1 U4355 ( .A1(n3557), .A2(n3681), .ZN(n3539) );
  NAND2_X1 U4356 ( .A1(n3541), .A2(n3058), .ZN(n3538) );
  NAND2_X1 U4357 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  XNOR2_X1 U4358 ( .A(n3540), .B(n3687), .ZN(n3548) );
  NAND2_X1 U4359 ( .A1(n3557), .A2(n3686), .ZN(n3543) );
  NAND2_X1 U4360 ( .A1(n3541), .A2(n3681), .ZN(n3542) );
  NAND2_X1 U4361 ( .A1(n3543), .A2(n3542), .ZN(n3549) );
  NAND2_X1 U4362 ( .A1(n3548), .A2(n3549), .ZN(n3566) );
  NAND2_X1 U4363 ( .A1(n3568), .A2(n3567), .ZN(n3544) );
  NAND2_X1 U4364 ( .A1(n3566), .A2(n3544), .ZN(n3545) );
  NOR2_X1 U4365 ( .A1(n3546), .A2(n3545), .ZN(n3553) );
  INV_X1 U4366 ( .A(n3568), .ZN(n3570) );
  NAND3_X1 U4367 ( .A1(n3566), .A2(n3547), .A3(n3570), .ZN(n3552) );
  INV_X1 U4368 ( .A(n3548), .ZN(n3551) );
  INV_X1 U4369 ( .A(n3549), .ZN(n3550) );
  NAND2_X1 U4370 ( .A1(n3551), .A2(n3550), .ZN(n3565) );
  OAI22_X1 U4371 ( .A1(n3824), .A2(n3691), .B1(n3560), .B2(n3689), .ZN(n3554)
         );
  XNOR2_X1 U4372 ( .A(n3554), .B(n3687), .ZN(n3606) );
  AOI22_X1 U4373 ( .A1(n3990), .A2(n3686), .B1(n3555), .B2(n3681), .ZN(n3608)
         );
  XNOR2_X1 U4374 ( .A(n3606), .B(n3608), .ZN(n3556) );
  XNOR2_X1 U4375 ( .A(n3607), .B(n3556), .ZN(n3564) );
  AOI22_X1 U4376 ( .A1(n3810), .A2(n3557), .B1(n3814), .B2(n3612), .ZN(n3559)
         );
  OAI211_X1 U4377 ( .C1(n3802), .C2(n3560), .A(n3559), .B(n3558), .ZN(n3561)
         );
  AOI21_X1 U4378 ( .B1(n3562), .B2(n3804), .A(n3561), .ZN(n3563) );
  OAI21_X1 U4379 ( .B1(n3564), .B2(n3816), .A(n3563), .ZN(U3212) );
  NAND2_X1 U4380 ( .A1(n3566), .A2(n3565), .ZN(n3573) );
  INV_X1 U4381 ( .A(n3546), .ZN(n3571) );
  OAI21_X1 U4382 ( .B1(n3546), .B2(n3568), .A(n3567), .ZN(n3569) );
  OAI21_X1 U4383 ( .B1(n3571), .B2(n3570), .A(n3569), .ZN(n3572) );
  XOR2_X1 U4384 ( .A(n3573), .B(n3572), .Z(n3580) );
  AOI22_X1 U4385 ( .A1(n3814), .A2(n3990), .B1(n3810), .B2(n4557), .ZN(n3575)
         );
  OAI211_X1 U4386 ( .C1(n3802), .C2(n3576), .A(n3575), .B(n3574), .ZN(n3577)
         );
  AOI21_X1 U4387 ( .B1(n3578), .B2(n3804), .A(n3577), .ZN(n3579) );
  OAI21_X1 U4388 ( .B1(n3580), .B2(n3816), .A(n3579), .ZN(U3231) );
  INV_X1 U4389 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4917) );
  OAI21_X1 U4390 ( .B1(n3582), .B2(n4552), .A(n3581), .ZN(n3583) );
  AOI21_X1 U4391 ( .B1(n4619), .B2(n3584), .A(n3583), .ZN(n3586) );
  MUX2_X1 U4392 ( .A(n4917), .B(n3586), .S(n4645), .Z(n3585) );
  OAI21_X1 U4393 ( .B1(n3589), .B2(n4417), .A(n3585), .ZN(U3491) );
  INV_X1 U4394 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3587) );
  MUX2_X1 U4395 ( .A(n3587), .B(n3586), .S(n4659), .Z(n3588) );
  OAI21_X1 U4396 ( .B1(n3589), .B2(n4358), .A(n3588), .ZN(U3530) );
  OAI21_X1 U4397 ( .B1(n3609), .B2(n4552), .A(n3590), .ZN(n3591) );
  AOI21_X1 U4398 ( .B1(n3592), .B2(n4619), .A(n3591), .ZN(n3594) );
  MUX2_X1 U4399 ( .A(n4788), .B(n3594), .S(n4645), .Z(n3593) );
  OAI21_X1 U4400 ( .B1(n3597), .B2(n4417), .A(n3593), .ZN(U3497) );
  INV_X1 U4401 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3595) );
  MUX2_X1 U4402 ( .A(n3595), .B(n3594), .S(n4659), .Z(n3596) );
  OAI21_X1 U4403 ( .B1(n4358), .B2(n3597), .A(n3596), .ZN(U3533) );
  NAND2_X1 U4404 ( .A1(n4228), .A2(n4227), .ZN(n3870) );
  XNOR2_X1 U4405 ( .A(n4230), .B(n3870), .ZN(n3599) );
  OAI22_X1 U4406 ( .A1(n3758), .A2(n4274), .B1(n3823), .B2(n4554), .ZN(n3598)
         );
  AOI21_X1 U4407 ( .B1(n3599), .B2(n4254), .A(n3598), .ZN(n4353) );
  XOR2_X1 U4408 ( .A(n3870), .B(n3600), .Z(n4356) );
  NAND2_X1 U4409 ( .A1(n4356), .A2(n5045), .ZN(n3605) );
  OAI21_X1 U4410 ( .B1(n4360), .B2(n4354), .A(n4283), .ZN(n4418) );
  INV_X1 U4411 ( .A(n4418), .ZN(n3603) );
  AOI22_X1 U4412 ( .A1(n5040), .A2(REG2_REG_17__SCAN_IN), .B1(n3761), .B2(
        n5034), .ZN(n3601) );
  OAI21_X1 U4413 ( .B1(n5039), .B2(n4354), .A(n3601), .ZN(n3602) );
  AOI21_X1 U4414 ( .B1(n3603), .B2(n5032), .A(n3602), .ZN(n3604) );
  OAI211_X1 U4415 ( .C1(n5040), .C2(n4353), .A(n3605), .B(n3604), .ZN(U3273)
         );
  OAI22_X1 U4416 ( .A1(n4433), .A2(n3691), .B1(n3689), .B2(n3609), .ZN(n3610)
         );
  XNOR2_X1 U4417 ( .A(n3610), .B(n3687), .ZN(n3613) );
  AND2_X1 U4418 ( .A1(n3826), .A2(n3681), .ZN(n3611) );
  AOI21_X1 U4419 ( .B1(n3612), .B2(n3686), .A(n3611), .ZN(n4440) );
  NOR2_X1 U4420 ( .A1(n3818), .A2(n4440), .ZN(n3622) );
  OR2_X1 U4421 ( .A1(n3823), .A2(n3671), .ZN(n3616) );
  NAND2_X1 U4422 ( .A1(n4439), .A2(n3681), .ZN(n3615) );
  NAND2_X1 U4423 ( .A1(n3616), .A2(n3615), .ZN(n3620) );
  OAI22_X1 U4424 ( .A1(n3823), .A2(n3691), .B1(n3617), .B2(n3689), .ZN(n3618)
         );
  XNOR2_X1 U4425 ( .A(n3618), .B(n3687), .ZN(n3619) );
  XOR2_X1 U4426 ( .A(n3620), .B(n3619), .Z(n4442) );
  NAND2_X1 U4427 ( .A1(n3819), .A2(n4442), .ZN(n3621) );
  OAI22_X1 U4428 ( .A1(n4436), .A2(n3691), .B1(n4354), .B2(n3689), .ZN(n3623)
         );
  XNOR2_X1 U4429 ( .A(n3623), .B(n3676), .ZN(n3756) );
  OR2_X1 U4430 ( .A1(n4436), .A2(n3671), .ZN(n3625) );
  OR2_X1 U4431 ( .A1(n3691), .A2(n4354), .ZN(n3624) );
  INV_X1 U4432 ( .A(n3756), .ZN(n3627) );
  INV_X1 U4433 ( .A(n3755), .ZN(n3626) );
  OAI22_X1 U4434 ( .A1(n3758), .A2(n3691), .B1(n4285), .B2(n3689), .ZN(n3628)
         );
  XNOR2_X1 U4435 ( .A(n3628), .B(n3687), .ZN(n3630) );
  OAI22_X1 U4436 ( .A1(n3758), .A2(n3671), .B1(n4285), .B2(n3691), .ZN(n3629)
         );
  NAND2_X1 U4437 ( .A1(n3630), .A2(n3629), .ZN(n3797) );
  NOR2_X1 U4438 ( .A1(n3630), .A2(n3629), .ZN(n3796) );
  AOI22_X1 U4439 ( .A1(n4235), .A2(n3686), .B1(n3681), .B2(n4256), .ZN(n3634)
         );
  NAND2_X1 U4440 ( .A1(n4235), .A2(n3681), .ZN(n3632) );
  NAND2_X1 U4441 ( .A1(n4256), .A2(n3058), .ZN(n3631) );
  NAND2_X1 U4442 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  XNOR2_X1 U4443 ( .A(n3633), .B(n3687), .ZN(n3636) );
  XOR2_X1 U4444 ( .A(n3634), .B(n3636), .Z(n3728) );
  INV_X1 U4445 ( .A(n3634), .ZN(n3635) );
  NAND2_X1 U4446 ( .A1(n4213), .A2(n3681), .ZN(n3639) );
  NAND2_X1 U4447 ( .A1(n3058), .A2(n4242), .ZN(n3638) );
  NAND2_X1 U4448 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  XNOR2_X1 U4449 ( .A(n3640), .B(n3687), .ZN(n3643) );
  NAND2_X1 U4450 ( .A1(n4213), .A2(n3686), .ZN(n3642) );
  NAND2_X1 U4451 ( .A1(n3681), .A2(n4242), .ZN(n3641) );
  NAND2_X1 U4452 ( .A1(n3642), .A2(n3641), .ZN(n3644) );
  NAND2_X1 U4453 ( .A1(n3643), .A2(n3644), .ZN(n3778) );
  INV_X1 U4454 ( .A(n3643), .ZN(n3646) );
  INV_X1 U4455 ( .A(n3644), .ZN(n3645) );
  NAND2_X1 U4456 ( .A1(n3646), .A2(n3645), .ZN(n3780) );
  NAND2_X1 U4457 ( .A1(n4236), .A2(n3681), .ZN(n3648) );
  NAND2_X1 U4458 ( .A1(n3058), .A2(n3650), .ZN(n3647) );
  NAND2_X1 U4459 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  XNOR2_X1 U4460 ( .A(n3649), .B(n3676), .ZN(n3736) );
  AND2_X1 U4461 ( .A1(n3681), .A2(n3650), .ZN(n3651) );
  AOI21_X1 U4462 ( .B1(n4236), .B2(n3686), .A(n3651), .ZN(n3735) );
  INV_X1 U4463 ( .A(n3736), .ZN(n3653) );
  INV_X1 U4464 ( .A(n3735), .ZN(n3652) );
  OAI22_X1 U4465 ( .A1(n3739), .A2(n3691), .B1(n4197), .B2(n3689), .ZN(n3654)
         );
  XNOR2_X1 U4466 ( .A(n3654), .B(n3687), .ZN(n3659) );
  AOI22_X1 U4467 ( .A1(n4214), .A2(n3686), .B1(n4203), .B2(n3681), .ZN(n3660)
         );
  XNOR2_X1 U4468 ( .A(n3659), .B(n3660), .ZN(n3790) );
  NAND2_X1 U4469 ( .A1(n3789), .A2(n3790), .ZN(n3718) );
  NAND2_X1 U4470 ( .A1(n4194), .A2(n3681), .ZN(n3656) );
  OR2_X1 U4471 ( .A1(n3689), .A2(n4186), .ZN(n3655) );
  NAND2_X1 U4472 ( .A1(n3656), .A2(n3655), .ZN(n3657) );
  XNOR2_X1 U4473 ( .A(n3657), .B(n3687), .ZN(n3666) );
  NOR2_X1 U4474 ( .A1(n3691), .A2(n4186), .ZN(n3658) );
  AOI21_X1 U4475 ( .B1(n4194), .B2(n3686), .A(n3658), .ZN(n3664) );
  XNOR2_X1 U4476 ( .A(n3666), .B(n3664), .ZN(n3719) );
  INV_X1 U4477 ( .A(n3659), .ZN(n3661) );
  NAND2_X1 U4478 ( .A1(n3661), .A2(n3660), .ZN(n3720) );
  NAND2_X1 U4479 ( .A1(n3718), .A2(n3662), .ZN(n3717) );
  NOR2_X1 U4480 ( .A1(n3691), .A2(n4166), .ZN(n3663) );
  AOI21_X1 U4481 ( .B1(n4141), .B2(n3686), .A(n3663), .ZN(n3668) );
  INV_X1 U4482 ( .A(n3664), .ZN(n3665) );
  NAND2_X1 U4483 ( .A1(n3666), .A2(n3665), .ZN(n3669) );
  NAND3_X1 U4484 ( .A1(n3717), .A2(n3668), .A3(n3669), .ZN(n3766) );
  OAI22_X1 U4485 ( .A1(n4183), .A2(n3691), .B1(n4166), .B2(n3689), .ZN(n3667)
         );
  XNOR2_X1 U4486 ( .A(n3667), .B(n3687), .ZN(n3768) );
  OAI22_X1 U4487 ( .A1(n4163), .A2(n3691), .B1(n4313), .B2(n3689), .ZN(n3670)
         );
  XNOR2_X1 U4488 ( .A(n3670), .B(n3687), .ZN(n3673) );
  OAI22_X1 U4489 ( .A1(n4163), .A2(n3671), .B1(n4313), .B2(n3691), .ZN(n3672)
         );
  NOR2_X1 U4490 ( .A1(n3673), .A2(n3672), .ZN(n3745) );
  NAND2_X1 U4491 ( .A1(n3673), .A2(n3672), .ZN(n3746) );
  NAND2_X1 U4492 ( .A1(n4142), .A2(n3681), .ZN(n3675) );
  OR2_X1 U4493 ( .A1(n3689), .A2(n4127), .ZN(n3674) );
  NAND2_X1 U4494 ( .A1(n3675), .A2(n3674), .ZN(n3677) );
  XNOR2_X1 U4495 ( .A(n3677), .B(n3676), .ZN(n3680) );
  NOR2_X1 U4496 ( .A1(n3691), .A2(n4127), .ZN(n3678) );
  AOI21_X1 U4497 ( .B1(n4142), .B2(n3686), .A(n3678), .ZN(n3679) );
  NOR2_X1 U4498 ( .A1(n3680), .A2(n3679), .ZN(n3807) );
  AOI22_X1 U4499 ( .A1(n3988), .A2(n3686), .B1(n3681), .B2(n4108), .ZN(n3685)
         );
  OAI22_X1 U4500 ( .A1(n4125), .A2(n3691), .B1(n3689), .B2(n4305), .ZN(n3682)
         );
  XNOR2_X1 U4501 ( .A(n3682), .B(n3687), .ZN(n3683) );
  XOR2_X1 U4502 ( .A(n3685), .B(n3683), .Z(n3711) );
  INV_X1 U4503 ( .A(n3683), .ZN(n3684) );
  AOI22_X1 U4504 ( .A1(n4102), .A2(n3686), .B1(n4092), .B2(n3681), .ZN(n3688)
         );
  XNOR2_X1 U4505 ( .A(n3688), .B(n3687), .ZN(n3694) );
  OAI22_X1 U4506 ( .A1(n3692), .A2(n3691), .B1(n3690), .B2(n3689), .ZN(n3693)
         );
  XNOR2_X1 U4507 ( .A(n3694), .B(n3693), .ZN(n3695) );
  XNOR2_X1 U4508 ( .A(n3696), .B(n3695), .ZN(n3703) );
  INV_X1 U4509 ( .A(n3697), .ZN(n4094) );
  NAND2_X1 U4510 ( .A1(n3988), .A2(n3810), .ZN(n3699) );
  AOI22_X1 U4511 ( .A1(n4438), .A2(n4092), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3698) );
  OAI211_X1 U4512 ( .C1(n4094), .C2(n4448), .A(n3699), .B(n3698), .ZN(n3700)
         );
  INV_X1 U4513 ( .A(n3700), .ZN(n3702) );
  NAND2_X1 U4514 ( .A1(n3987), .A2(n3814), .ZN(n3701) );
  OAI211_X1 U4515 ( .C1(n3703), .C2(n3816), .A(n3702), .B(n3701), .ZN(U3217)
         );
  NAND2_X1 U4516 ( .A1(n3704), .A2(n4443), .ZN(n3708) );
  AOI22_X1 U4517 ( .A1(REG3_REG_0__SCAN_IN), .A2(n3706), .B1(n4438), .B2(n3705), .ZN(n3707) );
  OAI211_X1 U4518 ( .C1(n3709), .C2(n4435), .A(n3708), .B(n3707), .ZN(U3229)
         );
  XNOR2_X1 U4519 ( .A(n3710), .B(n3711), .ZN(n3716) );
  NAND2_X1 U4520 ( .A1(n4142), .A2(n3810), .ZN(n3713) );
  AOI22_X1 U4521 ( .A1(n4438), .A2(n4108), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3712) );
  OAI211_X1 U4522 ( .C1(n4448), .C2(n4110), .A(n3713), .B(n3712), .ZN(n3714)
         );
  AOI21_X1 U4523 ( .B1(n4102), .B2(n3814), .A(n3714), .ZN(n3715) );
  OAI21_X1 U4524 ( .B1(n3716), .B2(n3816), .A(n3715), .ZN(U3211) );
  NAND2_X1 U4525 ( .A1(n3717), .A2(n4443), .ZN(n3727) );
  AOI21_X1 U4526 ( .B1(n3718), .B2(n3720), .A(n3719), .ZN(n3726) );
  INV_X1 U4527 ( .A(n3721), .ZN(n4187) );
  OAI22_X1 U4528 ( .A1(n3802), .A2(n4186), .B1(STATE_REG_SCAN_IN), .B2(n3722), 
        .ZN(n3724) );
  OAI22_X1 U4529 ( .A1(n4183), .A2(n4435), .B1(n3739), .B2(n4434), .ZN(n3723)
         );
  AOI211_X1 U4530 ( .C1(n4187), .C2(n3804), .A(n3724), .B(n3723), .ZN(n3725)
         );
  OAI21_X1 U4531 ( .B1(n3727), .B2(n3726), .A(n3725), .ZN(U3213) );
  XNOR2_X1 U4532 ( .A(n3729), .B(n3728), .ZN(n3730) );
  NAND2_X1 U4533 ( .A1(n3730), .A2(n4443), .ZN(n3733) );
  INV_X1 U4534 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4839) );
  NOR2_X1 U4535 ( .A1(n4839), .A2(STATE_REG_SCAN_IN), .ZN(n4067) );
  INV_X1 U4536 ( .A(n4213), .ZN(n4260) );
  OAI22_X1 U4537 ( .A1(n4260), .A2(n4435), .B1(n4434), .B2(n3758), .ZN(n3731)
         );
  AOI211_X1 U4538 ( .C1(n4256), .C2(n4438), .A(n4067), .B(n3731), .ZN(n3732)
         );
  OAI211_X1 U4539 ( .C1(n4448), .C2(n4265), .A(n3733), .B(n3732), .ZN(U3216)
         );
  XNOR2_X1 U4540 ( .A(n3736), .B(n3735), .ZN(n3737) );
  XNOR2_X1 U4541 ( .A(n3734), .B(n3737), .ZN(n3743) );
  OAI22_X1 U4542 ( .A1(n3802), .A2(n4335), .B1(STATE_REG_SCAN_IN), .B2(n3738), 
        .ZN(n3741) );
  OAI22_X1 U4543 ( .A1(n3739), .A2(n4435), .B1(n4260), .B2(n4434), .ZN(n3740)
         );
  AOI211_X1 U4544 ( .C1(n4220), .C2(n3804), .A(n3741), .B(n3740), .ZN(n3742)
         );
  OAI21_X1 U4545 ( .B1(n3743), .B2(n3816), .A(n3742), .ZN(U3220) );
  INV_X1 U4546 ( .A(n3745), .ZN(n3747) );
  NAND2_X1 U4547 ( .A1(n3747), .A2(n3746), .ZN(n3748) );
  XNOR2_X1 U4548 ( .A(n3744), .B(n3748), .ZN(n3753) );
  OAI22_X1 U4549 ( .A1(n3802), .A2(n4313), .B1(STATE_REG_SCAN_IN), .B2(n3749), 
        .ZN(n3750) );
  AOI21_X1 U4550 ( .B1(n4141), .B2(n3810), .A(n3750), .ZN(n3752) );
  AOI22_X1 U4551 ( .A1(n4142), .A2(n3814), .B1(n3804), .B2(n4146), .ZN(n3751)
         );
  OAI211_X1 U4552 ( .C1(n3753), .C2(n3816), .A(n3752), .B(n3751), .ZN(U3222)
         );
  XNOR2_X1 U4553 ( .A(n3756), .B(n3755), .ZN(n3757) );
  XNOR2_X1 U4554 ( .A(n3754), .B(n3757), .ZN(n3764) );
  NOR2_X1 U4555 ( .A1(STATE_REG_SCAN_IN), .A2(n2672), .ZN(n4540) );
  OAI22_X1 U4556 ( .A1(n3823), .A2(n4434), .B1(n4435), .B2(n3758), .ZN(n3759)
         );
  AOI211_X1 U4557 ( .C1(n3760), .C2(n4438), .A(n4540), .B(n3759), .ZN(n3763)
         );
  NAND2_X1 U4558 ( .A1(n3804), .A2(n3761), .ZN(n3762) );
  OAI211_X1 U4559 ( .C1(n3764), .C2(n3816), .A(n3763), .B(n3762), .ZN(U3225)
         );
  INV_X1 U4560 ( .A(n3766), .ZN(n3767) );
  NOR2_X1 U4561 ( .A1(n3765), .A2(n3767), .ZN(n3769) );
  XNOR2_X1 U4562 ( .A(n3769), .B(n3768), .ZN(n3775) );
  INV_X1 U4563 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3770) );
  OAI22_X1 U4564 ( .A1(n3802), .A2(n4166), .B1(STATE_REG_SCAN_IN), .B2(n3770), 
        .ZN(n3773) );
  OAI22_X1 U4565 ( .A1(n4163), .A2(n4435), .B1(n3771), .B2(n4434), .ZN(n3772)
         );
  AOI211_X1 U4566 ( .C1(n4167), .C2(n3804), .A(n3773), .B(n3772), .ZN(n3774)
         );
  OAI21_X1 U4567 ( .B1(n3775), .B2(n3816), .A(n3774), .ZN(U3226) );
  INV_X1 U4568 ( .A(n3776), .ZN(n3781) );
  AOI21_X1 U4569 ( .B1(n3780), .B2(n3778), .A(n3777), .ZN(n3779) );
  AOI21_X1 U4570 ( .B1(n3781), .B2(n3780), .A(n3779), .ZN(n3788) );
  INV_X1 U4571 ( .A(n4244), .ZN(n3786) );
  INV_X1 U4572 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4747) );
  OAI22_X1 U4573 ( .A1(n3802), .A2(n3782), .B1(STATE_REG_SCAN_IN), .B2(n4747), 
        .ZN(n3785) );
  INV_X1 U4574 ( .A(n4236), .ZN(n3783) );
  INV_X1 U4575 ( .A(n4235), .ZN(n4275) );
  OAI22_X1 U4576 ( .A1(n3783), .A2(n4435), .B1(n4434), .B2(n4275), .ZN(n3784)
         );
  AOI211_X1 U4577 ( .C1(n3786), .C2(n3804), .A(n3785), .B(n3784), .ZN(n3787)
         );
  OAI21_X1 U4578 ( .B1(n3788), .B2(n3816), .A(n3787), .ZN(U3230) );
  OAI21_X1 U4579 ( .B1(n3790), .B2(n3789), .A(n3718), .ZN(n3791) );
  NAND2_X1 U4580 ( .A1(n3791), .A2(n4443), .ZN(n3795) );
  AOI22_X1 U4581 ( .A1(n4438), .A2(n4203), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3794) );
  AOI22_X1 U4582 ( .A1(n4194), .A2(n3814), .B1(n3810), .B2(n4236), .ZN(n3793)
         );
  NAND2_X1 U4583 ( .A1(n3804), .A2(n4204), .ZN(n3792) );
  NAND4_X1 U4584 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(U3232)
         );
  NAND2_X1 U4585 ( .A1(n2462), .A2(n3797), .ZN(n3798) );
  XNOR2_X1 U4586 ( .A(n3799), .B(n3798), .ZN(n3806) );
  INV_X1 U4587 ( .A(n3800), .ZN(n4286) );
  AOI22_X1 U4588 ( .A1(n3810), .A2(n4281), .B1(n3814), .B2(n4235), .ZN(n3801)
         );
  NAND2_X1 U4589 ( .A1(REG3_REG_18__SCAN_IN), .A2(U3149), .ZN(n4038) );
  OAI211_X1 U4590 ( .C1(n3802), .C2(n4285), .A(n3801), .B(n4038), .ZN(n3803)
         );
  AOI21_X1 U4591 ( .B1(n4286), .B2(n3804), .A(n3803), .ZN(n3805) );
  OAI21_X1 U4592 ( .B1(n3806), .B2(n3816), .A(n3805), .ZN(U3235) );
  NOR2_X1 U4593 ( .A1(n3807), .A2(n2267), .ZN(n3808) );
  XNOR2_X1 U4594 ( .A(n3809), .B(n3808), .ZN(n3817) );
  NAND2_X1 U4595 ( .A1(n4122), .A2(n3810), .ZN(n3812) );
  AOI22_X1 U4596 ( .A1(n4438), .A2(n4121), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3811) );
  OAI211_X1 U4597 ( .C1(n4448), .C2(n4129), .A(n3812), .B(n3811), .ZN(n3813)
         );
  AOI21_X1 U4598 ( .B1(n3988), .B2(n3814), .A(n3813), .ZN(n3815) );
  OAI21_X1 U4599 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(U3237) );
  INV_X1 U4600 ( .A(n3819), .ZN(n3820) );
  NOR2_X1 U4601 ( .A1(n3818), .A2(n3820), .ZN(n3821) );
  XNOR2_X1 U4602 ( .A(n3821), .B(n4440), .ZN(n3822) );
  NAND2_X1 U4603 ( .A1(n3822), .A2(n4443), .ZN(n3828) );
  AND2_X1 U4604 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4521) );
  OAI22_X1 U4605 ( .A1(n3824), .A2(n4434), .B1(n4435), .B2(n3823), .ZN(n3825)
         );
  AOI211_X1 U4606 ( .C1(n3826), .C2(n4438), .A(n4521), .B(n3825), .ZN(n3827)
         );
  OAI211_X1 U4607 ( .C1(n4448), .C2(n3829), .A(n3828), .B(n3827), .ZN(U3238)
         );
  INV_X1 U4608 ( .A(n4076), .ZN(n3872) );
  AND2_X1 U4609 ( .A1(n2529), .A2(DATAI_30_), .ZN(n4299) );
  AOI211_X1 U4610 ( .C1(n3958), .C2(n3830), .A(n3866), .B(n3898), .ZN(n3964)
         );
  NAND2_X1 U4611 ( .A1(n3831), .A2(n3834), .ZN(n3948) );
  NAND2_X1 U4612 ( .A1(n3833), .A2(n3832), .ZN(n3931) );
  NAND2_X1 U4613 ( .A1(n3931), .A2(n3834), .ZN(n3947) );
  OAI21_X1 U4614 ( .B1(n3835), .B2(n3948), .A(n3947), .ZN(n3837) );
  AOI211_X1 U4615 ( .C1(n3837), .C2(n3952), .A(n2425), .B(n3953), .ZN(n3840)
         );
  INV_X1 U4616 ( .A(n3838), .ZN(n3839) );
  NOR2_X1 U4617 ( .A1(n3840), .A2(n3839), .ZN(n3842) );
  OAI21_X1 U4618 ( .B1(n3842), .B2(n3841), .A(n3958), .ZN(n3847) );
  OR2_X1 U4619 ( .A1(n3844), .A2(n3843), .ZN(n3853) );
  INV_X1 U4620 ( .A(n3845), .ZN(n3859) );
  AND2_X1 U4621 ( .A1(n2529), .A2(DATAI_31_), .ZN(n3873) );
  INV_X1 U4622 ( .A(n3873), .ZN(n4077) );
  NAND2_X1 U4623 ( .A1(n4076), .A2(n4077), .ZN(n3971) );
  INV_X1 U4624 ( .A(n3971), .ZN(n3846) );
  AOI21_X1 U4625 ( .B1(n4299), .B2(n3859), .A(n3846), .ZN(n3874) );
  OAI21_X1 U4626 ( .B1(n3987), .B2(n3848), .A(n3874), .ZN(n3852) );
  AOI211_X1 U4627 ( .C1(n3964), .C2(n3847), .A(n3853), .B(n3852), .ZN(n3857)
         );
  AND2_X1 U4628 ( .A1(n3987), .A2(n3848), .ZN(n3849) );
  OR2_X1 U4629 ( .A1(n3850), .A2(n3849), .ZN(n3965) );
  INV_X1 U4630 ( .A(n3965), .ZN(n3854) );
  NAND3_X1 U4631 ( .A1(n4105), .A2(n3854), .A3(n3851), .ZN(n3855) );
  AOI21_X1 U4632 ( .B1(n3854), .B2(n3853), .A(n3852), .ZN(n3969) );
  AOI22_X1 U4633 ( .A1(n3857), .A2(n3856), .B1(n3855), .B2(n3969), .ZN(n3858)
         );
  AOI21_X1 U4634 ( .B1(n3872), .B2(n4299), .A(n3858), .ZN(n3863) );
  NOR2_X1 U4635 ( .A1(n3859), .A2(n4299), .ZN(n3871) );
  INV_X1 U4636 ( .A(n3871), .ZN(n3860) );
  AOI21_X1 U4637 ( .B1(n3860), .B2(n4076), .A(n4077), .ZN(n3862) );
  OR3_X1 U4638 ( .A1(n3863), .A2(n3862), .A3(n3861), .ZN(n3978) );
  INV_X1 U4639 ( .A(n4116), .ZN(n3865) );
  OR2_X1 U4640 ( .A1(n3866), .A2(n3865), .ZN(n4137) );
  NAND2_X1 U4641 ( .A1(n4155), .A2(n3867), .ZN(n4178) );
  AND2_X1 U4642 ( .A1(n3869), .A2(n3868), .ZN(n4234) );
  XNOR2_X1 U4643 ( .A(n4235), .B(n4262), .ZN(n4252) );
  NOR4_X1 U4644 ( .A1(n4234), .A2(n4276), .A3(n4252), .A4(n3870), .ZN(n3878)
         );
  AOI21_X1 U4645 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3973) );
  AND4_X1 U4646 ( .A1(n3875), .A2(n4105), .A3(n3973), .A4(n3874), .ZN(n3876)
         );
  NAND4_X1 U4647 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3880)
         );
  NOR4_X1 U4648 ( .A1(n4178), .A2(n3881), .A3(n3880), .A4(n4604), .ZN(n3897)
         );
  NOR4_X1 U4649 ( .A1(n4550), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3896)
         );
  NOR4_X1 U4650 ( .A1(n2788), .A2(n2786), .A3(n3886), .A4(n3885), .ZN(n3895)
         );
  NAND4_X1 U4651 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3893)
         );
  NOR4_X1 U4652 ( .A1(n4200), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3894)
         );
  NAND4_X1 U4653 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3901)
         );
  NAND2_X1 U4654 ( .A1(n2385), .A2(n3899), .ZN(n4158) );
  INV_X1 U4655 ( .A(n3960), .ZN(n3900) );
  INV_X1 U4656 ( .A(n4212), .ZN(n4216) );
  NOR4_X1 U4657 ( .A1(n4137), .A2(n3901), .A3(n4158), .A4(n4216), .ZN(n3905)
         );
  INV_X1 U4658 ( .A(n3902), .ZN(n3904) );
  NAND2_X1 U4659 ( .A1(n3904), .A2(n3903), .ZN(n4118) );
  NAND3_X1 U4660 ( .A1(n2776), .A2(n3905), .A3(n4118), .ZN(n3976) );
  NOR2_X1 U4661 ( .A1(n4125), .A2(n4108), .ZN(n3968) );
  OAI211_X1 U4662 ( .C1(n2389), .C2(n4423), .A(n3908), .B(n3907), .ZN(n3911)
         );
  NAND3_X1 U4663 ( .A1(n3911), .A2(n3910), .A3(n3909), .ZN(n3914) );
  NAND3_X1 U4664 ( .A1(n3914), .A2(n3913), .A3(n3912), .ZN(n3917) );
  NAND3_X1 U4665 ( .A1(n3917), .A2(n3916), .A3(n3915), .ZN(n3920) );
  NAND4_X1 U4666 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3935), .ZN(n3923)
         );
  NAND3_X1 U4667 ( .A1(n3923), .A2(n3922), .A3(n3921), .ZN(n3930) );
  AND2_X1 U4668 ( .A1(n3925), .A2(n3924), .ZN(n3937) );
  INV_X1 U4669 ( .A(n3926), .ZN(n3929) );
  INV_X1 U4670 ( .A(n3927), .ZN(n3928) );
  AOI211_X1 U4671 ( .C1(n3930), .C2(n3937), .A(n3929), .B(n3928), .ZN(n3933)
         );
  NOR3_X1 U4672 ( .A1(n3933), .A2(n3932), .A3(n3931), .ZN(n3945) );
  INV_X1 U4673 ( .A(n3934), .ZN(n3938) );
  NAND4_X1 U4674 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3940)
         );
  INV_X1 U4675 ( .A(n3947), .ZN(n3939) );
  AOI21_X1 U4676 ( .B1(n3941), .B2(n3940), .A(n3939), .ZN(n3944) );
  OAI211_X1 U4677 ( .C1(n3945), .C2(n3944), .A(n3943), .B(n3942), .ZN(n3951)
         );
  INV_X1 U4678 ( .A(n3946), .ZN(n3949) );
  OAI21_X1 U4679 ( .B1(n3949), .B2(n3948), .A(n3947), .ZN(n3950) );
  AOI21_X1 U4680 ( .B1(n3951), .B2(n3950), .A(n2425), .ZN(n3956) );
  INV_X1 U4681 ( .A(n3952), .ZN(n3955) );
  INV_X1 U4682 ( .A(n3953), .ZN(n3954) );
  OAI21_X1 U4683 ( .B1(n3956), .B2(n3955), .A(n3954), .ZN(n3957) );
  AND2_X1 U4684 ( .A1(n3957), .A2(n4173), .ZN(n3961) );
  OAI211_X1 U4685 ( .C1(n3961), .C2(n3960), .A(n3959), .B(n3958), .ZN(n3963)
         );
  AOI21_X1 U4686 ( .B1(n3964), .B2(n3963), .A(n3962), .ZN(n3966) );
  NOR4_X1 U4687 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3974)
         );
  INV_X1 U4688 ( .A(n3973), .ZN(n3970) );
  AOI21_X1 U4689 ( .B1(n3971), .B2(n3970), .A(n3969), .ZN(n3972) );
  AOI21_X1 U4690 ( .B1(n3974), .B2(n3973), .A(n3972), .ZN(n3975) );
  MUX2_X1 U4691 ( .A(n3976), .B(n3975), .S(n2782), .Z(n3977) );
  NAND2_X1 U4692 ( .A1(n3978), .A2(n3977), .ZN(n3979) );
  XNOR2_X1 U4693 ( .A(n3979), .B(n4425), .ZN(n3986) );
  NOR2_X1 U4694 ( .A1(n3981), .A2(n3980), .ZN(n3984) );
  OAI21_X1 U4695 ( .B1(n3985), .B2(n3982), .A(B_REG_SCAN_IN), .ZN(n3983) );
  OAI22_X1 U4696 ( .A1(n3986), .A2(n3985), .B1(n3984), .B2(n3983), .ZN(U3239)
         );
  MUX2_X1 U4697 ( .A(DATAO_REG_29__SCAN_IN), .B(n3987), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4698 ( .A(DATAO_REG_28__SCAN_IN), .B(n4102), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4699 ( .A(DATAO_REG_27__SCAN_IN), .B(n3988), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4700 ( .A(DATAO_REG_24__SCAN_IN), .B(n4141), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4701 ( .A(DATAO_REG_22__SCAN_IN), .B(n4214), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4702 ( .A(DATAO_REG_21__SCAN_IN), .B(n4236), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4703 ( .A(DATAO_REG_19__SCAN_IN), .B(n4235), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4704 ( .A(DATAO_REG_18__SCAN_IN), .B(n4257), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4705 ( .A(DATAO_REG_17__SCAN_IN), .B(n4281), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4706 ( .A(DATAO_REG_16__SCAN_IN), .B(n3989), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4707 ( .A(DATAO_REG_14__SCAN_IN), .B(n3990), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4708 ( .A(DATAO_REG_12__SCAN_IN), .B(n4557), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4709 ( .A(DATAO_REG_11__SCAN_IN), .B(n3991), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4710 ( .A(DATAO_REG_10__SCAN_IN), .B(n3992), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4711 ( .A(DATAO_REG_9__SCAN_IN), .B(n3993), .S(U4043), .Z(U3559) );
  MUX2_X1 U4712 ( .A(DATAO_REG_7__SCAN_IN), .B(n3994), .S(U4043), .Z(U3557) );
  MUX2_X1 U4713 ( .A(DATAO_REG_6__SCAN_IN), .B(n3995), .S(U4043), .Z(U3556) );
  MUX2_X1 U4714 ( .A(DATAO_REG_5__SCAN_IN), .B(n3996), .S(U4043), .Z(U3555) );
  MUX2_X1 U4715 ( .A(DATAO_REG_3__SCAN_IN), .B(n3997), .S(U4043), .Z(U3553) );
  MUX2_X1 U4716 ( .A(DATAO_REG_2__SCAN_IN), .B(n2993), .S(U4043), .Z(U3552) );
  MUX2_X1 U4717 ( .A(DATAO_REG_1__SCAN_IN), .B(n2511), .S(U4043), .Z(U3551) );
  INV_X1 U4718 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4646) );
  NAND3_X1 U4719 ( .A1(n4542), .A2(IR_REG_0__SCAN_IN), .A3(n4646), .ZN(n4005)
         );
  AOI22_X1 U4720 ( .A1(n4541), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4004) );
  AOI21_X1 U4721 ( .B1(n4646), .B2(n3998), .A(n3999), .ZN(n4000) );
  MUX2_X1 U4722 ( .A(n4000), .B(n3999), .S(IR_REG_0__SCAN_IN), .Z(n4002) );
  NAND2_X1 U4723 ( .A1(n4002), .A2(n4001), .ZN(n4003) );
  NAND3_X1 U4724 ( .A1(n4005), .A2(n4004), .A3(n4003), .ZN(U3240) );
  OAI211_X1 U4725 ( .C1(n4008), .C2(n4007), .A(n4542), .B(n4006), .ZN(n4015)
         );
  OAI211_X1 U4726 ( .C1(n2918), .C2(n4011), .A(n4507), .B(n4010), .ZN(n4014)
         );
  INV_X1 U4727 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U4728 ( .A1(STATE_REG_SCAN_IN), .A2(n4940), .ZN(n4012) );
  AOI21_X1 U4729 ( .B1(n4541), .B2(ADDR_REG_1__SCAN_IN), .A(n4012), .ZN(n4013)
         );
  NAND4_X1 U4730 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(U3241)
         );
  NAND2_X1 U4731 ( .A1(n4017), .A2(n4429), .ZN(n4028) );
  OAI211_X1 U4732 ( .C1(n4020), .C2(n4019), .A(n4542), .B(n4018), .ZN(n4027)
         );
  OAI211_X1 U4733 ( .C1(n4023), .C2(n4022), .A(n4507), .B(n4021), .ZN(n4026)
         );
  AOI21_X1 U4734 ( .B1(n4541), .B2(ADDR_REG_5__SCAN_IN), .A(n4024), .ZN(n4025)
         );
  NAND4_X1 U4735 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(U3245)
         );
  XOR2_X1 U4736 ( .A(REG1_REG_18__SCAN_IN), .B(n4064), .Z(n4058) );
  NOR2_X1 U4737 ( .A1(n4051), .A2(REG1_REG_17__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U4738 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4047), .ZN(n4033) );
  INV_X1 U4739 ( .A(n4047), .ZN(n4587) );
  AOI22_X1 U4740 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4047), .B1(n4587), .B2(
        n3595), .ZN(n4524) );
  OR2_X1 U4741 ( .A1(n4030), .A2(n4029), .ZN(n4032) );
  NAND2_X1 U4742 ( .A1(n4032), .A2(n4031), .ZN(n4523) );
  NOR2_X1 U4743 ( .A1(n4048), .A2(n4034), .ZN(n4035) );
  INV_X1 U4744 ( .A(n4048), .ZN(n4586) );
  INV_X1 U4745 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4746 ( .A1(n4051), .A2(n4036), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4584), .ZN(n4543) );
  NOR2_X1 U4747 ( .A1(n4544), .A2(n4543), .ZN(n4545) );
  NOR2_X1 U4748 ( .A1(n4037), .A2(n4545), .ZN(n4059) );
  XOR2_X1 U4749 ( .A(n4058), .B(n4059), .Z(n4056) );
  INV_X1 U4750 ( .A(n4064), .ZN(n4041) );
  INV_X1 U4751 ( .A(n4038), .ZN(n4039) );
  AOI21_X1 U4752 ( .B1(n4541), .B2(ADDR_REG_18__SCAN_IN), .A(n4039), .ZN(n4040) );
  OAI21_X1 U4753 ( .B1(n4548), .B2(n4041), .A(n4040), .ZN(n4055) );
  INV_X1 U4754 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U4755 ( .A1(n4064), .A2(n4912), .ZN(n4042) );
  AOI21_X1 U4756 ( .B1(n4064), .B2(n4912), .A(n4042), .ZN(n4053) );
  NOR2_X1 U4757 ( .A1(n4051), .A2(REG2_REG_17__SCAN_IN), .ZN(n4043) );
  AOI21_X1 U4758 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4051), .A(n4043), .ZN(n4538) );
  NOR2_X1 U4759 ( .A1(n4045), .A2(n4044), .ZN(n4519) );
  NAND2_X1 U4760 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4047), .ZN(n4046) );
  OAI21_X1 U4761 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4047), .A(n4046), .ZN(n4518) );
  NOR2_X1 U4762 ( .A1(n4519), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U4763 ( .A1(n4049), .A2(n4586), .ZN(n4050) );
  AOI211_X1 U4764 ( .C1(n4053), .C2(n4052), .A(n4063), .B(n4535), .ZN(n4054)
         );
  AOI211_X1 U4765 ( .C1(n4056), .C2(n4542), .A(n4055), .B(n4054), .ZN(n4057)
         );
  INV_X1 U4766 ( .A(n4057), .ZN(U3258) );
  AOI22_X1 U4767 ( .A1(n4059), .A2(n4058), .B1(n4064), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n4062) );
  INV_X1 U4768 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4060) );
  MUX2_X1 U4769 ( .A(REG1_REG_19__SCAN_IN), .B(n4060), .S(n4069), .Z(n4061) );
  XNOR2_X1 U4770 ( .A(n4062), .B(n4061), .ZN(n4073) );
  INV_X1 U4771 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4065) );
  MUX2_X1 U4772 ( .A(n4065), .B(REG2_REG_19__SCAN_IN), .S(n4069), .Z(n4066) );
  AOI21_X1 U4773 ( .B1(n4541), .B2(ADDR_REG_19__SCAN_IN), .A(n4067), .ZN(n4068) );
  OAI21_X1 U4774 ( .B1(n4548), .B2(n4069), .A(n4068), .ZN(n4070) );
  OAI21_X1 U4775 ( .B1(n4074), .B2(n4073), .A(n4072), .ZN(U3259) );
  XNOR2_X1 U4776 ( .A(n4296), .B(n4077), .ZN(n4375) );
  NAND2_X1 U4777 ( .A1(n4076), .A2(n4075), .ZN(n4301) );
  OAI21_X1 U4778 ( .B1(n4077), .B2(n4552), .A(n4301), .ZN(n4373) );
  NAND2_X1 U4779 ( .A1(n4373), .A2(n4290), .ZN(n4079) );
  NAND2_X1 U4780 ( .A1(n5040), .A2(REG2_REG_31__SCAN_IN), .ZN(n4078) );
  OAI211_X1 U4781 ( .C1(n4375), .C2(n4263), .A(n4079), .B(n4078), .ZN(U3260)
         );
  INV_X1 U4782 ( .A(n4080), .ZN(n4089) );
  AOI22_X1 U4783 ( .A1(n4148), .A2(n4081), .B1(n5040), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n4088) );
  INV_X1 U4784 ( .A(n4082), .ZN(n4086) );
  OAI22_X1 U4785 ( .A1(n4084), .A2(n4263), .B1(n4083), .B2(n4264), .ZN(n4085)
         );
  OAI21_X1 U4786 ( .B1(n4086), .B2(n4085), .A(n4290), .ZN(n4087) );
  OAI211_X1 U4787 ( .C1(n4089), .C2(n4293), .A(n4088), .B(n4087), .ZN(U3354)
         );
  NAND2_X1 U4788 ( .A1(n4090), .A2(n5045), .ZN(n4098) );
  INV_X1 U4789 ( .A(n4091), .ZN(n4096) );
  AOI22_X1 U4790 ( .A1(n4148), .A2(n4092), .B1(n5040), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n4093) );
  OAI21_X1 U4791 ( .B1(n4094), .B2(n4264), .A(n4093), .ZN(n4095) );
  AOI21_X1 U4792 ( .B1(n4096), .B2(n5032), .A(n4095), .ZN(n4097) );
  OAI211_X1 U4793 ( .C1(n4099), .C2(n5040), .A(n4098), .B(n4097), .ZN(U3262)
         );
  OAI21_X1 U4794 ( .B1(n4105), .B2(n4101), .A(n4100), .ZN(n4103) );
  AOI222_X1 U4795 ( .A1(n4254), .A2(n4103), .B1(n4102), .B2(n4558), .C1(n4142), 
        .C2(n4282), .ZN(n4304) );
  XOR2_X1 U4796 ( .A(n4105), .B(n4104), .Z(n4307) );
  NAND2_X1 U4797 ( .A1(n4307), .A2(n5045), .ZN(n4114) );
  INV_X1 U4798 ( .A(n4126), .ZN(n4107) );
  INV_X1 U4799 ( .A(n4381), .ZN(n4112) );
  AOI22_X1 U4800 ( .A1(n4148), .A2(n4108), .B1(n5040), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4109) );
  OAI21_X1 U4801 ( .B1(n4110), .B2(n4264), .A(n4109), .ZN(n4111) );
  AOI21_X1 U4802 ( .B1(n4112), .B2(n5032), .A(n4111), .ZN(n4113) );
  OAI211_X1 U4803 ( .C1(n4304), .C2(n5040), .A(n4114), .B(n4113), .ZN(U3263)
         );
  XNOR2_X1 U4804 ( .A(n4115), .B(n4118), .ZN(n4311) );
  INV_X1 U4805 ( .A(n4311), .ZN(n4134) );
  NAND2_X1 U4806 ( .A1(n4117), .A2(n4116), .ZN(n4119) );
  XNOR2_X1 U4807 ( .A(n4119), .B(n4118), .ZN(n4120) );
  NAND2_X1 U4808 ( .A1(n4120), .A2(n4254), .ZN(n4124) );
  AOI22_X1 U4809 ( .A1(n4122), .A2(n4282), .B1(n4121), .B2(n4298), .ZN(n4123)
         );
  OAI211_X1 U4810 ( .C1(n4125), .C2(n4274), .A(n4124), .B(n4123), .ZN(n4310)
         );
  INV_X1 U4811 ( .A(n4145), .ZN(n4128) );
  OAI21_X1 U4812 ( .B1(n4128), .B2(n4127), .A(n4126), .ZN(n4385) );
  INV_X1 U4813 ( .A(n4129), .ZN(n4130) );
  AOI22_X1 U4814 ( .A1(n4130), .A2(n5034), .B1(REG2_REG_26__SCAN_IN), .B2(
        n5040), .ZN(n4131) );
  OAI21_X1 U4815 ( .B1(n4385), .B2(n4263), .A(n4131), .ZN(n4132) );
  AOI21_X1 U4816 ( .B1(n4310), .B2(n4290), .A(n4132), .ZN(n4133) );
  OAI21_X1 U4817 ( .B1(n4134), .B2(n4293), .A(n4133), .ZN(U3264) );
  XOR2_X1 U4818 ( .A(n4137), .B(n4136), .Z(n4316) );
  INV_X1 U4819 ( .A(n4316), .ZN(n4153) );
  INV_X1 U4820 ( .A(n4137), .ZN(n4138) );
  XNOR2_X1 U4821 ( .A(n4139), .B(n4138), .ZN(n4140) );
  NAND2_X1 U4822 ( .A1(n4140), .A2(n4254), .ZN(n4144) );
  AOI22_X1 U4823 ( .A1(n4142), .A2(n4558), .B1(n4282), .B2(n4141), .ZN(n4143)
         );
  NAND2_X1 U4824 ( .A1(n4144), .A2(n4143), .ZN(n4314) );
  OAI21_X1 U4825 ( .B1(n4164), .B2(n4313), .A(n4145), .ZN(n4389) );
  AOI22_X1 U4826 ( .A1(n4146), .A2(n5034), .B1(REG2_REG_25__SCAN_IN), .B2(
        n5040), .ZN(n4150) );
  NAND2_X1 U4827 ( .A1(n4148), .A2(n4147), .ZN(n4149) );
  OAI211_X1 U4828 ( .C1(n4389), .C2(n4263), .A(n4150), .B(n4149), .ZN(n4151)
         );
  AOI21_X1 U4829 ( .B1(n4314), .B2(n4290), .A(n4151), .ZN(n4152) );
  OAI21_X1 U4830 ( .B1(n4153), .B2(n4293), .A(n4152), .ZN(U3265) );
  XOR2_X1 U4831 ( .A(n4158), .B(n4154), .Z(n4320) );
  INV_X1 U4832 ( .A(n4320), .ZN(n4171) );
  NAND2_X1 U4833 ( .A1(n4156), .A2(n4155), .ZN(n4157) );
  XOR2_X1 U4834 ( .A(n4158), .B(n4157), .Z(n4159) );
  NAND2_X1 U4835 ( .A1(n4159), .A2(n4254), .ZN(n4162) );
  AOI22_X1 U4836 ( .A1(n4194), .A2(n4282), .B1(n4160), .B2(n4298), .ZN(n4161)
         );
  OAI211_X1 U4837 ( .C1(n4163), .C2(n4274), .A(n4162), .B(n4161), .ZN(n4319)
         );
  INV_X1 U4838 ( .A(n4164), .ZN(n4165) );
  OAI21_X1 U4839 ( .B1(n4184), .B2(n4166), .A(n4165), .ZN(n4393) );
  AOI22_X1 U4840 ( .A1(n4167), .A2(n5034), .B1(REG2_REG_24__SCAN_IN), .B2(
        n5040), .ZN(n4168) );
  OAI21_X1 U4841 ( .B1(n4393), .B2(n4263), .A(n4168), .ZN(n4169) );
  AOI21_X1 U4842 ( .B1(n4319), .B2(n4290), .A(n4169), .ZN(n4170) );
  OAI21_X1 U4843 ( .B1(n4171), .B2(n4293), .A(n4170), .ZN(U3266) );
  XNOR2_X1 U4844 ( .A(n4172), .B(n4178), .ZN(n4324) );
  INV_X1 U4845 ( .A(n4324), .ZN(n4191) );
  NAND2_X1 U4846 ( .A1(n4174), .A2(n4173), .ZN(n4211) );
  NAND2_X1 U4847 ( .A1(n4211), .A2(n4212), .ZN(n4210) );
  NAND2_X1 U4848 ( .A1(n4210), .A2(n4175), .ZN(n4193) );
  NAND2_X1 U4849 ( .A1(n4193), .A2(n2729), .ZN(n4192) );
  NAND2_X1 U4850 ( .A1(n4192), .A2(n4176), .ZN(n4177) );
  XOR2_X1 U4851 ( .A(n4178), .B(n4177), .Z(n4179) );
  NAND2_X1 U4852 ( .A1(n4179), .A2(n4254), .ZN(n4182) );
  AOI22_X1 U4853 ( .A1(n4214), .A2(n4282), .B1(n4298), .B2(n4180), .ZN(n4181)
         );
  OAI211_X1 U4854 ( .C1(n4183), .C2(n4274), .A(n4182), .B(n4181), .ZN(n4323)
         );
  INV_X1 U4855 ( .A(n4184), .ZN(n4185) );
  OAI21_X1 U4856 ( .B1(n2272), .B2(n4186), .A(n4185), .ZN(n4397) );
  AOI22_X1 U4857 ( .A1(n4187), .A2(n5034), .B1(REG2_REG_23__SCAN_IN), .B2(
        n5040), .ZN(n4188) );
  OAI21_X1 U4858 ( .B1(n4397), .B2(n4263), .A(n4188), .ZN(n4189) );
  AOI21_X1 U4859 ( .B1(n4323), .B2(n4290), .A(n4189), .ZN(n4190) );
  OAI21_X1 U4860 ( .B1(n4191), .B2(n4293), .A(n4190), .ZN(U3267) );
  OAI21_X1 U4861 ( .B1(n2729), .B2(n4193), .A(n4192), .ZN(n4199) );
  NAND2_X1 U4862 ( .A1(n4194), .A2(n4558), .ZN(n4196) );
  NAND2_X1 U4863 ( .A1(n4236), .A2(n4282), .ZN(n4195) );
  OAI211_X1 U4864 ( .C1(n4552), .C2(n4197), .A(n4196), .B(n4195), .ZN(n4198)
         );
  AOI21_X1 U4865 ( .B1(n4199), .B2(n4254), .A(n4198), .ZN(n4330) );
  INV_X1 U4866 ( .A(n4328), .ZN(n4202) );
  OR2_X1 U4867 ( .A1(n4201), .A2(n4200), .ZN(n4327) );
  NAND3_X1 U4868 ( .A1(n4202), .A2(n5045), .A3(n4327), .ZN(n4209) );
  AOI21_X1 U4869 ( .B1(n4203), .B2(n4218), .A(n2272), .ZN(n4398) );
  INV_X1 U4870 ( .A(n4204), .ZN(n4206) );
  INV_X1 U4871 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4205) );
  OAI22_X1 U4872 ( .A1(n4206), .A2(n4264), .B1(n4205), .B2(n4290), .ZN(n4207)
         );
  AOI21_X1 U4873 ( .B1(n4398), .B2(n5032), .A(n4207), .ZN(n4208) );
  OAI211_X1 U4874 ( .C1(n5040), .C2(n4330), .A(n4209), .B(n4208), .ZN(U3268)
         );
  OAI21_X1 U4875 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4215) );
  AOI222_X1 U4876 ( .A1(n4254), .A2(n4215), .B1(n4214), .B2(n4558), .C1(n4213), 
        .C2(n4282), .ZN(n4334) );
  XNOR2_X1 U4877 ( .A(n4217), .B(n4216), .ZN(n4337) );
  NAND2_X1 U4878 ( .A1(n4337), .A2(n5045), .ZN(n4225) );
  INV_X1 U4879 ( .A(n4341), .ZN(n4219) );
  OAI21_X1 U4880 ( .B1(n4219), .B2(n4335), .A(n4218), .ZN(n4407) );
  INV_X1 U4881 ( .A(n4407), .ZN(n4223) );
  AOI22_X1 U4882 ( .A1(n4220), .A2(n5034), .B1(n5040), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n4221) );
  OAI21_X1 U4883 ( .B1(n4335), .B2(n5039), .A(n4221), .ZN(n4222) );
  AOI21_X1 U4884 ( .B1(n4223), .B2(n5032), .A(n4222), .ZN(n4224) );
  OAI211_X1 U4885 ( .C1(n5040), .C2(n4334), .A(n4225), .B(n4224), .ZN(U3269)
         );
  XNOR2_X1 U4886 ( .A(n4226), .B(n4234), .ZN(n4340) );
  INV_X1 U4887 ( .A(n4227), .ZN(n4229) );
  OAI21_X1 U4888 ( .B1(n4230), .B2(n4229), .A(n4228), .ZN(n4277) );
  AOI21_X1 U4889 ( .B1(n4277), .B2(n4232), .A(n4231), .ZN(n4233) );
  XOR2_X1 U4890 ( .A(n4234), .B(n4233), .Z(n4239) );
  AOI22_X1 U4891 ( .A1(n4235), .A2(n4282), .B1(n4242), .B2(n4298), .ZN(n4238)
         );
  NAND2_X1 U4892 ( .A1(n4236), .A2(n4558), .ZN(n4237) );
  OAI211_X1 U4893 ( .C1(n4239), .C2(n4560), .A(n4238), .B(n4237), .ZN(n4240)
         );
  AOI21_X1 U4894 ( .B1(n4340), .B2(n4563), .A(n4240), .ZN(n4344) );
  INV_X1 U4895 ( .A(n4241), .ZN(n4261) );
  NAND2_X1 U4896 ( .A1(n4261), .A2(n4242), .ZN(n4342) );
  AND3_X1 U4897 ( .A1(n4342), .A2(n5032), .A3(n4341), .ZN(n4246) );
  INV_X1 U4898 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4243) );
  OAI22_X1 U4899 ( .A1(n4244), .A2(n4264), .B1(n4290), .B2(n4243), .ZN(n4245)
         );
  AOI211_X1 U4900 ( .C1(n4340), .C2(n4573), .A(n4246), .B(n4245), .ZN(n4247)
         );
  OAI21_X1 U4901 ( .B1(n4344), .B2(n5040), .A(n4247), .ZN(U3270) );
  XNOR2_X1 U4902 ( .A(n4248), .B(n4252), .ZN(n4348) );
  INV_X1 U4903 ( .A(n4348), .ZN(n4269) );
  INV_X1 U4904 ( .A(n4249), .ZN(n4251) );
  OAI21_X1 U4905 ( .B1(n4277), .B2(n4251), .A(n4250), .ZN(n4253) );
  XNOR2_X1 U4906 ( .A(n4253), .B(n4252), .ZN(n4255) );
  NAND2_X1 U4907 ( .A1(n4255), .A2(n4254), .ZN(n4259) );
  AOI22_X1 U4908 ( .A1(n4257), .A2(n4282), .B1(n4298), .B2(n4256), .ZN(n4258)
         );
  OAI211_X1 U4909 ( .C1(n4260), .C2(n4274), .A(n4259), .B(n4258), .ZN(n4347)
         );
  OAI21_X1 U4910 ( .B1(n2370), .B2(n4262), .A(n4261), .ZN(n4412) );
  NOR2_X1 U4911 ( .A1(n4412), .A2(n4263), .ZN(n4267) );
  OAI22_X1 U4912 ( .A1(n4290), .A2(n4065), .B1(n4265), .B2(n4264), .ZN(n4266)
         );
  AOI211_X1 U4913 ( .C1(n4347), .C2(n4290), .A(n4267), .B(n4266), .ZN(n4268)
         );
  OAI21_X1 U4914 ( .B1(n4269), .B2(n4293), .A(n4268), .ZN(U3271) );
  INV_X1 U4915 ( .A(n4270), .ZN(n4271) );
  AOI21_X1 U4916 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(n4352) );
  OAI22_X1 U4917 ( .A1(n4275), .A2(n4274), .B1(n4285), .B2(n4552), .ZN(n4280)
         );
  XNOR2_X1 U4918 ( .A(n4277), .B(n4276), .ZN(n4278) );
  NOR2_X1 U4919 ( .A1(n4278), .A2(n4560), .ZN(n4279) );
  AOI211_X1 U4920 ( .C1(n4282), .C2(n4281), .A(n4280), .B(n4279), .ZN(n4351)
         );
  INV_X1 U4921 ( .A(n4351), .ZN(n4291) );
  OAI211_X1 U4922 ( .C1(n2366), .C2(n4285), .A(n4638), .B(n4284), .ZN(n4350)
         );
  AOI22_X1 U4923 ( .A1(n5040), .A2(REG2_REG_18__SCAN_IN), .B1(n4286), .B2(
        n5034), .ZN(n4287) );
  OAI21_X1 U4924 ( .B1(n4350), .B2(n4288), .A(n4287), .ZN(n4289) );
  AOI21_X1 U4925 ( .B1(n4291), .B2(n4290), .A(n4289), .ZN(n4292) );
  OAI21_X1 U4926 ( .B1(n4352), .B2(n4293), .A(n4292), .ZN(U3272) );
  NAND2_X1 U4927 ( .A1(n4373), .A2(n4659), .ZN(n4295) );
  NAND2_X1 U4928 ( .A1(n4657), .A2(REG1_REG_31__SCAN_IN), .ZN(n4294) );
  OAI211_X1 U4929 ( .C1(n4375), .C2(n4358), .A(n4295), .B(n4294), .ZN(U3549)
         );
  AOI21_X1 U4930 ( .B1(n4299), .B2(n4297), .A(n4296), .ZN(n4449) );
  INV_X1 U4931 ( .A(n4449), .ZN(n4377) );
  NAND2_X1 U4932 ( .A1(n4299), .A2(n4298), .ZN(n4300) );
  AND2_X1 U4933 ( .A1(n4301), .A2(n4300), .ZN(n4451) );
  INV_X1 U4934 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U4935 ( .A(n4451), .B(n4302), .S(n4657), .Z(n4303) );
  OAI21_X1 U4936 ( .B1(n4377), .B2(n4358), .A(n4303), .ZN(U3548) );
  INV_X1 U4937 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4308) );
  OAI21_X1 U4938 ( .B1(n4305), .B2(n4552), .A(n4304), .ZN(n4306) );
  AOI21_X1 U4939 ( .B1(n4307), .B2(n4619), .A(n4306), .ZN(n4378) );
  MUX2_X1 U4940 ( .A(n4308), .B(n4378), .S(n4346), .Z(n4309) );
  OAI21_X1 U4941 ( .B1(n4358), .B2(n4381), .A(n4309), .ZN(U3545) );
  INV_X1 U4942 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4799) );
  AOI21_X1 U4943 ( .B1(n4311), .B2(n4619), .A(n4310), .ZN(n4382) );
  MUX2_X1 U4944 ( .A(n4799), .B(n4382), .S(n4659), .Z(n4312) );
  OAI21_X1 U4945 ( .B1(n4358), .B2(n4385), .A(n4312), .ZN(U3544) );
  INV_X1 U4946 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4317) );
  NOR2_X1 U4947 ( .A1(n4313), .A2(n4552), .ZN(n4315) );
  AOI211_X1 U4948 ( .C1(n4316), .C2(n4619), .A(n4315), .B(n4314), .ZN(n4386)
         );
  MUX2_X1 U4949 ( .A(n4317), .B(n4386), .S(n4346), .Z(n4318) );
  OAI21_X1 U4950 ( .B1(n4358), .B2(n4389), .A(n4318), .ZN(U3543) );
  INV_X1 U4951 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4321) );
  AOI21_X1 U4952 ( .B1(n4320), .B2(n4619), .A(n4319), .ZN(n4390) );
  MUX2_X1 U4953 ( .A(n4321), .B(n4390), .S(n4346), .Z(n4322) );
  OAI21_X1 U4954 ( .B1(n4358), .B2(n4393), .A(n4322), .ZN(U3542) );
  INV_X1 U4955 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4325) );
  AOI21_X1 U4956 ( .B1(n4324), .B2(n4619), .A(n4323), .ZN(n4394) );
  MUX2_X1 U4957 ( .A(n4325), .B(n4394), .S(n4346), .Z(n4326) );
  OAI21_X1 U4958 ( .B1(n4358), .B2(n4397), .A(n4326), .ZN(U3541) );
  NAND2_X1 U4959 ( .A1(n4327), .A2(n4619), .ZN(n4329) );
  OR2_X1 U4960 ( .A1(n4329), .A2(n4328), .ZN(n4331) );
  NAND2_X1 U4961 ( .A1(n4331), .A2(n4330), .ZN(n4399) );
  MUX2_X1 U4962 ( .A(REG1_REG_22__SCAN_IN), .B(n4399), .S(n4659), .Z(n4332) );
  AOI21_X1 U4963 ( .B1(n2879), .B2(n4398), .A(n4332), .ZN(n4333) );
  INV_X1 U4964 ( .A(n4333), .ZN(U3540) );
  INV_X1 U4965 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4338) );
  OAI21_X1 U4966 ( .B1(n4335), .B2(n4552), .A(n4334), .ZN(n4336) );
  AOI21_X1 U4967 ( .B1(n4337), .B2(n4619), .A(n4336), .ZN(n4404) );
  MUX2_X1 U4968 ( .A(n4338), .B(n4404), .S(n4346), .Z(n4339) );
  OAI21_X1 U4969 ( .B1(n4358), .B2(n4407), .A(n4339), .ZN(U3539) );
  INV_X1 U4970 ( .A(n4340), .ZN(n4345) );
  NAND3_X1 U4971 ( .A1(n4342), .A2(n4638), .A3(n4341), .ZN(n4343) );
  OAI211_X1 U4972 ( .C1(n4345), .C2(n4606), .A(n4344), .B(n4343), .ZN(n4408)
         );
  MUX2_X1 U4973 ( .A(REG1_REG_20__SCAN_IN), .B(n4408), .S(n4346), .Z(U3538) );
  AOI21_X1 U4974 ( .B1(n4348), .B2(n4619), .A(n4347), .ZN(n4410) );
  MUX2_X1 U4975 ( .A(n4410), .B(n4060), .S(n4657), .Z(n4349) );
  OAI21_X1 U4976 ( .B1(n4358), .B2(n4412), .A(n4349), .ZN(U3537) );
  INV_X1 U4977 ( .A(n4619), .ZN(n4363) );
  OAI211_X1 U4978 ( .C1(n4352), .C2(n4363), .A(n4351), .B(n4350), .ZN(n4413)
         );
  MUX2_X1 U4979 ( .A(REG1_REG_18__SCAN_IN), .B(n4413), .S(n4659), .Z(U3536) );
  OAI21_X1 U4980 ( .B1(n4354), .B2(n4552), .A(n4353), .ZN(n4355) );
  AOI21_X1 U4981 ( .B1(n4356), .B2(n4619), .A(n4355), .ZN(n4414) );
  MUX2_X1 U4982 ( .A(n4036), .B(n4414), .S(n4659), .Z(n4357) );
  OAI21_X1 U4983 ( .B1(n4358), .B2(n4418), .A(n4357), .ZN(U3535) );
  OR3_X1 U4984 ( .A1(n4360), .A2(n4359), .A3(n4631), .ZN(n4361) );
  OAI211_X1 U4985 ( .C1(n4364), .C2(n4363), .A(n4362), .B(n4361), .ZN(n4419)
         );
  MUX2_X1 U4986 ( .A(REG1_REG_16__SCAN_IN), .B(n4419), .S(n4659), .Z(U3534) );
  INV_X1 U4987 ( .A(n4365), .ZN(n4370) );
  NAND3_X1 U4988 ( .A1(n4367), .A2(n4638), .A3(n4366), .ZN(n4368) );
  OAI211_X1 U4989 ( .C1(n4370), .C2(n4606), .A(n4369), .B(n4368), .ZN(n4420)
         );
  MUX2_X1 U4990 ( .A(REG1_REG_14__SCAN_IN), .B(n4420), .S(n4659), .Z(U3532) );
  NOR2_X1 U4991 ( .A1(n4645), .A2(n4371), .ZN(n4372) );
  AOI21_X1 U4992 ( .B1(n4645), .B2(n4373), .A(n4372), .ZN(n4374) );
  OAI21_X1 U4993 ( .B1(n4375), .B2(n4417), .A(n4374), .ZN(U3517) );
  MUX2_X1 U4994 ( .A(n4451), .B(n2869), .S(n4643), .Z(n4376) );
  OAI21_X1 U4995 ( .B1(n4377), .B2(n4417), .A(n4376), .ZN(U3516) );
  MUX2_X1 U4996 ( .A(n4379), .B(n4378), .S(n4645), .Z(n4380) );
  OAI21_X1 U4997 ( .B1(n4381), .B2(n4417), .A(n4380), .ZN(U3513) );
  MUX2_X1 U4998 ( .A(n4383), .B(n4382), .S(n4645), .Z(n4384) );
  OAI21_X1 U4999 ( .B1(n4385), .B2(n4417), .A(n4384), .ZN(U3512) );
  MUX2_X1 U5000 ( .A(n4387), .B(n4386), .S(n4645), .Z(n4388) );
  OAI21_X1 U5001 ( .B1(n4389), .B2(n4417), .A(n4388), .ZN(U3511) );
  MUX2_X1 U5002 ( .A(n4391), .B(n4390), .S(n4645), .Z(n4392) );
  OAI21_X1 U5003 ( .B1(n4393), .B2(n4417), .A(n4392), .ZN(U3510) );
  MUX2_X1 U5004 ( .A(n4395), .B(n4394), .S(n4645), .Z(n4396) );
  OAI21_X1 U5005 ( .B1(n4397), .B2(n4417), .A(n4396), .ZN(U3509) );
  INV_X1 U5006 ( .A(n4398), .ZN(n4403) );
  INV_X1 U5007 ( .A(n4399), .ZN(n4400) );
  MUX2_X1 U5008 ( .A(n4401), .B(n4400), .S(n4645), .Z(n4402) );
  OAI21_X1 U5009 ( .B1(n4403), .B2(n4417), .A(n4402), .ZN(U3508) );
  MUX2_X1 U5010 ( .A(n4405), .B(n4404), .S(n4645), .Z(n4406) );
  OAI21_X1 U5011 ( .B1(n4407), .B2(n4417), .A(n4406), .ZN(U3507) );
  MUX2_X1 U5012 ( .A(REG0_REG_20__SCAN_IN), .B(n4408), .S(n4645), .Z(U3506) );
  INV_X1 U5013 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4409) );
  MUX2_X1 U5014 ( .A(n4410), .B(n4409), .S(n4643), .Z(n4411) );
  OAI21_X1 U5015 ( .B1(n4412), .B2(n4417), .A(n4411), .ZN(U3505) );
  MUX2_X1 U5016 ( .A(REG0_REG_18__SCAN_IN), .B(n4413), .S(n4645), .Z(U3503) );
  INV_X1 U5017 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4415) );
  MUX2_X1 U5018 ( .A(n4415), .B(n4414), .S(n4645), .Z(n4416) );
  OAI21_X1 U5019 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(U3501) );
  MUX2_X1 U5020 ( .A(REG0_REG_16__SCAN_IN), .B(n4419), .S(n4645), .Z(U3499) );
  MUX2_X1 U5021 ( .A(REG0_REG_14__SCAN_IN), .B(n4420), .S(n4645), .Z(U3495) );
  MUX2_X1 U5022 ( .A(n4421), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5023 ( .A(n4422), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5024 ( .A(n4423), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5025 ( .A(DATAI_20_), .B(n4424), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5026 ( .A(DATAI_19_), .B(n4425), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5027 ( .A(n4426), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5028 ( .A(n4427), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5029 ( .A(n4428), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5030 ( .A(n4429), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5031 ( .A(DATAI_4_), .B(n4430), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5032 ( .A(n4431), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5033 ( .A(n4432), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5034 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5035 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4749) );
  NOR2_X1 U5036 ( .A1(STATE_REG_SCAN_IN), .A2(n4749), .ZN(n4530) );
  OAI22_X1 U5037 ( .A1(n4436), .A2(n4435), .B1(n4434), .B2(n4433), .ZN(n4437)
         );
  AOI211_X1 U5038 ( .C1(n4439), .C2(n4438), .A(n4530), .B(n4437), .ZN(n4446)
         );
  AOI21_X1 U5039 ( .B1(n4440), .B2(n3819), .A(n3818), .ZN(n4441) );
  XOR2_X1 U5040 ( .A(n4442), .B(n4441), .Z(n4444) );
  NAND2_X1 U5041 ( .A1(n4444), .A2(n4443), .ZN(n4445) );
  OAI211_X1 U5042 ( .C1(n4448), .C2(n4447), .A(n4446), .B(n4445), .ZN(U3223)
         );
  AOI22_X1 U5043 ( .A1(n4449), .A2(n5032), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5040), .ZN(n4450) );
  OAI21_X1 U5044 ( .B1(n5040), .B2(n4451), .A(n4450), .ZN(U3261) );
  AOI22_X1 U5045 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4598), .B1(n4452), .B2(n4653), .ZN(n4454) );
  OAI21_X1 U5046 ( .B1(n4455), .B2(n4454), .A(n4542), .ZN(n4453) );
  AOI21_X1 U5047 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(n4456) );
  AOI211_X1 U5048 ( .C1(n4541), .C2(ADDR_REG_7__SCAN_IN), .A(n4457), .B(n4456), 
        .ZN(n4462) );
  OAI211_X1 U5049 ( .C1(n4460), .C2(n4459), .A(n4507), .B(n4458), .ZN(n4461)
         );
  OAI211_X1 U5050 ( .C1(n4548), .C2(n4598), .A(n4462), .B(n4461), .ZN(U3247)
         );
  OAI211_X1 U5051 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4464), .A(n4507), .B(n4463), 
        .ZN(n4466) );
  NAND2_X1 U5052 ( .A1(n4466), .A2(n4465), .ZN(n4467) );
  AOI21_X1 U5053 ( .B1(n4541), .B2(ADDR_REG_8__SCAN_IN), .A(n4467), .ZN(n4471)
         );
  OAI211_X1 U5054 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4469), .A(n4542), .B(n4468), 
        .ZN(n4470) );
  OAI211_X1 U5055 ( .C1(n4548), .C2(n4472), .A(n4471), .B(n4470), .ZN(U3248)
         );
  INV_X1 U5056 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4809) );
  OAI211_X1 U5057 ( .C1(n4475), .C2(n4474), .A(n4507), .B(n4473), .ZN(n4476)
         );
  OAI21_X1 U5058 ( .B1(n4477), .B2(n4809), .A(n4476), .ZN(n4478) );
  NOR2_X1 U5059 ( .A1(n4479), .A2(n4478), .ZN(n4484) );
  OAI211_X1 U5060 ( .C1(n4482), .C2(n4481), .A(n4542), .B(n4480), .ZN(n4483)
         );
  OAI211_X1 U5061 ( .C1(n4548), .C2(n4595), .A(n4484), .B(n4483), .ZN(U3249)
         );
  OAI211_X1 U5062 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4486), .A(n4542), .B(n4485), .ZN(n4490) );
  OAI211_X1 U5063 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4488), .A(n4507), .B(n4487), .ZN(n4489) );
  OAI211_X1 U5064 ( .C1(n4548), .C2(n4491), .A(n4490), .B(n4489), .ZN(n4492)
         );
  AOI211_X1 U5065 ( .C1(n4541), .C2(ADDR_REG_10__SCAN_IN), .A(n4493), .B(n4492), .ZN(n4494) );
  INV_X1 U5066 ( .A(n4494), .ZN(U3250) );
  OAI211_X1 U5067 ( .C1(n4497), .C2(n4496), .A(n4507), .B(n4495), .ZN(n4498)
         );
  NAND2_X1 U5068 ( .A1(n4499), .A2(n4498), .ZN(n4500) );
  AOI21_X1 U5069 ( .B1(n4541), .B2(ADDR_REG_11__SCAN_IN), .A(n4500), .ZN(n4505) );
  OAI211_X1 U5070 ( .C1(n4503), .C2(n4502), .A(n4542), .B(n4501), .ZN(n4504)
         );
  OAI211_X1 U5071 ( .C1(n4548), .C2(n4591), .A(n4505), .B(n4504), .ZN(U3251)
         );
  OAI211_X1 U5072 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4508), .A(n4507), .B(n4506), .ZN(n4510) );
  NAND2_X1 U5073 ( .A1(n4510), .A2(n4509), .ZN(n4511) );
  AOI21_X1 U5074 ( .B1(n4541), .B2(ADDR_REG_12__SCAN_IN), .A(n4511), .ZN(n4515) );
  OAI211_X1 U5075 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4513), .A(n4542), .B(n4512), .ZN(n4514) );
  OAI211_X1 U5076 ( .C1(n4548), .C2(n4516), .A(n4515), .B(n4514), .ZN(U3252)
         );
  AOI211_X1 U5077 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4535), .ZN(n4520)
         );
  AOI211_X1 U5078 ( .C1(n4541), .C2(ADDR_REG_15__SCAN_IN), .A(n4521), .B(n4520), .ZN(n4526) );
  OAI211_X1 U5079 ( .C1(n4524), .C2(n4523), .A(n4542), .B(n4522), .ZN(n4525)
         );
  OAI211_X1 U5080 ( .C1(n4548), .C2(n4587), .A(n4526), .B(n4525), .ZN(U3255)
         );
  AOI221_X1 U5081 ( .B1(n4528), .B2(n4527), .C1(n3531), .C2(n4527), .A(n4535), 
        .ZN(n4529) );
  AOI211_X1 U5082 ( .C1(n4541), .C2(ADDR_REG_16__SCAN_IN), .A(n4530), .B(n4529), .ZN(n4534) );
  OAI221_X1 U5083 ( .B1(n4532), .B2(REG1_REG_16__SCAN_IN), .C1(n4532), .C2(
        n4531), .A(n4542), .ZN(n4533) );
  OAI211_X1 U5084 ( .C1(n4548), .C2(n4586), .A(n4534), .B(n4533), .ZN(U3256)
         );
  AOI221_X1 U5085 ( .B1(n4538), .B2(n4537), .C1(n4536), .C2(n4537), .A(n4535), 
        .ZN(n4539) );
  AOI211_X1 U5086 ( .C1(n4541), .C2(ADDR_REG_17__SCAN_IN), .A(n4540), .B(n4539), .ZN(n4547) );
  OAI221_X1 U5087 ( .B1(n4545), .B2(n4544), .C1(n4545), .C2(n4543), .A(n4542), 
        .ZN(n4546) );
  OAI211_X1 U5088 ( .C1(n4548), .C2(n4584), .A(n4547), .B(n4546), .ZN(U3257)
         );
  XNOR2_X1 U5089 ( .A(n4549), .B(n4550), .ZN(n4640) );
  XNOR2_X1 U5090 ( .A(n4551), .B(n4550), .ZN(n4561) );
  OAI22_X1 U5091 ( .A1(n4555), .A2(n4554), .B1(n4553), .B2(n4552), .ZN(n4556)
         );
  AOI21_X1 U5092 ( .B1(n4558), .B2(n4557), .A(n4556), .ZN(n4559) );
  OAI21_X1 U5093 ( .B1(n4561), .B2(n4560), .A(n4559), .ZN(n4562) );
  AOI21_X1 U5094 ( .B1(n4563), .B2(n4640), .A(n4562), .ZN(n4642) );
  AOI22_X1 U5095 ( .A1(n4564), .A2(n5034), .B1(REG2_REG_11__SCAN_IN), .B2(
        n5040), .ZN(n4569) );
  AOI21_X1 U5096 ( .B1(n4567), .B2(n4566), .A(n4565), .ZN(n4637) );
  AOI22_X1 U5097 ( .A1(n4640), .A2(n4573), .B1(n5032), .B2(n4637), .ZN(n4568)
         );
  OAI211_X1 U5098 ( .C1(n5040), .C2(n4642), .A(n4569), .B(n4568), .ZN(U3279)
         );
  AOI22_X1 U5099 ( .A1(n5040), .A2(REG2_REG_3__SCAN_IN), .B1(n5034), .B2(n2532), .ZN(n4576) );
  INV_X1 U5100 ( .A(n4570), .ZN(n4574) );
  INV_X1 U5101 ( .A(n4571), .ZN(n4572) );
  AOI22_X1 U5102 ( .A1(n4574), .A2(n4573), .B1(n5032), .B2(n4572), .ZN(n4575)
         );
  OAI211_X1 U5103 ( .C1(n5040), .C2(n4577), .A(n4576), .B(n4575), .ZN(U3287)
         );
  AND2_X1 U5104 ( .A1(D_REG_31__SCAN_IN), .A2(n4582), .ZN(U3291) );
  AND2_X1 U5105 ( .A1(D_REG_30__SCAN_IN), .A2(n4582), .ZN(U3292) );
  AND2_X1 U5106 ( .A1(D_REG_29__SCAN_IN), .A2(n4582), .ZN(U3293) );
  AND2_X1 U5107 ( .A1(D_REG_28__SCAN_IN), .A2(n4582), .ZN(U3294) );
  NOR2_X1 U5108 ( .A1(n4581), .A2(n4769), .ZN(U3295) );
  NOR2_X1 U5109 ( .A1(n4581), .A2(n4579), .ZN(U3296) );
  AND2_X1 U5110 ( .A1(D_REG_25__SCAN_IN), .A2(n4582), .ZN(U3297) );
  INV_X1 U5111 ( .A(D_REG_24__SCAN_IN), .ZN(n4881) );
  NOR2_X1 U5112 ( .A1(n4581), .A2(n4881), .ZN(U3298) );
  AND2_X1 U5113 ( .A1(D_REG_23__SCAN_IN), .A2(n4582), .ZN(U3299) );
  AND2_X1 U5114 ( .A1(D_REG_22__SCAN_IN), .A2(n4582), .ZN(U3300) );
  INV_X1 U5115 ( .A(D_REG_21__SCAN_IN), .ZN(n4872) );
  NOR2_X1 U5116 ( .A1(n4581), .A2(n4872), .ZN(U3301) );
  AND2_X1 U5117 ( .A1(n4582), .A2(D_REG_20__SCAN_IN), .ZN(U3302) );
  AND2_X1 U5118 ( .A1(D_REG_19__SCAN_IN), .A2(n4582), .ZN(U3303) );
  AND2_X1 U5119 ( .A1(D_REG_18__SCAN_IN), .A2(n4582), .ZN(U3304) );
  NOR2_X1 U5120 ( .A1(n4581), .A2(n4580), .ZN(U3305) );
  AND2_X1 U5121 ( .A1(D_REG_16__SCAN_IN), .A2(n4582), .ZN(U3306) );
  INV_X1 U5122 ( .A(D_REG_15__SCAN_IN), .ZN(n4857) );
  NOR2_X1 U5123 ( .A1(n4581), .A2(n4857), .ZN(U3307) );
  INV_X1 U5124 ( .A(D_REG_14__SCAN_IN), .ZN(n4867) );
  NOR2_X1 U5125 ( .A1(n4581), .A2(n4867), .ZN(U3308) );
  NOR2_X1 U5126 ( .A1(n4581), .A2(n4773), .ZN(U3309) );
  AND2_X1 U5127 ( .A1(D_REG_12__SCAN_IN), .A2(n4582), .ZN(U3310) );
  AND2_X1 U5128 ( .A1(D_REG_11__SCAN_IN), .A2(n4582), .ZN(U3311) );
  AND2_X1 U5129 ( .A1(D_REG_10__SCAN_IN), .A2(n4582), .ZN(U3312) );
  INV_X1 U5130 ( .A(D_REG_9__SCAN_IN), .ZN(n4887) );
  NOR2_X1 U5131 ( .A1(n4581), .A2(n4887), .ZN(U3313) );
  AND2_X1 U5132 ( .A1(D_REG_8__SCAN_IN), .A2(n4582), .ZN(U3314) );
  AND2_X1 U5133 ( .A1(D_REG_7__SCAN_IN), .A2(n4582), .ZN(U3315) );
  AND2_X1 U5134 ( .A1(D_REG_6__SCAN_IN), .A2(n4582), .ZN(U3316) );
  INV_X1 U5135 ( .A(D_REG_5__SCAN_IN), .ZN(n4932) );
  NOR2_X1 U5136 ( .A1(n4581), .A2(n4932), .ZN(U3317) );
  AND2_X1 U5137 ( .A1(D_REG_4__SCAN_IN), .A2(n4582), .ZN(U3318) );
  INV_X1 U5138 ( .A(D_REG_3__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U5139 ( .A1(n4581), .A2(n4941), .ZN(U3319) );
  AND2_X1 U5140 ( .A1(D_REG_2__SCAN_IN), .A2(n4582), .ZN(U3320) );
  INV_X1 U5141 ( .A(DATAI_23_), .ZN(n4738) );
  AOI21_X1 U5142 ( .B1(U3149), .B2(n4738), .A(n4583), .ZN(U3329) );
  AOI22_X1 U5143 ( .A1(STATE_REG_SCAN_IN), .A2(n4584), .B1(n2687), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5144 ( .A(DATAI_16_), .ZN(n4585) );
  AOI22_X1 U5145 ( .A1(STATE_REG_SCAN_IN), .A2(n4586), .B1(n4585), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5146 ( .A(DATAI_15_), .ZN(n4751) );
  AOI22_X1 U5147 ( .A1(STATE_REG_SCAN_IN), .A2(n4587), .B1(n4751), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5148 ( .A1(U3149), .A2(n4588), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4589) );
  INV_X1 U5149 ( .A(n4589), .ZN(U3340) );
  INV_X1 U5150 ( .A(DATAI_11_), .ZN(n4590) );
  AOI22_X1 U5151 ( .A1(STATE_REG_SCAN_IN), .A2(n4591), .B1(n4590), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5152 ( .A1(U3149), .A2(n4592), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4593) );
  INV_X1 U5153 ( .A(n4593), .ZN(U3342) );
  INV_X1 U5154 ( .A(DATAI_9_), .ZN(n4594) );
  AOI22_X1 U5155 ( .A1(STATE_REG_SCAN_IN), .A2(n4595), .B1(n4594), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U5156 ( .A1(U3149), .A2(n4596), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4597) );
  INV_X1 U5157 ( .A(n4597), .ZN(U3344) );
  INV_X1 U5158 ( .A(DATAI_7_), .ZN(n4882) );
  AOI22_X1 U5159 ( .A1(STATE_REG_SCAN_IN), .A2(n4598), .B1(n4882), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5160 ( .A(n4599), .ZN(n4600) );
  NOR2_X1 U5161 ( .A1(n4601), .A2(n4600), .ZN(n4603) );
  AOI211_X1 U5162 ( .C1(n4639), .C2(n4604), .A(n4603), .B(n4602), .ZN(n4647)
         );
  AOI22_X1 U5163 ( .A1(n4645), .A2(n4647), .B1(n2506), .B2(n4643), .ZN(U3467)
         );
  OAI22_X1 U5164 ( .A1(n4607), .A2(n4606), .B1(n4631), .B2(n4605), .ZN(n4608)
         );
  NOR2_X1 U5165 ( .A1(n4609), .A2(n4608), .ZN(n4648) );
  AOI22_X1 U5166 ( .A1(n4645), .A2(n4648), .B1(n2496), .B2(n4643), .ZN(U3469)
         );
  NOR3_X1 U5167 ( .A1(n4611), .A2(n4610), .A3(n4631), .ZN(n4613) );
  AOI211_X1 U5168 ( .C1(n4639), .C2(n4614), .A(n4613), .B(n4612), .ZN(n4650)
         );
  INV_X1 U5169 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U5170 ( .A1(n4645), .A2(n4650), .B1(n4841), .B2(n4643), .ZN(U3471)
         );
  AOI211_X1 U5171 ( .C1(n4617), .C2(n4639), .A(n4616), .B(n4615), .ZN(n4652)
         );
  INV_X1 U5172 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4618) );
  AOI22_X1 U5173 ( .A1(n4645), .A2(n4652), .B1(n4618), .B2(n4643), .ZN(U3475)
         );
  NAND2_X1 U5174 ( .A1(n4620), .A2(n4619), .ZN(n4621) );
  INV_X1 U5175 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4624) );
  AOI22_X1 U5176 ( .A1(n4645), .A2(n4654), .B1(n4624), .B2(n4643), .ZN(U3481)
         );
  NOR3_X1 U5177 ( .A1(n4626), .A2(n4625), .A3(n4631), .ZN(n4628) );
  AOI211_X1 U5178 ( .C1(n4629), .C2(n4639), .A(n4628), .B(n4627), .ZN(n4655)
         );
  INV_X1 U5179 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5180 ( .A1(n4645), .A2(n4655), .B1(n4630), .B2(n4643), .ZN(U3483)
         );
  NOR3_X1 U5181 ( .A1(n4632), .A2(n2362), .A3(n4631), .ZN(n4634) );
  AOI211_X1 U5182 ( .C1(n4635), .C2(n4639), .A(n4634), .B(n4633), .ZN(n4656)
         );
  INV_X1 U5183 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5184 ( .A1(n4645), .A2(n4656), .B1(n4636), .B2(n4643), .ZN(U3487)
         );
  AOI22_X1 U5185 ( .A1(n4640), .A2(n4639), .B1(n4638), .B2(n4637), .ZN(n4641)
         );
  AND2_X1 U5186 ( .A1(n4642), .A2(n4641), .ZN(n4658) );
  INV_X1 U5187 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U5188 ( .A1(n4645), .A2(n4658), .B1(n4644), .B2(n4643), .ZN(U3489)
         );
  AOI22_X1 U5189 ( .A1(n4659), .A2(n4647), .B1(n4646), .B2(n4657), .ZN(U3518)
         );
  AOI22_X1 U5190 ( .A1(n4659), .A2(n4648), .B1(n2926), .B2(n4657), .ZN(U3519)
         );
  AOI22_X1 U5191 ( .A1(n4659), .A2(n4650), .B1(n4649), .B2(n4657), .ZN(U3520)
         );
  INV_X1 U5192 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4651) );
  AOI22_X1 U5193 ( .A1(n4659), .A2(n4652), .B1(n4651), .B2(n4657), .ZN(U3522)
         );
  AOI22_X1 U5194 ( .A1(n4659), .A2(n4654), .B1(n4653), .B2(n4657), .ZN(U3525)
         );
  INV_X1 U5195 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5196 ( .A1(n4659), .A2(n4655), .B1(n4791), .B2(n4657), .ZN(U3526)
         );
  INV_X1 U5197 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4928) );
  AOI22_X1 U5198 ( .A1(n4659), .A2(n4656), .B1(n4928), .B2(n4657), .ZN(U3528)
         );
  AOI22_X1 U5199 ( .A1(n4659), .A2(n4658), .B1(n4797), .B2(n4657), .ZN(U3529)
         );
  AOI22_X1 U5200 ( .A1(DATAI_26_), .A2(keyinput183), .B1(DATAI_29_), .B2(
        keyinput237), .ZN(n4660) );
  OAI221_X1 U5201 ( .B1(DATAI_26_), .B2(keyinput183), .C1(DATAI_29_), .C2(
        keyinput237), .A(n4660), .ZN(n4667) );
  AOI22_X1 U5202 ( .A1(DATAI_12_), .A2(keyinput251), .B1(DATAI_19_), .B2(
        keyinput140), .ZN(n4661) );
  OAI221_X1 U5203 ( .B1(DATAI_12_), .B2(keyinput251), .C1(DATAI_19_), .C2(
        keyinput140), .A(n4661), .ZN(n4666) );
  AOI22_X1 U5204 ( .A1(DATAI_5_), .A2(keyinput173), .B1(DATAI_4_), .B2(
        keyinput252), .ZN(n4662) );
  OAI221_X1 U5205 ( .B1(DATAI_5_), .B2(keyinput173), .C1(DATAI_4_), .C2(
        keyinput252), .A(n4662), .ZN(n4665) );
  AOI22_X1 U5206 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput203), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput172), .ZN(n4663) );
  OAI221_X1 U5207 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput203), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput172), .A(n4663), .ZN(n4664) );
  NOR4_X1 U5208 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4695)
         );
  AOI22_X1 U5209 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput141), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput182), .ZN(n4668) );
  OAI221_X1 U5210 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput141), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput182), .A(n4668), .ZN(n4675) );
  AOI22_X1 U5211 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput202), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput226), .ZN(n4669) );
  OAI221_X1 U5212 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput202), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput226), .A(n4669), .ZN(n4674) );
  AOI22_X1 U5213 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput149), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput241), .ZN(n4670) );
  OAI221_X1 U5214 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput149), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput241), .A(n4670), .ZN(n4673) );
  AOI22_X1 U5215 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput133), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput185), .ZN(n4671) );
  OAI221_X1 U5216 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput133), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput185), .A(n4671), .ZN(n4672) );
  NOR4_X1 U5217 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4694)
         );
  AOI22_X1 U5218 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput214), .B1(
        D_REG_3__SCAN_IN), .B2(keyinput205), .ZN(n4676) );
  OAI221_X1 U5219 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput214), .C1(
        D_REG_3__SCAN_IN), .C2(keyinput205), .A(n4676), .ZN(n4683) );
  AOI22_X1 U5220 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput169), .B1(
        D_REG_15__SCAN_IN), .B2(keyinput240), .ZN(n4677) );
  OAI221_X1 U5221 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput169), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput240), .A(n4677), .ZN(n4682) );
  AOI22_X1 U5222 ( .A1(D_REG_20__SCAN_IN), .A2(keyinput225), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput162), .ZN(n4678) );
  OAI221_X1 U5223 ( .B1(D_REG_20__SCAN_IN), .B2(keyinput225), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput162), .A(n4678), .ZN(n4681) );
  AOI22_X1 U5224 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput218), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput239), .ZN(n4679) );
  OAI221_X1 U5225 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput218), .C1(
        D_REG_21__SCAN_IN), .C2(keyinput239), .A(n4679), .ZN(n4680) );
  NOR4_X1 U5226 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4693)
         );
  AOI22_X1 U5227 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput242), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput238), .ZN(n4684) );
  OAI221_X1 U5228 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput242), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput238), .A(n4684), .ZN(n4691) );
  AOI22_X1 U5229 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput188), .B1(
        REG0_REG_2__SCAN_IN), .B2(keyinput253), .ZN(n4685) );
  OAI221_X1 U5230 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput188), .C1(
        REG0_REG_2__SCAN_IN), .C2(keyinput253), .A(n4685), .ZN(n4690) );
  AOI22_X1 U5231 ( .A1(REG0_REG_9__SCAN_IN), .A2(keyinput201), .B1(
        REG0_REG_12__SCAN_IN), .B2(keyinput158), .ZN(n4686) );
  OAI221_X1 U5232 ( .B1(REG0_REG_9__SCAN_IN), .B2(keyinput201), .C1(
        REG0_REG_12__SCAN_IN), .C2(keyinput158), .A(n4686), .ZN(n4689) );
  AOI22_X1 U5233 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput199), .B1(
        REG0_REG_29__SCAN_IN), .B2(keyinput179), .ZN(n4687) );
  OAI221_X1 U5234 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput199), .C1(
        REG0_REG_29__SCAN_IN), .C2(keyinput179), .A(n4687), .ZN(n4688) );
  NOR4_X1 U5235 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4692)
         );
  NAND4_X1 U5236 ( .A1(n4695), .A2(n4694), .A3(n4693), .A4(n4692), .ZN(n4836)
         );
  AOI22_X1 U5237 ( .A1(REG0_REG_30__SCAN_IN), .A2(keyinput219), .B1(
        REG1_REG_3__SCAN_IN), .B2(keyinput167), .ZN(n4696) );
  OAI221_X1 U5238 ( .B1(REG0_REG_30__SCAN_IN), .B2(keyinput219), .C1(
        REG1_REG_3__SCAN_IN), .C2(keyinput167), .A(n4696), .ZN(n4703) );
  AOI22_X1 U5239 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput255), .B1(
        REG1_REG_10__SCAN_IN), .B2(keyinput143), .ZN(n4697) );
  OAI221_X1 U5240 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput255), .C1(
        REG1_REG_10__SCAN_IN), .C2(keyinput143), .A(n4697), .ZN(n4702) );
  AOI22_X1 U5241 ( .A1(REG1_REG_24__SCAN_IN), .A2(keyinput148), .B1(
        REG1_REG_25__SCAN_IN), .B2(keyinput157), .ZN(n4698) );
  OAI221_X1 U5242 ( .B1(REG1_REG_24__SCAN_IN), .B2(keyinput148), .C1(
        REG1_REG_25__SCAN_IN), .C2(keyinput157), .A(n4698), .ZN(n4701) );
  AOI22_X1 U5243 ( .A1(REG1_REG_30__SCAN_IN), .A2(keyinput249), .B1(
        REG2_REG_1__SCAN_IN), .B2(keyinput186), .ZN(n4699) );
  OAI221_X1 U5244 ( .B1(REG1_REG_30__SCAN_IN), .B2(keyinput249), .C1(
        REG2_REG_1__SCAN_IN), .C2(keyinput186), .A(n4699), .ZN(n4700) );
  NOR4_X1 U5245 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(n4731)
         );
  AOI22_X1 U5246 ( .A1(REG2_REG_4__SCAN_IN), .A2(keyinput216), .B1(
        REG2_REG_6__SCAN_IN), .B2(keyinput231), .ZN(n4704) );
  OAI221_X1 U5247 ( .B1(REG2_REG_4__SCAN_IN), .B2(keyinput216), .C1(
        REG2_REG_6__SCAN_IN), .C2(keyinput231), .A(n4704), .ZN(n4711) );
  AOI22_X1 U5248 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput193), .B1(
        REG2_REG_9__SCAN_IN), .B2(keyinput195), .ZN(n4705) );
  OAI221_X1 U5249 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput193), .C1(
        REG2_REG_9__SCAN_IN), .C2(keyinput195), .A(n4705), .ZN(n4710) );
  AOI22_X1 U5250 ( .A1(REG2_REG_13__SCAN_IN), .A2(keyinput180), .B1(
        REG2_REG_17__SCAN_IN), .B2(keyinput204), .ZN(n4706) );
  OAI221_X1 U5251 ( .B1(REG2_REG_13__SCAN_IN), .B2(keyinput180), .C1(
        REG2_REG_17__SCAN_IN), .C2(keyinput204), .A(n4706), .ZN(n4709) );
  AOI22_X1 U5252 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput222), .B1(
        REG2_REG_22__SCAN_IN), .B2(keyinput156), .ZN(n4707) );
  OAI221_X1 U5253 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput222), .C1(
        REG2_REG_22__SCAN_IN), .C2(keyinput156), .A(n4707), .ZN(n4708) );
  NOR4_X1 U5254 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4730)
         );
  AOI22_X1 U5255 ( .A1(ADDR_REG_13__SCAN_IN), .A2(keyinput142), .B1(
        ADDR_REG_16__SCAN_IN), .B2(keyinput165), .ZN(n4712) );
  OAI221_X1 U5256 ( .B1(ADDR_REG_13__SCAN_IN), .B2(keyinput142), .C1(
        ADDR_REG_16__SCAN_IN), .C2(keyinput165), .A(n4712), .ZN(n4719) );
  AOI22_X1 U5257 ( .A1(ADDR_REG_4__SCAN_IN), .A2(keyinput228), .B1(
        ADDR_REG_6__SCAN_IN), .B2(keyinput170), .ZN(n4713) );
  OAI221_X1 U5258 ( .B1(ADDR_REG_4__SCAN_IN), .B2(keyinput228), .C1(
        ADDR_REG_6__SCAN_IN), .C2(keyinput170), .A(n4713), .ZN(n4718) );
  AOI22_X1 U5259 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput215), .B1(
        ADDR_REG_0__SCAN_IN), .B2(keyinput184), .ZN(n4714) );
  OAI221_X1 U5260 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput215), .C1(
        ADDR_REG_0__SCAN_IN), .C2(keyinput184), .A(n4714), .ZN(n4717) );
  AOI22_X1 U5261 ( .A1(DATAO_REG_15__SCAN_IN), .A2(keyinput196), .B1(
        DATAO_REG_11__SCAN_IN), .B2(keyinput171), .ZN(n4715) );
  OAI221_X1 U5262 ( .B1(DATAO_REG_15__SCAN_IN), .B2(keyinput196), .C1(
        DATAO_REG_11__SCAN_IN), .C2(keyinput171), .A(n4715), .ZN(n4716) );
  NOR4_X1 U5263 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4729)
         );
  AOI22_X1 U5264 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput243), .B1(
        DATAO_REG_19__SCAN_IN), .B2(keyinput192), .ZN(n4720) );
  OAI221_X1 U5265 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput243), .C1(
        DATAO_REG_19__SCAN_IN), .C2(keyinput192), .A(n4720), .ZN(n4727) );
  AOI22_X1 U5266 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput175), .B1(
        DATAO_REG_30__SCAN_IN), .B2(keyinput146), .ZN(n4721) );
  OAI221_X1 U5267 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput175), .C1(
        DATAO_REG_30__SCAN_IN), .C2(keyinput146), .A(n4721), .ZN(n4726) );
  AOI22_X1 U5268 ( .A1(ADDR_REG_11__SCAN_IN), .A2(keyinput254), .B1(
        ADDR_REG_19__SCAN_IN), .B2(keyinput247), .ZN(n4722) );
  OAI221_X1 U5269 ( .B1(ADDR_REG_11__SCAN_IN), .B2(keyinput254), .C1(
        ADDR_REG_19__SCAN_IN), .C2(keyinput247), .A(n4722), .ZN(n4725) );
  AOI22_X1 U5270 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput233), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput229), .ZN(n4723) );
  OAI221_X1 U5271 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput233), .C1(
        IR_REG_30__SCAN_IN), .C2(keyinput229), .A(n4723), .ZN(n4724) );
  NOR4_X1 U5272 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4728)
         );
  NAND4_X1 U5273 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4835)
         );
  AOI22_X1 U5274 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput147), .B1(n4733), 
        .B2(keyinput236), .ZN(n4732) );
  OAI221_X1 U5275 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput147), .C1(n4733), 
        .C2(keyinput236), .A(n4732), .ZN(n4745) );
  AOI22_X1 U5276 ( .A1(n4736), .A2(keyinput159), .B1(keyinput209), .B2(n4735), 
        .ZN(n4734) );
  OAI221_X1 U5277 ( .B1(n4736), .B2(keyinput159), .C1(n4735), .C2(keyinput209), 
        .A(n4734), .ZN(n4744) );
  AOI22_X1 U5278 ( .A1(n4739), .A2(keyinput197), .B1(n4738), .B2(keyinput212), 
        .ZN(n4737) );
  OAI221_X1 U5279 ( .B1(n4739), .B2(keyinput197), .C1(n4738), .C2(keyinput212), 
        .A(n4737), .ZN(n4743) );
  INV_X1 U5280 ( .A(DATAI_21_), .ZN(n4741) );
  AOI22_X1 U5281 ( .A1(n4902), .A2(keyinput191), .B1(keyinput232), .B2(n4741), 
        .ZN(n4740) );
  OAI221_X1 U5282 ( .B1(n4902), .B2(keyinput191), .C1(n4741), .C2(keyinput232), 
        .A(n4740), .ZN(n4742) );
  NOR4_X1 U5283 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4784)
         );
  AOI22_X1 U5284 ( .A1(n2672), .A2(keyinput155), .B1(n4747), .B2(keyinput130), 
        .ZN(n4746) );
  OAI221_X1 U5285 ( .B1(n2672), .B2(keyinput155), .C1(n4747), .C2(keyinput130), 
        .A(n4746), .ZN(n4757) );
  INV_X1 U5286 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5287 ( .A1(n4915), .A2(keyinput163), .B1(keyinput137), .B2(n4749), 
        .ZN(n4748) );
  OAI221_X1 U5288 ( .B1(n4915), .B2(keyinput163), .C1(n4749), .C2(keyinput137), 
        .A(n4748), .ZN(n4756) );
  AOI22_X1 U5289 ( .A1(n4751), .A2(keyinput144), .B1(n4882), .B2(keyinput223), 
        .ZN(n4750) );
  OAI221_X1 U5290 ( .B1(n4751), .B2(keyinput144), .C1(n4882), .C2(keyinput223), 
        .A(n4750), .ZN(n4755) );
  XNOR2_X1 U5291 ( .A(DATAI_0_), .B(keyinput176), .ZN(n4753) );
  XNOR2_X1 U5292 ( .A(DATAI_3_), .B(keyinput153), .ZN(n4752) );
  NAND2_X1 U5293 ( .A1(n4753), .A2(n4752), .ZN(n4754) );
  NOR4_X1 U5294 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n4783)
         );
  XNOR2_X1 U5295 ( .A(IR_REG_3__SCAN_IN), .B(keyinput160), .ZN(n4761) );
  XNOR2_X1 U5296 ( .A(IR_REG_0__SCAN_IN), .B(keyinput174), .ZN(n4760) );
  XNOR2_X1 U5297 ( .A(IR_REG_7__SCAN_IN), .B(keyinput194), .ZN(n4759) );
  XNOR2_X1 U5298 ( .A(IR_REG_1__SCAN_IN), .B(keyinput224), .ZN(n4758) );
  NAND4_X1 U5299 ( .A1(n4761), .A2(n4760), .A3(n4759), .A4(n4758), .ZN(n4767)
         );
  XNOR2_X1 U5300 ( .A(IR_REG_11__SCAN_IN), .B(keyinput235), .ZN(n4765) );
  XNOR2_X1 U5301 ( .A(IR_REG_6__SCAN_IN), .B(keyinput227), .ZN(n4764) );
  XNOR2_X1 U5302 ( .A(IR_REG_14__SCAN_IN), .B(keyinput129), .ZN(n4763) );
  XNOR2_X1 U5303 ( .A(IR_REG_13__SCAN_IN), .B(keyinput217), .ZN(n4762) );
  NAND4_X1 U5304 ( .A1(n4765), .A2(n4764), .A3(n4763), .A4(n4762), .ZN(n4766)
         );
  NOR2_X1 U5305 ( .A1(n4767), .A2(n4766), .ZN(n4782) );
  AOI22_X1 U5306 ( .A1(n4867), .A2(keyinput230), .B1(n4769), .B2(keyinput234), 
        .ZN(n4768) );
  OAI221_X1 U5307 ( .B1(n4867), .B2(keyinput230), .C1(n4769), .C2(keyinput234), 
        .A(n4768), .ZN(n4780) );
  AOI22_X1 U5308 ( .A1(n4772), .A2(keyinput248), .B1(n4771), .B2(keyinput161), 
        .ZN(n4770) );
  OAI221_X1 U5309 ( .B1(n4772), .B2(keyinput248), .C1(n4771), .C2(keyinput161), 
        .A(n4770), .ZN(n4779) );
  XNOR2_X1 U5310 ( .A(n4773), .B(keyinput134), .ZN(n4778) );
  XNOR2_X1 U5311 ( .A(IR_REG_22__SCAN_IN), .B(keyinput154), .ZN(n4776) );
  XNOR2_X1 U5312 ( .A(IR_REG_15__SCAN_IN), .B(keyinput206), .ZN(n4775) );
  XNOR2_X1 U5313 ( .A(IR_REG_18__SCAN_IN), .B(keyinput208), .ZN(n4774) );
  NAND3_X1 U5314 ( .A1(n4776), .A2(n4775), .A3(n4774), .ZN(n4777) );
  NOR4_X1 U5315 ( .A1(n4780), .A2(n4779), .A3(n4778), .A4(n4777), .ZN(n4781)
         );
  NAND4_X1 U5316 ( .A1(n4784), .A2(n4783), .A3(n4782), .A4(n4781), .ZN(n4834)
         );
  INV_X1 U5317 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4786) );
  AOI22_X1 U5318 ( .A1(n2533), .A2(keyinput164), .B1(n4786), .B2(keyinput181), 
        .ZN(n4785) );
  OAI221_X1 U5319 ( .B1(n2533), .B2(keyinput164), .C1(n4786), .C2(keyinput181), 
        .A(n4785), .ZN(n4795) );
  INV_X1 U5320 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U5321 ( .A1(n3495), .A2(keyinput139), .B1(keyinput189), .B2(n4788), 
        .ZN(n4787) );
  OAI221_X1 U5322 ( .B1(n3495), .B2(keyinput139), .C1(n4788), .C2(keyinput189), 
        .A(n4787), .ZN(n4794) );
  AOI22_X1 U5323 ( .A1(n4415), .A2(keyinput250), .B1(n4387), .B2(keyinput168), 
        .ZN(n4789) );
  OAI221_X1 U5324 ( .B1(n4415), .B2(keyinput250), .C1(n4387), .C2(keyinput168), 
        .A(n4789), .ZN(n4793) );
  AOI22_X1 U5325 ( .A1(n4371), .A2(keyinput198), .B1(n4791), .B2(keyinput136), 
        .ZN(n4790) );
  OAI221_X1 U5326 ( .B1(n4371), .B2(keyinput198), .C1(n4791), .C2(keyinput136), 
        .A(n4790), .ZN(n4792) );
  NOR4_X1 U5327 ( .A1(n4795), .A2(n4794), .A3(n4793), .A4(n4792), .ZN(n4832)
         );
  AOI22_X1 U5328 ( .A1(n3595), .A2(keyinput131), .B1(n4797), .B2(keyinput145), 
        .ZN(n4796) );
  OAI221_X1 U5329 ( .B1(n3595), .B2(keyinput131), .C1(n4797), .C2(keyinput145), 
        .A(n4796), .ZN(n4805) );
  INV_X1 U5330 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4916) );
  AOI22_X1 U5331 ( .A1(n4916), .A2(keyinput166), .B1(n4799), .B2(keyinput187), 
        .ZN(n4798) );
  OAI221_X1 U5332 ( .B1(n4916), .B2(keyinput166), .C1(n4799), .C2(keyinput187), 
        .A(n4798), .ZN(n4804) );
  INV_X1 U5333 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U5334 ( .A1(n4852), .A2(keyinput128), .B1(n3387), .B2(keyinput246), 
        .ZN(n4800) );
  OAI221_X1 U5335 ( .B1(n4852), .B2(keyinput128), .C1(n3387), .C2(keyinput246), 
        .A(n4800), .ZN(n4803) );
  AOI22_X1 U5336 ( .A1(n3531), .A2(keyinput221), .B1(keyinput150), .B2(n4912), 
        .ZN(n4801) );
  OAI221_X1 U5337 ( .B1(n3531), .B2(keyinput221), .C1(n4912), .C2(keyinput150), 
        .A(n4801), .ZN(n4802) );
  NOR4_X1 U5338 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4831)
         );
  INV_X1 U5339 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U5340 ( .A1(n4243), .A2(keyinput200), .B1(n4884), .B2(keyinput210), 
        .ZN(n4806) );
  OAI221_X1 U5341 ( .B1(n4243), .B2(keyinput200), .C1(n4884), .C2(keyinput210), 
        .A(n4806), .ZN(n4816) );
  INV_X1 U5342 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4927) );
  INV_X1 U5343 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4855) );
  AOI22_X1 U5344 ( .A1(n4927), .A2(keyinput138), .B1(keyinput220), .B2(n4855), 
        .ZN(n4807) );
  OAI221_X1 U5345 ( .B1(n4927), .B2(keyinput138), .C1(n4855), .C2(keyinput220), 
        .A(n4807), .ZN(n4815) );
  INV_X1 U5346 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U5347 ( .A1(n4809), .A2(keyinput207), .B1(keyinput177), .B2(n4930), 
        .ZN(n4808) );
  OAI221_X1 U5348 ( .B1(n4809), .B2(keyinput207), .C1(n4930), .C2(keyinput177), 
        .A(n4808), .ZN(n4814) );
  INV_X1 U5349 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4812) );
  AOI22_X1 U5350 ( .A1(n4812), .A2(keyinput151), .B1(keyinput132), .B2(n4811), 
        .ZN(n4810) );
  OAI221_X1 U5351 ( .B1(n4812), .B2(keyinput151), .C1(n4811), .C2(keyinput132), 
        .A(n4810), .ZN(n4813) );
  NOR4_X1 U5352 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4830)
         );
  AOI22_X1 U5353 ( .A1(n4858), .A2(keyinput244), .B1(keyinput190), .B2(n4818), 
        .ZN(n4817) );
  OAI221_X1 U5354 ( .B1(n4858), .B2(keyinput244), .C1(n4818), .C2(keyinput190), 
        .A(n4817), .ZN(n4828) );
  AOI22_X1 U5355 ( .A1(n4821), .A2(keyinput213), .B1(keyinput152), .B2(n4820), 
        .ZN(n4819) );
  OAI221_X1 U5356 ( .B1(n4821), .B2(keyinput213), .C1(n4820), .C2(keyinput152), 
        .A(n4819), .ZN(n4827) );
  AOI22_X1 U5357 ( .A1(n4823), .A2(keyinput135), .B1(keyinput245), .B2(n4842), 
        .ZN(n4822) );
  OAI221_X1 U5358 ( .B1(n4823), .B2(keyinput135), .C1(n4842), .C2(keyinput245), 
        .A(n4822), .ZN(n4826) );
  AOI22_X1 U5359 ( .A1(n4900), .A2(keyinput178), .B1(n4887), .B2(keyinput211), 
        .ZN(n4824) );
  OAI221_X1 U5360 ( .B1(n4900), .B2(keyinput178), .C1(n4887), .C2(keyinput211), 
        .A(n4824), .ZN(n4825) );
  NOR4_X1 U5361 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), .ZN(n4829)
         );
  NAND4_X1 U5362 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), .ZN(n4833)
         );
  NOR4_X1 U5363 ( .A1(n4836), .A2(n4835), .A3(n4834), .A4(n4833), .ZN(n5031)
         );
  AOI22_X1 U5364 ( .A1(n4839), .A2(keyinput105), .B1(n4838), .B2(keyinput113), 
        .ZN(n4837) );
  OAI221_X1 U5365 ( .B1(n4839), .B2(keyinput105), .C1(n4838), .C2(keyinput113), 
        .A(n4837), .ZN(n4850) );
  AOI22_X1 U5366 ( .A1(n4842), .A2(keyinput117), .B1(n4841), .B2(keyinput125), 
        .ZN(n4840) );
  OAI221_X1 U5367 ( .B1(n4842), .B2(keyinput117), .C1(n4841), .C2(keyinput125), 
        .A(n4840), .ZN(n4849) );
  AOI22_X1 U5368 ( .A1(n2533), .A2(keyinput36), .B1(n2506), .B2(keyinput60), 
        .ZN(n4843) );
  OAI221_X1 U5369 ( .B1(n2533), .B2(keyinput36), .C1(n2506), .C2(keyinput60), 
        .A(n4843), .ZN(n4848) );
  INV_X1 U5370 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5371 ( .A1(n4846), .A2(keyinput76), .B1(keyinput68), .B2(n4845), 
        .ZN(n4844) );
  OAI221_X1 U5372 ( .B1(n4846), .B2(keyinput76), .C1(n4845), .C2(keyinput68), 
        .A(n4844), .ZN(n4847) );
  NOR4_X1 U5373 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4897)
         );
  INV_X1 U5374 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4853) );
  AOI22_X1 U5375 ( .A1(n4853), .A2(keyinput126), .B1(n4852), .B2(keyinput0), 
        .ZN(n4851) );
  OAI221_X1 U5376 ( .B1(n4853), .B2(keyinput126), .C1(n4852), .C2(keyinput0), 
        .A(n4851), .ZN(n4865) );
  AOI22_X1 U5377 ( .A1(n4243), .A2(keyinput72), .B1(keyinput92), .B2(n4855), 
        .ZN(n4854) );
  OAI221_X1 U5378 ( .B1(n4243), .B2(keyinput72), .C1(n4855), .C2(keyinput92), 
        .A(n4854), .ZN(n4864) );
  AOI22_X1 U5379 ( .A1(n4858), .A2(keyinput116), .B1(n4857), .B2(keyinput112), 
        .ZN(n4856) );
  OAI221_X1 U5380 ( .B1(n4858), .B2(keyinput116), .C1(n4857), .C2(keyinput112), 
        .A(n4856), .ZN(n4863) );
  INV_X1 U5381 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4859) );
  XOR2_X1 U5382 ( .A(n4859), .B(keyinput100), .Z(n4861) );
  XNOR2_X1 U5383 ( .A(IR_REG_18__SCAN_IN), .B(keyinput80), .ZN(n4860) );
  NAND2_X1 U5384 ( .A1(n4861), .A2(n4860), .ZN(n4862) );
  NOR4_X1 U5385 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), .ZN(n4896)
         );
  AOI22_X1 U5386 ( .A1(n4868), .A2(keyinput107), .B1(keyinput102), .B2(n4867), 
        .ZN(n4866) );
  OAI221_X1 U5387 ( .B1(n4868), .B2(keyinput107), .C1(n4867), .C2(keyinput102), 
        .A(n4866), .ZN(n4879) );
  INV_X1 U5388 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U5389 ( .A1(n4870), .A2(keyinput127), .B1(n4415), .B2(keyinput122), 
        .ZN(n4869) );
  OAI221_X1 U5390 ( .B1(n4870), .B2(keyinput127), .C1(n4415), .C2(keyinput122), 
        .A(n4869), .ZN(n4878) );
  INV_X1 U5391 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4873) );
  AOI22_X1 U5392 ( .A1(n4873), .A2(keyinput119), .B1(n4872), .B2(keyinput111), 
        .ZN(n4871) );
  OAI221_X1 U5393 ( .B1(n4873), .B2(keyinput119), .C1(n4872), .C2(keyinput111), 
        .A(n4871), .ZN(n4877) );
  XNOR2_X1 U5394 ( .A(REG2_REG_24__SCAN_IN), .B(keyinput94), .ZN(n4875) );
  XNOR2_X1 U5395 ( .A(IR_REG_6__SCAN_IN), .B(keyinput99), .ZN(n4874) );
  NAND2_X1 U5396 ( .A1(n4875), .A2(n4874), .ZN(n4876) );
  NOR4_X1 U5397 ( .A1(n4879), .A2(n4878), .A3(n4877), .A4(n4876), .ZN(n4895)
         );
  AOI22_X1 U5398 ( .A1(n4882), .A2(keyinput95), .B1(n4881), .B2(keyinput90), 
        .ZN(n4880) );
  OAI221_X1 U5399 ( .B1(n4882), .B2(keyinput95), .C1(n4881), .C2(keyinput90), 
        .A(n4880), .ZN(n4893) );
  AOI22_X1 U5400 ( .A1(n2903), .A2(keyinput86), .B1(keyinput82), .B2(n4884), 
        .ZN(n4883) );
  OAI221_X1 U5401 ( .B1(n2903), .B2(keyinput86), .C1(n4884), .C2(keyinput82), 
        .A(n4883), .ZN(n4892) );
  INV_X1 U5402 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U5403 ( .A1(n4887), .A2(keyinput83), .B1(keyinput74), .B2(n4886), 
        .ZN(n4885) );
  OAI221_X1 U5404 ( .B1(n4887), .B2(keyinput83), .C1(n4886), .C2(keyinput74), 
        .A(n4885), .ZN(n4891) );
  AOI22_X1 U5405 ( .A1(n4889), .A2(keyinput78), .B1(keyinput71), .B2(n4379), 
        .ZN(n4888) );
  OAI221_X1 U5406 ( .B1(n4889), .B2(keyinput78), .C1(n4379), .C2(keyinput71), 
        .A(n4888), .ZN(n4890) );
  NOR4_X1 U5407 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n4890), .ZN(n4894)
         );
  NAND4_X1 U5408 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n5030)
         );
  AOI22_X1 U5409 ( .A1(n4900), .A2(keyinput50), .B1(n4899), .B2(keyinput47), 
        .ZN(n4898) );
  OAI221_X1 U5410 ( .B1(n4900), .B2(keyinput50), .C1(n4899), .C2(keyinput47), 
        .A(n4898), .ZN(n4910) );
  AOI22_X1 U5411 ( .A1(n4902), .A2(keyinput63), .B1(keyinput58), .B2(n2917), 
        .ZN(n4901) );
  OAI221_X1 U5412 ( .B1(n4902), .B2(keyinput63), .C1(n2917), .C2(keyinput58), 
        .A(n4901), .ZN(n4909) );
  AOI22_X1 U5413 ( .A1(n4371), .A2(keyinput70), .B1(n4904), .B2(keyinput66), 
        .ZN(n4903) );
  OAI221_X1 U5414 ( .B1(n4371), .B2(keyinput70), .C1(n4904), .C2(keyinput66), 
        .A(n4903), .ZN(n4908) );
  XNOR2_X1 U5415 ( .A(REG1_REG_26__SCAN_IN), .B(keyinput59), .ZN(n4906) );
  XNOR2_X1 U5416 ( .A(IR_REG_0__SCAN_IN), .B(keyinput46), .ZN(n4905) );
  NAND2_X1 U5417 ( .A1(n4906), .A2(n4905), .ZN(n4907) );
  NOR4_X1 U5418 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n4953)
         );
  AOI22_X1 U5419 ( .A1(n4912), .A2(keyinput22), .B1(n2672), .B2(keyinput27), 
        .ZN(n4911) );
  OAI221_X1 U5420 ( .B1(n4912), .B2(keyinput22), .C1(n2672), .C2(keyinput27), 
        .A(n4911), .ZN(n4923) );
  AOI22_X1 U5421 ( .A1(n2938), .A2(keyinput42), .B1(n3181), .B2(keyinput39), 
        .ZN(n4913) );
  OAI221_X1 U5422 ( .B1(n2938), .B2(keyinput42), .C1(n3181), .C2(keyinput39), 
        .A(n4913), .ZN(n4922) );
  AOI22_X1 U5423 ( .A1(n4916), .A2(keyinput38), .B1(n4915), .B2(keyinput35), 
        .ZN(n4914) );
  OAI221_X1 U5424 ( .B1(n4916), .B2(keyinput38), .C1(n4915), .C2(keyinput35), 
        .A(n4914), .ZN(n4921) );
  XOR2_X1 U5425 ( .A(n4917), .B(keyinput30), .Z(n4919) );
  XNOR2_X1 U5426 ( .A(IR_REG_22__SCAN_IN), .B(keyinput26), .ZN(n4918) );
  NAND2_X1 U5427 ( .A1(n4919), .A2(n4918), .ZN(n4920) );
  NOR4_X1 U5428 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(n4952)
         );
  AOI22_X1 U5429 ( .A1(n4925), .A2(keyinput18), .B1(n2586), .B2(keyinput19), 
        .ZN(n4924) );
  OAI221_X1 U5430 ( .B1(n4925), .B2(keyinput18), .C1(n2586), .C2(keyinput19), 
        .A(n4924), .ZN(n4936) );
  AOI22_X1 U5431 ( .A1(n4928), .A2(keyinput15), .B1(keyinput10), .B2(n4927), 
        .ZN(n4926) );
  OAI221_X1 U5432 ( .B1(n4928), .B2(keyinput15), .C1(n4927), .C2(keyinput10), 
        .A(n4926), .ZN(n4935) );
  AOI22_X1 U5433 ( .A1(n3495), .A2(keyinput11), .B1(keyinput49), .B2(n4930), 
        .ZN(n4929) );
  OAI221_X1 U5434 ( .B1(n3495), .B2(keyinput11), .C1(n4930), .C2(keyinput49), 
        .A(n4929), .ZN(n4934) );
  AOI22_X1 U5435 ( .A1(n4932), .A2(keyinput41), .B1(keyinput29), .B2(n4317), 
        .ZN(n4931) );
  OAI221_X1 U5436 ( .B1(n4932), .B2(keyinput41), .C1(n4317), .C2(keyinput29), 
        .A(n4931), .ZN(n4933) );
  NOR4_X1 U5437 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), .ZN(n4951)
         );
  INV_X1 U5438 ( .A(DATAI_3_), .ZN(n4938) );
  AOI22_X1 U5439 ( .A1(n4938), .A2(keyinput25), .B1(n3531), .B2(keyinput93), 
        .ZN(n4937) );
  OAI221_X1 U5440 ( .B1(n4938), .B2(keyinput25), .C1(n3531), .C2(keyinput93), 
        .A(n4937), .ZN(n4949) );
  AOI22_X1 U5441 ( .A1(n4941), .A2(keyinput77), .B1(keyinput13), .B2(n4940), 
        .ZN(n4939) );
  OAI221_X1 U5442 ( .B1(n4941), .B2(keyinput77), .C1(n4940), .C2(keyinput13), 
        .A(n4939), .ZN(n4948) );
  INV_X1 U5443 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4942) );
  XOR2_X1 U5444 ( .A(n4942), .B(keyinput73), .Z(n4946) );
  XNOR2_X1 U5445 ( .A(IR_REG_13__SCAN_IN), .B(keyinput89), .ZN(n4945) );
  XNOR2_X1 U5446 ( .A(IR_REG_14__SCAN_IN), .B(keyinput1), .ZN(n4944) );
  XNOR2_X1 U5447 ( .A(IR_REG_27__SCAN_IN), .B(keyinput5), .ZN(n4943) );
  NAND4_X1 U5448 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n4947)
         );
  NOR3_X1 U5449 ( .A1(n4949), .A2(n4948), .A3(n4947), .ZN(n4950) );
  NAND4_X1 U5450 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n5029)
         );
  OAI22_X1 U5451 ( .A1(DATAO_REG_0__SCAN_IN), .A2(keyinput4), .B1(
        DATAO_REG_23__SCAN_IN), .B2(keyinput7), .ZN(n4954) );
  AOI221_X1 U5452 ( .B1(DATAO_REG_0__SCAN_IN), .B2(keyinput4), .C1(keyinput7), 
        .C2(DATAO_REG_23__SCAN_IN), .A(n4954), .ZN(n4961) );
  OAI22_X1 U5453 ( .A1(REG1_REG_8__SCAN_IN), .A2(keyinput8), .B1(
        DATAO_REG_20__SCAN_IN), .B2(keyinput24), .ZN(n4955) );
  AOI221_X1 U5454 ( .B1(REG1_REG_8__SCAN_IN), .B2(keyinput8), .C1(keyinput24), 
        .C2(DATAO_REG_20__SCAN_IN), .A(n4955), .ZN(n4960) );
  OAI22_X1 U5455 ( .A1(DATAI_28_), .A2(keyinput31), .B1(REG1_REG_15__SCAN_IN), 
        .B2(keyinput3), .ZN(n4956) );
  AOI221_X1 U5456 ( .B1(DATAI_28_), .B2(keyinput31), .C1(keyinput3), .C2(
        REG1_REG_15__SCAN_IN), .A(n4956), .ZN(n4959) );
  OAI22_X1 U5457 ( .A1(DATAO_REG_11__SCAN_IN), .A2(keyinput43), .B1(keyinput23), .B2(ADDR_REG_2__SCAN_IN), .ZN(n4957) );
  AOI221_X1 U5458 ( .B1(DATAO_REG_11__SCAN_IN), .B2(keyinput43), .C1(
        ADDR_REG_2__SCAN_IN), .C2(keyinput23), .A(n4957), .ZN(n4958) );
  NAND4_X1 U5459 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4989)
         );
  OAI22_X1 U5460 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput44), .B1(keyinput48), 
        .B2(DATAI_0_), .ZN(n4962) );
  AOI221_X1 U5461 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput44), .C1(DATAI_0_), 
        .C2(keyinput48), .A(n4962), .ZN(n4969) );
  OAI22_X1 U5462 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput32), .B1(keyinput40), 
        .B2(REG0_REG_25__SCAN_IN), .ZN(n4963) );
  AOI221_X1 U5463 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput32), .C1(
        REG0_REG_25__SCAN_IN), .C2(keyinput40), .A(n4963), .ZN(n4968) );
  OAI22_X1 U5464 ( .A1(DATAI_15_), .A2(keyinput16), .B1(keyinput20), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n4964) );
  AOI221_X1 U5465 ( .B1(DATAI_15_), .B2(keyinput16), .C1(REG1_REG_24__SCAN_IN), 
        .C2(keyinput20), .A(n4964), .ZN(n4967) );
  OAI22_X1 U5466 ( .A1(REG2_REG_22__SCAN_IN), .A2(keyinput28), .B1(keyinput12), 
        .B2(DATAI_19_), .ZN(n4965) );
  AOI221_X1 U5467 ( .B1(REG2_REG_22__SCAN_IN), .B2(keyinput28), .C1(DATAI_19_), 
        .C2(keyinput12), .A(n4965), .ZN(n4966) );
  NAND4_X1 U5468 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n4988)
         );
  OAI22_X1 U5469 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput57), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput53), .ZN(n4970) );
  AOI221_X1 U5470 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput57), .C1(keyinput53), 
        .C2(REG0_REG_6__SCAN_IN), .A(n4970), .ZN(n4977) );
  OAI22_X1 U5471 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput33), .B1(keyinput61), 
        .B2(REG0_REG_15__SCAN_IN), .ZN(n4971) );
  AOI221_X1 U5472 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput33), .C1(
        REG0_REG_15__SCAN_IN), .C2(keyinput61), .A(n4971), .ZN(n4976) );
  OAI22_X1 U5473 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput21), .B1(keyinput37), 
        .B2(ADDR_REG_16__SCAN_IN), .ZN(n4972) );
  AOI221_X1 U5474 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput21), .C1(
        ADDR_REG_16__SCAN_IN), .C2(keyinput37), .A(n4972), .ZN(n4975) );
  OAI22_X1 U5475 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput9), .B1(keyinput17), 
        .B2(REG1_REG_11__SCAN_IN), .ZN(n4973) );
  AOI221_X1 U5476 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput9), .C1(
        REG1_REG_11__SCAN_IN), .C2(keyinput17), .A(n4973), .ZN(n4974) );
  NAND4_X1 U5477 ( .A1(n4977), .A2(n4976), .A3(n4975), .A4(n4974), .ZN(n4987)
         );
  OAI22_X1 U5478 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput65), .B1(keyinput69), 
        .B2(DATAI_24_), .ZN(n4978) );
  AOI221_X1 U5479 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput65), .C1(DATAI_24_), 
        .C2(keyinput69), .A(n4978), .ZN(n4985) );
  OAI22_X1 U5480 ( .A1(DATAI_27_), .A2(keyinput81), .B1(DATAO_REG_13__SCAN_IN), 
        .B2(keyinput85), .ZN(n4979) );
  AOI221_X1 U5481 ( .B1(DATAI_27_), .B2(keyinput81), .C1(keyinput85), .C2(
        DATAO_REG_13__SCAN_IN), .A(n4979), .ZN(n4984) );
  OAI22_X1 U5482 ( .A1(D_REG_20__SCAN_IN), .A2(keyinput97), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput101), .ZN(n4980) );
  AOI221_X1 U5483 ( .B1(D_REG_20__SCAN_IN), .B2(keyinput97), .C1(keyinput101), 
        .C2(IR_REG_30__SCAN_IN), .A(n4980), .ZN(n4983) );
  OAI22_X1 U5484 ( .A1(DATAI_29_), .A2(keyinput109), .B1(REG1_REG_30__SCAN_IN), 
        .B2(keyinput121), .ZN(n4981) );
  AOI221_X1 U5485 ( .B1(DATAI_29_), .B2(keyinput109), .C1(keyinput121), .C2(
        REG1_REG_30__SCAN_IN), .A(n4981), .ZN(n4982) );
  NAND4_X1 U5486 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n4986)
         );
  NOR4_X1 U5487 ( .A1(n4989), .A2(n4988), .A3(n4987), .A4(n4986), .ZN(n5027)
         );
  OAI22_X1 U5488 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput6), .B1(
        DATAO_REG_6__SCAN_IN), .B2(keyinput87), .ZN(n4990) );
  AOI221_X1 U5489 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput6), .C1(keyinput87), 
        .C2(DATAO_REG_6__SCAN_IN), .A(n4990), .ZN(n4997) );
  OAI22_X1 U5490 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput2), .B1(keyinput14), 
        .B2(ADDR_REG_13__SCAN_IN), .ZN(n4991) );
  AOI221_X1 U5491 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput2), .C1(
        ADDR_REG_13__SCAN_IN), .C2(keyinput14), .A(n4991), .ZN(n4996) );
  OAI22_X1 U5492 ( .A1(DATAI_26_), .A2(keyinput55), .B1(keyinput103), .B2(
        REG2_REG_6__SCAN_IN), .ZN(n4992) );
  AOI221_X1 U5493 ( .B1(DATAI_26_), .B2(keyinput55), .C1(REG2_REG_6__SCAN_IN), 
        .C2(keyinput103), .A(n4992), .ZN(n4995) );
  OAI22_X1 U5494 ( .A1(REG0_REG_30__SCAN_IN), .A2(keyinput91), .B1(keyinput79), 
        .B2(ADDR_REG_9__SCAN_IN), .ZN(n4993) );
  AOI221_X1 U5495 ( .B1(REG0_REG_30__SCAN_IN), .B2(keyinput91), .C1(
        ADDR_REG_9__SCAN_IN), .C2(keyinput79), .A(n4993), .ZN(n4994) );
  NAND4_X1 U5496 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), .ZN(n5025)
         );
  OAI22_X1 U5497 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput110), .B1(
        REG2_REG_10__SCAN_IN), .B2(keyinput118), .ZN(n4998) );
  AOI221_X1 U5498 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput110), .C1(keyinput118), 
        .C2(REG2_REG_10__SCAN_IN), .A(n4998), .ZN(n5005) );
  OAI22_X1 U5499 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput106), .B1(keyinput114), 
        .B2(REG0_REG_1__SCAN_IN), .ZN(n4999) );
  AOI221_X1 U5500 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput106), .C1(
        REG0_REG_1__SCAN_IN), .C2(keyinput114), .A(n4999), .ZN(n5004) );
  OAI22_X1 U5501 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput34), .B1(keyinput54), 
        .B2(REG3_REG_21__SCAN_IN), .ZN(n5000) );
  AOI221_X1 U5502 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput34), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput54), .A(n5000), .ZN(n5003) );
  OAI22_X1 U5503 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput98), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput62), .ZN(n5001) );
  AOI221_X1 U5504 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput98), .C1(keyinput62), .C2(DATAO_REG_8__SCAN_IN), .A(n5001), .ZN(n5002) );
  NAND4_X1 U5505 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n5024)
         );
  OAI22_X1 U5506 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput96), .B1(DATAI_23_), 
        .B2(keyinput84), .ZN(n5006) );
  AOI221_X1 U5507 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput96), .C1(keyinput84), 
        .C2(DATAI_23_), .A(n5006), .ZN(n5013) );
  OAI22_X1 U5508 ( .A1(DATAO_REG_19__SCAN_IN), .A2(keyinput64), .B1(
        keyinput115), .B2(DATAO_REG_21__SCAN_IN), .ZN(n5007) );
  AOI221_X1 U5509 ( .B1(DATAO_REG_19__SCAN_IN), .B2(keyinput64), .C1(
        DATAO_REG_21__SCAN_IN), .C2(keyinput115), .A(n5007), .ZN(n5012) );
  OAI22_X1 U5510 ( .A1(REG2_REG_13__SCAN_IN), .A2(keyinput52), .B1(DATAI_5_), 
        .B2(keyinput45), .ZN(n5008) );
  AOI221_X1 U5511 ( .B1(REG2_REG_13__SCAN_IN), .B2(keyinput52), .C1(keyinput45), .C2(DATAI_5_), .A(n5008), .ZN(n5011) );
  OAI22_X1 U5512 ( .A1(REG2_REG_4__SCAN_IN), .A2(keyinput88), .B1(keyinput56), 
        .B2(ADDR_REG_0__SCAN_IN), .ZN(n5009) );
  AOI221_X1 U5513 ( .B1(REG2_REG_4__SCAN_IN), .B2(keyinput88), .C1(
        ADDR_REG_0__SCAN_IN), .C2(keyinput56), .A(n5009), .ZN(n5010) );
  NAND4_X1 U5514 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n5023)
         );
  OAI22_X1 U5515 ( .A1(REG2_REG_9__SCAN_IN), .A2(keyinput67), .B1(DATAI_4_), 
        .B2(keyinput124), .ZN(n5014) );
  AOI221_X1 U5516 ( .B1(REG2_REG_9__SCAN_IN), .B2(keyinput67), .C1(keyinput124), .C2(DATAI_4_), .A(n5014), .ZN(n5021) );
  OAI22_X1 U5517 ( .A1(REG0_REG_29__SCAN_IN), .A2(keyinput51), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput75), .ZN(n5015) );
  AOI221_X1 U5518 ( .B1(REG0_REG_29__SCAN_IN), .B2(keyinput51), .C1(keyinput75), .C2(REG3_REG_10__SCAN_IN), .A(n5015), .ZN(n5020) );
  OAI22_X1 U5519 ( .A1(DATAI_12_), .A2(keyinput123), .B1(keyinput108), .B2(
        DATAI_30_), .ZN(n5016) );
  AOI221_X1 U5520 ( .B1(DATAI_12_), .B2(keyinput123), .C1(DATAI_30_), .C2(
        keyinput108), .A(n5016), .ZN(n5019) );
  OAI22_X1 U5521 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput120), .B1(DATAI_21_), 
        .B2(keyinput104), .ZN(n5017) );
  AOI221_X1 U5522 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput120), .C1(keyinput104), .C2(DATAI_21_), .A(n5017), .ZN(n5018) );
  NAND4_X1 U5523 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n5022)
         );
  NOR4_X1 U5524 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n5026)
         );
  NAND2_X1 U5525 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  NOR4_X1 U5526 ( .A1(n5031), .A2(n5030), .A3(n5029), .A4(n5028), .ZN(n5047)
         );
  NAND2_X1 U5527 ( .A1(n5033), .A2(n5032), .ZN(n5037) );
  AOI22_X1 U5528 ( .A1(n5040), .A2(REG2_REG_6__SCAN_IN), .B1(n5035), .B2(n5034), .ZN(n5036) );
  OAI211_X1 U5529 ( .C1(n5039), .C2(n5038), .A(n5037), .B(n5036), .ZN(n5043)
         );
  NOR2_X1 U5530 ( .A1(n5041), .A2(n5040), .ZN(n5042) );
  AOI211_X1 U5531 ( .C1(n5045), .C2(n5044), .A(n5043), .B(n5042), .ZN(n5046)
         );
  XNOR2_X1 U5532 ( .A(n5047), .B(n5046), .ZN(U3284) );
  INV_X2 U2498 ( .A(n2725), .ZN(n2702) );
endmodule

