

module b17_C_SARLock_k_64_5 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051;

  AOI21_X1 U11015 ( .B1(n12851), .B2(n12845), .A(n12850), .ZN(n14419) );
  INV_X2 U11016 ( .A(n17922), .ZN(n17893) );
  AND2_X1 U11017 ( .A1(n12906), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20104)
         );
  INV_X4 U11018 ( .A(n20101), .ZN(n12840) );
  OR2_X1 U11019 ( .A1(n10815), .A2(n10814), .ZN(n19724) );
  OR2_X1 U11020 ( .A1(n9857), .A2(n10813), .ZN(n10896) );
  OR2_X1 U11021 ( .A1(n9857), .A2(n10814), .ZN(n13440) );
  INV_X2 U11022 ( .A(n9583), .ZN(n9577) );
  NAND2_X1 U11023 ( .A1(n12740), .A2(n12739), .ZN(n12745) );
  CLKBUF_X2 U11024 ( .A(n10599), .Z(n11593) );
  CLKBUF_X2 U11025 ( .A(n9611), .Z(n9576) );
  AND2_X1 U11026 ( .A1(n9628), .A2(n16349), .ZN(n13886) );
  AND2_X1 U11027 ( .A1(n9628), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10912) );
  INV_X2 U11029 ( .A(n12858), .ZN(n12624) );
  CLKBUF_X2 U11030 ( .A(n11828), .Z(n12511) );
  INV_X1 U11031 ( .A(n9588), .ZN(n11809) );
  CLKBUF_X1 U11032 ( .A(n12510), .Z(n12487) );
  CLKBUF_X2 U11033 ( .A(n11665), .Z(n9580) );
  INV_X1 U11034 ( .A(n10713), .ZN(n10689) );
  AND2_X1 U11035 ( .A1(n11634), .A2(n14627), .ZN(n11790) );
  INV_X2 U11036 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10718) );
  AND2_X1 U11037 ( .A1(n9786), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11625) );
  CLKBUF_X1 U11038 ( .A(n20147), .Z(n9570) );
  NOR2_X1 U11039 ( .A1(n20104), .A2(n20106), .ZN(n20147) );
  CLKBUF_X1 U11040 ( .A(n20146), .Z(n9571) );
  NOR2_X1 U11041 ( .A1(n20106), .A2(n20105), .ZN(n20146) );
  CLKBUF_X1 U11042 ( .A(n18168), .Z(n9572) );
  NOR3_X1 U11043 ( .A1(n18700), .A2(n18254), .A3(n17427), .ZN(n18168) );
  INV_X4 U11044 ( .A(n18253), .ZN(n9587) );
  XNOR2_X1 U11045 ( .A(n20915), .B(keyinput47), .ZN(n20916) );
  AND2_X2 U11046 ( .A1(n11625), .A2(n9727), .ZN(n9619) );
  AND2_X2 U11047 ( .A1(n11625), .A2(n9727), .ZN(n9618) );
  INV_X1 U11048 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16349) );
  INV_X1 U11049 ( .A(n20109), .ZN(n13209) );
  BUF_X1 U11050 ( .A(n10462), .Z(n21040) );
  NAND2_X1 U11051 ( .A1(n14863), .A2(n13989), .ZN(n14011) );
  NOR2_X1 U11052 ( .A1(n14965), .A2(n13939), .ZN(n14869) );
  NAND2_X1 U11053 ( .A1(n15228), .A2(n15555), .ZN(n15229) );
  OR2_X1 U11054 ( .A1(n9857), .A2(n10807), .ZN(n10895) );
  OR2_X1 U11055 ( .A1(n10815), .A2(n10807), .ZN(n15615) );
  INV_X1 U11056 ( .A(n17148), .ZN(n17206) );
  BUF_X1 U11057 ( .A(n17226), .Z(n9622) );
  NOR2_X1 U11058 ( .A1(n14183), .A2(n14185), .ZN(n14167) );
  BUF_X1 U11059 ( .A(n11764), .Z(n13412) );
  CLKBUF_X2 U11060 ( .A(n11206), .Z(n11564) );
  NOR2_X1 U11061 ( .A1(n10716), .A2(n10705), .ZN(n10706) );
  OR2_X1 U11062 ( .A1(n9596), .A2(n9597), .ZN(n14845) );
  NOR2_X2 U11063 ( .A1(n15130), .A2(n10994), .ZN(n15120) );
  INV_X1 U11064 ( .A(n16949), .ZN(n16918) );
  INV_X1 U11065 ( .A(n18269), .ZN(n15632) );
  INV_X1 U11066 ( .A(n10231), .ZN(n10131) );
  NOR4_X2 U11067 ( .A1(n15632), .A2(n10403), .A3(n18291), .A4(n10393), .ZN(
        n17497) );
  INV_X1 U11068 ( .A(n19974), .ZN(n19987) );
  AOI21_X1 U11070 ( .B1(n14851), .B2(n14853), .A(n14852), .ZN(n14937) );
  BUF_X1 U11071 ( .A(n10711), .Z(n14062) );
  INV_X2 U11072 ( .A(n10102), .ZN(n17212) );
  INV_X1 U11073 ( .A(n17780), .ZN(n17758) );
  INV_X1 U11074 ( .A(n18716), .ZN(n18725) );
  OR3_X1 U11075 ( .A1(n11537), .A2(n15018), .A3(n19264), .ZN(n9573) );
  INV_X1 U11076 ( .A(n10086), .ZN(n17137) );
  NOR2_X1 U11077 ( .A1(n14964), .A2(n14966), .ZN(n14965) );
  AND2_X2 U11078 ( .A1(n12888), .A2(n11753), .ZN(n13401) );
  NOR2_X4 U11079 ( .A1(n10806), .A2(n13738), .ZN(n19284) );
  BUF_X1 U11080 ( .A(n10774), .Z(n11206) );
  AND2_X2 U11081 ( .A1(n11008), .A2(n11002), .ZN(n11016) );
  NOR2_X1 U11082 ( .A1(n18277), .A2(n16557), .ZN(n9574) );
  INV_X1 U11083 ( .A(n17911), .ZN(n17926) );
  AND2_X2 U11084 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13468) );
  INV_X2 U11085 ( .A(n10703), .ZN(n10609) );
  AND2_X4 U11086 ( .A1(n10726), .A2(n10599), .ZN(n10742) );
  NOR2_X2 U11087 ( .A1(n20126), .A2(n20130), .ZN(n13474) );
  AND2_X4 U11088 ( .A1(n13781), .A2(n10459), .ZN(n10622) );
  CLKBUF_X2 U11089 ( .A(n10622), .Z(n9623) );
  NAND2_X2 U11090 ( .A1(n9728), .A2(n12758), .ZN(n12763) );
  NAND2_X2 U11091 ( .A1(n9966), .A2(n9964), .ZN(n10726) );
  AOI21_X2 U11092 ( .B1(n11522), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11154), .ZN(n11161) );
  BUF_X1 U11093 ( .A(n15006), .Z(n9575) );
  OAI21_X2 U11094 ( .B1(n17918), .B2(n17702), .A(n18587), .ZN(n17763) );
  XNOR2_X2 U11095 ( .A(n12745), .B(n20080), .ZN(n13274) );
  NOR2_X2 U11096 ( .A1(n13520), .A2(n10059), .ZN(n14901) );
  NOR2_X1 U11097 ( .A1(n18731), .A2(n10090), .ZN(n10231) );
  INV_X4 U11098 ( .A(n10131), .ZN(n17250) );
  XNOR2_X2 U11099 ( .A(n13938), .B(n13937), .ZN(n14964) );
  NAND2_X2 U11100 ( .A1(n20079), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20080) );
  OR2_X1 U11101 ( .A1(n13151), .A2(n13673), .ZN(n10805) );
  AND2_X2 U11102 ( .A1(n15120), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15103) );
  NOR2_X1 U11103 ( .A1(n14857), .A2(n14859), .ZN(n14858) );
  AND2_X1 U11104 ( .A1(n9598), .A2(n10064), .ZN(n9597) );
  XOR2_X1 U11105 ( .A(n11614), .B(n14835), .Z(n15006) );
  INV_X1 U11106 ( .A(n17313), .ZN(n17309) );
  AND2_X1 U11107 ( .A1(n16245), .A2(n13937), .ZN(n13939) );
  AND3_X1 U11108 ( .A1(n17619), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17613), .ZN(n17603) );
  NOR2_X1 U11109 ( .A1(n17671), .A2(n10217), .ZN(n17614) );
  NOR2_X1 U11110 ( .A1(n17671), .A2(n17657), .ZN(n17658) );
  INV_X2 U11111 ( .A(n14579), .ZN(n15975) );
  BUF_X1 U11112 ( .A(n13503), .Z(n9615) );
  OR2_X1 U11113 ( .A1(n10805), .A2(n10788), .ZN(n19464) );
  OR2_X1 U11114 ( .A1(n10805), .A2(n10789), .ZN(n19347) );
  OR2_X1 U11115 ( .A1(n10815), .A2(n10813), .ZN(n13370) );
  NOR2_X1 U11116 ( .A1(n18722), .A2(n15828), .ZN(n17450) );
  OR3_X1 U11117 ( .A1(n11038), .A2(n11593), .A3(n11587), .ZN(n11130) );
  CLKBUF_X2 U11118 ( .A(n11712), .Z(n12835) );
  NOR2_X2 U11119 ( .A1(n10735), .A2(n10731), .ZN(n10717) );
  INV_X2 U11120 ( .A(n11284), .ZN(n11314) );
  NOR2_X2 U11121 ( .A1(n11757), .A2(n20109), .ZN(n13599) );
  CLKBUF_X2 U11122 ( .A(n11695), .Z(n20126) );
  CLKBUF_X2 U11123 ( .A(n11751), .Z(n20148) );
  CLKBUF_X2 U11124 ( .A(n11679), .Z(n20142) );
  INV_X4 U11125 ( .A(n10462), .ZN(n10722) );
  BUF_X1 U11126 ( .A(n10147), .Z(n17224) );
  CLKBUF_X2 U11127 ( .A(n13248), .Z(n21034) );
  INV_X4 U11128 ( .A(n17199), .ZN(n10142) );
  INV_X4 U11129 ( .A(n17156), .ZN(n17211) );
  INV_X1 U11130 ( .A(n11838), .ZN(n9588) );
  INV_X4 U11131 ( .A(n9722), .ZN(n17243) );
  INV_X4 U11132 ( .A(n15688), .ZN(n10178) );
  CLKBUF_X2 U11133 ( .A(n17249), .Z(n9616) );
  CLKBUF_X2 U11134 ( .A(n11789), .Z(n12302) );
  BUF_X2 U11135 ( .A(n11664), .Z(n12544) );
  INV_X2 U11136 ( .A(n9651), .ZN(n17245) );
  INV_X4 U11137 ( .A(n17142), .ZN(n10247) );
  CLKBUF_X1 U11138 ( .A(n14096), .Z(n9578) );
  INV_X1 U11139 ( .A(n12462), .ZN(n9579) );
  NOR2_X4 U11141 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11634) );
  NOR2_X2 U11143 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13488) );
  NOR2_X1 U11144 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16944) );
  NAND2_X1 U11145 ( .A1(n12846), .A2(n12845), .ZN(n14142) );
  AOI211_X1 U11146 ( .C1(n16027), .C2(n14443), .A(n14442), .B(n14441), .ZN(
        n14444) );
  XNOR2_X1 U11147 ( .A(n12850), .B(n12562), .ZN(n12896) );
  OAI21_X1 U11148 ( .B1(n14184), .B2(n14168), .A(n14152), .ZN(n14440) );
  OAI21_X1 U11149 ( .B1(n11617), .B2(n11618), .A(n11591), .ZN(n11599) );
  NOR2_X1 U11150 ( .A1(n14838), .A2(n14090), .ZN(n14108) );
  CLKBUF_X1 U11151 ( .A(n14167), .Z(n14184) );
  AOI211_X1 U11152 ( .C1(n15324), .C2(n16333), .A(n15323), .B(n15322), .ZN(
        n15325) );
  AND2_X1 U11153 ( .A1(n14454), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14466) );
  OR2_X1 U11154 ( .A1(n10002), .A2(n11142), .ZN(n11574) );
  NAND2_X1 U11155 ( .A1(n9814), .A2(n9813), .ZN(n14581) );
  OAI21_X1 U11156 ( .B1(n15192), .B2(n15081), .A(n15190), .ZN(n15175) );
  AOI21_X1 U11157 ( .B1(n15199), .B2(n15200), .A(n15080), .ZN(n15192) );
  AND2_X2 U11158 ( .A1(n14728), .A2(n9715), .ZN(n14835) );
  AND2_X1 U11159 ( .A1(n14741), .A2(n14726), .ZN(n14728) );
  AND2_X1 U11160 ( .A1(n14786), .A2(n9935), .ZN(n14741) );
  NOR2_X1 U11161 ( .A1(n14871), .A2(n13965), .ZN(n13986) );
  AND2_X1 U11162 ( .A1(n15220), .A2(n10986), .ZN(n10987) );
  NOR2_X1 U11163 ( .A1(n9995), .A2(n9724), .ZN(n9813) );
  OAI211_X1 U11164 ( .C1(n12827), .C2(n9997), .A(n12826), .B(n9992), .ZN(n9994) );
  NAND2_X1 U11165 ( .A1(n10046), .A2(n15526), .ZN(n15220) );
  OAI21_X1 U11166 ( .B1(n9629), .B2(n9872), .A(n9870), .ZN(n9869) );
  NAND2_X1 U11167 ( .A1(n12826), .A2(n9656), .ZN(n9995) );
  INV_X1 U11168 ( .A(n13759), .ZN(n9581) );
  INV_X1 U11169 ( .A(n14590), .ZN(n12826) );
  OR2_X1 U11170 ( .A1(n11035), .A2(n15526), .ZN(n9629) );
  OAI221_X1 U11171 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17729), 
        .C1(n20894), .C2(n17603), .A(n17602), .ZN(n17580) );
  NOR2_X1 U11172 ( .A1(n9667), .A2(n9736), .ZN(n9735) );
  AND2_X1 U11173 ( .A1(n14498), .A2(n12825), .ZN(n15987) );
  INV_X1 U11174 ( .A(n15541), .ZN(n10926) );
  NAND2_X1 U11175 ( .A1(n12818), .A2(n14511), .ZN(n14497) );
  AND2_X1 U11176 ( .A1(n14509), .A2(n9769), .ZN(n14498) );
  OAI21_X1 U11177 ( .B1(n17723), .B2(n18037), .A(n17722), .ZN(n17709) );
  AND2_X1 U11178 ( .A1(n10922), .A2(n11026), .ZN(n15541) );
  OR2_X1 U11179 ( .A1(n14918), .A2(n11486), .ZN(n14928) );
  NAND2_X1 U11180 ( .A1(n9862), .A2(n9864), .ZN(n15227) );
  NAND2_X1 U11181 ( .A1(n12833), .A2(n12824), .ZN(n9769) );
  NAND2_X1 U11182 ( .A1(n12008), .A2(n12007), .ZN(n13568) );
  XNOR2_X1 U11183 ( .A(n9947), .B(n12719), .ZN(n14542) );
  NAND2_X1 U11184 ( .A1(n9824), .A2(n9823), .ZN(n17671) );
  OR2_X1 U11185 ( .A1(n9825), .A2(n17833), .ZN(n9824) );
  NOR2_X1 U11186 ( .A1(n10213), .A2(n10212), .ZN(n17712) );
  INV_X1 U11187 ( .A(n10876), .ZN(n9742) );
  NAND2_X1 U11188 ( .A1(n12031), .A2(n12030), .ZN(n12807) );
  INV_X1 U11189 ( .A(n12028), .ZN(n12031) );
  NAND2_X1 U11190 ( .A1(n18965), .A2(n11596), .ZN(n11099) );
  NAND2_X1 U11191 ( .A1(n9827), .A2(n9641), .ZN(n9823) );
  NOR2_X1 U11192 ( .A1(n17893), .A2(n17676), .ZN(n17919) );
  OAI21_X1 U11193 ( .B1(n12759), .B2(n12093), .A(n11953), .ZN(n13510) );
  OAI21_X1 U11194 ( .B1(n12749), .B2(n12775), .A(n9632), .ZN(n13363) );
  NAND2_X1 U11195 ( .A1(n17915), .A2(n17427), .ZN(n17837) );
  OR2_X1 U11196 ( .A1(n11122), .A2(n11121), .ZN(n11129) );
  AND2_X1 U11197 ( .A1(n10959), .A2(n10958), .ZN(n15515) );
  NAND2_X1 U11198 ( .A1(n11997), .A2(n11996), .ZN(n12028) );
  NAND2_X1 U11199 ( .A1(n11979), .A2(n11947), .ZN(n12759) );
  NAND2_X1 U11200 ( .A1(n14289), .A2(n14210), .ZN(n14212) );
  NOR2_X2 U11201 ( .A1(n18277), .A2(n16557), .ZN(n17911) );
  OAI21_X2 U11202 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18909), .A(n16557), 
        .ZN(n17922) );
  AND3_X1 U11203 ( .A1(n9803), .A2(n13576), .A3(n11978), .ZN(n11997) );
  NOR2_X1 U11204 ( .A1(n17830), .A2(n18165), .ZN(n17829) );
  NAND2_X1 U11205 ( .A1(n18708), .A2(n18910), .ZN(n16557) );
  AND2_X1 U11206 ( .A1(n11896), .A2(n11895), .ZN(n9803) );
  NOR2_X1 U11207 ( .A1(n13194), .A2(n13282), .ZN(n13350) );
  NOR2_X1 U11208 ( .A1(n14310), .A2(n14299), .ZN(n14300) );
  OR3_X2 U11209 ( .A1(n11069), .A2(P2_EBX_REG_20__SCAN_IN), .A3(n11064), .ZN(
        n11117) );
  OR2_X1 U11210 ( .A1(n10888), .A2(n10887), .ZN(n10889) );
  OAI22_X1 U11211 ( .A1(n10832), .A2(n13440), .B1(n13370), .B2(n13948), .ZN(
        n10833) );
  NAND2_X1 U11212 ( .A1(n10818), .A2(n10817), .ZN(n19675) );
  NAND2_X1 U11213 ( .A1(n9804), .A2(n11945), .ZN(n13576) );
  NOR2_X1 U11214 ( .A1(n18177), .A2(n17845), .ZN(n17844) );
  NAND2_X1 U11215 ( .A1(n10798), .A2(n10797), .ZN(n9745) );
  OR2_X1 U11216 ( .A1(n10881), .A2(n10835), .ZN(n10837) );
  OAI22_X1 U11217 ( .A1(n13458), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12752), 
        .B2(n12804), .ZN(n11894) );
  NAND2_X1 U11218 ( .A1(n11862), .A2(n11850), .ZN(n11905) );
  XNOR2_X1 U11219 ( .A(n13491), .B(n20270), .ZN(n20415) );
  OAI211_X1 U11220 ( .C1(n20231), .C2(n9785), .A(n9784), .B(n11872), .ZN(
        n13491) );
  NAND2_X1 U11221 ( .A1(n11354), .A2(n11353), .ZN(n15504) );
  NAND2_X1 U11222 ( .A1(n12614), .A2(n12615), .ZN(n13390) );
  NOR2_X1 U11223 ( .A1(n19258), .A2(n10813), .ZN(n10797) );
  OR2_X1 U11224 ( .A1(n11849), .A2(n11848), .ZN(n11862) );
  AND2_X1 U11225 ( .A1(n11059), .A2(n9914), .ZN(n11089) );
  NOR2_X2 U11226 ( .A1(n19293), .A2(n19680), .ZN(n19294) );
  NOR2_X2 U11227 ( .A1(n19223), .A2(n19680), .ZN(n13380) );
  NOR2_X2 U11228 ( .A1(n14062), .A2(n19308), .ZN(n13381) );
  INV_X1 U11229 ( .A(n15732), .ZN(n15740) );
  NOR2_X2 U11230 ( .A1(n13453), .A2(n19680), .ZN(n13454) );
  NOR2_X2 U11231 ( .A1(n13448), .A2(n19680), .ZN(n13449) );
  AND2_X1 U11232 ( .A1(n16188), .A2(n9698), .ZN(n14361) );
  AND2_X1 U11233 ( .A1(n10785), .A2(n10790), .ZN(n13673) );
  NAND2_X1 U11234 ( .A1(n9750), .A2(n9749), .ZN(n10772) );
  AOI21_X1 U11235 ( .B1(n11866), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11867), .ZN(n11875) );
  NAND2_X1 U11236 ( .A1(n14674), .A2(n13650), .ZN(n19110) );
  NOR2_X1 U11237 ( .A1(n11334), .A2(n9969), .ZN(n9971) );
  INV_X2 U11238 ( .A(n17295), .ZN(n9582) );
  CLKBUF_X1 U11239 ( .A(n11865), .Z(n11866) );
  XNOR2_X1 U11240 ( .A(n11167), .B(n11165), .ZN(n11164) );
  NAND2_X1 U11241 ( .A1(n10767), .A2(n10768), .ZN(n10769) );
  NOR2_X1 U11242 ( .A1(n10325), .A2(n10324), .ZN(n10390) );
  AOI21_X1 U11243 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(n17886) );
  XNOR2_X1 U11244 ( .A(n13127), .B(n11326), .ZN(n13265) );
  NAND2_X1 U11245 ( .A1(n11016), .A2(n11015), .ZN(n11023) );
  AND2_X1 U11246 ( .A1(n10766), .A2(n10765), .ZN(n10767) );
  OR4_X1 U11247 ( .A1(n18284), .A2(n18287), .A3(n10395), .A4(n10326), .ZN(
        n10392) );
  INV_X1 U11248 ( .A(n13779), .ZN(n10741) );
  AND2_X1 U11249 ( .A1(n13130), .A2(n13129), .ZN(n13127) );
  INV_X1 U11250 ( .A(n17303), .ZN(n18295) );
  NAND2_X1 U11251 ( .A1(n12928), .A2(n10748), .ZN(n12939) );
  CLKBUF_X1 U11252 ( .A(n12889), .Z(n13220) );
  NAND2_X1 U11253 ( .A1(n9675), .A2(n11766), .ZN(n13211) );
  OAI211_X1 U11254 ( .C1(n10701), .C2(n11282), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n10700), .ZN(n10702) );
  NAND2_X1 U11255 ( .A1(n10999), .A2(n10998), .ZN(n11010) );
  INV_X1 U11256 ( .A(n10764), .ZN(n9583) );
  NAND2_X1 U11257 ( .A1(n13424), .A2(n11767), .ZN(n14623) );
  CLKBUF_X1 U11258 ( .A(n10691), .Z(n9591) );
  AND2_X1 U11259 ( .A1(n11286), .A2(n10728), .ZN(n10729) );
  OAI211_X1 U11260 ( .C1(n17199), .C2(n20973), .A(n10186), .B(n10185), .ZN(
        n17921) );
  INV_X1 U11261 ( .A(n11763), .ZN(n13424) );
  AND2_X1 U11262 ( .A1(n11765), .A2(n20148), .ZN(n11774) );
  MUX2_X1 U11263 ( .A(n11322), .B(n11000), .S(n11593), .Z(n11009) );
  NAND2_X1 U11264 ( .A1(n11162), .A2(n10725), .ZN(n11286) );
  MUX2_X1 U11265 ( .A(n11331), .B(n10648), .S(n11162), .Z(n10997) );
  OR2_X1 U11266 ( .A1(n11819), .A2(n11818), .ZN(n12810) );
  OR2_X1 U11267 ( .A1(n11803), .A2(n11802), .ZN(n12750) );
  AND2_X1 U11268 ( .A1(n13392), .A2(n20130), .ZN(n13204) );
  AOI211_X1 U11269 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n10112), .B(n10111), .ZN(n17434) );
  AND2_X2 U11270 ( .A1(n20109), .A2(n11757), .ZN(n13221) );
  NAND3_X2 U11271 ( .A1(n10075), .A2(n10155), .A3(n10154), .ZN(n17449) );
  AND4_X2 U11272 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n11587) );
  INV_X2 U11273 ( .A(n16494), .ZN(n16509) );
  NAND2_X2 U11274 ( .A1(n9589), .A2(n9590), .ZN(n20138) );
  CLKBUF_X3 U11275 ( .A(n10710), .Z(n21042) );
  INV_X1 U11276 ( .A(n11293), .ZN(n10714) );
  NAND2_X1 U11277 ( .A1(n10584), .A2(n10583), .ZN(n10713) );
  OR2_X1 U11278 ( .A1(n11709), .A2(n11708), .ZN(n11751) );
  NAND4_X1 U11279 ( .A1(n10082), .A2(n10081), .A3(n11662), .A4(n11661), .ZN(
        n11679) );
  NAND2_X2 U11280 ( .A1(n10455), .A2(n10454), .ZN(n10710) );
  AND4_X1 U11281 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11639) );
  AND4_X1 U11282 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11678) );
  AND4_X1 U11283 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n9589) );
  AND4_X1 U11284 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n10080) );
  NAND2_X1 U11285 ( .A1(n10545), .A2(n10544), .ZN(n11020) );
  INV_X4 U11286 ( .A(n10147), .ZN(n17244) );
  NAND2_X1 U11287 ( .A1(n10597), .A2(n10596), .ZN(n11293) );
  NOR2_X1 U11288 ( .A1(n9776), .A2(n9774), .ZN(n9773) );
  AND4_X1 U11289 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n9590) );
  NOR2_X1 U11290 ( .A1(n18868), .A2(n10084), .ZN(n10113) );
  AND3_X1 U11291 ( .A1(n9771), .A2(n11627), .A3(n9770), .ZN(n9775) );
  NAND2_X1 U11292 ( .A1(n9777), .A2(n9772), .ZN(n9774) );
  AND2_X2 U11293 ( .A1(n14096), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10850) );
  AND4_X1 U11294 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11749) );
  AND4_X1 U11295 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11748) );
  BUF_X2 U11296 ( .A(n11658), .Z(n12243) );
  NAND2_X2 U11297 ( .A1(n18925), .A2(n18789), .ZN(n18846) );
  NOR2_X1 U11298 ( .A1(n14016), .A2(n14015), .ZN(n10494) );
  AND2_X2 U11299 ( .A1(n10628), .A2(n16349), .ZN(n13907) );
  AND3_X1 U11300 ( .A1(n9671), .A2(n10490), .A3(n10489), .ZN(n10498) );
  AND2_X2 U11301 ( .A1(n9623), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10637) );
  INV_X2 U11302 ( .A(n16541), .ZN(U215) );
  INV_X2 U11303 ( .A(n12536), .ZN(n9585) );
  NAND2_X2 U11304 ( .A1(n19909), .A2(n19802), .ZN(n19857) );
  NOR2_X1 U11305 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16223), .ZN(n20044) );
  BUF_X4 U11306 ( .A(n10255), .Z(n9586) );
  INV_X2 U11308 ( .A(n12435), .ZN(n12543) );
  NAND2_X1 U11309 ( .A1(n16944), .A2(n9665), .ZN(n15688) );
  INV_X1 U11310 ( .A(n12482), .ZN(n9608) );
  AND2_X2 U11311 ( .A1(n11628), .A2(n13488), .ZN(n11828) );
  NAND2_X1 U11312 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18731) );
  INV_X2 U11313 ( .A(n16545), .ZN(n16547) );
  INV_X2 U11314 ( .A(n18926), .ZN(n18925) );
  OR2_X1 U11315 ( .A1(n10091), .A2(n10092), .ZN(n9652) );
  NOR2_X1 U11316 ( .A1(n10050), .A2(n18893), .ZN(n10093) );
  AND2_X2 U11317 ( .A1(n9609), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10855) );
  AND2_X1 U11318 ( .A1(n9998), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U11319 ( .A1(n18878), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10090) );
  AND2_X2 U11320 ( .A1(n13488), .A2(n13468), .ZN(n11665) );
  AND2_X1 U11321 ( .A1(n11902), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U11322 ( .A1(n9802), .A2(n11902), .ZN(n12482) );
  AND2_X2 U11323 ( .A1(n9787), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9727) );
  NAND2_X1 U11324 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18732) );
  NOR2_X4 U11325 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13781) );
  AND2_X1 U11326 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10522) );
  AND3_X1 U11327 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9802) );
  INV_X1 U11328 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14015) );
  INV_X1 U11329 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9786) );
  INV_X1 U11330 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9787) );
  INV_X1 U11331 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18885) );
  NAND4_X1 U11332 ( .A1(n9998), .A2(n11902), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12435) );
  INV_X1 U11333 ( .A(n10710), .ZN(n10711) );
  NOR2_X1 U11334 ( .A1(n10689), .A2(n10711), .ZN(n10690) );
  NAND2_X1 U11335 ( .A1(n10598), .A2(n10601), .ZN(n10691) );
  AND3_X2 U11336 ( .A1(n10718), .A2(n10430), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14099) );
  NOR2_X2 U11337 ( .A1(n20910), .A2(n17332), .ZN(n17327) );
  INV_X1 U11338 ( .A(n13054), .ZN(n9592) );
  NAND2_X1 U11339 ( .A1(n9593), .A2(n13055), .ZN(n13059) );
  NOR2_X1 U11340 ( .A1(n13057), .A2(n9592), .ZN(n9593) );
  AND2_X2 U11341 ( .A1(n12928), .A2(n10748), .ZN(n9594) );
  OR2_X1 U11342 ( .A1(n14871), .A2(n13965), .ZN(n9595) );
  NOR2_X1 U11343 ( .A1(n14857), .A2(n9599), .ZN(n9596) );
  INV_X1 U11344 ( .A(n14036), .ZN(n9598) );
  OR2_X1 U11345 ( .A1(n14859), .A2(n14036), .ZN(n9599) );
  NOR2_X1 U11347 ( .A1(n14858), .A2(n10064), .ZN(n14037) );
  NAND2_X1 U11348 ( .A1(n11281), .A2(n10722), .ZN(n10748) );
  AND2_X1 U11349 ( .A1(n10713), .A2(n11293), .ZN(n10601) );
  AND2_X1 U11350 ( .A1(n9602), .A2(n15537), .ZN(n9601) );
  NAND3_X1 U11351 ( .A1(n15229), .A2(n15538), .A3(n10926), .ZN(n9602) );
  NAND3_X1 U11352 ( .A1(n15229), .A2(n15538), .A3(n10926), .ZN(n9603) );
  NAND3_X1 U11353 ( .A1(n15229), .A2(n15538), .A3(n10926), .ZN(n15544) );
  NAND2_X2 U11354 ( .A1(n11756), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11854) );
  NAND2_X2 U11355 ( .A1(n11854), .A2(n11769), .ZN(n11865) );
  BUF_X1 U11356 ( .A(n11163), .Z(n9604) );
  NOR2_X1 U11357 ( .A1(n11572), .A2(n11580), .ZN(n9605) );
  OAI211_X1 U11358 ( .C1(n10763), .C2(n10456), .A(n10756), .B(n10755), .ZN(
        n9606) );
  INV_X1 U11359 ( .A(n11037), .ZN(n9607) );
  NOR2_X1 U11360 ( .A1(n11572), .A2(n11580), .ZN(n11153) );
  OAI211_X1 U11361 ( .C1(n10763), .C2(n10456), .A(n10756), .B(n10755), .ZN(
        n10761) );
  INV_X1 U11362 ( .A(n10704), .ZN(n10727) );
  NAND2_X2 U11363 ( .A1(n10747), .A2(n21040), .ZN(n12928) );
  INV_X2 U11364 ( .A(n10692), .ZN(n10747) );
  NAND2_X1 U11365 ( .A1(n11913), .A2(n20138), .ZN(n11763) );
  INV_X2 U11366 ( .A(n11679), .ZN(n11913) );
  OAI21_X1 U11367 ( .B1(n10928), .B2(n10927), .A(n9756), .ZN(n9754) );
  NAND2_X2 U11368 ( .A1(n10711), .A2(n10722), .ZN(n10725) );
  NOR2_X1 U11369 ( .A1(n14016), .A2(n10564), .ZN(n10565) );
  AND3_X2 U11370 ( .A1(n10718), .A2(n10430), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9609) );
  AND2_X1 U11371 ( .A1(n10747), .A2(n10736), .ZN(n10764) );
  NOR2_X2 U11372 ( .A1(n17521), .A2(n17323), .ZN(n17319) );
  BUF_X2 U11373 ( .A(n10240), .Z(n17303) );
  AOI211_X1 U11374 ( .C1(n10141), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n15694), .B(n15693), .ZN(n15695) );
  INV_X1 U11375 ( .A(n17137), .ZN(n9610) );
  INV_X1 U11376 ( .A(n17137), .ZN(n9611) );
  INV_X1 U11377 ( .A(n10086), .ZN(n9612) );
  INV_X4 U11378 ( .A(n10573), .ZN(n14096) );
  INV_X1 U11379 ( .A(n12431), .ZN(n9613) );
  INV_X1 U11380 ( .A(n12431), .ZN(n12545) );
  OR2_X4 U11381 ( .A1(n10805), .A2(n15566), .ZN(n10806) );
  INV_X1 U11382 ( .A(n12435), .ZN(n9614) );
  NAND2_X1 U11383 ( .A1(n10787), .A2(n10786), .ZN(n15566) );
  OR2_X1 U11384 ( .A1(n10791), .A2(n10786), .ZN(n10814) );
  AOI21_X2 U11385 ( .B1(n10774), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10759), .ZN(n10760) );
  NAND2_X2 U11386 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18893), .ZN(
        n10087) );
  INV_X1 U11387 ( .A(n11547), .ZN(n15018) );
  NOR2_X2 U11388 ( .A1(n13509), .A2(n13535), .ZN(n13536) );
  OR2_X1 U11389 ( .A1(n15077), .A2(n15076), .ZN(n15199) );
  NOR2_X2 U11390 ( .A1(n15077), .A2(n11097), .ZN(n11116) );
  NOR2_X2 U11391 ( .A1(n14869), .A2(n14872), .ZN(n14871) );
  XNOR2_X1 U11392 ( .A(n11905), .B(n12736), .ZN(n13503) );
  NAND2_X2 U11393 ( .A1(n12748), .A2(n12747), .ZN(n12757) );
  OR2_X1 U11394 ( .A1(n14570), .A2(n19920), .ZN(n12849) );
  NAND2_X2 U11395 ( .A1(n10003), .A2(n10004), .ZN(n15023) );
  XNOR2_X2 U11396 ( .A(n11912), .B(n11911), .ZN(n12741) );
  NAND3_X1 U11397 ( .A1(n18885), .A2(n18726), .A3(n10085), .ZN(n17249) );
  NOR2_X2 U11398 ( .A1(n10603), .A2(n10602), .ZN(n11281) );
  INV_X1 U11399 ( .A(n10113), .ZN(n10147) );
  BUF_X2 U11400 ( .A(n13052), .Z(n13738) );
  AND2_X1 U11401 ( .A1(n11628), .A2(n13488), .ZN(n9617) );
  INV_X2 U11402 ( .A(n11020), .ZN(n10599) );
  INV_X1 U11403 ( .A(n10551), .ZN(n9620) );
  INV_X2 U11404 ( .A(n9620), .ZN(n9621) );
  NOR2_X2 U11405 ( .A1(n13215), .A2(n13387), .ZN(n13413) );
  AOI21_X2 U11406 ( .B1(n15955), .B2(n14534), .A(n14421), .ZN(n14433) );
  XNOR2_X2 U11407 ( .A(n12763), .B(n13541), .ZN(n13525) );
  INV_X1 U11408 ( .A(n17249), .ZN(n17226) );
  OAI21_X2 U11409 ( .B1(n15065), .B2(n15066), .A(n15067), .ZN(n15058) );
  AOI21_X2 U11410 ( .B1(n11116), .B2(n11115), .A(n11114), .ZN(n15065) );
  XNOR2_X2 U11411 ( .A(n11027), .B(n11026), .ZN(n15535) );
  OR2_X1 U11412 ( .A1(n10394), .A2(n17497), .ZN(n9761) );
  OAI21_X2 U11413 ( .B1(n15827), .B2(n15826), .A(n18910), .ZN(n15828) );
  NOR3_X4 U11414 ( .A1(n16555), .A2(n18912), .A3(n15733), .ZN(n15827) );
  AND2_X2 U11415 ( .A1(n14896), .A2(n13861), .ZN(n14882) );
  NOR2_X2 U11416 ( .A1(n14895), .A2(n14898), .ZN(n14896) );
  NOR2_X4 U11417 ( .A1(n15044), .A2(n11491), .ZN(n15033) );
  NAND2_X2 U11418 ( .A1(n15103), .A2(n9725), .ZN(n15044) );
  XNOR2_X2 U11419 ( .A(n14011), .B(n10076), .ZN(n14857) );
  NAND2_X2 U11420 ( .A1(n13788), .A2(n9858), .ZN(n15130) );
  NAND2_X2 U11421 ( .A1(n10992), .A2(n10991), .ZN(n13788) );
  NAND2_X1 U11422 ( .A1(n9941), .A2(n10772), .ZN(n11163) );
  NAND2_X2 U11423 ( .A1(n10513), .A2(n10512), .ZN(n10704) );
  XNOR2_X2 U11424 ( .A(n9742), .B(n10878), .ZN(n13815) );
  NAND2_X1 U11425 ( .A1(n13120), .A2(n10717), .ZN(n9624) );
  NAND2_X1 U11426 ( .A1(n13120), .A2(n10717), .ZN(n11562) );
  AND2_X1 U11427 ( .A1(n9609), .A2(n16349), .ZN(n9625) );
  INV_X1 U11428 ( .A(n19913), .ZN(n13399) );
  OR2_X1 U11429 ( .A1(n10675), .A2(n10674), .ZN(n10877) );
  NOR2_X1 U11430 ( .A1(n21042), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11313) );
  AOI21_X1 U11431 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19874), .A(
        n10477), .ZN(n10482) );
  NOR2_X1 U11432 ( .A1(n10476), .A2(n10478), .ZN(n10477) );
  NOR2_X1 U11433 ( .A1(n20134), .A2(n20138), .ZN(n12854) );
  AND2_X1 U11434 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  INV_X1 U11435 ( .A(n14294), .ZN(n10026) );
  AND2_X1 U11436 ( .A1(n9684), .A2(n9953), .ZN(n9952) );
  INV_X1 U11437 ( .A(n13762), .ZN(n9953) );
  NAND2_X1 U11438 ( .A1(n13412), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12804) );
  CLKBUF_X1 U11439 ( .A(n11020), .Z(n11021) );
  NOR3_X1 U11440 ( .A1(n13964), .A2(n13963), .A3(n14874), .ZN(n13965) );
  OAI21_X1 U11441 ( .B1(n10010), .B2(n10037), .A(n10007), .ZN(n10006) );
  NAND2_X1 U11442 ( .A1(n9965), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9964) );
  NAND2_X1 U11443 ( .A1(n9967), .A2(n16349), .ZN(n9966) );
  INV_X1 U11444 ( .A(n16944), .ZN(n10092) );
  NAND2_X1 U11445 ( .A1(n18885), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10050) );
  AND2_X1 U11446 ( .A1(n10421), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9912) );
  NAND2_X1 U11447 ( .A1(n9761), .A2(n9760), .ZN(n9759) );
  INV_X1 U11448 ( .A(n18929), .ZN(n9760) );
  INV_X1 U11449 ( .A(n9759), .ZN(n16576) );
  INV_X1 U11450 ( .A(n11751), .ZN(n13810) );
  AND2_X1 U11451 ( .A1(n12525), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12526) );
  NAND2_X1 U11452 ( .A1(n12526), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12619) );
  INV_X1 U11453 ( .A(n13221), .ZN(n13101) );
  NAND2_X1 U11454 ( .A1(n9996), .A2(n14522), .ZN(n9814) );
  AOI21_X1 U11455 ( .B1(n12827), .B2(n14579), .A(n9997), .ZN(n9996) );
  INV_X1 U11456 ( .A(n9993), .ZN(n9992) );
  OAI21_X1 U11457 ( .B1(n9997), .B2(n14579), .A(n9656), .ZN(n9993) );
  AND2_X1 U11458 ( .A1(n13400), .A2(n13399), .ZN(n13416) );
  NAND2_X1 U11459 ( .A1(n9796), .A2(n9795), .ZN(n13398) );
  INV_X1 U11460 ( .A(n13390), .ZN(n13395) );
  AND2_X1 U11461 ( .A1(n9615), .A2(n12741), .ZN(n20632) );
  INV_X1 U11462 ( .A(n13692), .ZN(n9973) );
  NOR2_X1 U11463 ( .A1(n14649), .A2(n14703), .ZN(n11539) );
  OAI21_X1 U11464 ( .B1(n11579), .B2(n11580), .A(n10000), .ZN(n11617) );
  INV_X1 U11465 ( .A(n10001), .ZN(n10000) );
  OAI21_X1 U11466 ( .B1(n11578), .B2(n11580), .A(n15012), .ZN(n10001) );
  INV_X1 U11467 ( .A(n14837), .ZN(n9938) );
  AND2_X1 U11468 ( .A1(n11532), .A2(n11271), .ZN(n14699) );
  AND4_X1 U11469 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        n10979) );
  AND4_X1 U11470 ( .A1(n10966), .A2(n10965), .A3(n10964), .A4(n10963), .ZN(
        n10982) );
  INV_X1 U11471 ( .A(n13060), .ZN(n13117) );
  NAND2_X1 U11472 ( .A1(n12973), .A2(n19678), .ZN(n13155) );
  AND2_X1 U11473 ( .A1(n21039), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13150) );
  XNOR2_X1 U11474 ( .A(n13060), .B(n13061), .ZN(n12980) );
  AOI21_X1 U11475 ( .B1(n15738), .B2(n15737), .A(n15631), .ZN(n15825) );
  AND2_X1 U11476 ( .A1(n10420), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16410) );
  NOR2_X1 U11477 ( .A1(n16414), .A2(n16617), .ZN(n10420) );
  OR2_X1 U11478 ( .A1(n10207), .A2(n18165), .ZN(n17792) );
  INV_X1 U11479 ( .A(n18705), .ZN(n18104) );
  NOR2_X1 U11480 ( .A1(n10389), .A2(n10328), .ZN(n15734) );
  NAND2_X1 U11481 ( .A1(n18763), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18750) );
  NAND2_X1 U11482 ( .A1(n11501), .A2(n19777), .ZN(n12941) );
  INV_X1 U11483 ( .A(n14131), .ZN(n9962) );
  NAND2_X1 U11484 ( .A1(n14128), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14129) );
  INV_X1 U11485 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19900) );
  INV_X1 U11486 ( .A(n17708), .ZN(n17723) );
  INV_X1 U11487 ( .A(n12582), .ZN(n12594) );
  NAND2_X1 U11488 ( .A1(n11634), .A2(n13488), .ZN(n12431) );
  NAND2_X1 U11489 ( .A1(n12569), .A2(n12568), .ZN(n12573) );
  OR2_X1 U11490 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20103), .ZN(
        n12572) );
  NAND2_X1 U11491 ( .A1(n9794), .A2(n9793), .ZN(n9792) );
  NAND2_X1 U11492 ( .A1(n12604), .A2(n12605), .ZN(n9793) );
  NAND2_X1 U11493 ( .A1(n12603), .A2(n12602), .ZN(n9794) );
  NAND2_X1 U11494 ( .A1(n12606), .A2(n12605), .ZN(n9791) );
  NAND2_X1 U11495 ( .A1(n20777), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9789) );
  NAND2_X1 U11496 ( .A1(n11766), .A2(n11774), .ZN(n9734) );
  NAND2_X1 U11497 ( .A1(n13209), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11929) );
  NOR2_X1 U11498 ( .A1(n16284), .A2(n16282), .ZN(n11047) );
  INV_X1 U11499 ( .A(n15515), .ZN(n9756) );
  NAND2_X1 U11500 ( .A1(n16381), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10755) );
  OR2_X1 U11501 ( .A1(n10660), .A2(n10659), .ZN(n11335) );
  AND2_X1 U11502 ( .A1(n10727), .A2(n10726), .ZN(n10728) );
  AOI21_X1 U11503 ( .B1(n11284), .B2(n11293), .A(n10696), .ZN(n10697) );
  MUX2_X1 U11504 ( .A(n10727), .B(n10599), .S(n10703), .Z(n10698) );
  NAND2_X1 U11505 ( .A1(n11314), .A2(n10727), .ZN(n10610) );
  INV_X1 U11506 ( .A(n10199), .ZN(n10035) );
  NAND2_X1 U11507 ( .A1(n12844), .A2(n10032), .ZN(n10031) );
  INV_X1 U11508 ( .A(n14153), .ZN(n10032) );
  AND2_X1 U11509 ( .A1(n12324), .A2(n14315), .ZN(n10027) );
  OR2_X1 U11510 ( .A1(n14347), .A2(n14337), .ZN(n10016) );
  AND2_X1 U11511 ( .A1(n14240), .A2(n14353), .ZN(n12155) );
  INV_X1 U11512 ( .A(n13678), .ZN(n10019) );
  NAND2_X1 U11513 ( .A1(n20856), .A2(n20857), .ZN(n12559) );
  NAND2_X1 U11514 ( .A1(n11929), .A2(n12804), .ZN(n12583) );
  INV_X1 U11515 ( .A(n14169), .ZN(n9961) );
  OR2_X1 U11516 ( .A1(n14197), .A2(n14180), .ZN(n9959) );
  NAND2_X1 U11517 ( .A1(n9957), .A2(n14339), .ZN(n9956) );
  NOR2_X1 U11518 ( .A1(n14342), .A2(n14224), .ZN(n9957) );
  NAND2_X1 U11519 ( .A1(n9806), .A2(n9805), .ZN(n14489) );
  INV_X1 U11520 ( .A(n14497), .ZN(n9806) );
  NAND2_X1 U11521 ( .A1(n14519), .A2(n12819), .ZN(n9805) );
  OR2_X1 U11522 ( .A1(n12736), .A2(n13410), .ZN(n12740) );
  NAND2_X1 U11523 ( .A1(n11827), .A2(n11826), .ZN(n11849) );
  OAI21_X1 U11524 ( .B1(n11915), .B2(n9809), .A(n9670), .ZN(n11827) );
  INV_X1 U11525 ( .A(n11822), .ZN(n9809) );
  AND2_X2 U11526 ( .A1(n13468), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13476) );
  NAND2_X1 U11527 ( .A1(n11913), .A2(n20134), .ZN(n11680) );
  OAI21_X1 U11528 ( .B1(n16227), .B2(n13498), .A(n14639), .ZN(n20108) );
  INV_X1 U11529 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20476) );
  INV_X1 U11530 ( .A(n11582), .ZN(n11584) );
  AND2_X1 U11531 ( .A1(n11133), .A2(n14715), .ZN(n11147) );
  NOR2_X1 U11532 ( .A1(n11069), .A2(n11064), .ZN(n11065) );
  OR2_X1 U11533 ( .A1(n11072), .A2(n11067), .ZN(n11069) );
  NAND2_X1 U11534 ( .A1(n11074), .A2(n11130), .ZN(n11071) );
  NAND2_X1 U11535 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  NAND2_X1 U11536 ( .A1(n11085), .A2(n11058), .ZN(n9917) );
  NAND2_X1 U11537 ( .A1(n11056), .A2(n13591), .ZN(n11082) );
  NAND3_X1 U11538 ( .A1(n10763), .A2(n10753), .A3(n10752), .ZN(n10778) );
  NAND2_X1 U11539 ( .A1(n10774), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10752) );
  NOR2_X1 U11540 ( .A1(n9980), .A2(n9981), .ZN(n9979) );
  INV_X1 U11541 ( .A(n14917), .ZN(n9980) );
  INV_X1 U11542 ( .A(n13192), .ZN(n14034) );
  AND2_X1 U11543 ( .A1(n13935), .A2(n13934), .ZN(n13961) );
  INV_X1 U11544 ( .A(n16246), .ZN(n10061) );
  AND2_X1 U11545 ( .A1(n15504), .A2(n9697), .ZN(n15461) );
  INV_X1 U11546 ( .A(n15490), .ZN(n9982) );
  AND2_X1 U11547 ( .A1(n9686), .A2(n13796), .ZN(n9983) );
  NOR2_X1 U11548 ( .A1(n10918), .A2(n10917), .ZN(n11347) );
  NAND3_X1 U11549 ( .A1(n10609), .A2(n21042), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n13192) );
  NAND2_X1 U11550 ( .A1(n10714), .A2(n10713), .ZN(n10731) );
  NOR2_X1 U11551 ( .A1(n13803), .A2(n9856), .ZN(n9855) );
  INV_X1 U11552 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9856) );
  AND2_X1 U11553 ( .A1(n14737), .A2(n11139), .ZN(n11143) );
  INV_X1 U11554 ( .A(n14768), .ZN(n9975) );
  AND2_X1 U11555 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  INV_X1 U11556 ( .A(n14887), .ZN(n9944) );
  AND2_X1 U11557 ( .A1(n15133), .A2(n14892), .ZN(n9945) );
  INV_X1 U11558 ( .A(n15140), .ZN(n9877) );
  NOR2_X1 U11559 ( .A1(n9878), .A2(n9877), .ZN(n9876) );
  NOR2_X1 U11560 ( .A1(n9884), .A2(n15147), .ZN(n9882) );
  INV_X1 U11561 ( .A(n9871), .ZN(n9870) );
  OAI21_X1 U11562 ( .B1(n9872), .B2(n11047), .A(n10010), .ZN(n9871) );
  INV_X1 U11563 ( .A(n13790), .ZN(n10009) );
  NAND2_X1 U11564 ( .A1(n9757), .A2(n9755), .ZN(n10984) );
  AND2_X1 U11565 ( .A1(n10921), .A2(n15515), .ZN(n9755) );
  INV_X1 U11566 ( .A(n10928), .ZN(n9757) );
  NAND2_X1 U11567 ( .A1(n10984), .A2(n9754), .ZN(n11033) );
  AOI21_X1 U11568 ( .B1(n11206), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10777), .ZN(n11165) );
  INV_X1 U11569 ( .A(n13688), .ZN(n9934) );
  NOR2_X1 U11570 ( .A1(n9866), .A2(n11596), .ZN(n9863) );
  NOR2_X1 U11571 ( .A1(n13817), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9866) );
  AND4_X1 U11572 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(
        n10981) );
  NOR2_X2 U11573 ( .A1(n11010), .A2(n11009), .ZN(n11008) );
  AOI21_X1 U11574 ( .B1(n13155), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n15622), .ZN(n13156) );
  NAND2_X1 U11575 ( .A1(n13151), .A2(n13150), .ZN(n10053) );
  AND2_X1 U11576 ( .A1(n10522), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13178) );
  NAND2_X1 U11577 ( .A1(n10487), .A2(n21042), .ZN(n13071) );
  INV_X1 U11578 ( .A(n10815), .ZN(n10818) );
  NAND2_X1 U11579 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10499) );
  NOR2_X1 U11580 ( .A1(n10509), .A2(n10508), .ZN(n10510) );
  INV_X1 U11581 ( .A(n19894), .ZN(n19277) );
  AND2_X1 U11582 ( .A1(n10609), .A2(n10704), .ZN(n10600) );
  NOR3_X1 U11583 ( .A1(n18868), .A2(n18878), .A3(n10087), .ZN(n10086) );
  NAND2_X1 U11584 ( .A1(n18868), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10091) );
  AND2_X1 U11585 ( .A1(n10139), .A2(n10138), .ZN(n10140) );
  NAND2_X1 U11586 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n9835) );
  NOR2_X1 U11587 ( .A1(n17434), .A2(n10196), .ZN(n10201) );
  NOR2_X1 U11588 ( .A1(n17878), .A2(n10195), .ZN(n10198) );
  XNOR2_X1 U11589 ( .A(n9833), .B(n17449), .ZN(n10188) );
  AOI21_X1 U11590 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(n10349) );
  NOR2_X1 U11591 ( .A1(n10392), .A2(n10396), .ZN(n10394) );
  OAI21_X1 U11592 ( .B1(n10147), .B2(n18593), .A(n9765), .ZN(n9764) );
  AOI21_X1 U11593 ( .B1(n10247), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(n9766), .ZN(n9765) );
  NOR2_X1 U11594 ( .A1(n9616), .A2(n10308), .ZN(n9766) );
  INV_X1 U11595 ( .A(n10306), .ZN(n9767) );
  INV_X1 U11596 ( .A(n10313), .ZN(n9763) );
  AOI22_X1 U11597 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10313) );
  NOR2_X1 U11598 ( .A1(n14152), .A2(n10028), .ZN(n12850) );
  NAND2_X1 U11599 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  INV_X1 U11600 ( .A(n10031), .ZN(n10030) );
  INV_X1 U11601 ( .A(n12851), .ZN(n10029) );
  INV_X1 U11602 ( .A(n13356), .ZN(n11922) );
  INV_X1 U11603 ( .A(n14339), .ZN(n9955) );
  INV_X1 U11604 ( .A(n9721), .ZN(n9951) );
  NAND2_X1 U11605 ( .A1(n9737), .A2(n9735), .ZN(n9738) );
  NAND2_X1 U11606 ( .A1(n16188), .A2(n9684), .ZN(n16160) );
  NAND2_X1 U11607 ( .A1(n16188), .A2(n13700), .ZN(n16162) );
  OAI21_X1 U11608 ( .B1(n13363), .B2(n9731), .A(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9730) );
  NOR2_X1 U11609 ( .A1(n12759), .A2(n13575), .ZN(n20528) );
  INV_X1 U11610 ( .A(n12749), .ZN(n13575) );
  NOR2_X1 U11611 ( .A1(n20421), .A2(n20279), .ZN(n20650) );
  NAND2_X1 U11612 ( .A1(n11584), .A2(n11583), .ZN(n11592) );
  NAND2_X1 U11613 ( .A1(n14672), .A2(n9837), .ZN(n9839) );
  INV_X1 U11614 ( .A(n14702), .ZN(n9838) );
  AND2_X1 U11615 ( .A1(n11118), .A2(n9924), .ZN(n11133) );
  NOR2_X1 U11616 ( .A1(n9925), .A2(n9926), .ZN(n9924) );
  NAND2_X1 U11617 ( .A1(n9928), .A2(n9927), .ZN(n9926) );
  NOR2_X1 U11618 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n9927) );
  INV_X1 U11619 ( .A(n14672), .ZN(n14714) );
  OR2_X1 U11620 ( .A1(n14714), .A2(n15029), .ZN(n9840) );
  OR2_X1 U11621 ( .A1(n10678), .A2(n10519), .ZN(n12930) );
  AND2_X1 U11622 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NOR2_X1 U11623 ( .A1(n13829), .A2(n13521), .ZN(n10060) );
  NAND2_X1 U11624 ( .A1(n9676), .A2(n13828), .ZN(n13829) );
  OR2_X1 U11625 ( .A1(n11367), .A2(n11366), .ZN(n13519) );
  NAND2_X1 U11626 ( .A1(n9626), .A2(n14039), .ZN(n10057) );
  AND2_X1 U11627 ( .A1(n11471), .A2(n11470), .ZN(n14790) );
  NAND2_X1 U11628 ( .A1(n14806), .A2(n9693), .ZN(n15332) );
  INV_X1 U11629 ( .A(n15329), .ZN(n9986) );
  NOR2_X1 U11630 ( .A1(n15332), .A2(n14790), .ZN(n14789) );
  INV_X1 U11631 ( .A(n11334), .ZN(n9968) );
  AND2_X1 U11632 ( .A1(n13189), .A2(n13188), .ZN(n13190) );
  OR2_X1 U11633 ( .A1(n14651), .A2(n15026), .ZN(n14649) );
  NAND2_X1 U11634 ( .A1(n14669), .A2(n9846), .ZN(n14651) );
  AND2_X1 U11635 ( .A1(n9642), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9846) );
  NAND2_X1 U11636 ( .A1(n14669), .A2(n9642), .ZN(n14671) );
  NOR2_X1 U11637 ( .A1(n14656), .A2(n14654), .ZN(n14658) );
  NAND2_X1 U11638 ( .A1(n11586), .A2(n9932), .ZN(n11619) );
  NOR2_X1 U11639 ( .A1(n11587), .A2(n11613), .ZN(n9932) );
  AND2_X1 U11640 ( .A1(n9648), .A2(n10048), .ZN(n10047) );
  AND2_X1 U11641 ( .A1(n9707), .A2(n9936), .ZN(n9935) );
  INV_X1 U11642 ( .A(n14740), .ZN(n9936) );
  NOR2_X1 U11643 ( .A1(n15333), .A2(n11490), .ZN(n15306) );
  AOI21_X1 U11644 ( .B1(n9882), .B2(n9886), .A(n9879), .ZN(n9878) );
  INV_X1 U11645 ( .A(n15084), .ZN(n9879) );
  INV_X1 U11646 ( .A(n9882), .ZN(n9880) );
  AND2_X1 U11647 ( .A1(n9646), .A2(n10993), .ZN(n9858) );
  OAI21_X1 U11648 ( .B1(n9886), .B2(n15172), .A(n15163), .ZN(n9884) );
  OR2_X1 U11649 ( .A1(n11108), .A2(n15414), .ZN(n15173) );
  AND3_X1 U11650 ( .A1(n11344), .A2(n11343), .A3(n11342), .ZN(n13692) );
  NAND2_X1 U11651 ( .A1(n9972), .A2(n9703), .ZN(n13690) );
  AOI21_X1 U11652 ( .B1(n15566), .B2(n13150), .A(n12976), .ZN(n12979) );
  NOR2_X1 U11653 ( .A1(n19871), .A2(n19277), .ZN(n19462) );
  INV_X1 U11654 ( .A(n19720), .ZN(n19495) );
  NAND2_X1 U11655 ( .A1(n19871), .A2(n19894), .ZN(n19674) );
  NAND2_X1 U11656 ( .A1(n11503), .A2(n11502), .ZN(n19726) );
  NAND2_X1 U11657 ( .A1(n15594), .A2(n21039), .ZN(n11503) );
  NAND2_X1 U11658 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19726), .ZN(n19308) );
  NAND2_X1 U11659 ( .A1(n10348), .A2(n10350), .ZN(n18706) );
  NOR2_X1 U11660 ( .A1(n16615), .A2(n16616), .ZN(n16614) );
  OR2_X1 U11661 ( .A1(n16949), .A2(n17625), .ZN(n9902) );
  OR2_X1 U11662 ( .A1(n16693), .A2(n9903), .ZN(n9901) );
  OR2_X1 U11663 ( .A1(n17625), .A2(n17638), .ZN(n9903) );
  OR2_X1 U11664 ( .A1(n16693), .A2(n17638), .ZN(n9904) );
  NAND2_X1 U11665 ( .A1(n16723), .A2(n9892), .ZN(n9891) );
  INV_X1 U11666 ( .A(n17669), .ZN(n9892) );
  OR2_X1 U11667 ( .A1(n9893), .A2(n9891), .ZN(n9889) );
  NAND2_X1 U11668 ( .A1(n18914), .A2(n18269), .ZN(n16581) );
  NAND2_X1 U11669 ( .A1(n17271), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17242) );
  INV_X1 U11670 ( .A(n18291), .ZN(n17307) );
  INV_X1 U11671 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17050) );
  NOR2_X1 U11672 ( .A1(n18868), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10085) );
  NAND2_X1 U11673 ( .A1(n9820), .A2(n16944), .ZN(n17156) );
  INV_X1 U11674 ( .A(n10090), .ZN(n9820) );
  OAI21_X1 U11675 ( .B1(n10102), .B2(n17106), .A(n10151), .ZN(n10152) );
  NAND2_X1 U11676 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10151) );
  NOR2_X1 U11677 ( .A1(n10042), .A2(n10040), .ZN(n10039) );
  NAND2_X1 U11678 ( .A1(n16576), .A2(n16577), .ZN(n17457) );
  INV_X1 U11679 ( .A(n17564), .ZN(n9911) );
  AND2_X1 U11680 ( .A1(n17622), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17582) );
  NAND3_X1 U11681 ( .A1(n17731), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17679) );
  NOR2_X1 U11682 ( .A1(n16429), .A2(n9832), .ZN(n15744) );
  NAND2_X1 U11683 ( .A1(n16432), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9832) );
  AND2_X1 U11684 ( .A1(n10211), .A2(n9678), .ZN(n9825) );
  INV_X1 U11685 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U11686 ( .A1(n9827), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9826) );
  NAND2_X1 U11687 ( .A1(n10402), .A2(n10401), .ZN(n15732) );
  NAND2_X1 U11688 ( .A1(n9822), .A2(n9821), .ZN(n10045) );
  AOI21_X1 U11689 ( .B1(n10206), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n17729), .ZN(n9821) );
  NAND2_X1 U11690 ( .A1(n17844), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9822) );
  AND2_X1 U11691 ( .A1(n17792), .A2(n17724), .ZN(n17832) );
  XNOR2_X1 U11692 ( .A(n10198), .B(n10197), .ZN(n17860) );
  NOR2_X1 U11693 ( .A1(n17860), .A2(n17861), .ZN(n17859) );
  NOR2_X1 U11694 ( .A1(n10350), .A2(n10349), .ZN(n16555) );
  INV_X1 U11695 ( .A(n18706), .ZN(n15737) );
  NOR2_X1 U11696 ( .A1(n17303), .A2(n10351), .ZN(n10355) );
  INV_X1 U11697 ( .A(n17449), .ZN(n10365) );
  INV_X1 U11698 ( .A(n18917), .ZN(n18277) );
  AND2_X1 U11699 ( .A1(n13601), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13602) );
  INV_X1 U11700 ( .A(n19994), .ZN(n19962) );
  AND2_X2 U11701 ( .A1(n12856), .A2(n13399), .ZN(n20014) );
  AND2_X1 U11702 ( .A1(n14405), .A2(n13425), .ZN(n14409) );
  AND2_X1 U11703 ( .A1(n12619), .A2(n12528), .ZN(n14145) );
  OR2_X1 U11704 ( .A1(n20087), .A2(n12837), .ZN(n16033) );
  AND2_X1 U11705 ( .A1(n16033), .A2(n20084), .ZN(n16027) );
  AOI21_X1 U11706 ( .B1(n13813), .B2(n12624), .A(n9948), .ZN(n9947) );
  NOR2_X1 U11707 ( .A1(n13813), .A2(n9949), .ZN(n9948) );
  XNOR2_X1 U11708 ( .A(n12874), .B(n12873), .ZN(n14549) );
  NAND2_X1 U11709 ( .A1(n14567), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14551) );
  XNOR2_X1 U11710 ( .A(n9779), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14559) );
  NAND2_X1 U11711 ( .A1(n16047), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16035) );
  NOR2_X1 U11712 ( .A1(n16041), .A2(n16159), .ZN(n9811) );
  XNOR2_X1 U11713 ( .A(n14437), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16038) );
  AND2_X1 U11714 ( .A1(n13416), .A2(n13415), .ZN(n20093) );
  NAND2_X1 U11715 ( .A1(n9807), .A2(n11822), .ZN(n11912) );
  INV_X1 U11716 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20560) );
  CLKBUF_X1 U11717 ( .A(n13458), .Z(n20564) );
  INV_X1 U11718 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20559) );
  INV_X1 U11719 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20857) );
  INV_X1 U11720 ( .A(n19887), .ZN(n19278) );
  AOI21_X1 U11721 ( .B1(n14699), .B2(n16311), .A(n11542), .ZN(n11543) );
  INV_X1 U11722 ( .A(n16293), .ZN(n16306) );
  XNOR2_X1 U11723 ( .A(n11599), .B(n11598), .ZN(n9913) );
  AOI21_X1 U11724 ( .B1(n14686), .B2(n19261), .A(n15002), .ZN(n11612) );
  NOR2_X1 U11725 ( .A1(n11533), .A2(n10065), .ZN(n11534) );
  NAND2_X1 U11726 ( .A1(n11308), .A2(n11278), .ZN(n19257) );
  INV_X1 U11727 ( .A(n16338), .ZN(n19259) );
  AND2_X1 U11728 ( .A1(n11308), .A2(n19905), .ZN(n16338) );
  INV_X1 U11729 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19874) );
  NAND2_X1 U11730 ( .A1(n13673), .A2(n13150), .ZN(n12978) );
  AND2_X1 U11731 ( .A1(n19494), .A2(n19865), .ZN(n19429) );
  OR2_X1 U11732 ( .A1(n16614), .A2(n16918), .ZN(n9910) );
  NAND2_X1 U11733 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  INV_X1 U11734 ( .A(n16600), .ZN(n9907) );
  NAND2_X1 U11735 ( .A1(n16611), .A2(n16976), .ZN(n9908) );
  INV_X1 U11736 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17678) );
  INV_X1 U11737 ( .A(n16900), .ZN(n16947) );
  NOR2_X2 U11738 ( .A1(n17202), .A2(n15634), .ZN(n17170) );
  INV_X1 U11739 ( .A(n18299), .ZN(n17425) );
  NOR2_X1 U11740 ( .A1(n17342), .A2(n18299), .ZN(n17338) );
  NAND2_X1 U11741 ( .A1(n17338), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17337) );
  INV_X1 U11742 ( .A(n17837), .ZN(n17791) );
  NAND2_X1 U11743 ( .A1(n16410), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9899) );
  AND3_X1 U11744 ( .A1(n17635), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17622) );
  INV_X1 U11745 ( .A(n17834), .ZN(n17807) );
  INV_X1 U11746 ( .A(n12883), .ZN(n17820) );
  NOR2_X2 U11747 ( .A1(n17925), .A2(n17427), .ZN(n17834) );
  INV_X1 U11748 ( .A(n17915), .ZN(n17925) );
  OAI21_X1 U11749 ( .B1(n18032), .B2(n18031), .A(n18238), .ZN(n18156) );
  INV_X1 U11750 ( .A(n18210), .ZN(n18250) );
  INV_X1 U11751 ( .A(n12583), .ZN(n12601) );
  NAND2_X1 U11752 ( .A1(n9800), .A2(n9799), .ZN(n12582) );
  NAND2_X1 U11753 ( .A1(n12585), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U11754 ( .A1(n12583), .A2(n11757), .ZN(n9800) );
  AND3_X1 U11755 ( .A1(n11284), .A2(n10711), .A3(n10722), .ZN(n10699) );
  OAI21_X1 U11756 ( .B1(n10884), .B2(n10799), .A(n9743), .ZN(n10800) );
  NAND2_X1 U11757 ( .A1(n10798), .A2(n9744), .ZN(n9743) );
  XNOR2_X1 U11758 ( .A(n16349), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10478) );
  AOI22_X1 U11759 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10539) );
  OR2_X1 U11760 ( .A1(n12022), .A2(n12021), .ZN(n12796) );
  INV_X1 U11761 ( .A(n20138), .ZN(n12585) );
  NAND2_X1 U11762 ( .A1(n11822), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U11763 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U11764 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9771) );
  NAND2_X1 U11765 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9772) );
  NAND2_X1 U11766 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n9777) );
  OR2_X1 U11767 ( .A1(n11571), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10083) );
  INV_X1 U11768 ( .A(n15207), .ZN(n10007) );
  AND2_X1 U11769 ( .A1(n15481), .A2(n15479), .ZN(n10010) );
  AND2_X1 U11770 ( .A1(n19408), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U11771 ( .A1(n10798), .A2(n9631), .ZN(n10841) );
  OAI22_X1 U11772 ( .A1(n10810), .A2(n19724), .B1(n10896), .B2(n14001), .ZN(
        n10811) );
  AOI22_X1 U11773 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U11774 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10445) );
  AND2_X1 U11775 ( .A1(n10676), .A2(n10661), .ZN(n10515) );
  AOI22_X1 U11776 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U11777 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10548) );
  NOR2_X1 U11778 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18893), .ZN(
        n10335) );
  OR2_X1 U11779 ( .A1(n10322), .A2(n10317), .ZN(n10321) );
  NOR2_X1 U11780 ( .A1(n12320), .A2(n15867), .ZN(n12321) );
  INV_X1 U11781 ( .A(n12764), .ZN(n9990) );
  AND2_X1 U11782 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11949) );
  AND2_X1 U11783 ( .A1(n12192), .A2(n11924), .ZN(n10023) );
  NAND2_X1 U11784 ( .A1(n9732), .A2(n12834), .ZN(n12890) );
  AND2_X1 U11785 ( .A1(n12571), .A2(n12572), .ZN(n12581) );
  OR2_X1 U11786 ( .A1(n12573), .A2(n12570), .ZN(n12571) );
  AOI21_X1 U11787 ( .B1(n9790), .B2(n9688), .A(n9788), .ZN(n12612) );
  OAI21_X1 U11788 ( .B1(n12611), .B2(n12610), .A(n9789), .ZN(n9788) );
  NAND2_X1 U11789 ( .A1(n9792), .A2(n9791), .ZN(n9790) );
  INV_X1 U11790 ( .A(n12815), .ZN(n9997) );
  INV_X1 U11791 ( .A(n12802), .ZN(n9736) );
  INV_X1 U11792 ( .A(n16163), .ZN(n9954) );
  XNOR2_X1 U11793 ( .A(n12807), .B(n12034), .ZN(n12795) );
  NAND2_X1 U11794 ( .A1(n12624), .A2(n13221), .ZN(n12711) );
  OR2_X1 U11795 ( .A1(n11944), .A2(n11943), .ZN(n12766) );
  NOR2_X1 U11796 ( .A1(n11891), .A2(n11890), .ZN(n12752) );
  INV_X1 U11797 ( .A(n20134), .ZN(n11764) );
  NAND2_X1 U11798 ( .A1(n13390), .A2(n13391), .ZN(n9797) );
  NAND2_X1 U11799 ( .A1(n13393), .A2(n20126), .ZN(n9795) );
  INV_X1 U11800 ( .A(n11773), .ZN(n13208) );
  AND2_X1 U11801 ( .A1(n20138), .A2(n11757), .ZN(n12803) );
  AND3_X1 U11802 ( .A1(n20134), .A2(n20109), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12609) );
  INV_X1 U11803 ( .A(n12804), .ZN(n11860) );
  OR2_X1 U11804 ( .A1(n11844), .A2(n11843), .ZN(n12751) );
  OAI21_X1 U11805 ( .B1(n11905), .B2(n12736), .A(n11862), .ZN(n11897) );
  NOR2_X1 U11806 ( .A1(n11833), .A2(n11732), .ZN(n11733) );
  INV_X1 U11807 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11732) );
  NOR2_X1 U11808 ( .A1(n10073), .A2(n11641), .ZN(n11645) );
  OAI21_X1 U11809 ( .B1(n11782), .B2(n12481), .A(n11640), .ZN(n11641) );
  AOI22_X1 U11810 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11649) );
  NOR2_X1 U11811 ( .A1(n14702), .A2(n15029), .ZN(n9837) );
  INV_X1 U11812 ( .A(n11121), .ZN(n9928) );
  INV_X1 U11813 ( .A(n9917), .ZN(n9914) );
  NOR2_X1 U11814 ( .A1(n9918), .A2(n9916), .ZN(n11086) );
  INV_X1 U11815 ( .A(n11058), .ZN(n9916) );
  NOR2_X1 U11816 ( .A1(n11042), .A2(n9920), .ZN(n9919) );
  INV_X1 U11817 ( .A(n9922), .ZN(n9920) );
  INV_X1 U11818 ( .A(n11023), .ZN(n9921) );
  NOR2_X1 U11819 ( .A1(n11022), .A2(n9923), .ZN(n9922) );
  INV_X1 U11820 ( .A(n11030), .ZN(n9923) );
  NAND2_X1 U11821 ( .A1(n9595), .A2(n13988), .ZN(n13989) );
  AND2_X1 U11822 ( .A1(n14885), .A2(n16249), .ZN(n10062) );
  AND2_X1 U11823 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  INV_X1 U11824 ( .A(n14978), .ZN(n9988) );
  AND2_X1 U11825 ( .A1(n14987), .A2(n15356), .ZN(n9989) );
  INV_X1 U11826 ( .A(n11602), .ZN(n11606) );
  AND2_X1 U11827 ( .A1(n14827), .A2(n15431), .ZN(n9985) );
  INV_X1 U11828 ( .A(n13713), .ZN(n9984) );
  NAND2_X1 U11829 ( .A1(n13636), .A2(n9689), .ZN(n9969) );
  NAND2_X1 U11830 ( .A1(n10462), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10709) );
  NOR2_X1 U11831 ( .A1(n15059), .A2(n9848), .ZN(n9847) );
  INV_X1 U11832 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9848) );
  NOR2_X1 U11833 ( .A1(n18978), .A2(n9854), .ZN(n9853) );
  INV_X1 U11834 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U11835 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U11836 ( .A1(n11593), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10998) );
  AND2_X2 U11837 ( .A1(n10772), .A2(n10771), .ZN(n10782) );
  AND2_X1 U11838 ( .A1(n9708), .A2(n9940), .ZN(n9939) );
  INV_X1 U11839 ( .A(n11272), .ZN(n9940) );
  NAND2_X1 U11840 ( .A1(n11141), .A2(n11140), .ZN(n11142) );
  INV_X1 U11841 ( .A(n15025), .ZN(n11141) );
  INV_X1 U11842 ( .A(n15036), .ZN(n11140) );
  NOR2_X1 U11843 ( .A1(n15251), .A2(n15269), .ZN(n10049) );
  NAND2_X1 U11844 ( .A1(n15049), .A2(n9666), .ZN(n10003) );
  NAND2_X1 U11845 ( .A1(n10005), .A2(n11491), .ZN(n10004) );
  INV_X1 U11846 ( .A(n10735), .ZN(n10736) );
  INV_X1 U11847 ( .A(n14759), .ZN(n9937) );
  NAND2_X1 U11848 ( .A1(n12939), .A2(n10749), .ZN(n10750) );
  NOR2_X1 U11849 ( .A1(n15478), .A2(n11301), .ZN(n10036) );
  NAND2_X1 U11850 ( .A1(n9873), .A2(n9669), .ZN(n10012) );
  NAND2_X1 U11851 ( .A1(n9753), .A2(n19098), .ZN(n11034) );
  CLKBUF_X1 U11852 ( .A(n11562), .Z(n11258) );
  INV_X1 U11853 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13056) );
  AND2_X1 U11854 ( .A1(n10743), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12972) );
  NAND2_X1 U11855 ( .A1(n9594), .A2(n10754), .ZN(n11274) );
  NAND2_X1 U11856 ( .A1(n13151), .A2(n19258), .ZN(n9857) );
  NOR2_X1 U11857 ( .A1(n10573), .A2(n10561), .ZN(n10562) );
  NOR2_X1 U11858 ( .A1(n10581), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10582) );
  AND2_X1 U11859 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10581) );
  OR2_X1 U11860 ( .A1(n18711), .A2(n10398), .ZN(n15630) );
  NAND4_X1 U11861 ( .A1(n18868), .A2(n18878), .A3(n18885), .A4(n18726), .ZN(
        n17142) );
  NAND2_X1 U11862 ( .A1(n10181), .A2(n10043), .ZN(n10042) );
  NAND2_X1 U11863 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10043) );
  NOR2_X1 U11864 ( .A1(n10147), .A2(n10041), .ZN(n10040) );
  INV_X1 U11865 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10041) );
  INV_X1 U11866 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17107) );
  NOR2_X1 U11867 ( .A1(n15799), .A2(n15754), .ZN(n9831) );
  NOR2_X1 U11868 ( .A1(n18917), .A2(n17495), .ZN(n16574) );
  INV_X1 U11869 ( .A(n17792), .ZN(n18126) );
  OAI21_X1 U11870 ( .B1(n10034), .B2(n17859), .A(n10033), .ZN(n10205) );
  NAND2_X1 U11871 ( .A1(n17849), .A2(n9654), .ZN(n10033) );
  NAND2_X1 U11872 ( .A1(n10035), .A2(n9654), .ZN(n10034) );
  NOR2_X1 U11873 ( .A1(n10253), .A2(n10252), .ZN(n10396) );
  NOR2_X1 U11874 ( .A1(n18887), .A2(n18768), .ZN(n18268) );
  INV_X1 U11875 ( .A(n17497), .ZN(n17495) );
  OR2_X1 U11876 ( .A1(n20862), .A2(n12618), .ZN(n15872) );
  AND2_X1 U11877 ( .A1(n13359), .A2(n13358), .ZN(n13513) );
  NAND2_X1 U11878 ( .A1(n20148), .A2(n20142), .ZN(n13387) );
  AND2_X1 U11879 ( .A1(n13337), .A2(n13336), .ZN(n20015) );
  INV_X1 U11880 ( .A(n12098), .ZN(n12560) );
  NOR2_X1 U11881 ( .A1(n12471), .A2(n14186), .ZN(n12472) );
  AND2_X1 U11882 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12422), .ZN(
        n12423) );
  AND2_X1 U11883 ( .A1(n10025), .A2(n14291), .ZN(n10024) );
  CLKBUF_X1 U11884 ( .A(n14194), .Z(n14195) );
  NOR2_X1 U11885 ( .A1(n12376), .A2(n15840), .ZN(n12377) );
  NAND2_X1 U11886 ( .A1(n12377), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12381) );
  NAND2_X1 U11887 ( .A1(n12321), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12376) );
  NOR2_X1 U11888 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NAND2_X1 U11889 ( .A1(n12279), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12320) );
  NAND2_X1 U11890 ( .A1(n12257), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12278) );
  NOR2_X1 U11891 ( .A1(n20915), .A2(n12200), .ZN(n12257) );
  NOR2_X1 U11892 ( .A1(n10016), .A2(n10015), .ZN(n10014) );
  INV_X1 U11893 ( .A(n14223), .ZN(n10015) );
  CLKBUF_X1 U11894 ( .A(n14238), .Z(n14239) );
  AND2_X1 U11895 ( .A1(n12095), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12096) );
  NOR2_X1 U11896 ( .A1(n12090), .A2(n19941), .ZN(n12095) );
  NAND2_X1 U11897 ( .A1(n10019), .A2(n13743), .ZN(n10018) );
  AND3_X1 U11898 ( .A1(n12058), .A2(n12057), .A3(n12056), .ZN(n13678) );
  NAND2_X1 U11899 ( .A1(n12035), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12059) );
  AND2_X1 U11900 ( .A1(n12023), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U11901 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11949), .ZN(
        n12002) );
  NAND2_X1 U11902 ( .A1(n13354), .A2(n11924), .ZN(n13511) );
  AOI21_X1 U11903 ( .B1(n10022), .B2(n11946), .A(n10020), .ZN(n13357) );
  NOR2_X1 U11904 ( .A1(n11904), .A2(n10021), .ZN(n10020) );
  AND2_X1 U11905 ( .A1(n11899), .A2(n10023), .ZN(n10022) );
  INV_X1 U11906 ( .A(n11924), .ZN(n10021) );
  NAND2_X1 U11907 ( .A1(n11910), .A2(n11909), .ZN(n13201) );
  INV_X1 U11908 ( .A(n13205), .ZN(n12712) );
  INV_X1 U11909 ( .A(n12859), .ZN(n9949) );
  AND2_X1 U11910 ( .A1(n14519), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9782) );
  NOR2_X1 U11911 ( .A1(n14212), .A2(n9958), .ZN(n14156) );
  OR3_X1 U11912 ( .A1(n9959), .A2(n9961), .A3(n9960), .ZN(n9958) );
  NOR3_X1 U11913 ( .A1(n14212), .A2(n9959), .A3(n9961), .ZN(n14171) );
  NOR2_X1 U11914 ( .A1(n14212), .A2(n9959), .ZN(n14181) );
  AND2_X1 U11915 ( .A1(n14300), .A2(n12700), .ZN(n14289) );
  OR2_X1 U11916 ( .A1(n14317), .A2(n14308), .ZN(n14310) );
  OR2_X1 U11917 ( .A1(n14326), .A2(n14319), .ZN(n14317) );
  NOR3_X1 U11918 ( .A1(n14343), .A2(n14331), .A3(n9956), .ZN(n14333) );
  AOI21_X1 U11919 ( .B1(n14489), .B2(n12825), .A(n12822), .ZN(n14589) );
  AND2_X1 U11920 ( .A1(n12680), .A2(n12679), .ZN(n14224) );
  AND2_X1 U11921 ( .A1(n12675), .A2(n12674), .ZN(n14342) );
  NOR2_X1 U11922 ( .A1(n14343), .A2(n14342), .ZN(n14344) );
  XNOR2_X1 U11923 ( .A(n14579), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14511) );
  OR2_X1 U11924 ( .A1(n14352), .A2(n14245), .ZN(n14343) );
  AND2_X1 U11925 ( .A1(n13416), .A2(n13408), .ZN(n15810) );
  NAND2_X1 U11926 ( .A1(n14361), .A2(n14350), .ZN(n14352) );
  AND2_X1 U11927 ( .A1(n12666), .A2(n12665), .ZN(n13762) );
  NAND2_X1 U11928 ( .A1(n16012), .A2(n12801), .ZN(n9737) );
  NOR2_X1 U11929 ( .A1(n16184), .A2(n12657), .ZN(n16188) );
  OR2_X1 U11930 ( .A1(n13572), .A2(n13571), .ZN(n16184) );
  OR2_X1 U11931 ( .A1(n13533), .A2(n13532), .ZN(n13572) );
  NOR2_X1 U11932 ( .A1(n15810), .A2(n20098), .ZN(n14613) );
  AND2_X1 U11933 ( .A1(n15814), .A2(n14613), .ZN(n14600) );
  NAND2_X1 U11934 ( .A1(n13416), .A2(n13461), .ZN(n15814) );
  AND2_X1 U11935 ( .A1(n12624), .A2(n12642), .ZN(n13205) );
  XNOR2_X1 U11936 ( .A(n11857), .B(n11781), .ZN(n11915) );
  NAND2_X1 U11937 ( .A1(n11859), .A2(n20231), .ZN(n11876) );
  NAND2_X1 U11938 ( .A1(n9803), .A2(n13576), .ZN(n11979) );
  AND2_X1 U11939 ( .A1(n11727), .A2(n13214), .ZN(n12563) );
  INV_X1 U11940 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15761) );
  INV_X1 U11941 ( .A(n11874), .ZN(n9785) );
  NAND2_X1 U11942 ( .A1(n9783), .A2(n11874), .ZN(n9784) );
  AND3_X1 U11943 ( .A1(n13234), .A2(n13233), .A3(n13232), .ZN(n13494) );
  OR2_X1 U11944 ( .A1(n9615), .A2(n20107), .ZN(n20269) );
  OR2_X1 U11945 ( .A1(n9615), .A2(n12741), .ZN(n20318) );
  AND3_X1 U11946 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20777), .A3(n20108), 
        .ZN(n20149) );
  AND2_X1 U11947 ( .A1(n9615), .A2(n20107), .ZN(n20527) );
  NOR2_X1 U11948 ( .A1(n12749), .A2(n13577), .ZN(n20633) );
  AND2_X1 U11949 ( .A1(n10680), .A2(n10679), .ZN(n16362) );
  INV_X1 U11950 ( .A(n12930), .ZN(n16360) );
  NAND2_X1 U11951 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  NOR2_X1 U11952 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n9930) );
  INV_X1 U11953 ( .A(n11064), .ZN(n9931) );
  NAND2_X1 U11954 ( .A1(n11065), .A2(n11593), .ZN(n11061) );
  OR2_X1 U11955 ( .A1(n11065), .A2(n9711), .ZN(n11062) );
  AND2_X1 U11956 ( .A1(n11059), .A2(n9915), .ZN(n11077) );
  NOR2_X1 U11957 ( .A1(n9917), .A2(n9687), .ZN(n9915) );
  NAND2_X1 U11958 ( .A1(n11077), .A2(n11225), .ZN(n11074) );
  NOR2_X1 U11959 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16381) );
  NOR2_X1 U11960 ( .A1(n11023), .A2(n11022), .ZN(n11031) );
  NOR2_X1 U11961 ( .A1(n13632), .A2(n13822), .ZN(n13682) );
  NAND2_X1 U11962 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13632) );
  INV_X1 U11963 ( .A(n10779), .ZN(n10780) );
  NOR2_X1 U11964 ( .A1(n9627), .A2(n9977), .ZN(n14123) );
  NAND2_X1 U11965 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  NOR2_X1 U11966 ( .A1(n11525), .A2(n11608), .ZN(n9978) );
  NAND2_X1 U11967 ( .A1(n14845), .A2(n9643), .ZN(n10055) );
  INV_X1 U11968 ( .A(n9979), .ZN(n9976) );
  AND2_X1 U11969 ( .A1(n11484), .A2(n11485), .ZN(n14918) );
  NAND2_X1 U11970 ( .A1(n14806), .A2(n9987), .ZN(n15330) );
  NAND2_X1 U11971 ( .A1(n14806), .A2(n9989), .ZN(n15358) );
  AND2_X1 U11972 ( .A1(n11462), .A2(n11461), .ZN(n14807) );
  OR2_X1 U11973 ( .A1(n13840), .A2(n13839), .ZN(n19128) );
  AND2_X1 U11974 ( .A1(n14826), .A2(n9685), .ZN(n15419) );
  NAND2_X1 U11975 ( .A1(n15504), .A2(n9983), .ZN(n15489) );
  AND2_X1 U11976 ( .A1(n15504), .A2(n9686), .ZN(n13795) );
  NAND2_X1 U11977 ( .A1(n15504), .A2(n15503), .ZN(n15505) );
  OAI21_X1 U11978 ( .B1(n12926), .B2(n12925), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14109) );
  NOR2_X1 U11979 ( .A1(n10725), .A2(n10731), .ZN(n13121) );
  AND2_X1 U11980 ( .A1(n19196), .A2(n13126), .ZN(n14111) );
  AND2_X1 U11981 ( .A1(n13072), .A2(n21041), .ZN(n19224) );
  NOR2_X1 U11982 ( .A1(n12931), .A2(n12930), .ZN(n13649) );
  INV_X1 U11983 ( .A(n14109), .ZN(n14110) );
  AND2_X1 U11984 ( .A1(n11539), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14645) );
  AND2_X1 U11985 ( .A1(n11539), .A2(n9720), .ZN(n14647) );
  AND2_X1 U11986 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11507), .ZN(
        n14669) );
  NAND2_X1 U11987 ( .A1(n14669), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14668) );
  NAND2_X1 U11988 ( .A1(n14666), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14665) );
  NOR3_X1 U11989 ( .A1(n14657), .A2(n9851), .A3(n9850), .ZN(n14662) );
  NAND2_X1 U11990 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9850) );
  AND2_X1 U11991 ( .A1(n14662), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14666) );
  NOR2_X1 U11992 ( .A1(n14657), .A2(n15194), .ZN(n14659) );
  NAND2_X1 U11993 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n14658), .ZN(
        n14657) );
  INV_X1 U11994 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U11995 ( .A1(n13710), .A2(n9639), .ZN(n14656) );
  INV_X1 U11996 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13803) );
  NAND2_X1 U11997 ( .A1(n13710), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13802) );
  NOR2_X1 U11998 ( .A1(n19083), .A2(n13708), .ZN(n13710) );
  NAND2_X1 U11999 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n13709), .ZN(
        n13708) );
  NAND2_X1 U12000 ( .A1(n13682), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13706) );
  NOR2_X1 U12001 ( .A1(n13706), .A2(n16314), .ZN(n13709) );
  AND2_X1 U12002 ( .A1(n11174), .A2(n11179), .ZN(n9933) );
  INV_X1 U12003 ( .A(n11619), .ZN(n11590) );
  NAND2_X1 U12004 ( .A1(n11579), .A2(n11578), .ZN(n9999) );
  NAND2_X1 U12005 ( .A1(n14728), .A2(n9708), .ZN(n11271) );
  NAND2_X1 U12006 ( .A1(n14728), .A2(n9939), .ZN(n14836) );
  OR2_X1 U12007 ( .A1(n11144), .A2(n15269), .ZN(n15034) );
  INV_X1 U12008 ( .A(n14751), .ZN(n9974) );
  NAND2_X1 U12009 ( .A1(n14789), .A2(n9706), .ZN(n14766) );
  NAND2_X1 U12010 ( .A1(n14786), .A2(n9707), .ZN(n14761) );
  NAND2_X1 U12011 ( .A1(n14893), .A2(n9640), .ZN(n14787) );
  NOR2_X1 U12012 ( .A1(n14787), .A2(n14788), .ZN(n14786) );
  OR2_X1 U12013 ( .A1(n15402), .A2(n11489), .ZN(n15333) );
  NAND2_X1 U12014 ( .A1(n14893), .A2(n9943), .ZN(n15110) );
  INV_X1 U12015 ( .A(n9874), .ZN(n15129) );
  OAI21_X1 U12016 ( .B1(n15175), .B2(n9673), .A(n9875), .ZN(n9874) );
  NOR2_X1 U12017 ( .A1(n9876), .A2(n15087), .ZN(n9875) );
  AND2_X1 U12018 ( .A1(n14801), .A2(n11227), .ZN(n14893) );
  INV_X1 U12019 ( .A(n14802), .ZN(n11227) );
  NOR2_X1 U12020 ( .A1(n14818), .A2(n14913), .ZN(n15179) );
  NOR2_X1 U12021 ( .A1(n15486), .A2(n15487), .ZN(n15485) );
  NAND2_X1 U12022 ( .A1(n9868), .A2(n9758), .ZN(n15209) );
  INV_X1 U12023 ( .A(n9869), .ZN(n9868) );
  OR2_X1 U12024 ( .A1(n13515), .A2(n13516), .ZN(n15486) );
  OR2_X1 U12025 ( .A1(n16292), .A2(n16325), .ZN(n10988) );
  OAI21_X1 U12026 ( .B1(n9603), .B2(n11033), .A(n9859), .ZN(n15517) );
  NAND2_X1 U12027 ( .A1(n9603), .A2(n10960), .ZN(n9859) );
  NAND2_X1 U12028 ( .A1(n9604), .A2(n11164), .ZN(n11169) );
  CLKBUF_X1 U12029 ( .A(n15229), .Z(n15539) );
  AOI21_X1 U12030 ( .B1(n13817), .B2(n9691), .A(n9865), .ZN(n9864) );
  NOR2_X1 U12031 ( .A1(n13652), .A2(n16341), .ZN(n9865) );
  INV_X1 U12032 ( .A(n11300), .ZN(n15379) );
  NOR2_X1 U12033 ( .A1(n13261), .A2(n11334), .ZN(n13637) );
  CLKBUF_X1 U12034 ( .A(n11274), .Z(n11275) );
  NAND2_X1 U12035 ( .A1(n10053), .A2(n10051), .ZN(n13160) );
  AND2_X1 U12036 ( .A1(n10052), .A2(n13156), .ZN(n10051) );
  INV_X1 U12037 ( .A(n13158), .ZN(n10052) );
  NAND2_X1 U12038 ( .A1(n13149), .A2(n13148), .ZN(n13162) );
  NOR2_X1 U12039 ( .A1(n19871), .A2(n19467), .ZN(n19499) );
  INV_X1 U12040 ( .A(n19865), .ZN(n13444) );
  NAND2_X1 U12041 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  NOR2_X1 U12042 ( .A1(n10503), .A2(n9668), .ZN(n10511) );
  AND2_X1 U12043 ( .A1(n19871), .A2(n19277), .ZN(n19279) );
  NOR2_X2 U12044 ( .A1(n14110), .A2(n13376), .ZN(n19306) );
  NOR2_X2 U12045 ( .A1(n13375), .A2(n13376), .ZN(n19307) );
  INV_X1 U12046 ( .A(n10726), .ZN(n19309) );
  OR2_X1 U12047 ( .A1(n13642), .A2(n19676), .ZN(n16388) );
  AND2_X1 U12048 ( .A1(n9895), .A2(n9894), .ZN(n16637) );
  AND2_X1 U12049 ( .A1(n9896), .A2(n16949), .ZN(n9894) );
  OR2_X1 U12050 ( .A1(n16949), .A2(n16652), .ZN(n9896) );
  OR2_X1 U12051 ( .A1(n16659), .A2(n9897), .ZN(n9895) );
  NAND2_X1 U12052 ( .A1(n17586), .A2(n17598), .ZN(n9897) );
  OR2_X1 U12053 ( .A1(n16659), .A2(n16660), .ZN(n9898) );
  AND2_X1 U12054 ( .A1(n9901), .A2(n9900), .ZN(n16673) );
  AND2_X1 U12055 ( .A1(n9902), .A2(n16949), .ZN(n9900) );
  NOR2_X1 U12056 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16772), .ZN(n16757) );
  INV_X1 U12057 ( .A(n16964), .ZN(n16952) );
  NOR2_X1 U12058 ( .A1(n20919), .A2(n16756), .ZN(n9818) );
  NOR2_X1 U12059 ( .A1(n17205), .A2(n16843), .ZN(n9816) );
  NAND2_X1 U12060 ( .A1(n10140), .A2(n9835), .ZN(n9834) );
  INV_X1 U12061 ( .A(n10150), .ZN(n10102) );
  NOR2_X1 U12062 ( .A1(n18750), .A2(n16555), .ZN(n17496) );
  INV_X1 U12063 ( .A(n10420), .ZN(n10422) );
  NAND2_X1 U12064 ( .A1(n17622), .A2(n9912), .ZN(n12879) );
  NOR2_X1 U12065 ( .A1(n17679), .A2(n16591), .ZN(n17635) );
  NOR2_X1 U12066 ( .A1(n17742), .A2(n17741), .ZN(n17731) );
  AND3_X1 U12067 ( .A1(n9905), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17855) );
  NAND2_X1 U12068 ( .A1(n15744), .A2(n9831), .ZN(n9830) );
  AND2_X1 U12069 ( .A1(n15745), .A2(n10220), .ZN(n15795) );
  NAND2_X1 U12070 ( .A1(n15744), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15794) );
  AOI21_X1 U12071 ( .B1(n17603), .B2(n17930), .A(n17729), .ZN(n10218) );
  OAI21_X1 U12072 ( .B1(n17712), .B2(n17600), .A(n10215), .ZN(n10216) );
  NOR2_X1 U12073 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17659), .ZN(
        n17647) );
  NOR2_X1 U12074 ( .A1(n17712), .A2(n17642), .ZN(n17657) );
  INV_X1 U12075 ( .A(n18723), .ZN(n18081) );
  NOR2_X1 U12076 ( .A1(n18725), .A2(n18707), .ZN(n18057) );
  AND2_X1 U12077 ( .A1(n9759), .A2(n10403), .ZN(n10405) );
  XNOR2_X1 U12078 ( .A(n10205), .B(n10204), .ZN(n17845) );
  XNOR2_X1 U12079 ( .A(n10188), .B(n18235), .ZN(n17903) );
  NAND2_X1 U12080 ( .A1(n18929), .A2(n15738), .ZN(n18736) );
  NOR2_X2 U12081 ( .A1(n10404), .A2(n10392), .ZN(n16575) );
  NOR3_X1 U12082 ( .A1(n9767), .A2(n9764), .A3(n9763), .ZN(n9762) );
  NOR2_X1 U12083 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18268), .ZN(n18564) );
  AOI211_X1 U12084 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n10303), .B(n10302), .ZN(n10304) );
  AOI211_X1 U12085 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n10272), .B(n10271), .ZN(n10273) );
  OAI211_X1 U12086 ( .C1(n9651), .C2(n17050), .A(n10285), .B(n10284), .ZN(
        n18291) );
  AOI22_X1 U12087 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10285) );
  AOI211_X1 U12088 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n10283), .B(n10282), .ZN(n10284) );
  OAI21_X1 U12089 ( .B1(n18104), .B2(n18706), .A(n9692), .ZN(n18708) );
  AOI211_X1 U12090 ( .C1(n15738), .C2(n15737), .A(n15827), .B(n15736), .ZN(
        n18738) );
  INV_X1 U12091 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15867) );
  INV_X1 U12092 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14247) );
  NOR2_X2 U12093 ( .A1(n13614), .A2(n12721), .ZN(n19977) );
  INV_X1 U12094 ( .A(n19949), .ZN(n19989) );
  NAND2_X1 U12095 ( .A1(n15872), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19949) );
  NAND2_X1 U12096 ( .A1(n20862), .A2(n12723), .ZN(n19994) );
  INV_X1 U12097 ( .A(n20014), .ZN(n14362) );
  INV_X1 U12098 ( .A(n15953), .ZN(n14399) );
  AND2_X1 U12099 ( .A1(n12895), .A2(n13399), .ZN(n14405) );
  INV_X1 U12100 ( .A(n14409), .ZN(n14404) );
  NOR2_X2 U12102 ( .A1(n20075), .A2(n13410), .ZN(n20061) );
  XNOR2_X1 U12103 ( .A(n12621), .B(n12620), .ZN(n13601) );
  OR2_X1 U12104 ( .A1(n12619), .A2(n14133), .ZN(n12621) );
  OR2_X1 U12105 ( .A1(n12844), .A2(n12843), .ZN(n12846) );
  INV_X1 U12106 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20915) );
  INV_X1 U12107 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19948) );
  NOR2_X1 U12108 ( .A1(n16035), .A2(n14548), .ZN(n14567) );
  NOR2_X1 U12109 ( .A1(n16045), .A2(n16057), .ZN(n16047) );
  NOR2_X1 U12110 ( .A1(n16088), .A2(n16079), .ZN(n16068) );
  NAND2_X1 U12111 ( .A1(n16092), .A2(n14546), .ZN(n16088) );
  AND2_X1 U12112 ( .A1(n16100), .A2(n9798), .ZN(n16092) );
  INV_X1 U12113 ( .A(n14545), .ZN(n9798) );
  NAND2_X1 U12114 ( .A1(n9814), .A2(n9812), .ZN(n14482) );
  INV_X1 U12115 ( .A(n9995), .ZN(n9812) );
  NAND2_X1 U12116 ( .A1(n13525), .A2(n13526), .ZN(n9991) );
  AND2_X1 U12117 ( .A1(n13416), .A2(n9801), .ZN(n20098) );
  CLKBUF_X1 U12118 ( .A(n11915), .Z(n11916) );
  INV_X1 U12119 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20601) );
  INV_X1 U12120 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20103) );
  OAI21_X1 U12121 ( .B1(n13497), .B2(n16228), .A(n20279), .ZN(n20102) );
  CLKBUF_X1 U12122 ( .A(n13488), .Z(n13489) );
  INV_X1 U12123 ( .A(n15785), .ZN(n14639) );
  OR2_X1 U12124 ( .A1(n20227), .A2(n20190), .ZN(n20263) );
  OAI221_X1 U12125 ( .B1(n20281), .B2(n20566), .C1(n20281), .C2(n20280), .A(
        n20650), .ZN(n20306) );
  OAI211_X1 U12126 ( .C1(n20443), .C2(n20566), .A(n20484), .B(n20427), .ZN(
        n20445) );
  INV_X1 U12127 ( .A(n20414), .ZN(n20444) );
  OAI22_X1 U12128 ( .A1(n20489), .A2(n20488), .B1(n20487), .B2(n20637), .ZN(
        n20513) );
  AND2_X1 U12129 ( .A1(n20521), .A2(n20520), .ZN(n20550) );
  OAI211_X1 U12130 ( .C1(n20694), .C2(n20651), .A(n20650), .B(n20649), .ZN(
        n20698) );
  AND2_X1 U12131 ( .A1(n20707), .A2(n20706), .ZN(n20765) );
  NAND2_X1 U12132 ( .A1(n15781), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19913) );
  INV_X1 U12133 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20776) );
  INV_X1 U12134 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20566) );
  XNOR2_X1 U12135 ( .A(n11592), .B(n11585), .ZN(n11586) );
  AND2_X1 U12136 ( .A1(n9840), .A2(n19118), .ZN(n14701) );
  AND2_X1 U12137 ( .A1(n11595), .A2(n11134), .ZN(n14724) );
  INV_X1 U12138 ( .A(n9840), .ZN(n14713) );
  AND2_X1 U12139 ( .A1(n13656), .A2(n13646), .ZN(n19086) );
  INV_X1 U12140 ( .A(n19127), .ZN(n14829) );
  INV_X1 U12141 ( .A(n19086), .ZN(n19112) );
  AND2_X1 U12142 ( .A1(n13656), .A2(n13655), .ZN(n19122) );
  XNOR2_X1 U12143 ( .A(n11566), .B(n11565), .ZN(n14130) );
  INV_X1 U12144 ( .A(n14699), .ZN(n14856) );
  OR2_X1 U12145 ( .A1(n11530), .A2(n14712), .ZN(n15250) );
  NAND2_X1 U12146 ( .A1(n10060), .A2(n14903), .ZN(n10059) );
  OR2_X1 U12147 ( .A1(n11408), .A2(n11407), .ZN(n13826) );
  NOR2_X1 U12148 ( .A1(n11395), .A2(n11394), .ZN(n19142) );
  INV_X1 U12149 ( .A(n19148), .ZN(n19156) );
  NAND2_X1 U12150 ( .A1(n14039), .A2(n10057), .ZN(n10056) );
  CLKBUF_X1 U12151 ( .A(n14863), .Z(n14864) );
  CLKBUF_X1 U12152 ( .A(n14869), .Z(n14870) );
  AND2_X1 U12153 ( .A1(n14111), .A2(n14110), .ZN(n19166) );
  AND2_X1 U12154 ( .A1(n19196), .A2(n10742), .ZN(n19164) );
  NOR2_X1 U12155 ( .A1(n13261), .A2(n9970), .ZN(n15546) );
  NAND2_X1 U12156 ( .A1(n9703), .A2(n9973), .ZN(n9970) );
  AND2_X1 U12157 ( .A1(n19196), .A2(n19309), .ZN(n19214) );
  INV_X1 U12158 ( .A(n19196), .ZN(n19213) );
  NAND2_X1 U12159 ( .A1(n19196), .A2(n11314), .ZN(n19218) );
  NOR2_X1 U12160 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13073), .ZN(n13248) );
  INV_X1 U12161 ( .A(n13137), .ZN(n13091) );
  NAND2_X1 U12162 ( .A1(n9845), .A2(n11567), .ZN(n9841) );
  INV_X1 U12163 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19083) );
  INV_X1 U12164 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13822) );
  NAND2_X1 U12165 ( .A1(n12941), .A2(n11504), .ZN(n16315) );
  INV_X1 U12166 ( .A(n16315), .ZN(n16297) );
  AND2_X1 U12167 ( .A1(n11516), .A2(n10710), .ZN(n16293) );
  OAI21_X1 U12168 ( .B1(n15175), .B2(n9880), .A(n9878), .ZN(n15141) );
  NAND2_X1 U12169 ( .A1(n9883), .A2(n9881), .ZN(n15148) );
  INV_X1 U12170 ( .A(n9884), .ZN(n9881) );
  NAND2_X1 U12171 ( .A1(n15175), .A2(n9885), .ZN(n9883) );
  OAI21_X1 U12172 ( .B1(n15175), .B2(n15082), .A(n15173), .ZN(n15164) );
  CLKBUF_X1 U12173 ( .A(n13151), .Z(n13164) );
  NAND2_X1 U12174 ( .A1(n9867), .A2(n13652), .ZN(n13819) );
  INV_X1 U12175 ( .A(n16331), .ZN(n19261) );
  INV_X1 U12176 ( .A(n19257), .ZN(n16333) );
  NAND2_X1 U12177 ( .A1(n15379), .A2(n15378), .ZN(n15565) );
  NAND2_X1 U12178 ( .A1(n13117), .A2(n13116), .ZN(n19894) );
  INV_X1 U12179 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19891) );
  INV_X1 U12180 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19881) );
  NAND2_X1 U12181 ( .A1(n13149), .A2(n13068), .ZN(n19877) );
  NAND2_X1 U12182 ( .A1(n13063), .A2(n12981), .ZN(n19887) );
  AND2_X1 U12183 ( .A1(n13163), .A2(n13191), .ZN(n19871) );
  OR2_X1 U12184 ( .A1(n13162), .A2(n13161), .ZN(n13163) );
  AND2_X1 U12185 ( .A1(n19462), .A2(n19865), .ZN(n19396) );
  INV_X1 U12186 ( .A(n19412), .ZN(n19430) );
  OR3_X1 U12187 ( .A1(n19471), .A2(n19680), .A3(n19470), .ZN(n19490) );
  NOR2_X2 U12188 ( .A1(n19674), .A2(n13444), .ZN(n19623) );
  INV_X1 U12189 ( .A(n19731), .ZN(n19652) );
  NOR2_X2 U12190 ( .A1(n19674), .A2(n13377), .ZN(n19670) );
  INV_X1 U12191 ( .A(n19735), .ZN(n19689) );
  INV_X1 U12192 ( .A(n19751), .ZN(n19697) );
  OR3_X1 U12193 ( .A1(n19681), .A2(n19680), .A3(n19679), .ZN(n19710) );
  OAI21_X1 U12194 ( .B1(n19686), .B2(n19685), .A(n19684), .ZN(n19709) );
  AND2_X1 U12195 ( .A1(n19279), .A2(n19433), .ZN(n19707) );
  INV_X1 U12196 ( .A(n19776), .ZN(n19708) );
  INV_X1 U12197 ( .A(n19634), .ZN(n19737) );
  INV_X1 U12198 ( .A(n19643), .ZN(n19754) );
  NOR2_X1 U12199 ( .A1(n19674), .A2(n19720), .ZN(n19755) );
  INV_X1 U12200 ( .A(n19620), .ZN(n19762) );
  INV_X1 U12201 ( .A(n19758), .ZN(n19771) );
  INV_X1 U12202 ( .A(n16388), .ZN(n19777) );
  INV_X1 U12203 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n21039) );
  XNOR2_X1 U12204 ( .A(n18917), .B(n15632), .ZN(n18929) );
  INV_X1 U12205 ( .A(n9761), .ZN(n16556) );
  INV_X1 U12206 ( .A(n17496), .ZN(n17458) );
  INV_X1 U12207 ( .A(n9910), .ZN(n16605) );
  AND2_X1 U12208 ( .A1(n9898), .A2(n16949), .ZN(n16651) );
  AND2_X1 U12209 ( .A1(n9904), .A2(n16949), .ZN(n16681) );
  AND2_X1 U12210 ( .A1(n9888), .A2(n9887), .ZN(n16702) );
  NOR2_X2 U12211 ( .A1(n16578), .A2(n16581), .ZN(n16920) );
  OR2_X1 U12212 ( .A1(n9893), .A2(n9890), .ZN(n16712) );
  INV_X1 U12213 ( .A(n9889), .ZN(n16711) );
  INV_X1 U12214 ( .A(n16920), .ZN(n16959) );
  NOR2_X1 U12215 ( .A1(n16976), .A2(n16975), .ZN(n17003) );
  NOR3_X1 U12216 ( .A1(n17016), .A2(n16969), .A3(n16968), .ZN(n17009) );
  NAND2_X1 U12217 ( .A1(n17024), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17016) );
  NOR2_X1 U12218 ( .A1(n17027), .A2(n9819), .ZN(n17024) );
  NAND2_X1 U12219 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .ZN(n9819) );
  NAND2_X1 U12220 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17046), .ZN(n17027) );
  INV_X1 U12221 ( .A(n17027), .ZN(n17032) );
  NOR2_X1 U12222 ( .A1(n17061), .A2(n17062), .ZN(n17033) );
  AND2_X1 U12223 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17033), .ZN(n17046) );
  NAND2_X1 U12224 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17074), .ZN(n17062) );
  NAND2_X1 U12225 ( .A1(n17135), .A2(n9647), .ZN(n17090) );
  NAND2_X1 U12226 ( .A1(n17135), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n17119) );
  NOR2_X1 U12227 ( .A1(n17121), .A2(n17151), .ZN(n17135) );
  NAND2_X1 U12228 ( .A1(n17170), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n17151) );
  NAND2_X1 U12229 ( .A1(n17240), .A2(n9645), .ZN(n17202) );
  NOR2_X1 U12230 ( .A1(n17242), .A2(n17262), .ZN(n17240) );
  NAND2_X1 U12231 ( .A1(n17240), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17239) );
  INV_X1 U12232 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17269) );
  NOR2_X1 U12233 ( .A1(n17272), .A2(n17267), .ZN(n17271) );
  AND2_X1 U12234 ( .A1(n17291), .A2(n9815), .ZN(n17273) );
  INV_X1 U12235 ( .A(n17278), .ZN(n9815) );
  NAND2_X1 U12236 ( .A1(n17273), .A2(P3_EBX_REG_5__SCAN_IN), .ZN(n17272) );
  NOR2_X1 U12237 ( .A1(n15825), .A2(n15633), .ZN(n17291) );
  OR3_X1 U12238 ( .A1(n18917), .A2(n15632), .A3(n18750), .ZN(n15633) );
  INV_X1 U12239 ( .A(n17291), .ZN(n17294) );
  NAND2_X1 U12240 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17327), .ZN(n17323) );
  INV_X1 U12241 ( .A(n17337), .ZN(n17333) );
  NAND2_X1 U12242 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17333), .ZN(n17332) );
  NOR2_X1 U12243 ( .A1(n17380), .A2(n17302), .ZN(n17343) );
  OAI211_X2 U12244 ( .C1(n15688), .C2(n17264), .A(n10295), .B(n10294), .ZN(
        n18299) );
  AOI22_X1 U12245 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10247), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10295) );
  AOI211_X1 U12246 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n10293), .B(n10292), .ZN(n10294) );
  INV_X1 U12247 ( .A(n17373), .ZN(n17369) );
  NAND2_X1 U12248 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17369), .ZN(n17368) );
  INV_X1 U12249 ( .A(n17383), .ZN(n17372) );
  NAND2_X1 U12250 ( .A1(n17384), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17380) );
  NOR2_X1 U12251 ( .A1(n17546), .A2(n17408), .ZN(n17407) );
  NOR2_X1 U12252 ( .A1(n15828), .A2(n17425), .ZN(n17414) );
  AND2_X1 U12253 ( .A1(n10121), .A2(n10120), .ZN(n10126) );
  NAND2_X1 U12254 ( .A1(n17414), .A2(n18722), .ZN(n17448) );
  INV_X1 U12255 ( .A(n17450), .ZN(n17447) );
  NOR2_X1 U12256 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  INV_X1 U12257 ( .A(n17414), .ZN(n17453) );
  NOR2_X1 U12258 ( .A1(n10184), .A2(n10038), .ZN(n10185) );
  INV_X1 U12259 ( .A(n17448), .ZN(n17451) );
  NOR2_X1 U12260 ( .A1(n17458), .A2(n17457), .ZN(n17476) );
  NOR2_X1 U12261 ( .A1(n18917), .A2(n17559), .ZN(n17549) );
  OAI211_X1 U12262 ( .C1(n18917), .C2(n18918), .A(n17497), .B(n17496), .ZN(
        n17552) );
  BUF_X1 U12263 ( .A(n17552), .Z(n17559) );
  NAND2_X1 U12265 ( .A1(n17573), .A2(n17574), .ZN(n17572) );
  INV_X1 U12266 ( .A(n17582), .ZN(n17595) );
  NOR2_X1 U12267 ( .A1(n17820), .A2(n18046), .ZN(n17708) );
  NAND3_X1 U12268 ( .A1(n17786), .A2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17742) );
  NOR3_X1 U12269 ( .A1(n16857), .A2(n17784), .A3(n10419), .ZN(n17786) );
  INV_X1 U12270 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10419) );
  INV_X1 U12271 ( .A(n18587), .ZN(n18648) );
  INV_X1 U12272 ( .A(n17797), .ZN(n17821) );
  NAND2_X1 U12273 ( .A1(n9905), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17866) );
  NOR2_X2 U12274 ( .A1(n16575), .A2(n15732), .ZN(n18716) );
  AND2_X1 U12275 ( .A1(n10211), .A2(n9658), .ZN(n9829) );
  NAND2_X1 U12276 ( .A1(n18057), .A2(n18723), .ZN(n18162) );
  AND2_X1 U12277 ( .A1(n18710), .A2(n9768), .ZN(n18723) );
  OR2_X1 U12278 ( .A1(n15732), .A2(n18711), .ZN(n9768) );
  NAND2_X1 U12279 ( .A1(n10044), .A2(n17724), .ZN(n17831) );
  INV_X1 U12280 ( .A(n10045), .ZN(n10044) );
  INV_X1 U12281 ( .A(n17832), .ZN(n18173) );
  NOR2_X1 U12282 ( .A1(n17859), .A2(n10199), .ZN(n17850) );
  INV_X1 U12283 ( .A(n18736), .ZN(n18707) );
  NAND2_X1 U12284 ( .A1(n10355), .A2(n10327), .ZN(n18700) );
  AOI21_X2 U12285 ( .B1(n15734), .B2(n10356), .A(n18750), .ZN(n18238) );
  INV_X1 U12286 ( .A(n18238), .ZN(n18254) );
  NOR2_X1 U12287 ( .A1(n18700), .A2(n18254), .ZN(n18252) );
  INV_X1 U12288 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18271) );
  INV_X1 U12289 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18266) );
  OAI211_X1 U12290 ( .C1(n18750), .C2(n18738), .A(n18267), .B(n15739), .ZN(
        n18891) );
  INV_X1 U12291 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18593) );
  INV_X1 U12292 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18597) );
  INV_X1 U12293 ( .A(n18750), .ZN(n18910) );
  NOR2_X1 U12294 ( .A1(n18859), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18763) );
  INV_X1 U12295 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18859) );
  INV_X1 U12296 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18862) );
  NAND2_X1 U12297 ( .A1(n18787), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18926) );
  AOI21_X1 U12299 ( .B1(n12864), .B2(n12863), .A(n12862), .ZN(n12865) );
  NOR2_X1 U12300 ( .A1(n20014), .A2(n12861), .ZN(n12862) );
  OAI21_X1 U12301 ( .B1(n14559), .B2(n19920), .A(n14420), .ZN(P1_U2969) );
  AND2_X1 U12302 ( .A1(n9950), .A2(n9946), .ZN(n9778) );
  NAND2_X1 U12303 ( .A1(n14542), .A2(n20093), .ZN(n9946) );
  NOR3_X1 U12304 ( .A1(n14540), .A2(n14541), .A3(n9663), .ZN(n9950) );
  OAI211_X1 U12305 ( .C1(n16038), .C2(n16204), .A(n16040), .B(n9810), .ZN(
        P1_U3004) );
  AOI21_X1 U12306 ( .B1(n16039), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9811), .ZN(n9810) );
  INV_X1 U12307 ( .A(n11545), .ZN(n11546) );
  OAI211_X1 U12308 ( .C1(n14132), .C2(n19264), .A(n9963), .B(n9860), .ZN(
        P2_U3015) );
  AND2_X1 U12309 ( .A1(n9962), .A2(n9861), .ZN(n9860) );
  INV_X1 U12310 ( .A(n14126), .ZN(n9861) );
  NOR2_X1 U12311 ( .A1(n11616), .A2(n11615), .ZN(n11624) );
  INV_X1 U12312 ( .A(n11535), .ZN(n11536) );
  AOI21_X1 U12313 ( .B1(n9910), .B2(n9909), .A(n9906), .ZN(n16601) );
  AND2_X1 U12314 ( .A1(n10427), .A2(n10426), .ZN(n10428) );
  AOI22_X1 U12315 ( .A1(n17709), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n18040), .B2(n17834), .ZN(n17699) );
  AND2_X1 U12316 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  NOR2_X1 U12317 ( .A1(n10091), .A2(n18731), .ZN(n10150) );
  OR2_X2 U12318 ( .A1(n10087), .A2(n10090), .ZN(n9722) );
  NAND2_X1 U12319 ( .A1(n13788), .A2(n9644), .ZN(n15176) );
  AND2_X1 U12320 ( .A1(n14038), .A2(n10058), .ZN(n9626) );
  NAND2_X1 U12321 ( .A1(n19147), .A2(n13522), .ZN(n13830) );
  NOR2_X2 U12322 ( .A1(n17427), .A2(n16436), .ZN(n17833) );
  INV_X1 U12323 ( .A(n17833), .ZN(n17729) );
  INV_X1 U12324 ( .A(n11788), .ZN(n12536) );
  OR2_X1 U12325 ( .A1(n14719), .A2(n14718), .ZN(n9627) );
  OR3_X2 U12326 ( .A1(n18868), .A2(n18893), .A3(n18732), .ZN(n9649) );
  OR3_X2 U12327 ( .A1(n18868), .A2(n18878), .A3(n10092), .ZN(n9651) );
  NAND2_X1 U12328 ( .A1(n15103), .A2(n9723), .ZN(n15055) );
  AND2_X4 U12329 ( .A1(n10431), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9628) );
  NAND2_X1 U12330 ( .A1(n13788), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13787) );
  NAND2_X1 U12331 ( .A1(n9661), .A2(n13790), .ZN(n13789) );
  NAND2_X1 U12332 ( .A1(n10721), .A2(n11020), .ZN(n11284) );
  AND2_X1 U12333 ( .A1(n14314), .A2(n10025), .ZN(n14290) );
  AND2_X1 U12334 ( .A1(n13681), .A2(n10066), .ZN(n9630) );
  INV_X2 U12335 ( .A(n10627), .ZN(n10628) );
  AND2_X1 U12336 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9631) );
  AND2_X1 U12337 ( .A1(n14789), .A2(n9719), .ZN(n14734) );
  AND2_X1 U12338 ( .A1(n12755), .A2(n12756), .ZN(n9632) );
  INV_X1 U12339 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17865) );
  AND2_X1 U12340 ( .A1(n9830), .A2(n9714), .ZN(n9633) );
  OR2_X1 U12341 ( .A1(n15480), .A2(n10009), .ZN(n9634) );
  NAND2_X1 U12342 ( .A1(n12774), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9635) );
  AND2_X1 U12343 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9636)
         );
  NAND2_X1 U12344 ( .A1(n13680), .A2(n13681), .ZN(n13280) );
  NAND2_X1 U12345 ( .A1(n14882), .A2(n9681), .ZN(n14877) );
  AND2_X1 U12346 ( .A1(n17135), .A2(n9818), .ZN(n9637) );
  OR3_X1 U12347 ( .A1(n14657), .A2(n9852), .A3(n15194), .ZN(n9638) );
  AND2_X1 U12348 ( .A1(n9855), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9639) );
  AND2_X1 U12349 ( .A1(n9943), .A2(n9942), .ZN(n9640) );
  AND2_X1 U12350 ( .A1(n17729), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9641) );
  NOR2_X1 U12351 ( .A1(n16918), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9893) );
  AND2_X1 U12352 ( .A1(n9847), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9642) );
  NOR2_X1 U12353 ( .A1(n14840), .A2(n14846), .ZN(n9643) );
  INV_X1 U12354 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15166) );
  AND2_X1 U12355 ( .A1(n10036), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9644) );
  AND2_X1 U12356 ( .A1(n9816), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n9645) );
  AND2_X1 U12357 ( .A1(n9644), .A2(n11488), .ZN(n9646) );
  AND2_X1 U12358 ( .A1(n9818), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n9647) );
  AND2_X1 U12359 ( .A1(n10049), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9648) );
  AND2_X2 U12360 ( .A1(n9621), .A2(n16349), .ZN(n10669) );
  NAND2_X1 U12361 ( .A1(n14522), .A2(n12815), .ZN(n14488) );
  AND2_X2 U12362 ( .A1(n9623), .A2(n16349), .ZN(n10662) );
  AND2_X2 U12363 ( .A1(n13410), .A2(n20109), .ZN(n11773) );
  AND4_X1 U12364 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n9650) );
  AND2_X1 U12365 ( .A1(n14314), .A2(n14315), .ZN(n14302) );
  AND2_X1 U12366 ( .A1(n9873), .A2(n9629), .ZN(n15213) );
  NAND2_X1 U12367 ( .A1(n11633), .A2(n13468), .ZN(n11713) );
  OR2_X1 U12368 ( .A1(n14152), .A2(n10031), .ZN(n12845) );
  OR2_X1 U12369 ( .A1(n11069), .A2(n9929), .ZN(n9653) );
  INV_X1 U12370 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U12371 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10202), .ZN(
        n9654) );
  OR2_X1 U12372 ( .A1(n11098), .A2(n15319), .ZN(n9655) );
  OR2_X1 U12373 ( .A1(n14579), .A2(n12816), .ZN(n9656) );
  NAND2_X1 U12374 ( .A1(n10055), .A2(n10054), .ZN(n14838) );
  AND4_X1 U12375 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n9657) );
  NAND2_X1 U12376 ( .A1(n10013), .A2(n12178), .ZN(n14336) );
  NOR2_X1 U12377 ( .A1(n14238), .A2(n10016), .ZN(n14221) );
  NAND2_X1 U12378 ( .A1(n14314), .A2(n10027), .ZN(n14293) );
  AND2_X1 U12379 ( .A1(n11857), .A2(n11856), .ZN(n11859) );
  OR2_X1 U12380 ( .A1(n13151), .A2(n10796), .ZN(n10884) );
  NAND2_X1 U12381 ( .A1(n9921), .A2(n9922), .ZN(n11038) );
  NAND2_X1 U12383 ( .A1(n9738), .A2(n12813), .ZN(n13769) );
  NAND2_X1 U12384 ( .A1(n9737), .A2(n12802), .ZN(n13721) );
  OR2_X1 U12385 ( .A1(n17729), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9658) );
  OR3_X1 U12386 ( .A1(n11537), .A2(n15018), .A3(n16308), .ZN(n9659) );
  OR3_X1 U12387 ( .A1(n11122), .A2(n11121), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n9660) );
  AND2_X1 U12388 ( .A1(n10012), .A2(n10011), .ZN(n9661) );
  OR2_X1 U12389 ( .A1(n14142), .A2(n20106), .ZN(n9662) );
  NOR3_X1 U12390 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14552), .ZN(n9663) );
  NAND2_X1 U12391 ( .A1(n12978), .A2(n12977), .ZN(n13060) );
  OR2_X1 U12392 ( .A1(n10091), .A2(n10087), .ZN(n17148) );
  AND2_X1 U12393 ( .A1(n10008), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9664) );
  XNOR2_X1 U12394 ( .A(n10599), .B(n10721), .ZN(n10608) );
  NAND2_X1 U12395 ( .A1(n10920), .A2(n10919), .ZN(n10927) );
  INV_X1 U12396 ( .A(n10927), .ZN(n10921) );
  INV_X1 U12397 ( .A(n10057), .ZN(n14852) );
  AND2_X1 U12398 ( .A1(n18878), .A2(n18868), .ZN(n9665) );
  XNOR2_X1 U12399 ( .A(n10760), .B(n10761), .ZN(n10784) );
  NAND2_X1 U12400 ( .A1(n10056), .A2(n14061), .ZN(n14839) );
  OR2_X1 U12401 ( .A1(n10005), .A2(n11491), .ZN(n9666) );
  AND2_X1 U12402 ( .A1(n13722), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9667) );
  NOR2_X1 U12403 ( .A1(n10573), .A2(n10502), .ZN(n9668) );
  NAND2_X1 U12404 ( .A1(n10779), .A2(n10778), .ZN(n10785) );
  INV_X1 U12405 ( .A(n9886), .ZN(n9885) );
  NAND2_X1 U12406 ( .A1(n15173), .A2(n15162), .ZN(n9886) );
  AND2_X1 U12407 ( .A1(n9629), .A2(n11047), .ZN(n9669) );
  AND2_X1 U12408 ( .A1(n9808), .A2(n11911), .ZN(n9670) );
  AND2_X1 U12409 ( .A1(n11051), .A2(n11199), .ZN(n11056) );
  AND2_X1 U12410 ( .A1(n13788), .A2(n9646), .ZN(n15149) );
  OR2_X1 U12411 ( .A1(n10573), .A2(n10488), .ZN(n9671) );
  AND4_X1 U12412 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n9672) );
  INV_X1 U12413 ( .A(n18284), .ZN(n10397) );
  OAI211_X1 U12414 ( .C1(n9651), .C2(n17189), .A(n10305), .B(n10304), .ZN(
        n18284) );
  INV_X1 U12415 ( .A(n9833), .ZN(n17446) );
  OR3_X1 U12416 ( .A1(n9834), .A2(n10137), .A3(n10136), .ZN(n9833) );
  INV_X1 U12417 ( .A(n11046), .ZN(n10011) );
  OR2_X1 U12418 ( .A1(n16285), .A2(n15214), .ZN(n11046) );
  OR2_X1 U12419 ( .A1(n9880), .A2(n9877), .ZN(n9673) );
  AND2_X1 U12420 ( .A1(n15103), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9674) );
  AND2_X1 U12421 ( .A1(n11774), .A2(n13412), .ZN(n9675) );
  NAND2_X1 U12422 ( .A1(n9999), .A2(n11581), .ZN(n15013) );
  AND2_X1 U12423 ( .A1(n13827), .A2(n13826), .ZN(n9676) );
  AND2_X1 U12424 ( .A1(n15033), .A2(n10047), .ZN(n15019) );
  INV_X1 U12425 ( .A(n10703), .ZN(n10721) );
  OAI21_X1 U12426 ( .B1(n14581), .B2(n12829), .A(n12833), .ZN(n14473) );
  NOR2_X1 U12427 ( .A1(n9634), .A2(n11046), .ZN(n10008) );
  INV_X1 U12428 ( .A(n10008), .ZN(n9872) );
  AND2_X1 U12429 ( .A1(n13788), .A2(n10036), .ZN(n9677) );
  AND2_X1 U12430 ( .A1(n9658), .A2(n9828), .ZN(n9678) );
  NAND2_X1 U12431 ( .A1(n10712), .A2(n21042), .ZN(n10735) );
  AND2_X2 U12432 ( .A1(n11313), .A2(n10742), .ZN(n11602) );
  AND2_X1 U12433 ( .A1(n14826), .A2(n14827), .ZN(n14825) );
  AND2_X1 U12434 ( .A1(n14826), .A2(n9985), .ZN(n15416) );
  AND2_X1 U12435 ( .A1(n14882), .A2(n14885), .ZN(n14883) );
  NOR2_X1 U12436 ( .A1(n13662), .A2(n13678), .ZN(n13677) );
  NAND2_X1 U12437 ( .A1(n14893), .A2(n9945), .ZN(n14886) );
  AND2_X1 U12438 ( .A1(n14666), .A2(n9853), .ZN(n9679) );
  AND2_X1 U12439 ( .A1(n13710), .A2(n9855), .ZN(n9680) );
  AND2_X1 U12440 ( .A1(n10062), .A2(n14878), .ZN(n9681) );
  AND2_X1 U12441 ( .A1(n14882), .A2(n10062), .ZN(n14876) );
  AND2_X1 U12442 ( .A1(n13536), .A2(n13568), .ZN(n9682) );
  AND2_X1 U12443 ( .A1(n14669), .A2(n9847), .ZN(n9683) );
  AND2_X1 U12444 ( .A1(n13700), .A2(n9954), .ZN(n9684) );
  NAND2_X1 U12445 ( .A1(n12794), .A2(n16018), .ZN(n16012) );
  NAND2_X1 U12446 ( .A1(n9991), .A2(n12764), .ZN(n13547) );
  AND2_X1 U12447 ( .A1(n9985), .A2(n15417), .ZN(n9685) );
  NOR2_X1 U12448 ( .A1(n13662), .A2(n10018), .ZN(n13742) );
  AND2_X1 U12449 ( .A1(n14806), .A2(n14987), .ZN(n14986) );
  NOR2_X1 U12450 ( .A1(n15397), .A2(n14807), .ZN(n14806) );
  NAND2_X1 U12451 ( .A1(n10207), .A2(n18165), .ZN(n17724) );
  NOR2_X1 U12452 ( .A1(n11328), .A2(n11327), .ZN(n11332) );
  NAND2_X1 U12453 ( .A1(n14789), .A2(n14781), .ZN(n14765) );
  NOR2_X1 U12454 ( .A1(n15181), .A2(n14904), .ZN(n14801) );
  AND2_X1 U12455 ( .A1(n13160), .A2(n13189), .ZN(n13161) );
  AND2_X1 U12456 ( .A1(n9984), .A2(n15503), .ZN(n9686) );
  NAND2_X1 U12457 ( .A1(n10611), .A2(n10610), .ZN(n10695) );
  AND2_X1 U12458 ( .A1(n11593), .A2(n11060), .ZN(n9687) );
  OR2_X1 U12459 ( .A1(n12609), .A2(n12607), .ZN(n9688) );
  AND2_X1 U12460 ( .A1(n9973), .A2(n15547), .ZN(n9689) );
  NAND2_X1 U12461 ( .A1(n11082), .A2(n11130), .ZN(n11059) );
  INV_X1 U12462 ( .A(n11059), .ZN(n9918) );
  AND2_X1 U12463 ( .A1(n11315), .A2(n11330), .ZN(n9690) );
  NAND2_X1 U12464 ( .A1(n13652), .A2(n16341), .ZN(n9691) );
  INV_X1 U12465 ( .A(n9849), .ZN(n14661) );
  NOR3_X1 U12466 ( .A1(n14657), .A2(n9851), .A3(n9852), .ZN(n9849) );
  OR2_X1 U12467 ( .A1(n18700), .A2(n10416), .ZN(n9692) );
  AND2_X1 U12468 ( .A1(n9987), .A2(n9986), .ZN(n9693) );
  INV_X1 U12469 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20777) );
  OR2_X1 U12470 ( .A1(n11457), .A2(n11456), .ZN(n14903) );
  OR2_X1 U12471 ( .A1(n14212), .A2(n14197), .ZN(n9694) );
  AND2_X2 U12472 ( .A1(n11628), .A2(n11625), .ZN(n11838) );
  INV_X1 U12473 ( .A(n11792), .ZN(n11833) );
  NAND2_X1 U12474 ( .A1(n14786), .A2(n14775), .ZN(n14758) );
  OR2_X1 U12475 ( .A1(n14343), .A2(n9956), .ZN(n9695) );
  INV_X1 U12476 ( .A(n15975), .ZN(n14519) );
  AND2_X1 U12477 ( .A1(n14893), .A2(n14892), .ZN(n14891) );
  INV_X1 U12478 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U12479 ( .A1(n11913), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12093) );
  AND2_X1 U12480 ( .A1(n9685), .A2(n15398), .ZN(n9696) );
  NAND2_X1 U12481 ( .A1(n18284), .A2(n18299), .ZN(n10403) );
  AND2_X1 U12482 ( .A1(n9983), .A2(n9982), .ZN(n9697) );
  AND2_X1 U12483 ( .A1(n9952), .A2(n9951), .ZN(n9698) );
  AND2_X1 U12484 ( .A1(n9681), .A2(n10061), .ZN(n9699) );
  AND2_X1 U12485 ( .A1(n9912), .A2(n9911), .ZN(n9700) );
  AND2_X1 U12486 ( .A1(n9826), .A2(n9825), .ZN(n9701) );
  INV_X1 U12487 ( .A(n13376), .ZN(n16311) );
  NAND3_X2 U12488 ( .A1(n19869), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19726), 
        .ZN(n13376) );
  INV_X2 U12489 ( .A(n19159), .ZN(n19153) );
  OR2_X1 U12490 ( .A1(n20148), .A2(n20856), .ZN(n9702) );
  AND2_X1 U12491 ( .A1(n9968), .A2(n13636), .ZN(n9703) );
  INV_X1 U12492 ( .A(n13261), .ZN(n9972) );
  NOR2_X1 U12493 ( .A1(n16189), .A2(n16188), .ZN(n9704) );
  NAND2_X1 U12494 ( .A1(n13416), .A2(n13404), .ZN(n16204) );
  NAND2_X1 U12495 ( .A1(n13680), .A2(n9630), .ZN(n13518) );
  INV_X1 U12496 ( .A(n16723), .ZN(n9890) );
  NAND2_X1 U12497 ( .A1(n16188), .A2(n9952), .ZN(n9705) );
  AND2_X1 U12498 ( .A1(n9975), .A2(n14781), .ZN(n9706) );
  INV_X1 U12499 ( .A(n15760), .ZN(n9801) );
  NAND2_X1 U12500 ( .A1(n9934), .A2(n11174), .ZN(n13193) );
  AND2_X1 U12501 ( .A1(n14775), .A2(n9937), .ZN(n9707) );
  AND2_X1 U12502 ( .A1(n14711), .A2(n11531), .ZN(n9708) );
  NAND2_X1 U12503 ( .A1(n11350), .A2(n11349), .ZN(n15522) );
  INV_X1 U12504 ( .A(n11587), .ZN(n11596) );
  OR2_X1 U12505 ( .A1(n17833), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9709) );
  AND2_X1 U12506 ( .A1(n15461), .A2(n15460), .ZN(n14826) );
  INV_X1 U12507 ( .A(n19118), .ZN(n19102) );
  OAI22_X2 U12508 ( .A1(n21039), .A2(n11548), .B1(n13633), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19118) );
  AND3_X1 U12509 ( .A1(n13743), .A2(n10019), .A3(n13760), .ZN(n9710) );
  INV_X1 U12510 ( .A(n11119), .ZN(n9925) );
  NAND2_X1 U12511 ( .A1(n13191), .A2(n13190), .ZN(n13680) );
  NAND2_X1 U12512 ( .A1(n11858), .A2(n9783), .ZN(n20157) );
  AND2_X1 U12513 ( .A1(n11593), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9711) );
  OR3_X1 U12514 ( .A1(n14343), .A2(n14342), .A3(n9955), .ZN(n9712) );
  AND2_X1 U12515 ( .A1(n19147), .A2(n10060), .ZN(n9713) );
  AND2_X1 U12516 ( .A1(n10224), .A2(n9709), .ZN(n9714) );
  AND2_X1 U12517 ( .A1(n9939), .A2(n9938), .ZN(n9715) );
  AND2_X1 U12518 ( .A1(n13680), .A2(n9636), .ZN(n19146) );
  AND2_X1 U12519 ( .A1(n9889), .A2(n16949), .ZN(n9716) );
  NOR2_X1 U12520 ( .A1(n17850), .A2(n17849), .ZN(n9717) );
  NAND2_X1 U12521 ( .A1(n17240), .A2(n9816), .ZN(n9817) );
  INV_X1 U12522 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17918) );
  INV_X1 U12523 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15194) );
  AND2_X1 U12524 ( .A1(n9853), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9718) );
  AND2_X1 U12525 ( .A1(n12177), .A2(n12176), .ZN(n14347) );
  AND2_X1 U12526 ( .A1(n9706), .A2(n9974), .ZN(n9719) );
  AND2_X1 U12527 ( .A1(n20377), .A2(n12847), .ZN(n16029) );
  INV_X1 U12528 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16217) );
  INV_X1 U12529 ( .A(n15109), .ZN(n9942) );
  AND2_X1 U12530 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9720) );
  AND3_X1 U12531 ( .A1(n13104), .A2(n13399), .A3(n13390), .ZN(n20087) );
  INV_X1 U12532 ( .A(n10590), .ZN(n10627) );
  NAND2_X1 U12533 ( .A1(n12668), .A2(n12667), .ZN(n9721) );
  INV_X1 U12534 ( .A(n9845), .ZN(n9844) );
  NAND2_X1 U12535 ( .A1(n9720), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9845) );
  INV_X1 U12536 ( .A(n11494), .ZN(n19115) );
  AND2_X1 U12537 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9723) );
  INV_X1 U12538 ( .A(n16905), .ZN(n9905) );
  NAND2_X1 U12539 ( .A1(n16101), .A2(n16091), .ZN(n9724) );
  INV_X1 U12540 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10037) );
  AND2_X1 U12541 ( .A1(n10995), .A2(n9723), .ZN(n9725) );
  INV_X1 U12542 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9852) );
  INV_X1 U12543 ( .A(n11610), .ZN(n10048) );
  INV_X1 U12544 ( .A(n16029), .ZN(n20106) );
  AOI22_X2 U12545 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9571), .B1(DATAI_28_), 
        .B2(n9570), .ZN(n20749) );
  AOI22_X2 U12546 ( .A1(DATAI_23_), .A2(n9570), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n9571), .ZN(n20701) );
  AOI22_X2 U12547 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9571), .B1(DATAI_27_), 
        .B2(n9570), .ZN(n20742) );
  AOI22_X2 U12548 ( .A1(DATAI_21_), .A2(n9570), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n9571), .ZN(n20685) );
  NOR3_X2 U12549 ( .A1(n18589), .A2(n18397), .A3(n18396), .ZN(n18366) );
  AOI22_X2 U12550 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9571), .B1(DATAI_30_), 
        .B2(n9570), .ZN(n20763) );
  AOI22_X2 U12551 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9571), .B1(DATAI_18_), 
        .B2(n9570), .ZN(n20667) );
  NOR3_X2 U12552 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18589), .A3(
        n18490), .ZN(n18460) );
  NOR3_X2 U12553 ( .A1(n18589), .A2(n18562), .A3(n18536), .ZN(n18530) );
  NOR2_X2 U12554 ( .A1(n18862), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18589) );
  AOI22_X2 U12555 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9571), .B1(DATAI_24_), 
        .B2(n9570), .ZN(n20721) );
  AOI22_X2 U12556 ( .A1(DATAI_17_), .A2(n9570), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9571), .ZN(n20661) );
  CLKBUF_X1 U12557 ( .A(n15948), .Z(n9726) );
  AND2_X2 U12558 ( .A1(n9727), .A2(n14627), .ZN(n11743) );
  AND2_X2 U12559 ( .A1(n9727), .A2(n13488), .ZN(n11664) );
  AND2_X1 U12560 ( .A1(n9727), .A2(n11633), .ZN(n11788) );
  NAND2_X1 U12561 ( .A1(n13364), .A2(n13363), .ZN(n9728) );
  OR2_X1 U12562 ( .A1(n9730), .A2(n9729), .ZN(n12764) );
  NOR2_X1 U12563 ( .A1(n13364), .A2(n9731), .ZN(n9729) );
  INV_X1 U12564 ( .A(n12758), .ZN(n9731) );
  XNOR2_X2 U12565 ( .A(n12757), .B(n13420), .ZN(n13364) );
  AND2_X1 U12566 ( .A1(n9734), .A2(n12858), .ZN(n13207) );
  NOR2_X1 U12567 ( .A1(n9734), .A2(n9733), .ZN(n9732) );
  INV_X1 U12568 ( .A(n13204), .ZN(n9733) );
  NAND2_X2 U12569 ( .A1(n13769), .A2(n12814), .ZN(n14522) );
  NAND2_X1 U12570 ( .A1(n9739), .A2(n12783), .ZN(n16017) );
  NAND2_X1 U12571 ( .A1(n16024), .A2(n16025), .ZN(n9739) );
  NAND3_X1 U12572 ( .A1(n9741), .A2(n9740), .A3(n9635), .ZN(n16024) );
  NAND3_X1 U12573 ( .A1(n13525), .A2(n13548), .A3(n13526), .ZN(n9740) );
  NAND2_X1 U12574 ( .A1(n9990), .A2(n13548), .ZN(n9741) );
  OAI21_X2 U12575 ( .B1(n14265), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11861), 
        .ZN(n12736) );
  NAND2_X2 U12576 ( .A1(n20157), .A2(n11876), .ZN(n14265) );
  OAI21_X1 U12577 ( .B1(n14549), .B2(n16204), .A(n9778), .ZN(P1_U3000) );
  OAI21_X1 U12578 ( .B1(n14549), .B2(n19920), .A(n12875), .ZN(P1_U2968) );
  AND2_X2 U12579 ( .A1(n10863), .A2(n10862), .ZN(n10876) );
  AND2_X1 U12580 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U12581 ( .A1(n9745), .A2(n19434), .ZN(n19438) );
  OAI22_X1 U12582 ( .A1(n10881), .A2(n10929), .B1(n14064), .B2(n9745), .ZN(
        n10933) );
  OAI22_X1 U12583 ( .A1(n10881), .A2(n10883), .B1(n10882), .B2(n9745), .ZN(
        n10888) );
  NAND3_X1 U12584 ( .A1(n9748), .A2(n10782), .A3(n9746), .ZN(n9941) );
  NAND2_X1 U12585 ( .A1(n9747), .A2(n9751), .ZN(n9746) );
  INV_X1 U12586 ( .A(n10785), .ZN(n9747) );
  NAND2_X1 U12587 ( .A1(n10792), .A2(n9751), .ZN(n9748) );
  NAND2_X1 U12588 ( .A1(n9752), .A2(n10760), .ZN(n9751) );
  INV_X1 U12589 ( .A(n10770), .ZN(n9749) );
  INV_X1 U12590 ( .A(n10769), .ZN(n9750) );
  NAND2_X1 U12591 ( .A1(n10786), .A2(n9751), .ZN(n10783) );
  NAND2_X1 U12592 ( .A1(n10784), .A2(n10785), .ZN(n10786) );
  INV_X1 U12593 ( .A(n9606), .ZN(n9752) );
  NAND3_X1 U12594 ( .A1(n10984), .A2(n9754), .A3(n11587), .ZN(n9753) );
  NOR2_X2 U12595 ( .A1(n15023), .A2(n11142), .ZN(n11572) );
  AOI21_X2 U12596 ( .B1(n15058), .B2(n15057), .A(n11126), .ZN(n15049) );
  NOR2_X2 U12597 ( .A1(n15209), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15076) );
  NAND3_X1 U12598 ( .A1(n11037), .A2(n10008), .A3(n11036), .ZN(n9758) );
  NAND3_X1 U12599 ( .A1(n9672), .A2(n10307), .A3(n9762), .ZN(n18269) );
  NOR2_X2 U12600 ( .A1(n18917), .A2(n16557), .ZN(n17915) );
  INV_X4 U12601 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18893) );
  NOR2_X2 U12602 ( .A1(n18162), .A2(n18277), .ZN(n18705) );
  INV_X1 U12603 ( .A(n9769), .ZN(n14507) );
  NAND3_X1 U12604 ( .A1(n11639), .A2(n9775), .A3(n9773), .ZN(n11695) );
  INV_X1 U12605 ( .A(n11626), .ZN(n9776) );
  NAND2_X1 U12606 ( .A1(n9781), .A2(n9780), .ZN(n9779) );
  NAND2_X1 U12607 ( .A1(n14415), .A2(n15975), .ZN(n9780) );
  NAND2_X1 U12608 ( .A1(n12868), .A2(n9782), .ZN(n9781) );
  INV_X1 U12609 ( .A(n11859), .ZN(n9783) );
  NAND2_X1 U12610 ( .A1(n9797), .A2(n13392), .ZN(n9796) );
  AND2_X2 U12611 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14627) );
  NAND2_X1 U12612 ( .A1(n20415), .A2(n20777), .ZN(n9804) );
  NAND2_X1 U12613 ( .A1(n11896), .A2(n11895), .ZN(n11946) );
  NAND2_X1 U12614 ( .A1(n11915), .A2(n20777), .ZN(n9807) );
  NOR3_X2 U12615 ( .A1(n10071), .A2(n18712), .A3(n10403), .ZN(n15738) );
  INV_X1 U12616 ( .A(n9817), .ZN(n17204) );
  NOR2_X2 U12617 ( .A1(n17090), .A2(n18299), .ZN(n17074) );
  INV_X2 U12618 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18878) );
  NOR2_X1 U12619 ( .A1(n17844), .A2(n10206), .ZN(n10207) );
  NAND2_X1 U12620 ( .A1(n9826), .A2(n9829), .ZN(n17701) );
  INV_X1 U12621 ( .A(n10212), .ZN(n9827) );
  NOR2_X2 U12622 ( .A1(n16429), .A2(n17928), .ZN(n16435) );
  NAND2_X1 U12623 ( .A1(n19102), .A2(n9838), .ZN(n9836) );
  NAND2_X1 U12624 ( .A1(n9839), .A2(n9836), .ZN(n14700) );
  OR2_X1 U12625 ( .A1(n11539), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9843) );
  NAND3_X1 U12626 ( .A1(n9843), .A2(n9842), .A3(n9841), .ZN(n13633) );
  NAND3_X1 U12627 ( .A1(n11539), .A2(n9844), .A3(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U12628 ( .A1(n14666), .A2(n9718), .ZN(n14667) );
  INV_X1 U12629 ( .A(n14667), .ZN(n11507) );
  NAND2_X1 U12631 ( .A1(n13815), .A2(n11587), .ZN(n9867) );
  NAND2_X1 U12632 ( .A1(n13815), .A2(n9863), .ZN(n9862) );
  NAND2_X1 U12633 ( .A1(n11037), .A2(n11036), .ZN(n9873) );
  AOI21_X1 U12634 ( .B1(n16949), .B2(n9891), .A(n16703), .ZN(n9887) );
  NAND2_X1 U12635 ( .A1(n16949), .A2(n9893), .ZN(n9888) );
  NAND2_X1 U12636 ( .A1(n9895), .A2(n9896), .ZN(n16650) );
  INV_X1 U12637 ( .A(n9898), .ZN(n16658) );
  XNOR2_X2 U12638 ( .A(n9899), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16949) );
  NAND2_X1 U12639 ( .A1(n9901), .A2(n9902), .ZN(n16680) );
  INV_X1 U12640 ( .A(n9904), .ZN(n16692) );
  NAND4_X1 U12641 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n9905), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16857) );
  NOR3_X1 U12642 ( .A1(n16918), .A2(n16606), .A3(n18767), .ZN(n9909) );
  NAND2_X1 U12643 ( .A1(n17622), .A2(n9700), .ZN(n16414) );
  NAND2_X1 U12644 ( .A1(n9913), .A2(n16293), .ZN(n11600) );
  NAND2_X1 U12645 ( .A1(n9913), .A2(n16338), .ZN(n9963) );
  NAND2_X1 U12646 ( .A1(n9921), .A2(n9919), .ZN(n11044) );
  NAND2_X1 U12647 ( .A1(n11118), .A2(n11119), .ZN(n11122) );
  NAND2_X1 U12648 ( .A1(n9934), .A2(n9933), .ZN(n13194) );
  AND2_X1 U12649 ( .A1(n14728), .A2(n14711), .ZN(n11530) );
  INV_X1 U12650 ( .A(n14154), .ZN(n9960) );
  INV_X2 U12651 ( .A(n11713), .ZN(n11658) );
  NAND4_X1 U12652 ( .A1(n10532), .A2(n10533), .A3(n10530), .A4(n10531), .ZN(
        n9965) );
  NAND4_X1 U12653 ( .A1(n10528), .A2(n10529), .A3(n10526), .A4(n10527), .ZN(
        n9967) );
  NAND2_X1 U12654 ( .A1(n9971), .A2(n9972), .ZN(n11350) );
  NOR2_X1 U12655 ( .A1(n9627), .A2(n11525), .ZN(n11484) );
  OR3_X1 U12656 ( .A1(n9627), .A2(n9976), .A3(n11525), .ZN(n11607) );
  INV_X1 U12657 ( .A(n11485), .ZN(n9981) );
  NAND2_X1 U12658 ( .A1(n14826), .A2(n9696), .ZN(n15397) );
  NAND2_X2 U12659 ( .A1(n9657), .A2(n11678), .ZN(n20134) );
  OAI211_X2 U12660 ( .C1(n14522), .C2(n9995), .A(n9994), .B(n14481), .ZN(
        n14480) );
  INV_X1 U12661 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11902) );
  NAND3_X1 U12662 ( .A1(n10003), .A2(n10004), .A3(n10083), .ZN(n10002) );
  INV_X1 U12663 ( .A(n15047), .ZN(n10005) );
  AOI21_X2 U12664 ( .B1(n10012), .B2(n9664), .A(n10006), .ZN(n15077) );
  NAND3_X2 U12665 ( .A1(n10876), .A2(n10878), .A3(n10877), .ZN(n10928) );
  INV_X1 U12666 ( .A(n13608), .ZN(n12040) );
  NAND3_X1 U12667 ( .A1(n13536), .A2(n13568), .A3(n13609), .ZN(n13608) );
  INV_X1 U12668 ( .A(n14238), .ZN(n10013) );
  NAND2_X1 U12669 ( .A1(n10013), .A2(n10014), .ZN(n14222) );
  INV_X1 U12670 ( .A(n13662), .ZN(n10017) );
  NAND2_X1 U12671 ( .A1(n10017), .A2(n9710), .ZN(n13759) );
  NAND2_X1 U12672 ( .A1(n11946), .A2(n11899), .ZN(n12749) );
  NAND2_X1 U12673 ( .A1(n14314), .A2(n10024), .ZN(n14208) );
  NOR2_X1 U12674 ( .A1(n14152), .A2(n14153), .ZN(n12843) );
  NAND3_X1 U12675 ( .A1(n13214), .A2(n11727), .A3(n13410), .ZN(n12888) );
  NAND2_X2 U12676 ( .A1(n10557), .A2(n10558), .ZN(n10703) );
  NAND3_X1 U12677 ( .A1(n10182), .A2(n10183), .A3(n10039), .ZN(n10038) );
  NAND2_X1 U12678 ( .A1(n10045), .A2(n17724), .ZN(n17726) );
  OR2_X2 U12679 ( .A1(n17579), .A2(n10218), .ZN(n16429) );
  NAND2_X1 U12680 ( .A1(n10962), .A2(n10961), .ZN(n10046) );
  NAND2_X1 U12681 ( .A1(n15544), .A2(n15537), .ZN(n10962) );
  NAND2_X1 U12682 ( .A1(n15033), .A2(n9648), .ZN(n11547) );
  AND2_X1 U12683 ( .A1(n15033), .A2(n10049), .ZN(n11521) );
  NAND2_X1 U12684 ( .A1(n15033), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15030) );
  NAND2_X2 U12685 ( .A1(n10443), .A2(n10442), .ZN(n10462) );
  NAND2_X1 U12686 ( .A1(n10053), .A2(n13156), .ZN(n13159) );
  XNOR2_X2 U12687 ( .A(n11163), .B(n11164), .ZN(n13151) );
  NAND3_X1 U12688 ( .A1(n9626), .A2(n14039), .A3(n9643), .ZN(n10054) );
  NAND2_X1 U12689 ( .A1(n14039), .A2(n14038), .ZN(n14851) );
  INV_X1 U12690 ( .A(n14853), .ZN(n10058) );
  AND2_X2 U12691 ( .A1(n14882), .A2(n9699), .ZN(n13938) );
  NAND2_X1 U12692 ( .A1(n11763), .A2(n20130), .ZN(n11772) );
  AOI21_X1 U12693 ( .B1(n9576), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n10248), .ZN(n10249) );
  AOI22_X1 U12694 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U12695 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  NAND2_X1 U12696 ( .A1(n15485), .A2(n13586), .ZN(n14820) );
  INV_X1 U12697 ( .A(n14820), .ZN(n11212) );
  INV_X1 U12698 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10456) );
  NOR3_X1 U12699 ( .A1(n15946), .A2(n13810), .A3(n20138), .ZN(n15948) );
  NAND2_X1 U12700 ( .A1(n11212), .A2(n11211), .ZN(n14818) );
  XNOR2_X1 U12701 ( .A(n11549), .B(n11548), .ZN(n14132) );
  INV_X1 U12702 ( .A(n13066), .ZN(n13064) );
  NAND2_X1 U12703 ( .A1(n10695), .A2(n13125), .ZN(n11279) );
  BUF_X1 U12704 ( .A(n15044), .Z(n15056) );
  NAND2_X1 U12705 ( .A1(n12896), .A2(n10063), .ZN(n12913) );
  NAND2_X1 U12706 ( .A1(n13065), .A2(n13064), .ZN(n13149) );
  INV_X1 U12707 ( .A(n13067), .ZN(n13065) );
  INV_X1 U12708 ( .A(n13151), .ZN(n10798) );
  AOI22_X1 U12709 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U12710 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U12711 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U12712 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10438) );
  OR2_X1 U12713 ( .A1(n12980), .A2(n12979), .ZN(n12981) );
  NAND2_X1 U12714 ( .A1(n12979), .A2(n12980), .ZN(n13063) );
  NOR2_X1 U12715 ( .A1(n15106), .A2(n15105), .ZN(n15107) );
  AOI21_X2 U12716 ( .B1(n15536), .B2(n15535), .A(n11028), .ZN(n15531) );
  OR2_X1 U12717 ( .A1(n18871), .A2(n18771), .ZN(n18911) );
  INV_X1 U12718 ( .A(n17556), .ZN(n17558) );
  AND2_X1 U12719 ( .A1(n18299), .A2(n17291), .ZN(n17295) );
  AND2_X1 U12720 ( .A1(n14405), .A2(n13810), .ZN(n10063) );
  NOR2_X1 U12721 ( .A1(n14613), .A2(n13427), .ZN(n16171) );
  OR2_X1 U12722 ( .A1(n13614), .A2(n12730), .ZN(n15883) );
  INV_X1 U12723 ( .A(n12741), .ZN(n20107) );
  AND2_X1 U12724 ( .A1(n14011), .A2(n10076), .ZN(n10064) );
  AND2_X1 U12725 ( .A1(n14699), .A2(n16333), .ZN(n10065) );
  INV_X1 U12726 ( .A(n13704), .ZN(n11192) );
  INV_X1 U12727 ( .A(n11318), .ZN(n11383) );
  AND2_X1 U12728 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10066) );
  AND2_X1 U12729 ( .A1(n10580), .A2(n10579), .ZN(n10067) );
  AND4_X1 U12730 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10068) );
  OR2_X1 U12731 ( .A1(n12712), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10069) );
  AND4_X1 U12732 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10070) );
  OR2_X1 U12733 ( .A1(n18280), .A2(n17307), .ZN(n10071) );
  INV_X1 U12734 ( .A(n13705), .ZN(n11191) );
  OR2_X1 U12735 ( .A1(n14848), .A2(n13376), .ZN(n10072) );
  AND2_X1 U12736 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10073) );
  INV_X1 U12737 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20856) );
  OR2_X1 U12738 ( .A1(n12712), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10074) );
  INV_X1 U12739 ( .A(n14411), .ZN(n15950) );
  AND4_X1 U12740 ( .A1(n10146), .A2(n10145), .A3(n10144), .A4(n10143), .ZN(
        n10075) );
  AND2_X1 U12741 ( .A1(n14010), .A2(n14034), .ZN(n10076) );
  INV_X1 U12742 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19941) );
  INV_X1 U12743 ( .A(n20869), .ZN(n20868) );
  INV_X1 U12744 ( .A(n10128), .ZN(n10357) );
  OR2_X1 U12745 ( .A1(n12712), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10077) );
  INV_X1 U12746 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U12747 ( .A1(n11516), .A2(n14062), .ZN(n16308) );
  INV_X1 U12748 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12386) );
  OR2_X1 U12749 ( .A1(n13287), .A2(n11757), .ZN(n13334) );
  NAND2_X1 U12750 ( .A1(n10730), .A2(n10729), .ZN(n13779) );
  INV_X1 U12751 ( .A(n20716), .ZN(n20635) );
  AND2_X1 U12752 ( .A1(n10745), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10078) );
  NOR3_X1 U12753 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18731), .ZN(n10255) );
  NAND2_X1 U12754 ( .A1(n20014), .A2(n13810), .ZN(n14358) );
  AND3_X1 U12755 ( .A1(n20559), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10079) );
  INV_X1 U12756 ( .A(n11033), .ZN(n10961) );
  INV_X1 U12757 ( .A(n11664), .ZN(n12480) );
  AND2_X1 U12758 ( .A1(n11660), .A2(n11659), .ZN(n10081) );
  AND4_X1 U12759 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n10082) );
  OR3_X1 U12760 ( .A1(n12601), .A2(n12600), .A3(n12599), .ZN(n12602) );
  NAND2_X1 U12761 ( .A1(n13392), .A2(n20138), .ZN(n11663) );
  INV_X1 U12762 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11672) );
  INV_X1 U12763 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10508) );
  INV_X1 U12764 ( .A(n11789), .ZN(n12534) );
  OR2_X1 U12765 ( .A1(n11993), .A2(n11992), .ZN(n12785) );
  INV_X1 U12766 ( .A(n13987), .ZN(n13988) );
  INV_X1 U12767 ( .A(n12584), .ZN(n12577) );
  INV_X1 U12768 ( .A(n14360), .ZN(n12117) );
  INV_X1 U12769 ( .A(n14236), .ZN(n12101) );
  AOI21_X1 U12770 ( .B1(n11712), .B2(n20126), .A(n13810), .ZN(n11710) );
  NAND2_X1 U12771 ( .A1(n11335), .A2(n14062), .ZN(n10826) );
  INV_X1 U12772 ( .A(n10731), .ZN(n10745) );
  NOR2_X1 U12773 ( .A1(n9649), .A2(n17282), .ZN(n10119) );
  NAND2_X1 U12774 ( .A1(n10395), .A2(n10397), .ZN(n10319) );
  NOR2_X1 U12775 ( .A1(n12573), .A2(n12572), .ZN(n12608) );
  INV_X1 U12776 ( .A(n14330), .ZN(n12237) );
  INV_X1 U12777 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11948) );
  INV_X1 U12778 ( .A(n12029), .ZN(n12030) );
  OR2_X1 U12779 ( .A1(n11968), .A2(n11967), .ZN(n12777) );
  OR2_X1 U12780 ( .A1(n11854), .A2(n11864), .ZN(n11874) );
  INV_X1 U12781 ( .A(n19142), .ZN(n13828) );
  INV_X1 U12782 ( .A(n13964), .ZN(n13937) );
  OR2_X1 U12783 ( .A1(n10957), .A2(n10956), .ZN(n11029) );
  INV_X1 U12784 ( .A(n13196), .ZN(n11179) );
  NAND2_X1 U12785 ( .A1(n10925), .A2(n10924), .ZN(n15538) );
  NAND2_X1 U12786 ( .A1(n19258), .A2(n10795), .ZN(n10796) );
  OAI21_X1 U12787 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18878), .A(
        n10330), .ZN(n10331) );
  AOI21_X1 U12788 ( .B1(n17250), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n10119), .ZN(n10120) );
  AND2_X1 U12789 ( .A1(n12609), .A2(n12803), .ZN(n12606) );
  INV_X1 U12790 ( .A(n14347), .ZN(n12178) );
  INV_X1 U12791 ( .A(n12520), .ZN(n12556) );
  NAND2_X1 U12792 ( .A1(n20138), .A2(n11764), .ZN(n11712) );
  OR2_X1 U12793 ( .A1(n10464), .A2(n10463), .ZN(n10465) );
  NAND2_X1 U12794 ( .A1(n10448), .A2(n16349), .ZN(n10455) );
  XNOR2_X1 U12795 ( .A(n13986), .B(n13987), .ZN(n14862) );
  INV_X1 U12796 ( .A(n15011), .ZN(n11589) );
  AND4_X1 U12797 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10980) );
  INV_X1 U12798 ( .A(n15221), .ZN(n16288) );
  INV_X1 U12799 ( .A(n11317), .ZN(n11382) );
  OR2_X1 U12800 ( .A1(n11299), .A2(n11298), .ZN(n13181) );
  INV_X1 U12801 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15678) );
  INV_X1 U12802 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17157) );
  INV_X1 U12803 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20941) );
  INV_X1 U12804 ( .A(n10124), .ZN(n10125) );
  INV_X1 U12805 ( .A(n16433), .ZN(n10219) );
  NOR2_X1 U12806 ( .A1(n10357), .A2(n10192), .ZN(n10177) );
  OAI21_X1 U12807 ( .B1(n10397), .B2(n10391), .A(n10390), .ZN(n10404) );
  INV_X1 U12808 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17225) );
  INV_X1 U12809 ( .A(n12706), .ZN(n12717) );
  OR2_X1 U12810 ( .A1(n12150), .A2(n15914), .ZN(n12157) );
  INV_X1 U12811 ( .A(n12381), .ZN(n12422) );
  NOR2_X1 U12812 ( .A1(n14623), .A2(n20777), .ZN(n12520) );
  INV_X1 U12813 ( .A(n12093), .ZN(n12192) );
  AND2_X1 U12814 ( .A1(n20376), .A2(n20408), .ZN(n20382) );
  AND2_X1 U12815 ( .A1(n20519), .A2(n20551), .ZN(n20523) );
  AND2_X1 U12816 ( .A1(n13485), .A2(n13484), .ZN(n15758) );
  INV_X1 U12817 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15155) );
  INV_X1 U12818 ( .A(n14819), .ZN(n11211) );
  AND2_X1 U12819 ( .A1(n11477), .A2(n11476), .ZN(n14751) );
  AND2_X1 U12820 ( .A1(n11469), .A2(n11468), .ZN(n15329) );
  INV_X1 U12821 ( .A(n11382), .ZN(n11357) );
  NOR2_X1 U12822 ( .A1(n9605), .A2(n11152), .ZN(n11154) );
  INV_X1 U12823 ( .A(n15293), .ZN(n10995) );
  OR2_X1 U12824 ( .A1(n15565), .A2(n15567), .ZN(n15411) );
  NOR2_X1 U12825 ( .A1(n15467), .A2(n15491), .ZN(n15445) );
  OAI21_X1 U12826 ( .B1(n11321), .B2(n11316), .A(n9690), .ZN(n13129) );
  AND2_X1 U12827 ( .A1(n10678), .A2(n10712), .ZN(n10486) );
  INV_X1 U12828 ( .A(n10216), .ZN(n10217) );
  AOI211_X1 U12829 ( .C1(n18287), .C2(n18722), .A(n10403), .B(n10315), .ZN(
        n10327) );
  AOI21_X1 U12830 ( .B1(n15740), .B2(n16575), .A(n16574), .ZN(n15733) );
  INV_X2 U12831 ( .A(n9649), .ZN(n17258) );
  AND2_X1 U12832 ( .A1(n12179), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12199) );
  NOR2_X1 U12833 ( .A1(n12157), .A2(n14247), .ZN(n12179) );
  NAND2_X1 U12834 ( .A1(n11928), .A2(n11927), .ZN(n20270) );
  INV_X1 U12835 ( .A(n20862), .ZN(n13614) );
  NAND2_X1 U12836 ( .A1(n12472), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12524) );
  NAND2_X1 U12837 ( .A1(n12423), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12471) );
  INV_X1 U12838 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U12839 ( .A1(n12199), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12200) );
  INV_X1 U12840 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15914) );
  OR2_X1 U12841 ( .A1(n12059), .A2(n19948), .ZN(n12090) );
  NOR2_X1 U12842 ( .A1(n12002), .A2(n12001), .ZN(n12023) );
  INV_X1 U12843 ( .A(n20635), .ZN(n20377) );
  CLKBUF_X3 U12844 ( .A(n12831), .Z(n15955) );
  AND2_X1 U12845 ( .A1(n12692), .A2(n12691), .ZN(n14308) );
  NOR2_X1 U12846 ( .A1(n20566), .A2(n13395), .ZN(n15785) );
  AND2_X1 U12847 ( .A1(n20236), .A2(n20235), .ZN(n20240) );
  AND2_X1 U12848 ( .A1(n20274), .A2(n20273), .ZN(n20302) );
  AND2_X1 U12849 ( .A1(n20380), .A2(n20379), .ZN(n20407) );
  NOR2_X1 U12850 ( .A1(n20639), .A2(n20279), .ZN(n20484) );
  AOI21_X1 U12851 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20601), .A(n20279), 
        .ZN(n20715) );
  OAI22_X1 U12852 ( .A1(n16375), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n10483), .B2(n10482), .ZN(n10678) );
  OR2_X1 U12853 ( .A1(n21033), .A2(n13644), .ZN(n19096) );
  AND3_X1 U12854 ( .A1(n11370), .A2(n11369), .A3(n11368), .ZN(n13713) );
  INV_X1 U12855 ( .A(n19115), .ZN(n19088) );
  NOR2_X1 U12856 ( .A1(n11099), .A2(n15339), .ZN(n15093) );
  OR2_X1 U12857 ( .A1(n19016), .A2(n11105), .ZN(n15162) );
  OR2_X1 U12858 ( .A1(n10984), .A2(n11041), .ZN(n10991) );
  NOR2_X1 U12859 ( .A1(n10514), .A2(n10486), .ZN(n16367) );
  INV_X1 U12860 ( .A(n19318), .ZN(n15609) );
  OR2_X1 U12861 ( .A1(n19877), .A2(n19887), .ZN(n13377) );
  INV_X1 U12862 ( .A(n13377), .ZN(n19433) );
  OR2_X1 U12863 ( .A1(n19877), .A2(n19278), .ZN(n19720) );
  AOI21_X1 U12864 ( .B1(n10343), .B2(n10347), .A(n10342), .ZN(n10350) );
  NOR2_X1 U12865 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16727), .ZN(n16714) );
  NOR2_X1 U12866 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16749), .ZN(n16736) );
  NOR2_X1 U12867 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16800), .ZN(n16783) );
  NOR2_X1 U12868 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16872), .ZN(n16850) );
  INV_X1 U12869 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15687) );
  NAND2_X1 U12870 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10138) );
  INV_X1 U12871 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17741) );
  NAND2_X1 U12872 ( .A1(n17755), .A2(n17922), .ZN(n17702) );
  NAND2_X1 U12873 ( .A1(n17614), .A2(n17974), .ZN(n17613) );
  NOR2_X1 U12874 ( .A1(n18078), .A2(n17749), .ZN(n18065) );
  INV_X1 U12875 ( .A(n18203), .ZN(n18222) );
  INV_X1 U12876 ( .A(n18101), .ZN(n18125) );
  OAI21_X1 U12877 ( .B1(n10193), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n17885), .ZN(n17879) );
  NOR2_X1 U12878 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20716) );
  INV_X1 U12879 ( .A(n19954), .ZN(n12623) );
  INV_X1 U12880 ( .A(n14142), .ZN(n14143) );
  NAND2_X1 U12881 ( .A1(n14333), .A2(n14324), .ZN(n14326) );
  INV_X1 U12882 ( .A(n14358), .ZN(n12863) );
  AND2_X1 U12883 ( .A1(n12524), .A2(n12474), .ZN(n14443) );
  INV_X1 U12884 ( .A(n14384), .ZN(n15848) );
  INV_X1 U12885 ( .A(n14394), .ZN(n15887) );
  NAND2_X1 U12886 ( .A1(n12096), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12150) );
  INV_X1 U12887 ( .A(n16033), .ZN(n20085) );
  INV_X1 U12888 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12873) );
  INV_X1 U12889 ( .A(n15814), .ZN(n16063) );
  INV_X1 U12890 ( .A(n16204), .ZN(n20094) );
  NAND2_X1 U12891 ( .A1(n20777), .A2(n20108), .ZN(n20279) );
  NOR2_X1 U12892 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16214) );
  OAI22_X1 U12893 ( .A1(n20120), .A2(n20119), .B1(n20487), .B2(n20118), .ZN(
        n20152) );
  OAI22_X1 U12894 ( .A1(n20198), .A2(n20197), .B1(n20487), .B2(n20345), .ZN(
        n20221) );
  NAND2_X1 U12895 ( .A1(n12759), .A2(n12749), .ZN(n20227) );
  INV_X1 U12896 ( .A(n20276), .ZN(n20305) );
  INV_X1 U12897 ( .A(n20369), .ZN(n20335) );
  NOR2_X1 U12898 ( .A1(n12749), .A2(n13576), .ZN(n20385) );
  INV_X1 U12899 ( .A(n20511), .ZN(n20479) );
  INV_X1 U12900 ( .A(n20318), .ZN(n20611) );
  INV_X1 U12901 ( .A(n20557), .ZN(n20544) );
  OAI22_X1 U12902 ( .A1(n20572), .A2(n20571), .B1(n20570), .B2(n20569), .ZN(
        n20595) );
  INV_X1 U12903 ( .A(n20269), .ZN(n20558) );
  AND2_X1 U12904 ( .A1(n20633), .A2(n20611), .ZN(n20697) );
  AND2_X1 U12905 ( .A1(n20633), .A2(n20527), .ZN(n20770) );
  AND2_X1 U12906 ( .A1(n20776), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15781) );
  INV_X1 U12907 ( .A(n20839), .ZN(n20833) );
  INV_X1 U12908 ( .A(n19084), .ZN(n19109) );
  AND2_X1 U12909 ( .A1(n14111), .A2(n14109), .ZN(n19165) );
  AND3_X1 U12910 ( .A1(n11398), .A2(n11397), .A3(n11396), .ZN(n15490) );
  OR2_X1 U12911 ( .A1(n14111), .A2(n19164), .ZN(n19198) );
  INV_X1 U12912 ( .A(n13647), .ZN(n13078) );
  INV_X1 U12913 ( .A(n16308), .ZN(n11517) );
  AND2_X1 U12914 ( .A1(n16315), .A2(n12993), .ZN(n16305) );
  AND2_X1 U12915 ( .A1(n15085), .A2(n15086), .ZN(n15140) );
  AND2_X1 U12916 ( .A1(n19087), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16282) );
  AND2_X1 U12917 ( .A1(n10688), .A2(n19777), .ZN(n11308) );
  AND2_X1 U12918 ( .A1(n11308), .A2(n11296), .ZN(n11300) );
  INV_X1 U12919 ( .A(n19264), .ZN(n16319) );
  NOR2_X2 U12920 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19869) );
  NOR2_X1 U12921 ( .A1(n16367), .A2(n19678), .ZN(n15594) );
  INV_X1 U12922 ( .A(n19323), .ZN(n19340) );
  AND2_X1 U12923 ( .A1(n19877), .A2(n19278), .ZN(n19318) );
  OAI21_X1 U12924 ( .B1(n19383), .B2(n19382), .A(n19381), .ZN(n19401) );
  AND2_X1 U12925 ( .A1(n19462), .A2(n19433), .ZN(n19457) );
  AND2_X1 U12926 ( .A1(n19494), .A2(n19433), .ZN(n19489) );
  INV_X1 U12927 ( .A(n19493), .ZN(n19521) );
  NOR2_X1 U12928 ( .A1(n19871), .A2(n19894), .ZN(n19494) );
  NOR2_X2 U12929 ( .A1(n19674), .A2(n15609), .ZN(n19572) );
  AND2_X1 U12930 ( .A1(n19279), .A2(n19318), .ZN(n19584) );
  INV_X1 U12931 ( .A(n19726), .ZN(n19680) );
  AND2_X1 U12932 ( .A1(n19877), .A2(n19887), .ZN(n19865) );
  AND2_X1 U12933 ( .A1(n13379), .A2(n13378), .ZN(n19669) );
  INV_X1 U12934 ( .A(n19564), .ZN(n19742) );
  INV_X1 U12935 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19676) );
  AND3_X1 U12936 ( .A1(n19791), .A2(n19855), .A3(n19796), .ZN(n21041) );
  INV_X1 U12937 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19791) );
  NOR2_X1 U12938 ( .A1(n18703), .A2(n17458), .ZN(n18914) );
  NOR2_X1 U12939 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16704), .ZN(n16691) );
  NOR2_X1 U12940 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16821), .ZN(n16809) );
  NOR2_X1 U12941 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16842), .ZN(n16827) );
  NOR2_X1 U12942 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16892), .ZN(n16876) );
  NOR2_X2 U12943 ( .A1(n18862), .A2(n16961), .ZN(n16900) );
  NOR2_X1 U12944 ( .A1(n17505), .A2(n17368), .ZN(n17362) );
  NOR2_X1 U12945 ( .A1(n18299), .A2(n17380), .ZN(n17374) );
  AOI21_X1 U12947 ( .B1(n17578), .B2(n17928), .A(n17563), .ZN(n12885) );
  NOR2_X1 U12948 ( .A1(n10385), .A2(n17829), .ZN(n18123) );
  NAND2_X1 U12949 ( .A1(n17702), .A2(n17780), .ZN(n17914) );
  NOR2_X1 U12950 ( .A1(n17580), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17579) );
  INV_X1 U12951 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18113) );
  NOR2_X1 U12952 ( .A1(n9587), .A2(n18238), .ZN(n18211) );
  INV_X1 U12953 ( .A(n18564), .ZN(n18372) );
  NOR2_X1 U12954 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18862), .ZN(
        n18887) );
  INV_X1 U12955 ( .A(n18395), .ZN(n18461) );
  INV_X1 U12956 ( .A(n18442), .ZN(n18508) );
  INV_X1 U12957 ( .A(n18487), .ZN(n18554) );
  AND2_X1 U12958 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18648), .ZN(n18679) );
  INV_X1 U12959 ( .A(n14110), .ZN(n13375) );
  NOR2_X1 U12960 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12927), .ZN(n16533)
         );
  NAND3_X1 U12961 ( .A1(n13390), .A2(n13411), .A3(n13399), .ZN(n13287) );
  NAND2_X1 U12962 ( .A1(n12957), .A2(n13287), .ZN(n20862) );
  NAND2_X1 U12963 ( .A1(n14143), .A2(n12623), .ZN(n14151) );
  NAND2_X1 U12964 ( .A1(n15872), .A2(n13602), .ZN(n19974) );
  NAND2_X1 U12965 ( .A1(n15872), .A2(n12622), .ZN(n19954) );
  INV_X1 U12966 ( .A(n19977), .ZN(n20005) );
  AND2_X1 U12967 ( .A1(n13600), .A2(n19954), .ZN(n19990) );
  OR2_X1 U12968 ( .A1(n15946), .A2(n12908), .ZN(n15953) );
  OR2_X1 U12969 ( .A1(n14356), .A2(n14355), .ZN(n15999) );
  INV_X1 U12970 ( .A(n20015), .ZN(n20046) );
  NOR2_X1 U12971 ( .A1(n13287), .A2(n13286), .ZN(n13330) );
  INV_X1 U12972 ( .A(n16027), .ZN(n16023) );
  INV_X1 U12973 ( .A(n20087), .ZN(n19920) );
  INV_X1 U12974 ( .A(n20093), .ZN(n16159) );
  OR2_X1 U12975 ( .A1(n20227), .A2(n20269), .ZN(n20183) );
  OR2_X1 U12976 ( .A1(n20227), .A2(n20318), .ZN(n20225) );
  OR2_X1 U12977 ( .A1(n20227), .A2(n20226), .ZN(n20276) );
  NAND2_X1 U12978 ( .A1(n20385), .A2(n20558), .ZN(n20339) );
  NAND2_X1 U12979 ( .A1(n20385), .A2(n20611), .ZN(n20369) );
  NAND2_X1 U12980 ( .A1(n20385), .A2(n20632), .ZN(n20406) );
  NAND2_X1 U12981 ( .A1(n20528), .A2(n20558), .ZN(n20475) );
  NAND2_X1 U12982 ( .A1(n20528), .A2(n20611), .ZN(n20511) );
  NAND2_X1 U12983 ( .A1(n20528), .A2(n20632), .ZN(n20557) );
  NAND2_X1 U12984 ( .A1(n20528), .A2(n20527), .ZN(n20599) );
  NAND2_X1 U12985 ( .A1(n20633), .A2(n20558), .ZN(n20631) );
  NAND2_X1 U12986 ( .A1(n20633), .A2(n20632), .ZN(n20774) );
  INV_X1 U12987 ( .A(n20845), .ZN(n20780) );
  INV_X1 U12988 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20970) );
  OR2_X1 U12989 ( .A1(n20794), .A2(n20869), .ZN(n20835) );
  AND2_X1 U12990 ( .A1(n12934), .A2(n16360), .ZN(n21033) );
  INV_X1 U12991 ( .A(n19122), .ZN(n19090) );
  NAND2_X1 U12992 ( .A1(n21033), .A2(n13640), .ZN(n19127) );
  INV_X1 U12993 ( .A(n19214), .ZN(n19173) );
  AND2_X1 U12994 ( .A1(n13124), .A2(n19777), .ZN(n19196) );
  AND2_X1 U12995 ( .A1(n19173), .A2(n19218), .ZN(n19205) );
  INV_X1 U12996 ( .A(n19198), .ZN(n19222) );
  INV_X1 U12997 ( .A(n19224), .ZN(n19254) );
  NAND2_X1 U12998 ( .A1(n13649), .A2(n14062), .ZN(n13647) );
  INV_X1 U12999 ( .A(n16305), .ZN(n16304) );
  INV_X1 U13000 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16314) );
  NAND2_X1 U13001 ( .A1(n11308), .A2(n16359), .ZN(n19264) );
  INV_X1 U13002 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16375) );
  NAND2_X1 U13003 ( .A1(n19318), .A2(n19462), .ZN(n19323) );
  NAND2_X1 U13004 ( .A1(n19318), .A2(n19494), .ZN(n19373) );
  INV_X1 U13005 ( .A(n19429), .ZN(n19399) );
  INV_X1 U13006 ( .A(n19457), .ZN(n19456) );
  INV_X1 U13007 ( .A(n19489), .ZN(n19486) );
  NAND2_X1 U13008 ( .A1(n19495), .A2(n19494), .ZN(n19555) );
  INV_X1 U13009 ( .A(n19584), .ZN(n19606) );
  INV_X1 U13010 ( .A(n19617), .ZN(n19627) );
  NAND2_X1 U13011 ( .A1(n19279), .A2(n19865), .ZN(n19651) );
  INV_X1 U13012 ( .A(n19670), .ZN(n19668) );
  INV_X1 U13013 ( .A(n19707), .ZN(n19705) );
  INV_X1 U13014 ( .A(n19755), .ZN(n19775) );
  INV_X1 U13015 ( .A(n19864), .ZN(n19785) );
  NAND2_X1 U13016 ( .A1(n19791), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19910) );
  NOR2_X1 U13017 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16687), .ZN(n16678) );
  INV_X1 U13018 ( .A(n16965), .ZN(n16953) );
  INV_X1 U13019 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17264) );
  INV_X1 U13020 ( .A(n16439), .ZN(n17427) );
  NAND2_X1 U13021 ( .A1(n17476), .A2(n18269), .ZN(n17474) );
  INV_X1 U13022 ( .A(n17476), .ZN(n17494) );
  AOI21_X1 U13023 ( .B1(n16639), .B2(n17565), .A(n12885), .ZN(n12886) );
  OR2_X1 U13024 ( .A1(n17723), .A2(n17989), .ZN(n17690) );
  NAND2_X1 U13025 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17919), .ZN(n17780) );
  INV_X1 U13026 ( .A(n17914), .ZN(n17905) );
  OR2_X1 U13027 ( .A1(n18372), .A2(n18513), .ZN(n18587) );
  INV_X1 U13028 ( .A(n9572), .ZN(n18144) );
  INV_X1 U13029 ( .A(n18211), .ZN(n18239) );
  INV_X1 U13030 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18397) );
  INV_X1 U13031 ( .A(n18693), .ZN(n18584) );
  INV_X1 U13032 ( .A(n18858), .ZN(n18772) );
  INV_X1 U13033 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18787) );
  OAI21_X1 U13034 ( .B1(n14367), .B2(n14364), .A(n12865), .ZN(P1_U2842) );
  OAI211_X1 U13035 ( .C1(n15010), .C2(n19264), .A(n11624), .B(n11623), .ZN(
        P2_U3016) );
  NAND2_X1 U13036 ( .A1(n12887), .A2(n12886), .ZN(P3_U2803) );
  INV_X2 U13037 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18868) );
  INV_X1 U13038 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20949) );
  INV_X1 U13039 ( .A(n10093), .ZN(n10084) );
  AOI22_X1 U13040 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U13041 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10089) );
  NOR3_X2 U13042 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n10087), .ZN(n10141) );
  BUF_X4 U13043 ( .A(n10141), .Z(n17251) );
  AOI22_X1 U13044 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10088) );
  OAI211_X1 U13045 ( .C1(n9649), .C2(n17264), .A(n10089), .B(n10088), .ZN(
        n10099) );
  AOI22_X1 U13046 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10097) );
  INV_X2 U13047 ( .A(n9652), .ZN(n17171) );
  AOI22_X1 U13048 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10096) );
  NAND2_X2 U13049 ( .A1(n18868), .A2(n10093), .ZN(n17199) );
  AOI22_X1 U13050 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10142), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U13051 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10094) );
  NAND4_X1 U13052 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n10098) );
  AOI211_X1 U13053 ( .C1(n9622), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n10099), .B(n10098), .ZN(n10100) );
  OAI211_X1 U13054 ( .C1(n17148), .C2(n20949), .A(n10101), .B(n10100), .ZN(
        n16439) );
  INV_X1 U13055 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15700) );
  INV_X2 U13056 ( .A(n17148), .ZN(n17108) );
  AOI22_X1 U13057 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10103) );
  OAI21_X1 U13058 ( .B1(n17156), .B2(n15700), .A(n10103), .ZN(n10112) );
  INV_X1 U13059 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U13060 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10110) );
  INV_X1 U13061 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U13062 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10104) );
  OAI21_X1 U13063 ( .B1(n9616), .B2(n17059), .A(n10104), .ZN(n10108) );
  INV_X1 U13064 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U13065 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U13066 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10105) );
  OAI211_X1 U13067 ( .C1(n9649), .C2(n17275), .A(n10106), .B(n10105), .ZN(
        n10107) );
  AOI211_X1 U13068 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n10108), .B(n10107), .ZN(n10109) );
  OAI211_X1 U13069 ( .C1(n17224), .C2(n15699), .A(n10110), .B(n10109), .ZN(
        n10111) );
  INV_X1 U13070 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18605) );
  AOI22_X1 U13071 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10114) );
  OAI21_X1 U13072 ( .B1(n9651), .B2(n18605), .A(n10114), .ZN(n10118) );
  INV_X1 U13073 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U13074 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U13075 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10115) );
  OAI211_X1 U13076 ( .C1(n9616), .C2(n17079), .A(n10116), .B(n10115), .ZN(
        n10117) );
  AOI211_X1 U13077 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n10118), .B(n10117), .ZN(n10127) );
  AOI22_X1 U13078 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10142), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10121) );
  INV_X1 U13079 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17282) );
  INV_X1 U13080 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U13081 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10122) );
  OAI21_X1 U13082 ( .B1(n9652), .B2(n10123), .A(n10122), .ZN(n10124) );
  NAND3_X1 U13083 ( .A1(n10127), .A2(n10126), .A3(n10125), .ZN(n10128) );
  INV_X1 U13084 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U13085 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10130) );
  OAI211_X1 U13086 ( .C1(n9649), .C2(n17289), .A(n10130), .B(n10129), .ZN(
        n10137) );
  AOI22_X1 U13087 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U13088 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U13089 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U13090 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10132) );
  NAND4_X1 U13091 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10136) );
  INV_X2 U13092 ( .A(n9652), .ZN(n17207) );
  AOI22_X1 U13093 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U13094 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10231), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17211), .ZN(n10146) );
  AOI22_X1 U13095 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10141), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10178), .ZN(n10145) );
  AOI22_X1 U13096 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10142), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U13097 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10143) );
  AOI22_X1 U13098 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17244), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10155) );
  INV_X1 U13099 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17290) );
  AOI22_X1 U13100 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17108), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17243), .ZN(n10149) );
  AOI22_X1 U13101 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17171), .ZN(n10148) );
  OAI211_X1 U13102 ( .C1(n9649), .C2(n17290), .A(n10149), .B(n10148), .ZN(
        n10153) );
  INV_X1 U13104 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17106) );
  NAND2_X1 U13105 ( .A1(n9833), .A2(n17449), .ZN(n10192) );
  INV_X1 U13106 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U13107 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10165) );
  INV_X1 U13108 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U13109 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13110 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10156) );
  OAI211_X1 U13111 ( .C1(n9649), .C2(n17279), .A(n10157), .B(n10156), .ZN(
        n10163) );
  AOI22_X1 U13112 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13113 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13114 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10142), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U13115 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10158) );
  NAND4_X1 U13116 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        n10162) );
  AOI211_X1 U13117 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n10163), .B(n10162), .ZN(n10164) );
  OAI211_X1 U13118 ( .C1(n9612), .C2(n17182), .A(n10165), .B(n10164), .ZN(
        n10176) );
  NAND2_X1 U13119 ( .A1(n10177), .A2(n10176), .ZN(n10196) );
  AOI22_X1 U13120 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10175) );
  INV_X1 U13121 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U13122 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13123 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10166) );
  OAI211_X1 U13124 ( .C1(n9616), .C2(n17155), .A(n10167), .B(n10166), .ZN(
        n10173) );
  AOI22_X1 U13125 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13126 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13127 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U13128 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10168) );
  NAND4_X1 U13129 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10172) );
  AOI211_X1 U13130 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10173), .B(n10172), .ZN(n10174) );
  OAI211_X1 U13131 ( .C1(n9649), .C2(n17269), .A(n10175), .B(n10174), .ZN(
        n10200) );
  NAND2_X1 U13132 ( .A1(n10201), .A2(n10200), .ZN(n16436) );
  INV_X1 U13133 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17928) );
  INV_X1 U13134 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20894) );
  INV_X1 U13135 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18059) );
  INV_X1 U13136 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18177) );
  INV_X1 U13137 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17861) );
  INV_X1 U13138 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18204) );
  INV_X1 U13139 ( .A(n10176), .ZN(n17438) );
  XNOR2_X1 U13140 ( .A(n17438), .B(n10177), .ZN(n10194) );
  XOR2_X1 U13141 ( .A(n18204), .B(n10194), .Z(n17880) );
  INV_X1 U13142 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18872) );
  NOR2_X1 U13143 ( .A1(n17449), .A2(n18872), .ZN(n10187) );
  XNOR2_X1 U13144 ( .A(n18872), .B(n17449), .ZN(n17913) );
  INV_X1 U13145 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20973) );
  AOI22_X1 U13146 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10186) );
  INV_X1 U13147 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20925) );
  AOI22_X1 U13148 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13149 ( .A1(n10178), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10179) );
  OAI211_X1 U13150 ( .C1(n9649), .C2(n20925), .A(n10180), .B(n10179), .ZN(
        n10184) );
  AOI22_X1 U13151 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13152 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10231), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13153 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U13154 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17921), .ZN(
        n17920) );
  NOR2_X1 U13155 ( .A1(n17913), .A2(n17920), .ZN(n17912) );
  NOR2_X1 U13156 ( .A1(n10187), .A2(n17912), .ZN(n17902) );
  INV_X1 U13157 ( .A(n17902), .ZN(n10191) );
  INV_X1 U13158 ( .A(n17903), .ZN(n10190) );
  INV_X1 U13159 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18235) );
  NOR2_X1 U13160 ( .A1(n18235), .A2(n10188), .ZN(n10189) );
  XNOR2_X1 U13161 ( .A(n10357), .B(n10192), .ZN(n17887) );
  NOR2_X1 U13162 ( .A1(n17886), .A2(n17887), .ZN(n10193) );
  NAND2_X1 U13163 ( .A1(n17886), .A2(n17887), .ZN(n17885) );
  NOR2_X1 U13164 ( .A1(n17880), .A2(n17879), .ZN(n17878) );
  AND2_X1 U13165 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10194), .ZN(
        n10195) );
  XNOR2_X1 U13166 ( .A(n17434), .B(n10196), .ZN(n10197) );
  NOR2_X1 U13167 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  INV_X1 U13168 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18178) );
  INV_X1 U13169 ( .A(n10200), .ZN(n17430) );
  XNOR2_X1 U13170 ( .A(n17430), .B(n10201), .ZN(n10202) );
  XOR2_X1 U13171 ( .A(n18178), .B(n10202), .Z(n17849) );
  AOI21_X1 U13172 ( .B1(n16436), .B2(n17427), .A(n17833), .ZN(n10203) );
  INV_X1 U13173 ( .A(n10203), .ZN(n10204) );
  NOR2_X1 U13174 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  INV_X1 U13175 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18165) );
  INV_X1 U13176 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18078) );
  INV_X1 U13177 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18155) );
  INV_X1 U13178 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18138) );
  NOR2_X1 U13179 ( .A1(n18155), .A2(n18138), .ZN(n17790) );
  NAND2_X1 U13180 ( .A1(n17790), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18114) );
  NOR2_X1 U13181 ( .A1(n18114), .A2(n18113), .ZN(n18083) );
  NAND3_X1 U13182 ( .A1(n18083), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18066) );
  NOR2_X1 U13183 ( .A1(n18078), .A2(n18066), .ZN(n17988) );
  INV_X1 U13184 ( .A(n17988), .ZN(n18046) );
  NOR2_X1 U13185 ( .A1(n17726), .A2(n18046), .ZN(n10212) );
  INV_X1 U13186 ( .A(n17724), .ZN(n10209) );
  NAND2_X1 U13187 ( .A1(n18155), .A2(n18138), .ZN(n17802) );
  INV_X1 U13188 ( .A(n17802), .ZN(n17725) );
  NOR4_X1 U13189 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U13190 ( .A1(n10209), .A2(n17725), .A3(n10208), .A4(n18078), .ZN(
        n10210) );
  NAND2_X1 U13191 ( .A1(n17729), .A2(n10210), .ZN(n10211) );
  INV_X1 U13192 ( .A(n10211), .ZN(n10213) );
  NAND2_X1 U13193 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17642) );
  INV_X1 U13194 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18001) );
  INV_X1 U13195 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20969) );
  NAND2_X1 U13196 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18005) );
  NOR2_X1 U13197 ( .A1(n20969), .A2(n18005), .ZN(n17987) );
  INV_X1 U13198 ( .A(n17987), .ZN(n17643) );
  NOR2_X1 U13199 ( .A1(n18001), .A2(n17643), .ZN(n17994) );
  NAND2_X1 U13200 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17994), .ZN(
        n16427) );
  NOR2_X1 U13201 ( .A1(n17658), .A2(n16427), .ZN(n17619) );
  NOR2_X1 U13202 ( .A1(n17642), .A2(n16427), .ZN(n17589) );
  NAND2_X1 U13203 ( .A1(n17589), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17600) );
  NAND2_X1 U13204 ( .A1(n18001), .A2(n17729), .ZN(n17696) );
  NOR2_X1 U13205 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17696), .ZN(
        n10214) );
  INV_X1 U13206 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17984) );
  NAND2_X1 U13207 ( .A1(n10214), .A2(n17984), .ZN(n17659) );
  INV_X1 U13208 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17649) );
  INV_X1 U13209 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17967) );
  NAND3_X1 U13210 ( .A1(n17647), .A2(n17649), .A3(n17967), .ZN(n10215) );
  INV_X1 U13211 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17974) );
  NAND2_X1 U13212 ( .A1(n17729), .A2(n17613), .ZN(n17602) );
  AND2_X1 U13213 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17930) );
  NAND2_X1 U13214 ( .A1(n17928), .A2(n16429), .ZN(n16434) );
  INV_X1 U13215 ( .A(n16434), .ZN(n15745) );
  NOR2_X1 U13216 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17833), .ZN(
        n16433) );
  NOR2_X1 U13217 ( .A1(n10219), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10220) );
  NOR2_X1 U13218 ( .A1(n17833), .A2(n15795), .ZN(n10225) );
  INV_X1 U13219 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15799) );
  INV_X1 U13220 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17562) );
  NOR2_X1 U13221 ( .A1(n17562), .A2(n17729), .ZN(n16432) );
  OAI21_X1 U13222 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n15799), .A(
        n15794), .ZN(n10223) );
  NAND2_X1 U13223 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17833), .ZN(
        n10221) );
  OAI22_X1 U13224 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17833), .B1(
        n10221), .B2(n15799), .ZN(n10222) );
  OAI21_X1 U13225 ( .B1(n10225), .B2(n10223), .A(n10222), .ZN(n10228) );
  OAI21_X1 U13226 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17833), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10224) );
  INV_X1 U13227 ( .A(n10225), .ZN(n10226) );
  NAND2_X1 U13228 ( .A1(n9633), .A2(n10226), .ZN(n10227) );
  NAND2_X1 U13229 ( .A1(n10228), .A2(n10227), .ZN(n10429) );
  AOI22_X1 U13230 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10229) );
  OAI21_X1 U13231 ( .B1(n9651), .B2(n17157), .A(n10229), .ZN(n10239) );
  INV_X1 U13232 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U13233 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13234 ( .A1(n10113), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17226), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10230) );
  OAI21_X1 U13235 ( .B1(n15688), .B2(n17269), .A(n10230), .ZN(n10235) );
  INV_X1 U13236 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U13237 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10231), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U13238 ( .A1(n10150), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10232) );
  OAI211_X1 U13239 ( .C1(n9649), .C2(n17158), .A(n10233), .B(n10232), .ZN(
        n10234) );
  AOI211_X1 U13240 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10235), .B(n10234), .ZN(n10236) );
  OAI211_X1 U13241 ( .C1(n17199), .C2(n16989), .A(n10237), .B(n10236), .ZN(
        n10238) );
  AOI211_X1 U13242 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n10239), .B(n10238), .ZN(n10240) );
  AOI22_X1 U13243 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10241) );
  OAI21_X1 U13244 ( .B1(n9652), .B2(n15687), .A(n10241), .ZN(n10253) );
  INV_X1 U13245 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17095) );
  OAI22_X1 U13246 ( .A1(n9651), .A2(n17095), .B1(n15688), .B2(n17289), .ZN(
        n10246) );
  AOI22_X1 U13247 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13248 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10231), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13249 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10242) );
  NAND3_X1 U13250 ( .A1(n10244), .A2(n10243), .A3(n10242), .ZN(n10245) );
  AOI211_X1 U13251 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n10246), .B(n10245), .ZN(n10251) );
  AOI22_X1 U13252 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10250) );
  NOR2_X1 U13253 ( .A1(n17199), .A2(n15678), .ZN(n10248) );
  NAND3_X1 U13254 ( .A1(n10251), .A2(n10250), .A3(n10249), .ZN(n10252) );
  AOI22_X1 U13255 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10254) );
  OAI21_X1 U13256 ( .B1(n9651), .B2(n17107), .A(n10254), .ZN(n10264) );
  AOI22_X1 U13257 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13258 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U13259 ( .B1(n10147), .B2(n18597), .A(n10256), .ZN(n10260) );
  AOI22_X1 U13260 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13261 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10257) );
  OAI211_X1 U13262 ( .C1(n20941), .C2(n9649), .A(n10258), .B(n10257), .ZN(
        n10259) );
  AOI211_X1 U13263 ( .C1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .C2(n9622), .A(
        n10260), .B(n10259), .ZN(n10261) );
  OAI211_X1 U13264 ( .C1(n17148), .C2(n17225), .A(n10262), .B(n10261), .ZN(
        n10263) );
  AOI211_X4 U13265 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n10264), .B(n10263), .ZN(n18917) );
  NAND2_X1 U13266 ( .A1(n10396), .A2(n18277), .ZN(n10351) );
  INV_X1 U13267 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13268 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10274) );
  INV_X1 U13269 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U13270 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13271 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10265) );
  OAI211_X1 U13272 ( .C1(n9616), .C2(n17173), .A(n10266), .B(n10265), .ZN(
        n10272) );
  AOI22_X1 U13273 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13274 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U13275 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10142), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U13276 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10267) );
  NAND4_X1 U13277 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        n10271) );
  OAI211_X1 U13278 ( .C1(n9612), .C2(n10275), .A(n10274), .B(n10273), .ZN(
        n18287) );
  AOI22_X1 U13279 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13280 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10276) );
  OAI211_X1 U13281 ( .C1(n9616), .C2(n15700), .A(n10277), .B(n10276), .ZN(
        n10283) );
  AOI22_X1 U13282 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13283 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13284 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U13285 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10278) );
  NAND4_X1 U13286 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NAND2_X1 U13287 ( .A1(n17303), .A2(n18291), .ZN(n18722) );
  INV_X1 U13288 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U13289 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13290 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10286) );
  OAI211_X1 U13291 ( .C1(n9616), .C2(n16988), .A(n10287), .B(n10286), .ZN(
        n10293) );
  AOI22_X1 U13292 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13293 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13294 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U13295 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10288) );
  NAND4_X1 U13296 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10292) );
  INV_X1 U13297 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U13298 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10305) );
  INV_X1 U13299 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U13300 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13301 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10296) );
  OAI211_X1 U13302 ( .C1(n9649), .C2(n17087), .A(n10297), .B(n10296), .ZN(
        n10303) );
  AOI22_X1 U13303 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13304 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13305 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U13306 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10298) );
  NAND4_X1 U13307 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10302) );
  INV_X1 U13308 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13309 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13310 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13311 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13312 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13313 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U13314 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10309) );
  NOR2_X1 U13315 ( .A1(n18917), .A2(n18269), .ZN(n10314) );
  INV_X1 U13316 ( .A(n10396), .ZN(n18280) );
  NOR2_X1 U13317 ( .A1(n10314), .A2(n18280), .ZN(n10317) );
  NAND2_X1 U13318 ( .A1(n17307), .A2(n18295), .ZN(n10398) );
  NAND2_X1 U13319 ( .A1(n10317), .A2(n10398), .ZN(n10315) );
  NAND2_X1 U13320 ( .A1(n18917), .A2(n18269), .ZN(n10316) );
  AOI21_X1 U13321 ( .B1(n18299), .B2(n18722), .A(n10316), .ZN(n10389) );
  NAND2_X1 U13322 ( .A1(n18291), .A2(n18295), .ZN(n10326) );
  INV_X1 U13323 ( .A(n10326), .ZN(n10322) );
  NOR2_X2 U13324 ( .A1(n18287), .A2(n18295), .ZN(n10388) );
  OAI21_X1 U13325 ( .B1(n18280), .B2(n18269), .A(n18722), .ZN(n10318) );
  OAI21_X1 U13326 ( .B1(n10322), .B2(n10388), .A(n10318), .ZN(n10320) );
  NAND2_X1 U13327 ( .A1(n18299), .A2(n15632), .ZN(n10395) );
  NAND3_X1 U13328 ( .A1(n10321), .A2(n10320), .A3(n10319), .ZN(n10325) );
  OAI21_X1 U13329 ( .B1(n17425), .B2(n10322), .A(n18287), .ZN(n10323) );
  INV_X1 U13330 ( .A(n10323), .ZN(n10324) );
  AOI21_X1 U13331 ( .B1(n10327), .B2(n10390), .A(n10394), .ZN(n10328) );
  OAI22_X1 U13332 ( .A1(n18885), .A2(n18397), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10345) );
  INV_X1 U13333 ( .A(n10345), .ZN(n10334) );
  AOI22_X1 U13334 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18271), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18878), .ZN(n10337) );
  NAND2_X1 U13335 ( .A1(n10345), .A2(n10335), .ZN(n10329) );
  OAI21_X1 U13336 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18885), .A(
        n10329), .ZN(n10336) );
  NAND2_X1 U13337 ( .A1(n10337), .A2(n10336), .ZN(n10330) );
  NAND2_X1 U13338 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10331), .ZN(
        n10338) );
  OAI22_X1 U13339 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18266), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10331), .ZN(n10340) );
  AOI21_X1 U13340 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10338), .A(
        n10340), .ZN(n10332) );
  AOI21_X1 U13341 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18266), .A(
        n10332), .ZN(n10341) );
  OAI21_X1 U13342 ( .B1(n10335), .B2(n10334), .A(n10341), .ZN(n10333) );
  AOI21_X1 U13343 ( .B1(n18893), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n10335), .ZN(n10346) );
  INV_X1 U13344 ( .A(n10346), .ZN(n10344) );
  XOR2_X1 U13345 ( .A(n10337), .B(n10336), .Z(n10343) );
  NOR2_X1 U13346 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18266), .ZN(
        n10339) );
  AOI22_X1 U13347 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10340), .B1(
        n10339), .B2(n10338), .ZN(n10347) );
  INV_X1 U13348 ( .A(n10341), .ZN(n10342) );
  AOI21_X1 U13349 ( .B1(n10349), .B2(n10344), .A(n10350), .ZN(n10416) );
  INV_X1 U13350 ( .A(n10416), .ZN(n18701) );
  NAND3_X1 U13351 ( .A1(n10347), .A2(n10346), .A3(n10345), .ZN(n10348) );
  NAND2_X1 U13352 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18918) );
  NAND2_X2 U13353 ( .A1(n18925), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18850) );
  OAI211_X1 U13354 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18787), .B(n18850), .ZN(n18915) );
  OAI211_X1 U13355 ( .C1(n10396), .C2(n18277), .A(n10351), .B(n18915), .ZN(
        n10352) );
  NAND2_X1 U13356 ( .A1(n18918), .A2(n10352), .ZN(n16553) );
  NOR2_X1 U13357 ( .A1(n16555), .A2(n16553), .ZN(n10353) );
  MUX2_X1 U13358 ( .A(n15737), .B(n10353), .S(n10071), .Z(n10354) );
  AOI21_X1 U13359 ( .B1(n10355), .B2(n18701), .A(n10354), .ZN(n10356) );
  INV_X1 U13360 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18873) );
  NAND2_X1 U13361 ( .A1(n17921), .A2(n17449), .ZN(n10362) );
  NAND2_X1 U13362 ( .A1(n17446), .A2(n10362), .ZN(n10361) );
  NAND2_X1 U13363 ( .A1(n10361), .A2(n10128), .ZN(n10371) );
  NOR2_X1 U13364 ( .A1(n17438), .A2(n10371), .ZN(n10359) );
  INV_X1 U13365 ( .A(n17434), .ZN(n10358) );
  NAND2_X1 U13366 ( .A1(n10359), .A2(n10358), .ZN(n10374) );
  NOR2_X1 U13367 ( .A1(n17430), .A2(n10374), .ZN(n10378) );
  NAND2_X1 U13368 ( .A1(n10378), .A2(n16439), .ZN(n10379) );
  XNOR2_X1 U13369 ( .A(n10359), .B(n17434), .ZN(n10360) );
  AND2_X1 U13370 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10360), .ZN(
        n10373) );
  XOR2_X1 U13371 ( .A(n17861), .B(n10360), .Z(n17864) );
  XNOR2_X1 U13372 ( .A(n10361), .B(n10128), .ZN(n10369) );
  INV_X1 U13373 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18213) );
  NOR2_X1 U13374 ( .A1(n10369), .A2(n18213), .ZN(n10370) );
  XOR2_X1 U13375 ( .A(n17446), .B(n10362), .Z(n10363) );
  NOR2_X1 U13376 ( .A1(n10363), .A2(n18235), .ZN(n10368) );
  XOR2_X1 U13377 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10363), .Z(
        n17901) );
  INV_X1 U13378 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18890) );
  NOR2_X1 U13379 ( .A1(n10365), .A2(n18890), .ZN(n10367) );
  INV_X1 U13380 ( .A(n17921), .ZN(n10366) );
  NAND3_X1 U13381 ( .A1(n10366), .A2(n10365), .A3(n18890), .ZN(n10364) );
  OAI221_X1 U13382 ( .B1(n10367), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n10366), .C2(n10365), .A(n10364), .ZN(n17900) );
  NOR2_X1 U13383 ( .A1(n17901), .A2(n17900), .ZN(n17899) );
  NOR2_X1 U13384 ( .A1(n10368), .A2(n17899), .ZN(n17891) );
  XOR2_X1 U13385 ( .A(n10369), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n17890) );
  NOR2_X1 U13386 ( .A1(n17891), .A2(n17890), .ZN(n17889) );
  NOR2_X1 U13387 ( .A1(n10370), .A2(n17889), .ZN(n17873) );
  XNOR2_X1 U13388 ( .A(n10371), .B(n17438), .ZN(n17874) );
  NOR2_X1 U13389 ( .A1(n17873), .A2(n17874), .ZN(n10372) );
  NAND2_X1 U13390 ( .A1(n17873), .A2(n17874), .ZN(n17872) );
  OAI21_X1 U13391 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n10372), .A(
        n17872), .ZN(n17863) );
  NOR2_X1 U13392 ( .A1(n17864), .A2(n17863), .ZN(n17862) );
  NOR2_X1 U13393 ( .A1(n10373), .A2(n17862), .ZN(n10375) );
  XNOR2_X1 U13394 ( .A(n10374), .B(n17430), .ZN(n10376) );
  NOR2_X1 U13395 ( .A1(n10375), .A2(n10376), .ZN(n10377) );
  XNOR2_X1 U13396 ( .A(n10376), .B(n10375), .ZN(n17854) );
  NOR2_X1 U13397 ( .A1(n17854), .A2(n18178), .ZN(n17853) );
  NOR2_X1 U13398 ( .A1(n10377), .A2(n17853), .ZN(n10380) );
  XNOR2_X1 U13399 ( .A(n10378), .B(n16439), .ZN(n10381) );
  NAND2_X1 U13400 ( .A1(n10380), .A2(n10381), .ZN(n17838) );
  NAND2_X1 U13401 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17838), .ZN(
        n10383) );
  NOR2_X1 U13402 ( .A1(n10379), .A2(n10383), .ZN(n10385) );
  INV_X1 U13403 ( .A(n10379), .ZN(n10384) );
  OR2_X1 U13404 ( .A1(n10381), .A2(n10380), .ZN(n17839) );
  OAI21_X1 U13405 ( .B1(n10384), .B2(n10383), .A(n17839), .ZN(n10382) );
  AOI21_X1 U13406 ( .B1(n10384), .B2(n10383), .A(n10382), .ZN(n17830) );
  INV_X1 U13407 ( .A(n18083), .ZN(n18082) );
  INV_X1 U13408 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18106) );
  NOR2_X1 U13409 ( .A1(n18082), .A2(n18106), .ZN(n18079) );
  INV_X1 U13410 ( .A(n18079), .ZN(n18088) );
  NOR2_X1 U13411 ( .A1(n18123), .A2(n18088), .ZN(n17748) );
  NAND2_X1 U13412 ( .A1(n17748), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17747) );
  NOR2_X2 U13413 ( .A1(n17747), .A2(n18078), .ZN(n18064) );
  INV_X1 U13414 ( .A(n17589), .ZN(n10386) );
  NAND2_X1 U13415 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17950) );
  INV_X1 U13416 ( .A(n17950), .ZN(n17952) );
  NAND3_X1 U13417 ( .A1(n17952), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10410) );
  NOR2_X1 U13418 ( .A1(n10386), .A2(n10410), .ZN(n12884) );
  NAND2_X1 U13419 ( .A1(n18064), .A2(n12884), .ZN(n16407) );
  NAND2_X1 U13420 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16419) );
  INV_X1 U13421 ( .A(n16419), .ZN(n15755) );
  NAND2_X1 U13422 ( .A1(n15755), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15798) );
  NOR2_X1 U13423 ( .A1(n16407), .A2(n15798), .ZN(n16406) );
  NAND2_X1 U13424 ( .A1(n16406), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10387) );
  XOR2_X1 U13425 ( .A(n18873), .B(n10387), .Z(n10418) );
  NAND2_X1 U13426 ( .A1(n10396), .A2(n10388), .ZN(n10393) );
  AOI21_X1 U13427 ( .B1(n10071), .B2(n10393), .A(n10389), .ZN(n10391) );
  NOR2_X1 U13428 ( .A1(n16576), .A2(n16574), .ZN(n10402) );
  INV_X1 U13429 ( .A(n10395), .ZN(n10400) );
  NAND2_X1 U13430 ( .A1(n10397), .A2(n10396), .ZN(n18711) );
  INV_X1 U13431 ( .A(n15630), .ZN(n10399) );
  NAND3_X1 U13432 ( .A1(n10400), .A2(n18917), .A3(n10399), .ZN(n10401) );
  NAND2_X1 U13433 ( .A1(n17303), .A2(n18287), .ZN(n18712) );
  AOI21_X1 U13434 ( .B1(n10405), .B2(n18277), .A(n10404), .ZN(n18710) );
  NAND2_X1 U13435 ( .A1(n18705), .A2(n18238), .ZN(n18210) );
  INV_X1 U13436 ( .A(n18066), .ZN(n18056) );
  NAND2_X1 U13437 ( .A1(n18126), .A2(n18056), .ZN(n17749) );
  NAND2_X1 U13438 ( .A1(n12884), .A2(n18065), .ZN(n16418) );
  NOR2_X1 U13439 ( .A1(n15798), .A2(n16418), .ZN(n16420) );
  NAND2_X1 U13440 ( .A1(n16420), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10406) );
  XOR2_X1 U13441 ( .A(n10406), .B(n18873), .Z(n10417) );
  NAND2_X1 U13442 ( .A1(n17427), .A2(n18252), .ZN(n18172) );
  INV_X1 U13443 ( .A(n18172), .ZN(n15751) );
  AOI22_X1 U13444 ( .A1(n10418), .A2(n18250), .B1(n10417), .B2(n15751), .ZN(
        n10414) );
  NAND2_X1 U13445 ( .A1(n18238), .A2(n18162), .ZN(n18240) );
  NAND2_X1 U13446 ( .A1(n18716), .A2(n18723), .ZN(n18203) );
  NOR2_X1 U13447 ( .A1(n18177), .A2(n18178), .ZN(n18157) );
  NAND2_X1 U13448 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18157), .ZN(
        n10407) );
  INV_X1 U13449 ( .A(n10407), .ZN(n18030) );
  NAND3_X1 U13450 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18029) );
  NAND2_X1 U13451 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18202) );
  NOR2_X1 U13452 ( .A1(n18029), .A2(n18202), .ZN(n18161) );
  NAND2_X1 U13453 ( .A1(n18030), .A2(n18161), .ZN(n18097) );
  INV_X1 U13454 ( .A(n18097), .ZN(n18135) );
  NAND2_X1 U13455 ( .A1(n17988), .A2(n18135), .ZN(n18034) );
  INV_X1 U13456 ( .A(n18034), .ZN(n17983) );
  AOI21_X1 U13457 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18227) );
  OR2_X1 U13458 ( .A1(n18029), .A2(n18227), .ZN(n18159) );
  NOR2_X1 U13459 ( .A1(n18159), .A2(n10407), .ZN(n18052) );
  NOR2_X1 U13460 ( .A1(n17642), .A2(n18046), .ZN(n17691) );
  NAND2_X1 U13461 ( .A1(n18052), .A2(n17691), .ZN(n18039) );
  OR2_X1 U13462 ( .A1(n16427), .A2(n18039), .ZN(n17968) );
  OAI21_X1 U13463 ( .B1(n10410), .B2(n17968), .A(n18707), .ZN(n10408) );
  INV_X1 U13464 ( .A(n10408), .ZN(n17935) );
  NOR2_X1 U13465 ( .A1(n18723), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18224) );
  AOI211_X1 U13466 ( .C1(n18081), .C2(n17928), .A(n17935), .B(n18224), .ZN(
        n10409) );
  OAI221_X1 U13467 ( .B1(n18222), .B2(n12884), .C1(n18222), .C2(n17983), .A(
        n10409), .ZN(n15747) );
  OAI211_X1 U13468 ( .C1(n15747), .C2(n15798), .A(n18162), .B(n18238), .ZN(
        n15800) );
  INV_X1 U13469 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18871) );
  NAND2_X1 U13470 ( .A1(n18871), .A2(n18862), .ZN(n18928) );
  OR3_X2 U13471 ( .A1(n18928), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18253) );
  OAI211_X1 U13472 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18240), .A(
        n15800), .B(n18239), .ZN(n10412) );
  INV_X1 U13473 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18847) );
  NOR2_X1 U13474 ( .A1(n18847), .A2(n18253), .ZN(n10425) );
  NOR2_X1 U13475 ( .A1(n10410), .A2(n18254), .ZN(n16428) );
  AOI21_X1 U13476 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18081), .A(
        n18725), .ZN(n18220) );
  NAND2_X1 U13477 ( .A1(n17589), .A2(n17983), .ZN(n17929) );
  OAI22_X1 U13478 ( .A1(n18736), .A2(n17968), .B1(n18220), .B2(n17929), .ZN(
        n17951) );
  NAND2_X1 U13479 ( .A1(n16428), .A2(n17951), .ZN(n15752) );
  NOR4_X1 U13480 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15798), .A3(
        n15799), .A4(n15752), .ZN(n10411) );
  AOI211_X1 U13481 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n10412), .A(
        n10425), .B(n10411), .ZN(n10413) );
  OAI21_X1 U13482 ( .B1(n10429), .B2(n18144), .A(n10415), .ZN(P3_U2831) );
  AOI22_X1 U13483 ( .A1(n9574), .A2(n10418), .B1(n17791), .B2(n10417), .ZN(
        n10427) );
  INV_X1 U13484 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18753) );
  NAND2_X1 U13485 ( .A1(n18753), .A2(n18862), .ZN(n16550) );
  NAND2_X1 U13486 ( .A1(n18928), .A2(n16550), .ZN(n18259) );
  INV_X1 U13487 ( .A(n18259), .ZN(n18909) );
  INV_X1 U13488 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18916) );
  NOR2_X1 U13489 ( .A1(n18871), .A2(n18916), .ZN(n17676) );
  INV_X1 U13490 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16603) );
  NAND2_X1 U13491 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16905) );
  NAND2_X1 U13492 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17797) );
  NAND3_X1 U13493 ( .A1(n17821), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17784) );
  NAND2_X1 U13494 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17681) );
  NOR2_X1 U13495 ( .A1(n17678), .A2(n17681), .ZN(n17664) );
  NAND2_X1 U13496 ( .A1(n17664), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16591) );
  NAND2_X1 U13497 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17596) );
  INV_X1 U13498 ( .A(n17596), .ZN(n17581) );
  NAND2_X1 U13499 ( .A1(n17581), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12882) );
  INV_X1 U13500 ( .A(n12882), .ZN(n10421) );
  NAND2_X1 U13501 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17564) );
  INV_X1 U13502 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16617) );
  NAND2_X1 U13503 ( .A1(n18859), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18771) );
  INV_X1 U13504 ( .A(n18771), .ZN(n17755) );
  NOR2_X1 U13505 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18920) );
  AOI21_X1 U13506 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18920), .ZN(n18768) );
  NAND3_X1 U13507 ( .A1(n18753), .A2(n18862), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18513) );
  NAND2_X1 U13508 ( .A1(n10420), .A2(n17763), .ZN(n16398) );
  XNOR2_X1 U13509 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10423) );
  NOR2_X1 U13510 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17702), .ZN(
        n16411) );
  NAND2_X1 U13511 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17582), .ZN(
        n16589) );
  INV_X1 U13512 ( .A(n16589), .ZN(n12877) );
  NAND2_X1 U13513 ( .A1(n10421), .A2(n12877), .ZN(n16584) );
  NOR2_X1 U13514 ( .A1(n17564), .A2(n16584), .ZN(n16409) );
  NAND2_X1 U13515 ( .A1(n18648), .A2(n10422), .ZN(n16415) );
  OAI211_X1 U13516 ( .C1(n16409), .C2(n18771), .A(n17922), .B(n16415), .ZN(
        n16408) );
  NOR2_X1 U13517 ( .A1(n16411), .A2(n16408), .ZN(n16397) );
  OAI22_X1 U13518 ( .A1(n16398), .A2(n10423), .B1(n16397), .B2(n16603), .ZN(
        n10424) );
  AOI211_X1 U13519 ( .C1(n17758), .C2(n16949), .A(n10425), .B(n10424), .ZN(
        n10426) );
  OAI21_X1 U13520 ( .B1(n10429), .B2(n17807), .A(n10428), .ZN(P3_U2799) );
  NAND2_X2 U13521 ( .A1(n13781), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10573) );
  INV_X2 U13522 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13523 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10435) );
  AND3_X4 U13524 ( .A1(n10456), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13525 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10434) );
  AND2_X4 U13526 ( .A1(n10522), .A2(n10718), .ZN(n10621) );
  AOI22_X1 U13527 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10433) );
  AND2_X2 U13528 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13182) );
  AND2_X4 U13529 ( .A1(n13182), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10619) );
  AND2_X4 U13530 ( .A1(n13182), .A2(n10459), .ZN(n10590) );
  AOI22_X1 U13531 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10432) );
  NAND4_X1 U13532 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10436) );
  NAND2_X1 U13533 ( .A1(n10436), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10443) );
  AOI22_X1 U13534 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13535 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9609), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13536 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13537 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  NAND2_X1 U13538 ( .A1(n10441), .A2(n10508), .ZN(n10442) );
  AOI22_X1 U13539 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13540 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14099), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13541 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10444) );
  NAND4_X1 U13542 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10448) );
  AOI22_X1 U13543 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13544 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13545 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14099), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13546 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10453) );
  NAND2_X1 U13547 ( .A1(n10453), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10454) );
  NAND2_X2 U13548 ( .A1(n10462), .A2(n10710), .ZN(n11162) );
  NAND2_X1 U13549 ( .A1(n10709), .A2(n21042), .ZN(n10461) );
  NAND2_X1 U13550 ( .A1(n19891), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U13551 ( .A1(n10456), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13552 ( .A1(n10458), .A2(n10457), .ZN(n10464) );
  NAND2_X1 U13553 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19900), .ZN(
        n10463) );
  NAND2_X1 U13554 ( .A1(n10465), .A2(n10458), .ZN(n10473) );
  NAND2_X1 U13555 ( .A1(n19881), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10474) );
  NAND2_X1 U13556 ( .A1(n10459), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13557 ( .A1(n10474), .A2(n10460), .ZN(n10471) );
  XNOR2_X1 U13558 ( .A(n10473), .B(n10471), .ZN(n10516) );
  MUX2_X1 U13559 ( .A(n10461), .B(n11162), .S(n10516), .Z(n10470) );
  INV_X1 U13560 ( .A(n10516), .ZN(n10648) );
  OAI21_X1 U13561 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19900), .A(
        n10463), .ZN(n10635) );
  INV_X1 U13562 ( .A(n11162), .ZN(n13645) );
  OAI21_X1 U13563 ( .B1(n10635), .B2(n10464), .A(n13645), .ZN(n10468) );
  INV_X1 U13564 ( .A(n10635), .ZN(n10466) );
  NAND2_X1 U13565 ( .A1(n10464), .A2(n10463), .ZN(n10636) );
  AND2_X1 U13566 ( .A1(n10465), .A2(n10636), .ZN(n10518) );
  OAI211_X1 U13567 ( .C1(n21042), .C2(n10466), .A(n10722), .B(n10518), .ZN(
        n10467) );
  OAI211_X1 U13568 ( .C1(n10648), .C2(n10725), .A(n10468), .B(n10467), .ZN(
        n10469) );
  NAND2_X1 U13569 ( .A1(n10470), .A2(n10469), .ZN(n10480) );
  INV_X1 U13570 ( .A(n10471), .ZN(n10472) );
  NAND2_X1 U13571 ( .A1(n10473), .A2(n10472), .ZN(n10475) );
  NAND2_X1 U13572 ( .A1(n10475), .A2(n10474), .ZN(n10479) );
  INV_X1 U13573 ( .A(n10479), .ZN(n10476) );
  NAND3_X1 U13574 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10482), .A3(
        n16375), .ZN(n10676) );
  XNOR2_X1 U13575 ( .A(n10479), .B(n10478), .ZN(n10661) );
  MUX2_X1 U13576 ( .A(n11162), .B(n10480), .S(n10515), .Z(n10481) );
  INV_X1 U13577 ( .A(n10481), .ZN(n10484) );
  AND2_X1 U13578 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16375), .ZN(
        n10483) );
  NOR2_X1 U13579 ( .A1(n10484), .A2(n10678), .ZN(n10485) );
  MUX2_X1 U13580 ( .A(n10485), .B(n16375), .S(n21039), .Z(n10514) );
  INV_X1 U13581 ( .A(n16367), .ZN(n10487) );
  INV_X1 U13582 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U13583 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13584 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10489) );
  NAND2_X1 U13585 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10493) );
  NAND2_X1 U13586 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10492) );
  NAND2_X1 U13587 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10491) );
  NAND4_X1 U13588 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10508), .ZN(
        n10495) );
  INV_X1 U13589 ( .A(n10622), .ZN(n14016) );
  NOR2_X1 U13590 ( .A1(n10495), .A2(n10494), .ZN(n10497) );
  NAND2_X1 U13591 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10496) );
  NAND3_X1 U13592 ( .A1(n10498), .A2(n10497), .A3(n10496), .ZN(n10513) );
  NAND2_X1 U13593 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10501) );
  NAND2_X1 U13594 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10500) );
  NAND3_X1 U13595 ( .A1(n10501), .A2(n10500), .A3(n10499), .ZN(n10503) );
  INV_X1 U13596 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10502) );
  NAND2_X1 U13597 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10507) );
  NAND2_X1 U13598 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13599 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10505) );
  NAND2_X1 U13600 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10504) );
  NAND4_X1 U13601 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10509) );
  OAI211_X1 U13602 ( .C1(n21040), .C2(n10514), .A(n13071), .B(n10727), .ZN(
        n10687) );
  NAND2_X1 U13603 ( .A1(n10516), .A2(n10515), .ZN(n10520) );
  INV_X1 U13604 ( .A(n10520), .ZN(n10517) );
  OAI21_X1 U13605 ( .B1(n10635), .B2(n10520), .A(n16360), .ZN(n10521) );
  INV_X1 U13606 ( .A(n10521), .ZN(n10525) );
  AND2_X2 U13607 ( .A1(n9621), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10668) );
  INV_X1 U13608 ( .A(n10668), .ZN(n10523) );
  NOR2_X1 U13609 ( .A1(n13178), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12952) );
  NAND2_X1 U13610 ( .A1(n10523), .A2(n12952), .ZN(n10524) );
  INV_X1 U13611 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12950) );
  NAND2_X1 U13612 ( .A1(n10524), .A2(n12950), .ZN(n19896) );
  MUX2_X1 U13613 ( .A(n10525), .B(n19896), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n15823) );
  AOI22_X1 U13614 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13615 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13616 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10621), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13617 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13618 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13619 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13620 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13621 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13622 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13623 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13624 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13625 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10538) );
  NAND2_X1 U13626 ( .A1(n10538), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10545) );
  AOI22_X1 U13627 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13628 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13629 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10543) );
  NAND2_X1 U13630 ( .A1(n10543), .A2(n10508), .ZN(n10544) );
  AOI22_X1 U13631 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13632 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13633 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10546) );
  NAND4_X1 U13634 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10550) );
  NAND2_X1 U13635 ( .A1(n10550), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10558) );
  AOI22_X1 U13636 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13637 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13638 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13639 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10552) );
  NAND4_X1 U13640 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10556) );
  NAND2_X1 U13641 ( .A1(n10556), .A2(n16349), .ZN(n10557) );
  NAND4_X1 U13642 ( .A1(n10704), .A2(n10726), .A3(n11020), .A4(n10703), .ZN(
        n10602) );
  INV_X1 U13643 ( .A(n10602), .ZN(n10598) );
  NAND2_X1 U13644 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U13645 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10559) );
  NAND2_X1 U13646 ( .A1(n10560), .A2(n10559), .ZN(n10563) );
  INV_X1 U13647 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U13648 ( .A1(n10563), .A2(n10562), .ZN(n10571) );
  INV_X1 U13649 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10564) );
  NOR2_X1 U13650 ( .A1(n10565), .A2(n10508), .ZN(n10570) );
  NAND2_X1 U13651 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10569) );
  NAND2_X1 U13652 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10568) );
  NAND2_X1 U13653 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10567) );
  NAND2_X1 U13654 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10566) );
  NAND3_X1 U13655 ( .A1(n10571), .A2(n10570), .A3(n10070), .ZN(n10584) );
  INV_X1 U13656 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10572) );
  OR2_X1 U13657 ( .A1(n10573), .A2(n10572), .ZN(n10574) );
  NAND2_X1 U13658 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10578) );
  NAND2_X1 U13659 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13660 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13661 ( .A1(n10551), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10575) );
  NAND2_X1 U13662 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13663 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10579) );
  NAND4_X1 U13664 ( .A1(n10574), .A2(n10068), .A3(n10067), .A4(n10582), .ZN(
        n10583) );
  AOI22_X1 U13665 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13666 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10551), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13667 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9609), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13668 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10585) );
  NAND4_X1 U13669 ( .A1(n10588), .A2(n10587), .A3(n10586), .A4(n10585), .ZN(
        n10589) );
  NAND2_X1 U13670 ( .A1(n10589), .A2(n10508), .ZN(n10597) );
  AOI22_X1 U13671 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13672 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13673 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10595) );
  NAND2_X1 U13674 ( .A1(n10595), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10596) );
  NOR2_X1 U13675 ( .A1(n9591), .A2(n14062), .ZN(n10618) );
  NAND2_X1 U13676 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n21038) );
  INV_X1 U13677 ( .A(n21038), .ZN(n19786) );
  NOR2_X1 U13678 ( .A1(n12930), .A2(n19786), .ZN(n12943) );
  INV_X1 U13679 ( .A(n12943), .ZN(n10616) );
  NAND3_X2 U13680 ( .A1(n10601), .A2(n10600), .A3(n10742), .ZN(n10692) );
  MUX2_X1 U13681 ( .A(n10692), .B(n10713), .S(n14062), .Z(n10615) );
  INV_X2 U13682 ( .A(n19910), .ZN(n19909) );
  NAND2_X2 U13683 ( .A1(n19909), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19855) );
  NOR2_X1 U13684 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n18940) );
  INV_X1 U13685 ( .A(n18940), .ZN(n19796) );
  NAND2_X1 U13686 ( .A1(n21038), .A2(n21041), .ZN(n13639) );
  INV_X1 U13687 ( .A(n13639), .ZN(n10683) );
  NAND2_X1 U13688 ( .A1(n10683), .A2(n10747), .ZN(n10613) );
  NAND2_X1 U13689 ( .A1(n10714), .A2(n10689), .ZN(n10603) );
  NOR2_X1 U13690 ( .A1(n21042), .A2(n10704), .ZN(n11297) );
  NAND2_X1 U13691 ( .A1(n10713), .A2(n10726), .ZN(n10696) );
  NOR2_X1 U13692 ( .A1(n10696), .A2(n10714), .ZN(n10604) );
  OAI21_X1 U13693 ( .B1(n11297), .B2(n21040), .A(n10604), .ZN(n10605) );
  NAND2_X1 U13694 ( .A1(n10748), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U13695 ( .A1(n10608), .A2(n13125), .ZN(n10606) );
  AND2_X1 U13696 ( .A1(n14062), .A2(n21040), .ZN(n16379) );
  NAND2_X1 U13697 ( .A1(n10606), .A2(n16379), .ZN(n11280) );
  NAND2_X1 U13698 ( .A1(n10607), .A2(n11280), .ZN(n11299) );
  INV_X1 U13699 ( .A(n11299), .ZN(n10612) );
  NAND2_X1 U13700 ( .A1(n10704), .A2(n10608), .ZN(n10611) );
  OAI211_X1 U13701 ( .C1(n12930), .C2(n10613), .A(n10612), .B(n10695), .ZN(
        n10614) );
  INV_X1 U13702 ( .A(n10614), .ZN(n12947) );
  OAI21_X1 U13703 ( .B1(n10616), .B2(n10615), .A(n12947), .ZN(n10617) );
  AOI21_X1 U13704 ( .B1(n15823), .B2(n10618), .A(n10617), .ZN(n10682) );
  INV_X1 U13705 ( .A(n10619), .ZN(n10620) );
  INV_X2 U13706 ( .A(n10620), .ZN(n15584) );
  AND2_X2 U13707 ( .A1(n15584), .A2(n16349), .ZN(n11371) );
  AND2_X1 U13708 ( .A1(n9609), .A2(n16349), .ZN(n10911) );
  AOI22_X1 U13709 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13710 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10625) );
  AND2_X2 U13711 ( .A1(n13178), .A2(n10718), .ZN(n13913) );
  AND2_X1 U13712 ( .A1(n10621), .A2(n16349), .ZN(n10663) );
  AOI22_X1 U13713 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10624) );
  AND2_X1 U13714 ( .A1(n14096), .A2(n16349), .ZN(n10650) );
  AOI22_X1 U13715 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10637), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10623) );
  NAND4_X1 U13716 ( .A1(n10626), .A2(n10625), .A3(n10624), .A4(n10623), .ZN(
        n10634) );
  AOI22_X1 U13717 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13718 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10631) );
  AND2_X2 U13719 ( .A1(n13178), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13912) );
  AOI22_X1 U13720 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10630) );
  AND2_X2 U13721 ( .A1(n10628), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10906) );
  AOI22_X1 U13722 ( .A1(n10906), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10855), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10629) );
  NAND4_X1 U13723 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10633) );
  NOR2_X1 U13724 ( .A1(n10634), .A2(n10633), .ZN(n11316) );
  MUX2_X1 U13725 ( .A(n11316), .B(n10635), .S(n11162), .Z(n11004) );
  INV_X1 U13726 ( .A(n10636), .ZN(n10649) );
  AOI22_X1 U13727 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10662), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13728 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13729 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U13730 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13907), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10638) );
  NAND4_X1 U13731 ( .A1(n10641), .A2(n10640), .A3(n10639), .A4(n10638), .ZN(
        n10647) );
  AOI22_X1 U13732 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10911), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13733 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13886), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13734 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n13913), .B1(
        n10855), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n13912), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10642) );
  NAND4_X1 U13736 ( .A1(n10645), .A2(n10644), .A3(n10643), .A4(n10642), .ZN(
        n10646) );
  NOR2_X1 U13737 ( .A1(n10647), .A2(n10646), .ZN(n11331) );
  OAI21_X1 U13738 ( .B1(n11004), .B2(n10649), .A(n10997), .ZN(n10677) );
  AOI22_X1 U13739 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10650), .B1(
        n10637), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13740 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13741 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13742 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U13743 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10660) );
  AOI22_X1 U13744 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10911), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13745 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n13913), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13746 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n13912), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13747 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10655) );
  NAND4_X1 U13748 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  MUX2_X1 U13749 ( .A(n11335), .B(n10661), .S(n11162), .Z(n10996) );
  AOI22_X1 U13750 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10662), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13751 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13752 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11371), .B1(
        n13907), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13754 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10675) );
  AOI22_X1 U13755 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13756 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13757 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13758 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13759 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  MUX2_X1 U13760 ( .A(n10676), .B(n10877), .S(n13645), .Z(n11014) );
  NAND3_X1 U13761 ( .A1(n10677), .A2(n10996), .A3(n11014), .ZN(n10680) );
  INV_X1 U13762 ( .A(n10678), .ZN(n10679) );
  INV_X1 U13763 ( .A(n16379), .ZN(n10681) );
  NOR2_X1 U13764 ( .A1(n9591), .A2(n10681), .ZN(n16359) );
  NAND2_X1 U13765 ( .A1(n16362), .A2(n16359), .ZN(n16370) );
  AND2_X1 U13766 ( .A1(n10682), .A2(n16370), .ZN(n10686) );
  INV_X1 U13767 ( .A(n13071), .ZN(n10684) );
  NAND3_X1 U13768 ( .A1(n10684), .A2(n10689), .A3(n10683), .ZN(n10685) );
  NAND3_X1 U13769 ( .A1(n10687), .A2(n10686), .A3(n10685), .ZN(n10688) );
  NAND2_X1 U13770 ( .A1(n16384), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13642) );
  INV_X1 U13771 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13993) );
  NAND2_X1 U13772 ( .A1(n10691), .A2(n10690), .ZN(n10693) );
  NAND2_X1 U13773 ( .A1(n10693), .A2(n10692), .ZN(n11306) );
  AND2_X1 U13774 ( .A1(n11293), .A2(n21040), .ZN(n10694) );
  NAND2_X1 U13775 ( .A1(n11306), .A2(n10694), .ZN(n10708) );
  INV_X1 U13776 ( .A(n10699), .ZN(n10701) );
  NAND2_X1 U13777 ( .A1(n10698), .A2(n10697), .ZN(n11282) );
  NAND2_X1 U13778 ( .A1(n10699), .A2(n11281), .ZN(n10700) );
  INV_X1 U13779 ( .A(n10702), .ZN(n10707) );
  NAND4_X1 U13780 ( .A1(n10743), .A2(n10599), .A3(n10704), .A4(n19309), .ZN(
        n10716) );
  NAND2_X1 U13781 ( .A1(n21040), .A2(n10714), .ZN(n10705) );
  NAND2_X2 U13782 ( .A1(n11306), .A2(n10706), .ZN(n11295) );
  OAI211_X2 U13783 ( .C1(n10708), .C2(n11279), .A(n10707), .B(n11295), .ZN(
        n10763) );
  INV_X1 U13784 ( .A(n10709), .ZN(n10712) );
  INV_X1 U13785 ( .A(n10717), .ZN(n10715) );
  NAND2_X1 U13786 ( .A1(n10763), .A2(n10715), .ZN(n10720) );
  INV_X1 U13787 ( .A(n10716), .ZN(n13120) );
  NAND2_X1 U13788 ( .A1(n11562), .A2(n10718), .ZN(n10719) );
  NAND2_X1 U13789 ( .A1(n10720), .A2(n10719), .ZN(n10734) );
  NAND3_X1 U13790 ( .A1(n10599), .A2(n10609), .A3(n10722), .ZN(n10724) );
  NAND2_X1 U13791 ( .A1(n11314), .A2(n11293), .ZN(n10723) );
  OAI21_X1 U13792 ( .B1(n10724), .B2(n11293), .A(n10723), .ZN(n10730) );
  AND2_X1 U13793 ( .A1(n10741), .A2(n10745), .ZN(n11276) );
  INV_X1 U13794 ( .A(n16381), .ZN(n10773) );
  NOR2_X1 U13795 ( .A1(n10773), .A2(n19900), .ZN(n10732) );
  AOI21_X1 U13796 ( .B1(n11276), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10732), 
        .ZN(n10733) );
  NAND2_X1 U13797 ( .A1(n10734), .A2(n10733), .ZN(n10779) );
  INV_X1 U13798 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11003) );
  NOR2_X1 U13799 ( .A1(n11562), .A2(n11003), .ZN(n10740) );
  INV_X1 U13800 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13801 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10737) );
  OAI211_X1 U13802 ( .C1(n9583), .C2(n10738), .A(n10773), .B(n10737), .ZN(
        n10739) );
  NOR2_X1 U13803 ( .A1(n10740), .A2(n10739), .ZN(n10753) );
  NAND2_X1 U13804 ( .A1(n10741), .A2(n10078), .ZN(n10751) );
  INV_X1 U13805 ( .A(n10725), .ZN(n10744) );
  NAND4_X1 U13806 ( .A1(n10745), .A2(n10744), .A3(n10742), .A4(n12972), .ZN(
        n10746) );
  NOR2_X1 U13807 ( .A1(n21042), .A2(n21039), .ZN(n10749) );
  NAND3_X2 U13808 ( .A1(n10751), .A2(n10746), .A3(n10750), .ZN(n10774) );
  NAND3_X1 U13809 ( .A1(n13121), .A2(n10742), .A3(n10743), .ZN(n10754) );
  NAND2_X1 U13810 ( .A1(n11274), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10756) );
  NAND2_X1 U13811 ( .A1(n10764), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U13812 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10757) );
  OAI211_X1 U13813 ( .C1(n9624), .C2(n12983), .A(n10758), .B(n10757), .ZN(
        n10759) );
  AOI21_X1 U13814 ( .B1(n21039), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10762) );
  OAI21_X1 U13815 ( .B1(n10763), .B2(n10459), .A(n10762), .ZN(n10770) );
  NAND2_X1 U13816 ( .A1(n10774), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10768) );
  AOI22_X1 U13817 ( .A1(n10764), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10766) );
  NAND2_X1 U13818 ( .A1(n11201), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U13819 ( .A1(n10770), .A2(n10769), .ZN(n10771) );
  OAI22_X1 U13820 ( .A1(n10763), .A2(n16349), .B1(n10773), .B2(n19874), .ZN(
        n11167) );
  INV_X1 U13821 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13651) );
  NAND2_X1 U13822 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13823 ( .A1(n10764), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U13824 ( .C1(n11562), .C2(n13651), .A(n10776), .B(n10775), .ZN(
        n10777) );
  INV_X1 U13825 ( .A(n10778), .ZN(n10781) );
  NAND2_X1 U13826 ( .A1(n10781), .A2(n10780), .ZN(n10790) );
  XNOR2_X2 U13827 ( .A(n10783), .B(n10782), .ZN(n13052) );
  INV_X1 U13828 ( .A(n10784), .ZN(n10792) );
  NAND2_X1 U13829 ( .A1(n10792), .A2(n9747), .ZN(n10787) );
  NAND2_X1 U13830 ( .A1(n13738), .A2(n15566), .ZN(n10788) );
  INV_X1 U13831 ( .A(n15566), .ZN(n13784) );
  OR2_X1 U13832 ( .A1(n13738), .A2(n13784), .ZN(n10789) );
  INV_X1 U13833 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13991) );
  OAI22_X1 U13834 ( .A1(n13993), .A2(n19464), .B1(n19347), .B2(n13991), .ZN(
        n10804) );
  INV_X1 U13835 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10793) );
  INV_X2 U13836 ( .A(n13052), .ZN(n19258) );
  INV_X1 U13837 ( .A(n10790), .ZN(n10791) );
  OR3_X2 U13838 ( .A1(n13151), .A2(n19258), .A3(n10814), .ZN(n10881) );
  NAND2_X1 U13839 ( .A1(n10792), .A2(n13673), .ZN(n10813) );
  OR3_X1 U13840 ( .A1(n13151), .A2(n13738), .A3(n10813), .ZN(n10930) );
  INV_X1 U13841 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13992) );
  OAI22_X1 U13842 ( .A1(n10793), .A2(n10881), .B1(n10930), .B2(n13992), .ZN(
        n10794) );
  INV_X1 U13843 ( .A(n10794), .ZN(n10802) );
  INV_X1 U13844 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10799) );
  INV_X1 U13845 ( .A(n10814), .ZN(n10795) );
  INV_X1 U13846 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13990) );
  INV_X1 U13847 ( .A(n10800), .ZN(n10801) );
  NAND2_X1 U13848 ( .A1(n10802), .A2(n10801), .ZN(n10803) );
  NOR2_X1 U13849 ( .A1(n10804), .A2(n10803), .ZN(n10824) );
  NOR2_X4 U13850 ( .A1(n10806), .A2(n19258), .ZN(n19408) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19284), .B1(
        n19408), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10823) );
  INV_X1 U13852 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10809) );
  OR2_X1 U13853 ( .A1(n13673), .A2(n15566), .ZN(n10807) );
  NAND2_X1 U13854 ( .A1(n13151), .A2(n13738), .ZN(n10815) );
  INV_X1 U13855 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10808) );
  OAI22_X1 U13856 ( .A1(n10809), .A2(n10895), .B1(n15615), .B2(n10808), .ZN(
        n10812) );
  INV_X1 U13857 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10810) );
  INV_X1 U13858 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14001) );
  NOR2_X1 U13859 ( .A1(n10812), .A2(n10811), .ZN(n10822) );
  INV_X1 U13860 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13999) );
  INV_X1 U13861 ( .A(n13673), .ZN(n15579) );
  NAND2_X1 U13862 ( .A1(n15566), .A2(n15579), .ZN(n10816) );
  INV_X1 U13863 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14000) );
  OAI22_X1 U13864 ( .A1(n13999), .A2(n13370), .B1(n10892), .B2(n14000), .ZN(
        n10820) );
  INV_X1 U13865 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20876) );
  INV_X1 U13866 ( .A(n10816), .ZN(n10817) );
  INV_X1 U13867 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14002) );
  OAI22_X1 U13868 ( .A1(n20876), .A2(n13440), .B1(n19675), .B2(n14002), .ZN(
        n10819) );
  NOR2_X1 U13869 ( .A1(n10820), .A2(n10819), .ZN(n10821) );
  NAND4_X1 U13870 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10825) );
  NAND2_X1 U13871 ( .A1(n10825), .A2(n21042), .ZN(n10827) );
  NAND2_X2 U13872 ( .A1(n10827), .A2(n10826), .ZN(n10878) );
  INV_X1 U13873 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10828) );
  INV_X1 U13874 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15613) );
  OAI22_X1 U13875 ( .A1(n10828), .A2(n15615), .B1(n10896), .B2(n15613), .ZN(
        n10831) );
  INV_X1 U13876 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10829) );
  INV_X1 U13877 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13949) );
  OAI22_X1 U13878 ( .A1(n10829), .A2(n19724), .B1(n10892), .B2(n13949), .ZN(
        n10830) );
  NOR2_X1 U13879 ( .A1(n10831), .A2(n10830), .ZN(n10849) );
  INV_X1 U13880 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10832) );
  INV_X1 U13881 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13948) );
  AOI21_X1 U13882 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n19284), .A(
        n10833), .ZN(n10848) );
  INV_X1 U13883 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13940) );
  INV_X1 U13884 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10834) );
  OAI22_X1 U13885 ( .A1(n13940), .A2(n19347), .B1(n10895), .B2(n10834), .ZN(
        n10839) );
  INV_X1 U13886 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13942) );
  INV_X1 U13887 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10835) );
  INV_X1 U13888 ( .A(n10884), .ZN(n19380) );
  NAND2_X1 U13889 ( .A1(n19380), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10836) );
  OAI211_X1 U13890 ( .C1(n19464), .C2(n13942), .A(n10837), .B(n10836), .ZN(
        n10838) );
  NOR2_X1 U13891 ( .A1(n10839), .A2(n10838), .ZN(n10847) );
  INV_X1 U13892 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13950) );
  OR2_X1 U13893 ( .A1(n19675), .A2(n13950), .ZN(n10843) );
  INV_X1 U13894 ( .A(n10930), .ZN(n19317) );
  NAND2_X1 U13895 ( .A1(n19317), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10842) );
  INV_X1 U13896 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10840) );
  NAND4_X1 U13897 ( .A1(n10843), .A2(n21042), .A3(n10842), .A4(n10841), .ZN(
        n10845) );
  NOR2_X1 U13898 ( .A1(n10845), .A2(n10844), .ZN(n10846) );
  NAND4_X1 U13899 ( .A1(n10846), .A2(n10848), .A3(n10847), .A4(n10849), .ZN(
        n10863) );
  OR2_X1 U13900 ( .A1(n11316), .A2(n21042), .ZN(n10864) );
  INV_X1 U13901 ( .A(n10864), .ZN(n12988) );
  AOI22_X1 U13902 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10911), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13903 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13904 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10906), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11371), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13906 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10861) );
  AOI22_X1 U13907 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13907), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13909 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10855), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13910 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13911 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10860) );
  NOR2_X1 U13912 ( .A1(n10861), .A2(n10860), .ZN(n11322) );
  INV_X1 U13913 ( .A(n11322), .ZN(n10865) );
  NAND2_X1 U13914 ( .A1(n12988), .A2(n10865), .ZN(n10869) );
  NAND2_X1 U13915 ( .A1(n10869), .A2(n11331), .ZN(n10862) );
  INV_X1 U13916 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19255) );
  AND2_X1 U13917 ( .A1(n10864), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12987) );
  XNOR2_X1 U13918 ( .A(n11316), .B(n10865), .ZN(n10866) );
  NAND2_X1 U13919 ( .A1(n12987), .A2(n10866), .ZN(n10868) );
  XOR2_X1 U13920 ( .A(n10866), .B(n12987), .Z(n13002) );
  NAND2_X1 U13921 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13002), .ZN(
        n10867) );
  NAND2_X1 U13922 ( .A1(n10868), .A2(n10867), .ZN(n10870) );
  XNOR2_X1 U13923 ( .A(n19255), .B(n10870), .ZN(n12964) );
  XNOR2_X1 U13924 ( .A(n11331), .B(n10869), .ZN(n12963) );
  NAND2_X1 U13925 ( .A1(n12964), .A2(n12963), .ZN(n12962) );
  NAND2_X1 U13926 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10870), .ZN(
        n10871) );
  NAND2_X1 U13927 ( .A1(n12962), .A2(n10871), .ZN(n10872) );
  INV_X1 U13928 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16341) );
  XNOR2_X1 U13929 ( .A(n10872), .B(n16341), .ZN(n13816) );
  NAND2_X1 U13930 ( .A1(n13815), .A2(n13816), .ZN(n10874) );
  NAND2_X1 U13931 ( .A1(n10872), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U13932 ( .A1(n10874), .A2(n10873), .ZN(n10923) );
  NAND2_X1 U13933 ( .A1(n10878), .A2(n10876), .ZN(n10875) );
  INV_X1 U13934 ( .A(n10877), .ZN(n11341) );
  XNOR2_X1 U13935 ( .A(n10875), .B(n11341), .ZN(n10924) );
  XNOR2_X1 U13936 ( .A(n10923), .B(n10924), .ZN(n15228) );
  INV_X1 U13937 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15555) );
  AOI22_X1 U13938 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19284), .B1(
        n19408), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10905) );
  INV_X1 U13939 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10880) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10879) );
  OAI22_X1 U13941 ( .A1(n10880), .A2(n19464), .B1(n19347), .B2(n10879), .ZN(
        n10890) );
  INV_X1 U13942 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10883) );
  INV_X1 U13943 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10882) );
  INV_X1 U13944 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10886) );
  INV_X1 U13945 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10885) );
  OAI22_X1 U13946 ( .A1(n10886), .A2(n10884), .B1(n10930), .B2(n10885), .ZN(
        n10887) );
  NOR2_X1 U13947 ( .A1(n10890), .A2(n10889), .ZN(n10904) );
  INV_X1 U13948 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10891) );
  INV_X1 U13949 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14042) );
  OAI22_X1 U13950 ( .A1(n10891), .A2(n19724), .B1(n13370), .B2(n14042), .ZN(
        n10894) );
  INV_X1 U13951 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14045) );
  INV_X1 U13952 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14043) );
  OAI22_X1 U13953 ( .A1(n14045), .A2(n19675), .B1(n10892), .B2(n14043), .ZN(
        n10893) );
  NOR2_X1 U13954 ( .A1(n10894), .A2(n10893), .ZN(n10903) );
  INV_X1 U13955 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10897) );
  INV_X1 U13956 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14044) );
  OAI22_X1 U13957 ( .A1(n10897), .A2(n10895), .B1(n10896), .B2(n14044), .ZN(
        n10901) );
  INV_X1 U13958 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10899) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10898) );
  OAI22_X1 U13960 ( .A1(n10899), .A2(n15615), .B1(n13440), .B2(n10898), .ZN(
        n10900) );
  NOR2_X1 U13961 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  NAND4_X1 U13962 ( .A1(n10905), .A2(n10904), .A3(n10903), .A4(n10902), .ZN(
        n10920) );
  AOI22_X1 U13963 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13964 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13965 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13966 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10907) );
  NAND4_X1 U13967 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n10918) );
  AOI22_X1 U13968 ( .A1(n10911), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13969 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13970 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13971 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10913) );
  NAND4_X1 U13972 ( .A1(n10916), .A2(n10915), .A3(n10914), .A4(n10913), .ZN(
        n10917) );
  NAND2_X1 U13973 ( .A1(n11347), .A2(n14062), .ZN(n10919) );
  XNOR2_X2 U13974 ( .A(n10928), .B(n10921), .ZN(n11019) );
  INV_X1 U13975 ( .A(n11019), .ZN(n10922) );
  INV_X1 U13976 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11026) );
  INV_X1 U13977 ( .A(n10923), .ZN(n10925) );
  NAND2_X1 U13978 ( .A1(n11019), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15537) );
  AOI22_X1 U13979 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19284), .B1(
        n19408), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10947) );
  INV_X1 U13980 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14067) );
  INV_X1 U13981 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14065) );
  OAI22_X1 U13982 ( .A1(n14067), .A2(n19464), .B1(n19347), .B2(n14065), .ZN(
        n10935) );
  INV_X1 U13983 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10929) );
  INV_X1 U13984 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14064) );
  INV_X1 U13985 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10931) );
  INV_X1 U13986 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14066) );
  OAI22_X1 U13987 ( .A1(n10931), .A2(n10884), .B1(n10930), .B2(n14066), .ZN(
        n10932) );
  OR2_X1 U13988 ( .A1(n10933), .A2(n10932), .ZN(n10934) );
  NOR2_X1 U13989 ( .A1(n10935), .A2(n10934), .ZN(n10946) );
  INV_X1 U13990 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14077) );
  INV_X1 U13991 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14078) );
  OAI22_X1 U13992 ( .A1(n14077), .A2(n10896), .B1(n13370), .B2(n14078), .ZN(
        n10938) );
  INV_X1 U13993 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10936) );
  INV_X1 U13994 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14075) );
  OAI22_X1 U13995 ( .A1(n10936), .A2(n19724), .B1(n10892), .B2(n14075), .ZN(
        n10937) );
  NOR2_X1 U13996 ( .A1(n10938), .A2(n10937), .ZN(n10945) );
  INV_X1 U13997 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10940) );
  INV_X1 U13998 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10939) );
  OAI22_X1 U13999 ( .A1(n10940), .A2(n15615), .B1(n13440), .B2(n10939), .ZN(
        n10943) );
  INV_X1 U14000 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10941) );
  INV_X1 U14001 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14073) );
  OAI22_X1 U14002 ( .A1(n10941), .A2(n10895), .B1(n19675), .B2(n14073), .ZN(
        n10942) );
  NOR2_X1 U14003 ( .A1(n10943), .A2(n10942), .ZN(n10944) );
  NAND4_X1 U14004 ( .A1(n10947), .A2(n10946), .A3(n10945), .A4(n10944), .ZN(
        n10959) );
  AOI22_X1 U14005 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10662), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U14006 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U14007 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U14008 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10948) );
  NAND4_X1 U14009 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .ZN(
        n10957) );
  AOI22_X1 U14010 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10911), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U14011 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14013 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U14014 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10956) );
  INV_X1 U14015 ( .A(n11029), .ZN(n11348) );
  NAND2_X1 U14016 ( .A1(n11348), .A2(n14062), .ZN(n10958) );
  NAND2_X1 U14017 ( .A1(n10961), .A2(n15537), .ZN(n10960) );
  NAND2_X1 U14018 ( .A1(n15517), .A2(n9601), .ZN(n15219) );
  NAND3_X1 U14019 ( .A1(n15220), .A2(n15219), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10983) );
  NAND2_X1 U14020 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10966) );
  NAND2_X1 U14021 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10965) );
  NAND2_X1 U14022 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10964) );
  NAND2_X1 U14023 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10963) );
  NAND2_X1 U14024 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U14025 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10969) );
  NAND2_X1 U14026 ( .A1(n10906), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10968) );
  NAND2_X1 U14027 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10967) );
  NAND2_X1 U14028 ( .A1(n10668), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10974) );
  NAND2_X1 U14029 ( .A1(n13886), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10973) );
  NAND2_X1 U14030 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10972) );
  NAND2_X1 U14031 ( .A1(n10669), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14032 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10978) );
  NAND2_X1 U14033 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10977) );
  NAND2_X1 U14034 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10976) );
  NAND2_X1 U14035 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10975) );
  XNOR2_X1 U14036 ( .A(n10984), .B(n11587), .ZN(n15222) );
  NAND2_X1 U14037 ( .A1(n10983), .A2(n15222), .ZN(n16290) );
  INV_X1 U14038 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16324) );
  OAI21_X1 U14039 ( .B1(n10984), .B2(n11587), .A(n16324), .ZN(n10985) );
  NAND2_X1 U14040 ( .A1(n11596), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11041) );
  NAND2_X1 U14041 ( .A1(n10985), .A2(n10991), .ZN(n16292) );
  INV_X1 U14042 ( .A(n16292), .ZN(n10986) );
  NAND2_X1 U14043 ( .A1(n15219), .A2(n10987), .ZN(n10989) );
  INV_X1 U14044 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16325) );
  NAND2_X1 U14045 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  NAND2_X1 U14046 ( .A1(n16290), .A2(n10990), .ZN(n10992) );
  INV_X1 U14047 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15478) );
  NAND2_X1 U14048 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15436) );
  INV_X1 U14049 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15414) );
  NOR2_X1 U14050 ( .A1(n15436), .A2(n15414), .ZN(n11488) );
  INV_X1 U14051 ( .A(n11488), .ZN(n11302) );
  NAND2_X1 U14052 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15372) );
  INV_X1 U14053 ( .A(n15372), .ZN(n10993) );
  NAND2_X1 U14054 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U14055 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15293) );
  INV_X1 U14056 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11491) );
  INV_X1 U14057 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15251) );
  INV_X1 U14058 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11576) );
  XNOR2_X1 U14059 ( .A(n11547), .B(n11576), .ZN(n11515) );
  MUX2_X1 U14060 ( .A(n10996), .B(n13651), .S(n11593), .Z(n11002) );
  NAND2_X1 U14061 ( .A1(n10997), .A2(n11021), .ZN(n10999) );
  OR2_X1 U14062 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(
        n11000) );
  INV_X1 U14063 ( .A(n11016), .ZN(n11001) );
  OAI21_X1 U14064 ( .B1(n11002), .B2(n11008), .A(n11001), .ZN(n13652) );
  MUX2_X1 U14065 ( .A(n11004), .B(n11003), .S(n11593), .Z(n13670) );
  INV_X1 U14066 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12986) );
  NOR2_X1 U14067 ( .A1(n13670), .A2(n12986), .ZN(n12985) );
  INV_X1 U14068 ( .A(n12985), .ZN(n11006) );
  INV_X1 U14069 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12983) );
  NAND3_X1 U14070 ( .A1(n11593), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U14071 ( .A1(n11009), .A2(n11005), .ZN(n13747) );
  NOR2_X1 U14072 ( .A1(n11006), .A2(n13747), .ZN(n11007) );
  INV_X1 U14073 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13776) );
  XNOR2_X1 U14074 ( .A(n13747), .B(n11006), .ZN(n13001) );
  NOR2_X1 U14075 ( .A1(n13776), .A2(n13001), .ZN(n13000) );
  NOR2_X1 U14076 ( .A1(n11007), .A2(n13000), .ZN(n12960) );
  INV_X1 U14077 ( .A(n11008), .ZN(n11012) );
  NAND2_X1 U14078 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  NAND2_X1 U14079 ( .A1(n11012), .A2(n11011), .ZN(n13736) );
  OAI21_X1 U14080 ( .B1(n12960), .B2(n13736), .A(n19255), .ZN(n11013) );
  NAND2_X1 U14081 ( .A1(n12960), .A2(n13736), .ZN(n12959) );
  AND2_X1 U14082 ( .A1(n11013), .A2(n12959), .ZN(n13817) );
  INV_X1 U14083 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11172) );
  MUX2_X1 U14084 ( .A(n11014), .B(n11172), .S(n11593), .Z(n11015) );
  OAI21_X1 U14085 ( .B1(n11016), .B2(n11015), .A(n11023), .ZN(n13696) );
  XNOR2_X1 U14086 ( .A(n13696), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15226) );
  NAND2_X1 U14087 ( .A1(n15227), .A2(n15226), .ZN(n11018) );
  OR2_X1 U14088 ( .A1(n13696), .A2(n15555), .ZN(n11017) );
  NAND2_X1 U14089 ( .A1(n11018), .A2(n11017), .ZN(n15536) );
  NAND2_X1 U14090 ( .A1(n11019), .A2(n11587), .ZN(n11025) );
  MUX2_X1 U14091 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n11347), .S(n11021), .Z(
        n11022) );
  AND2_X1 U14092 ( .A1(n11023), .A2(n11022), .ZN(n11024) );
  OR2_X1 U14093 ( .A1(n11024), .A2(n11031), .ZN(n19113) );
  NAND2_X1 U14094 ( .A1(n11025), .A2(n19113), .ZN(n11027) );
  AND2_X1 U14095 ( .A1(n11027), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11028) );
  INV_X1 U14096 ( .A(n15531), .ZN(n11037) );
  INV_X1 U14097 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11182) );
  MUX2_X1 U14098 ( .A(n11029), .B(n11182), .S(n11593), .Z(n11030) );
  OR2_X1 U14099 ( .A1(n11031), .A2(n11030), .ZN(n11032) );
  NAND2_X1 U14100 ( .A1(n11038), .A2(n11032), .ZN(n19098) );
  XNOR2_X1 U14101 ( .A(n11034), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15532) );
  INV_X1 U14102 ( .A(n15532), .ZN(n11036) );
  INV_X1 U14103 ( .A(n11034), .ZN(n11035) );
  INV_X1 U14104 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15526) );
  MUX2_X1 U14105 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n11587), .S(n11021), .Z(
        n11042) );
  INV_X1 U14106 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11189) );
  NOR2_X1 U14107 ( .A1(n11021), .A2(n11189), .ZN(n11039) );
  OR2_X2 U14108 ( .A1(n11044), .A2(n11039), .ZN(n11049) );
  NAND2_X1 U14109 ( .A1(n11044), .A2(n11039), .ZN(n11040) );
  NAND2_X1 U14110 ( .A1(n11049), .A2(n11040), .ZN(n13716) );
  NOR2_X1 U14111 ( .A1(n13716), .A2(n11041), .ZN(n16284) );
  NAND2_X1 U14112 ( .A1(n11038), .A2(n11042), .ZN(n11043) );
  AND2_X1 U14113 ( .A1(n11044), .A2(n11043), .ZN(n19087) );
  INV_X1 U14114 ( .A(n13716), .ZN(n11045) );
  AOI21_X1 U14115 ( .B1(n11045), .B2(n11596), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16285) );
  NOR2_X1 U14116 ( .A1(n19087), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15214) );
  NAND2_X1 U14117 ( .A1(n11593), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11048) );
  XNOR2_X1 U14118 ( .A(n11049), .B(n11048), .ZN(n19073) );
  NAND2_X1 U14119 ( .A1(n19073), .A2(n11596), .ZN(n11054) );
  INV_X1 U14120 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U14121 ( .A1(n11054), .A2(n11301), .ZN(n13790) );
  NOR2_X2 U14122 ( .A1(n11049), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11051) );
  INV_X1 U14123 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U14124 ( .A1(n11593), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11050) );
  OAI21_X1 U14125 ( .B1(n11051), .B2(n11050), .A(n11130), .ZN(n11052) );
  OR2_X1 U14126 ( .A1(n11056), .A2(n11052), .ZN(n19061) );
  INV_X1 U14127 ( .A(n19061), .ZN(n11053) );
  AOI21_X1 U14128 ( .B1(n11053), .B2(n11596), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15480) );
  NAND3_X1 U14129 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n11596), .ZN(n15481) );
  INV_X1 U14130 ( .A(n11054), .ZN(n11055) );
  NAND2_X1 U14131 ( .A1(n11055), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15479) );
  NAND2_X1 U14132 ( .A1(n11593), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11057) );
  INV_X1 U14133 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U14134 ( .B1(n11056), .B2(n11057), .A(n9918), .ZN(n19052) );
  NOR2_X1 U14135 ( .A1(n19052), .A2(n11587), .ZN(n15207) );
  NAND2_X1 U14136 ( .A1(n11593), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11058) );
  NAND2_X1 U14137 ( .A1(n11593), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11085) );
  INV_X1 U14138 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11219) );
  INV_X1 U14139 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19015) );
  NAND2_X1 U14140 ( .A1(n11219), .A2(n19015), .ZN(n11060) );
  INV_X1 U14141 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11225) );
  NAND2_X1 U14142 ( .A1(n11593), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11070) );
  INV_X1 U14143 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16256) );
  NOR2_X1 U14144 ( .A1(n11021), .A2(n16256), .ZN(n11067) );
  INV_X1 U14145 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11236) );
  NOR2_X1 U14146 ( .A1(n11021), .A2(n11236), .ZN(n11064) );
  NAND2_X1 U14147 ( .A1(n11062), .A2(n11061), .ZN(n11063) );
  INV_X1 U14148 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11240) );
  AND2_X1 U14149 ( .A1(n11063), .A2(n11117), .ZN(n18965) );
  INV_X1 U14150 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15339) );
  NAND2_X1 U14151 ( .A1(n11099), .A2(n15339), .ZN(n15091) );
  AND2_X1 U14152 ( .A1(n11069), .A2(n11064), .ZN(n11066) );
  OR2_X1 U14153 ( .A1(n11066), .A2(n11065), .ZN(n18979) );
  INV_X1 U14154 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15348) );
  OAI21_X1 U14155 ( .B1(n18979), .B2(n11587), .A(n15348), .ZN(n15117) );
  NAND2_X1 U14156 ( .A1(n11072), .A2(n11067), .ZN(n11068) );
  AND2_X1 U14157 ( .A1(n11069), .A2(n11068), .ZN(n18990) );
  NAND2_X1 U14158 ( .A1(n18990), .A2(n11596), .ZN(n11109) );
  INV_X1 U14159 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U14160 ( .A1(n11109), .A2(n15355), .ZN(n15126) );
  NAND2_X1 U14161 ( .A1(n15117), .A2(n15126), .ZN(n15088) );
  OR2_X1 U14162 ( .A1(n11071), .A2(n11070), .ZN(n11073) );
  AND2_X1 U14163 ( .A1(n11073), .A2(n11072), .ZN(n19000) );
  NAND2_X1 U14164 ( .A1(n19000), .A2(n11596), .ZN(n11102) );
  INV_X1 U14165 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15376) );
  NAND2_X1 U14166 ( .A1(n11102), .A2(n15376), .ZN(n15085) );
  NAND2_X1 U14167 ( .A1(n11593), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11075) );
  OAI211_X1 U14168 ( .C1(n11077), .C2(n11075), .A(n11130), .B(n11074), .ZN(
        n14812) );
  OR2_X1 U14169 ( .A1(n14812), .A2(n11587), .ZN(n11076) );
  XNOR2_X1 U14170 ( .A(n11076), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15083) );
  INV_X1 U14171 ( .A(n11077), .ZN(n11080) );
  AND2_X1 U14172 ( .A1(n11089), .A2(n11219), .ZN(n11091) );
  INV_X1 U14173 ( .A(n11091), .ZN(n11078) );
  NAND3_X1 U14174 ( .A1(n11078), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n11593), 
        .ZN(n11079) );
  NAND2_X1 U14175 ( .A1(n11080), .A2(n11079), .ZN(n19016) );
  OR2_X1 U14176 ( .A1(n19016), .A2(n11587), .ZN(n11081) );
  INV_X1 U14177 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15403) );
  NAND2_X1 U14178 ( .A1(n11081), .A2(n15403), .ZN(n15163) );
  NAND2_X1 U14179 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n11082), .ZN(n11083) );
  NOR2_X1 U14180 ( .A1(n11021), .A2(n11083), .ZN(n11084) );
  NOR2_X1 U14181 ( .A1(n11086), .A2(n11084), .ZN(n14822) );
  NAND2_X1 U14182 ( .A1(n14822), .A2(n11596), .ZN(n15078) );
  INV_X1 U14183 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15447) );
  NAND2_X1 U14184 ( .A1(n15078), .A2(n15447), .ZN(n15079) );
  NOR2_X1 U14185 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  NOR2_X1 U14186 ( .A1(n11089), .A2(n11087), .ZN(n19038) );
  NAND2_X1 U14187 ( .A1(n19038), .A2(n11596), .ZN(n11088) );
  INV_X1 U14188 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11106) );
  NAND2_X1 U14189 ( .A1(n11088), .A2(n11106), .ZN(n15190) );
  AND3_X1 U14190 ( .A1(n15163), .A2(n15079), .A3(n15190), .ZN(n11093) );
  NOR2_X1 U14191 ( .A1(n11089), .A2(n11219), .ZN(n11090) );
  MUX2_X1 U14192 ( .A(n11090), .B(n11089), .S(n11021), .Z(n11092) );
  NOR2_X1 U14193 ( .A1(n11092), .A2(n11091), .ZN(n19029) );
  NAND2_X1 U14194 ( .A1(n19029), .A2(n11596), .ZN(n11108) );
  NAND2_X1 U14195 ( .A1(n11108), .A2(n15414), .ZN(n15172) );
  NAND4_X1 U14196 ( .A1(n15085), .A2(n15083), .A3(n11093), .A4(n15172), .ZN(
        n11094) );
  NOR2_X1 U14197 ( .A1(n15088), .A2(n11094), .ZN(n11096) );
  NAND3_X1 U14198 ( .A1(n11117), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11593), 
        .ZN(n11095) );
  OAI211_X1 U14199 ( .C1(n11117), .C2(P2_EBX_REG_21__SCAN_IN), .A(n11095), .B(
        n11130), .ZN(n14793) );
  OR2_X1 U14200 ( .A1(n14793), .A2(n11587), .ZN(n11098) );
  INV_X1 U14201 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15319) );
  NAND2_X1 U14202 ( .A1(n11098), .A2(n15319), .ZN(n15094) );
  NAND3_X1 U14203 ( .A1(n15091), .A2(n11096), .A3(n15094), .ZN(n11097) );
  NAND2_X1 U14204 ( .A1(n15076), .A2(n15447), .ZN(n11115) );
  INV_X1 U14205 ( .A(n18979), .ZN(n11101) );
  NOR2_X1 U14206 ( .A1(n11587), .A2(n15348), .ZN(n11100) );
  NAND2_X1 U14207 ( .A1(n11101), .A2(n11100), .ZN(n15116) );
  INV_X1 U14208 ( .A(n11102), .ZN(n11103) );
  NAND2_X1 U14209 ( .A1(n11103), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15086) );
  INV_X1 U14210 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15388) );
  OR2_X1 U14211 ( .A1(n11587), .A2(n15388), .ZN(n11104) );
  OR2_X1 U14212 ( .A1(n14812), .A2(n11104), .ZN(n15084) );
  OR2_X1 U14213 ( .A1(n11587), .A2(n15403), .ZN(n11105) );
  NOR2_X1 U14214 ( .A1(n11587), .A2(n11106), .ZN(n11107) );
  NAND2_X1 U14215 ( .A1(n19038), .A2(n11107), .ZN(n15189) );
  AND4_X1 U14216 ( .A1(n15086), .A2(n15084), .A3(n15162), .A4(n15189), .ZN(
        n11111) );
  INV_X1 U14217 ( .A(n11109), .ZN(n11110) );
  NAND2_X1 U14218 ( .A1(n11110), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15127) );
  NAND4_X1 U14219 ( .A1(n15116), .A2(n11111), .A3(n15173), .A4(n15127), .ZN(
        n11112) );
  NOR2_X1 U14220 ( .A1(n15093), .A2(n11112), .ZN(n11113) );
  NAND2_X1 U14221 ( .A1(n9655), .A2(n11113), .ZN(n11114) );
  NAND2_X1 U14222 ( .A1(n11130), .A2(n9653), .ZN(n11118) );
  NAND2_X1 U14223 ( .A1(n11593), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U14224 ( .A1(n9925), .A2(n9653), .ZN(n11120) );
  AND2_X1 U14225 ( .A1(n11122), .A2(n11120), .ZN(n14783) );
  AOI21_X1 U14226 ( .B1(n14783), .B2(n11596), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15066) );
  NAND3_X1 U14227 ( .A1(n14783), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11596), .ZN(n15067) );
  INV_X1 U14228 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11250) );
  NOR2_X1 U14229 ( .A1(n11021), .A2(n11250), .ZN(n11121) );
  NAND2_X1 U14230 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  AND2_X1 U14231 ( .A1(n11129), .A2(n11123), .ZN(n14772) );
  NAND2_X1 U14232 ( .A1(n14772), .A2(n11596), .ZN(n11124) );
  XNOR2_X1 U14233 ( .A(n11124), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15057) );
  INV_X1 U14234 ( .A(n14772), .ZN(n11125) );
  INV_X1 U14235 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15296) );
  NOR3_X1 U14236 ( .A1(n11125), .A2(n11587), .A3(n15296), .ZN(n11126) );
  INV_X1 U14237 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14747) );
  NOR2_X1 U14238 ( .A1(n11021), .A2(n14747), .ZN(n11128) );
  INV_X1 U14239 ( .A(n11129), .ZN(n11127) );
  MUX2_X1 U14240 ( .A(n11128), .B(n14747), .S(n11127), .Z(n14750) );
  NAND2_X1 U14241 ( .A1(n11130), .A2(n11596), .ZN(n11138) );
  NOR2_X1 U14242 ( .A1(n14750), .A2(n11138), .ZN(n15047) );
  INV_X1 U14243 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11257) );
  INV_X1 U14244 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n14715) );
  INV_X1 U14245 ( .A(n11130), .ZN(n11131) );
  NOR2_X1 U14246 ( .A1(n11147), .A2(n11131), .ZN(n11595) );
  NAND2_X1 U14247 ( .A1(n11593), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11132) );
  OR2_X1 U14248 ( .A1(n11133), .A2(n11132), .ZN(n11134) );
  INV_X1 U14249 ( .A(n14724), .ZN(n11135) );
  NOR2_X1 U14250 ( .A1(n11135), .A2(n11587), .ZN(n11136) );
  NAND3_X1 U14251 ( .A1(n14724), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11596), .ZN(n11145) );
  OAI21_X1 U14252 ( .B1(n11136), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11145), .ZN(n15025) );
  NAND2_X1 U14253 ( .A1(n11593), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11137) );
  MUX2_X1 U14254 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n11137), .S(n9660), .Z(
        n14737) );
  INV_X1 U14255 ( .A(n11138), .ZN(n11139) );
  NOR2_X1 U14256 ( .A1(n11143), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15036) );
  INV_X1 U14257 ( .A(n11143), .ZN(n11144) );
  INV_X1 U14258 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U14259 ( .A1(n11145), .A2(n15034), .ZN(n11580) );
  INV_X1 U14260 ( .A(n11595), .ZN(n11146) );
  NAND2_X1 U14261 ( .A1(n11593), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U14262 ( .A1(n11146), .A2(n11148), .ZN(n11155) );
  INV_X1 U14263 ( .A(n11147), .ZN(n11150) );
  INV_X1 U14264 ( .A(n11148), .ZN(n11149) );
  NAND2_X1 U14265 ( .A1(n11150), .A2(n11149), .ZN(n11151) );
  NAND2_X1 U14266 ( .A1(n11155), .A2(n11151), .ZN(n14707) );
  NOR2_X1 U14267 ( .A1(n14707), .A2(n11587), .ZN(n11571) );
  XNOR2_X1 U14268 ( .A(n11153), .B(n11571), .ZN(n11522) );
  INV_X1 U14269 ( .A(n11571), .ZN(n11152) );
  INV_X1 U14270 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U14271 ( .A1(n11593), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11157) );
  NAND2_X1 U14272 ( .A1(n11156), .A2(n11157), .ZN(n11582) );
  INV_X1 U14273 ( .A(n11157), .ZN(n11158) );
  NAND2_X1 U14274 ( .A1(n11155), .A2(n11158), .ZN(n11159) );
  NAND2_X1 U14275 ( .A1(n11582), .A2(n11159), .ZN(n14695) );
  NOR2_X1 U14276 ( .A1(n14695), .A2(n11587), .ZN(n11575) );
  XNOR2_X1 U14277 ( .A(n11575), .B(n11576), .ZN(n11160) );
  XNOR2_X1 U14278 ( .A(n11161), .B(n11160), .ZN(n11514) );
  NOR2_X1 U14279 ( .A1(n9591), .A2(n11162), .ZN(n19905) );
  NAND2_X1 U14280 ( .A1(n11514), .A2(n16338), .ZN(n11499) );
  INV_X1 U14281 ( .A(n11165), .ZN(n11166) );
  OR2_X1 U14282 ( .A1(n11167), .A2(n11166), .ZN(n11168) );
  NAND2_X1 U14283 ( .A1(n11169), .A2(n11168), .ZN(n13688) );
  NAND2_X1 U14284 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U14285 ( .A1(n9577), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11170) );
  OAI211_X1 U14286 ( .C1(n11258), .C2(n11172), .A(n11171), .B(n11170), .ZN(
        n11173) );
  AOI21_X1 U14287 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11173), .ZN(n13687) );
  INV_X1 U14288 ( .A(n13687), .ZN(n11174) );
  INV_X1 U14289 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14290 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11176) );
  NAND2_X1 U14291 ( .A1(n9577), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U14292 ( .C1(n11258), .C2(n11177), .A(n11176), .B(n11175), .ZN(
        n11178) );
  AOI21_X1 U14293 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11178), .ZN(n13196) );
  NAND2_X1 U14294 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U14295 ( .A1(n9577), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11180) );
  OAI211_X1 U14296 ( .C1(n11258), .C2(n11182), .A(n11181), .B(n11180), .ZN(
        n11183) );
  AOI21_X1 U14297 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11183), .ZN(n13282) );
  INV_X1 U14298 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U14299 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11185) );
  AOI22_X1 U14300 ( .A1(n9577), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11184) );
  OAI211_X1 U14301 ( .C1(n11258), .C2(n11186), .A(n11185), .B(n11184), .ZN(
        n13349) );
  NAND2_X1 U14302 ( .A1(n13350), .A2(n13349), .ZN(n13704) );
  NAND2_X1 U14303 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U14304 ( .A1(n9577), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11187) );
  OAI211_X1 U14305 ( .C1(n11258), .C2(n11189), .A(n11188), .B(n11187), .ZN(
        n11190) );
  AOI21_X1 U14306 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11190), .ZN(n13705) );
  NAND2_X1 U14307 ( .A1(n11192), .A2(n11191), .ZN(n13515) );
  INV_X1 U14308 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11195) );
  NAND2_X1 U14309 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11194) );
  NAND2_X1 U14310 ( .A1(n9577), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11193) );
  OAI211_X1 U14311 ( .C1(n11258), .C2(n11195), .A(n11194), .B(n11193), .ZN(
        n11196) );
  AOI21_X1 U14312 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11196), .ZN(n13516) );
  NAND2_X1 U14313 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U14314 ( .A1(n9577), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11197) );
  OAI211_X1 U14315 ( .C1(n11258), .C2(n11199), .A(n11198), .B(n11197), .ZN(
        n11200) );
  AOI21_X1 U14316 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11200), .ZN(n15487) );
  NAND2_X1 U14317 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11205) );
  AOI22_X1 U14318 ( .A1(n9577), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11203) );
  NAND2_X1 U14319 ( .A1(n11201), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11202) );
  AND2_X1 U14320 ( .A1(n11203), .A2(n11202), .ZN(n11204) );
  NAND2_X1 U14321 ( .A1(n11205), .A2(n11204), .ZN(n13586) );
  INV_X1 U14322 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U14323 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14324 ( .A1(n9577), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11207) );
  OAI211_X1 U14325 ( .C1(n11258), .C2(n11209), .A(n11208), .B(n11207), .ZN(
        n11210) );
  AOI21_X1 U14326 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11210), .ZN(n14819) );
  INV_X1 U14327 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U14328 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U14329 ( .A1(n9577), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11213) );
  OAI211_X1 U14330 ( .C1(n11258), .C2(n11215), .A(n11214), .B(n11213), .ZN(
        n11216) );
  AOI21_X1 U14331 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11216), .ZN(n14913) );
  NAND2_X1 U14332 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11218) );
  AOI22_X1 U14333 ( .A1(n9577), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11217) );
  OAI211_X1 U14334 ( .C1(n11258), .C2(n11219), .A(n11218), .B(n11217), .ZN(
        n15178) );
  NAND2_X1 U14335 ( .A1(n15179), .A2(n15178), .ZN(n15181) );
  NAND2_X1 U14336 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11221) );
  NAND2_X1 U14337 ( .A1(n9577), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11220) );
  OAI211_X1 U14338 ( .C1(n11258), .C2(n19015), .A(n11221), .B(n11220), .ZN(
        n11222) );
  AOI21_X1 U14339 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11222), .ZN(n14904) );
  NAND2_X1 U14340 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14341 ( .A1(n9577), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11223) );
  OAI211_X1 U14342 ( .C1(n11258), .C2(n11225), .A(n11224), .B(n11223), .ZN(
        n11226) );
  AOI21_X1 U14343 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11226), .ZN(n14802) );
  NAND2_X1 U14344 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11231) );
  AOI22_X1 U14345 ( .A1(n9577), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11229) );
  NAND2_X1 U14346 ( .A1(n11201), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11228) );
  AND2_X1 U14347 ( .A1(n11229), .A2(n11228), .ZN(n11230) );
  NAND2_X1 U14348 ( .A1(n11231), .A2(n11230), .ZN(n14892) );
  NAND2_X1 U14349 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11233) );
  AOI22_X1 U14350 ( .A1(n9577), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11232) );
  OAI211_X1 U14351 ( .C1(n11258), .C2(n16256), .A(n11233), .B(n11232), .ZN(
        n15133) );
  NAND2_X1 U14352 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U14353 ( .A1(n9577), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11234) );
  OAI211_X1 U14354 ( .C1(n11258), .C2(n11236), .A(n11235), .B(n11234), .ZN(
        n11237) );
  AOI21_X1 U14355 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11237), .ZN(n14887) );
  NAND2_X1 U14356 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14357 ( .A1(n9577), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11238) );
  OAI211_X1 U14358 ( .C1(n11258), .C2(n11240), .A(n11239), .B(n11238), .ZN(
        n11241) );
  AOI21_X1 U14359 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11241), .ZN(n15109) );
  INV_X1 U14360 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U14361 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U14362 ( .A1(n9577), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11242) );
  OAI211_X1 U14363 ( .C1(n11258), .C2(n14879), .A(n11243), .B(n11242), .ZN(
        n11244) );
  AOI21_X1 U14364 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11244), .ZN(n14788) );
  INV_X1 U14365 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11247) );
  NAND2_X1 U14366 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11246) );
  AOI22_X1 U14367 ( .A1(n9577), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11245) );
  OAI211_X1 U14368 ( .C1(n11258), .C2(n11247), .A(n11246), .B(n11245), .ZN(
        n14775) );
  NAND2_X1 U14369 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U14370 ( .A1(n9577), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11248) );
  OAI211_X1 U14371 ( .C1(n11258), .C2(n11250), .A(n11249), .B(n11248), .ZN(
        n11251) );
  AOI21_X1 U14372 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11251), .ZN(n14759) );
  NAND2_X1 U14373 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U14374 ( .A1(n9577), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11252) );
  OAI211_X1 U14375 ( .C1(n11258), .C2(n14747), .A(n11253), .B(n11252), .ZN(
        n11254) );
  AOI21_X1 U14376 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11254), .ZN(n14740) );
  NAND2_X1 U14377 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11256) );
  AOI22_X1 U14378 ( .A1(n9577), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11255) );
  OAI211_X1 U14379 ( .C1(n11258), .C2(n11257), .A(n11256), .B(n11255), .ZN(
        n14726) );
  NAND2_X1 U14380 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11262) );
  AOI22_X1 U14381 ( .A1(n9577), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11260) );
  NAND2_X1 U14382 ( .A1(n11201), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11259) );
  AND2_X1 U14383 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  NAND2_X1 U14384 ( .A1(n11262), .A2(n11261), .ZN(n14711) );
  NAND2_X1 U14385 ( .A1(n11564), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11266) );
  AOI22_X1 U14386 ( .A1(n9577), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11264) );
  NAND2_X1 U14387 ( .A1(n11201), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11263) );
  AND2_X1 U14388 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  NAND2_X1 U14389 ( .A1(n11266), .A2(n11265), .ZN(n11531) );
  INV_X1 U14390 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14391 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U14392 ( .A1(n9577), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11267) );
  OAI211_X1 U14393 ( .C1(n11258), .C2(n11269), .A(n11268), .B(n11267), .ZN(
        n11270) );
  AOI21_X1 U14394 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11270), .ZN(n11272) );
  NAND2_X1 U14395 ( .A1(n11271), .A2(n11272), .ZN(n11273) );
  NAND2_X1 U14396 ( .A1(n14836), .A2(n11273), .ZN(n14848) );
  NAND2_X1 U14397 ( .A1(n11275), .A2(n14062), .ZN(n11277) );
  INV_X1 U14398 ( .A(n11276), .ZN(n13175) );
  NAND2_X1 U14399 ( .A1(n11277), .A2(n13175), .ZN(n11278) );
  NAND2_X1 U14400 ( .A1(n11279), .A2(n21042), .ZN(n13780) );
  NAND2_X1 U14401 ( .A1(n13780), .A2(n11280), .ZN(n11294) );
  INV_X1 U14402 ( .A(n11281), .ZN(n11283) );
  NAND3_X1 U14403 ( .A1(n11283), .A2(n10722), .A3(n11282), .ZN(n11291) );
  NAND2_X1 U14404 ( .A1(n11284), .A2(n14062), .ZN(n11285) );
  NAND2_X1 U14405 ( .A1(n10716), .A2(n11285), .ZN(n11287) );
  AOI21_X1 U14406 ( .B1(n11287), .B2(n11286), .A(n10731), .ZN(n11289) );
  OAI22_X1 U14407 ( .A1(n11286), .A2(n10704), .B1(n10713), .B2(n10722), .ZN(
        n11288) );
  NOR2_X1 U14408 ( .A1(n11289), .A2(n11288), .ZN(n11290) );
  NAND2_X1 U14409 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  AOI21_X1 U14410 ( .B1(n11294), .B2(n11293), .A(n11292), .ZN(n15593) );
  NAND2_X1 U14411 ( .A1(n15593), .A2(n11295), .ZN(n11296) );
  NAND2_X1 U14412 ( .A1(n11297), .A2(n11314), .ZN(n11298) );
  INV_X1 U14413 ( .A(n13181), .ZN(n16358) );
  NAND2_X1 U14414 ( .A1(n11308), .A2(n16358), .ZN(n15378) );
  NAND2_X1 U14415 ( .A1(n19869), .A2(n16381), .ZN(n11494) );
  INV_X1 U14416 ( .A(n11494), .ZN(n16322) );
  NOR2_X1 U14417 ( .A1(n11308), .A2(n16322), .ZN(n15567) );
  NAND3_X1 U14418 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15528) );
  NOR2_X1 U14419 ( .A1(n15526), .A2(n15528), .ZN(n15500) );
  NAND3_X1 U14420 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n15500), .ZN(n11487) );
  NAND2_X1 U14421 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19275) );
  NAND2_X1 U14422 ( .A1(n19255), .A2(n19275), .ZN(n19269) );
  AOI21_X1 U14423 ( .B1(n11300), .B2(n19275), .A(n15567), .ZN(n19256) );
  NAND2_X1 U14424 ( .A1(n11300), .A2(n19255), .ZN(n19276) );
  OAI211_X1 U14425 ( .C1(n15378), .C2(n19269), .A(n19256), .B(n19276), .ZN(
        n15520) );
  AOI211_X1 U14426 ( .C1(n15411), .C2(n11487), .A(n15520), .B(n11301), .ZN(
        n15459) );
  NAND3_X1 U14427 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n15459), .ZN(n15412) );
  NOR2_X1 U14428 ( .A1(n15412), .A2(n11302), .ZN(n15363) );
  NOR2_X1 U14429 ( .A1(n15376), .A2(n15372), .ZN(n15364) );
  NAND3_X1 U14430 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15363), .A3(
        n15364), .ZN(n15328) );
  NOR2_X1 U14431 ( .A1(n15348), .A2(n15339), .ZN(n15334) );
  NAND2_X1 U14432 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15334), .ZN(
        n11490) );
  OAI21_X1 U14433 ( .B1(n15328), .B2(n11490), .A(n15411), .ZN(n15320) );
  NAND2_X1 U14434 ( .A1(n15411), .A2(n15293), .ZN(n11303) );
  AND2_X1 U14435 ( .A1(n11303), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14436 ( .A1(n15320), .A2(n11304), .ZN(n15281) );
  NAND2_X1 U14437 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11493) );
  INV_X1 U14438 ( .A(n15565), .ZN(n15382) );
  NAND2_X1 U14439 ( .A1(n15320), .A2(n15382), .ZN(n15271) );
  OAI21_X1 U14440 ( .B1(n15281), .B2(n11493), .A(n15271), .ZN(n11305) );
  AND2_X1 U14441 ( .A1(n11305), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11529) );
  INV_X1 U14442 ( .A(n15271), .ZN(n15253) );
  NOR2_X1 U14443 ( .A1(n11529), .A2(n15253), .ZN(n15236) );
  AND2_X1 U14444 ( .A1(n11306), .A2(n10741), .ZN(n12946) );
  INV_X1 U14445 ( .A(n12946), .ZN(n16366) );
  OAI21_X1 U14446 ( .B1(n14062), .B2(n9594), .A(n16366), .ZN(n11307) );
  NAND2_X1 U14447 ( .A1(n11308), .A2(n11307), .ZN(n16331) );
  NAND2_X1 U14448 ( .A1(n11602), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11312) );
  INV_X1 U14449 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13135) );
  NAND2_X1 U14450 ( .A1(n21042), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11309) );
  OAI211_X1 U14451 ( .C1(n13125), .C2(n13135), .A(n11309), .B(n19678), .ZN(
        n11310) );
  INV_X1 U14452 ( .A(n11310), .ZN(n11311) );
  NAND2_X1 U14453 ( .A1(n11312), .A2(n11311), .ZN(n13130) );
  NAND2_X1 U14454 ( .A1(n11313), .A2(n11021), .ZN(n11321) );
  MUX2_X1 U14455 ( .A(n13125), .B(n19900), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11315) );
  AND2_X2 U14456 ( .A1(n21042), .A2(n19678), .ZN(n11318) );
  NAND2_X1 U14457 ( .A1(n11314), .A2(n11318), .ZN(n11330) );
  NAND2_X1 U14458 ( .A1(n11602), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11320) );
  NOR2_X1 U14459 ( .A1(n13125), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14460 ( .A1(n11317), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11319) );
  NAND2_X1 U14461 ( .A1(n11320), .A2(n11319), .ZN(n11326) );
  OR2_X1 U14462 ( .A1(n11322), .A2(n11321), .ZN(n11325) );
  NAND2_X1 U14463 ( .A1(n11284), .A2(n13125), .ZN(n11323) );
  MUX2_X1 U14464 ( .A(n11323), .B(n19891), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11324) );
  NAND2_X1 U14465 ( .A1(n11325), .A2(n11324), .ZN(n13264) );
  NOR2_X1 U14466 ( .A1(n13265), .A2(n13264), .ZN(n11328) );
  NOR2_X1 U14467 ( .A1(n13127), .A2(n11326), .ZN(n11327) );
  NAND2_X1 U14468 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11329) );
  OAI211_X1 U14469 ( .C1(n11321), .C2(n11331), .A(n11330), .B(n11329), .ZN(
        n11333) );
  XNOR2_X1 U14470 ( .A(n11332), .B(n11333), .ZN(n13263) );
  INV_X1 U14471 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19250) );
  INV_X1 U14472 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19804) );
  OAI222_X1 U14473 ( .A1(n11383), .A2(n19255), .B1(n11382), .B2(n19250), .C1(
        n11606), .C2(n19804), .ZN(n13262) );
  NOR2_X1 U14474 ( .A1(n13263), .A2(n13262), .ZN(n13261) );
  NOR2_X1 U14475 ( .A1(n11332), .A2(n11333), .ZN(n11334) );
  INV_X1 U14476 ( .A(n11335), .ZN(n11340) );
  AOI22_X1 U14477 ( .A1(n11318), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11337) );
  NAND2_X1 U14478 ( .A1(n11357), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11336) );
  AND2_X1 U14479 ( .A1(n11337), .A2(n11336), .ZN(n11339) );
  NAND2_X1 U14480 ( .A1(n11602), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11338) );
  OAI211_X1 U14481 ( .C1(n11321), .C2(n11340), .A(n11339), .B(n11338), .ZN(
        n13636) );
  NAND2_X1 U14482 ( .A1(n11602), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14483 ( .A1(n11357), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11343) );
  OR2_X1 U14484 ( .A1(n11321), .A2(n11341), .ZN(n11342) );
  NAND2_X1 U14485 ( .A1(n11602), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14486 ( .A1(n11357), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11345) );
  OAI211_X1 U14487 ( .C1(n11321), .C2(n11347), .A(n11346), .B(n11345), .ZN(
        n15547) );
  OR2_X1 U14488 ( .A1(n11321), .A2(n11348), .ZN(n11349) );
  NAND2_X1 U14489 ( .A1(n11602), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14490 ( .A1(n11357), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U14491 ( .A1(n11352), .A2(n11351), .ZN(n15523) );
  NAND2_X1 U14492 ( .A1(n15522), .A2(n15523), .ZN(n11354) );
  OR2_X1 U14493 ( .A1(n11321), .A2(n11587), .ZN(n11353) );
  NAND2_X1 U14494 ( .A1(n11602), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14495 ( .A1(n11357), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14496 ( .A1(n11356), .A2(n11355), .ZN(n15503) );
  NAND2_X1 U14497 ( .A1(n11602), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14498 ( .A1(n11357), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14499 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10637), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14500 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14501 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14502 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11358) );
  NAND4_X1 U14503 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n11367) );
  AOI22_X1 U14504 ( .A1(n13886), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14505 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10855), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14506 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14507 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11362) );
  NAND4_X1 U14508 ( .A1(n11365), .A2(n11364), .A3(n11363), .A4(n11362), .ZN(
        n11366) );
  INV_X1 U14509 ( .A(n13519), .ZN(n19150) );
  OR2_X1 U14510 ( .A1(n11321), .A2(n19150), .ZN(n11368) );
  AOI22_X1 U14511 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14512 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14513 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14515 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11381) );
  AOI22_X1 U14516 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14517 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14518 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14519 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14520 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11380) );
  NOR2_X1 U14521 ( .A1(n11381), .A2(n11380), .ZN(n13521) );
  AOI22_X1 U14522 ( .A1(n11357), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11318), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U14523 ( .A1(n11602), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11384) );
  OAI211_X1 U14524 ( .C1(n11321), .C2(n13521), .A(n11385), .B(n11384), .ZN(
        n13796) );
  NAND2_X1 U14525 ( .A1(n11602), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14526 ( .A1(n11357), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14527 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10850), .B1(
        n10637), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14528 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14529 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11386) );
  NAND4_X1 U14531 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11395) );
  AOI22_X1 U14532 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n13912), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14533 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n13913), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14534 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n9625), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14535 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11390) );
  NAND4_X1 U14536 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11394) );
  OR2_X1 U14537 ( .A1(n11321), .A2(n19142), .ZN(n11396) );
  AOI22_X1 U14538 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14539 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14540 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14541 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U14542 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11408) );
  AOI22_X1 U14543 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14544 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14545 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14546 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14547 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  INV_X1 U14548 ( .A(n13826), .ZN(n11411) );
  NAND2_X1 U14549 ( .A1(n11602), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14550 ( .A1(n11357), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11409) );
  OAI211_X1 U14551 ( .C1(n11321), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        n15460) );
  AOI22_X1 U14552 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10650), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14553 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14554 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14555 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13907), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14556 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11421) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14558 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13886), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14559 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10855), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14560 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13912), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14561 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11420) );
  NOR2_X1 U14562 ( .A1(n11421), .A2(n11420), .ZN(n19138) );
  NAND2_X1 U14563 ( .A1(n11602), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14564 ( .A1(n11357), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11422) );
  OAI211_X1 U14565 ( .C1(n11321), .C2(n19138), .A(n11423), .B(n11422), .ZN(
        n14827) );
  AOI22_X1 U14566 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14567 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14568 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14569 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14570 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11433) );
  AOI22_X1 U14571 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14572 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14573 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14574 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11428) );
  NAND4_X1 U14575 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(
        n11432) );
  NOR2_X1 U14576 ( .A1(n11433), .A2(n11432), .ZN(n14909) );
  NAND2_X1 U14577 ( .A1(n11602), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14578 ( .A1(n11357), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11434) );
  OAI211_X1 U14579 ( .C1(n11321), .C2(n14909), .A(n11435), .B(n11434), .ZN(
        n15431) );
  AOI22_X1 U14580 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14581 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14582 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14583 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13907), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11436) );
  NAND4_X1 U14584 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n11445) );
  AOI22_X1 U14585 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9625), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14586 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13913), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14587 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13912), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14588 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11440) );
  NAND4_X1 U14589 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11444) );
  NOR2_X1 U14590 ( .A1(n11445), .A2(n11444), .ZN(n19133) );
  NAND2_X1 U14591 ( .A1(n11602), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14592 ( .A1(n11357), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11446) );
  OAI211_X1 U14593 ( .C1(n11321), .C2(n19133), .A(n11447), .B(n11446), .ZN(
        n15417) );
  INV_X1 U14594 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19827) );
  INV_X1 U14595 ( .A(n11321), .ZN(n11458) );
  AOI22_X1 U14596 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14597 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14598 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14599 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U14600 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11457) );
  AOI22_X1 U14601 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14602 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14603 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14604 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U14605 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11456) );
  NAND2_X1 U14606 ( .A1(n11458), .A2(n14903), .ZN(n11460) );
  AOI22_X1 U14607 ( .A1(n11317), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11459) );
  OAI211_X1 U14608 ( .C1(n11606), .C2(n19827), .A(n11460), .B(n11459), .ZN(
        n15398) );
  NAND2_X1 U14609 ( .A1(n11602), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14610 ( .A1(n11317), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11461) );
  INV_X1 U14611 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U14612 ( .A1(n11317), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11463) );
  OAI21_X1 U14613 ( .B1(n11606), .B2(n19830), .A(n11463), .ZN(n14987) );
  NAND2_X1 U14614 ( .A1(n11602), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14615 ( .A1(n11317), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11464) );
  NAND2_X1 U14616 ( .A1(n11465), .A2(n11464), .ZN(n15356) );
  NAND2_X1 U14617 ( .A1(n11602), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U14618 ( .A1(n11317), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11466) );
  AND2_X1 U14619 ( .A1(n11467), .A2(n11466), .ZN(n14978) );
  NAND2_X1 U14620 ( .A1(n11602), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14621 ( .A1(n11317), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U14622 ( .A1(n11602), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14623 ( .A1(n11357), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14624 ( .A1(n11602), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14625 ( .A1(n11317), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14626 ( .A1(n11473), .A2(n11472), .ZN(n14781) );
  NAND2_X1 U14627 ( .A1(n11602), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14628 ( .A1(n11317), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11474) );
  AND2_X1 U14629 ( .A1(n11475), .A2(n11474), .ZN(n14768) );
  NAND2_X1 U14630 ( .A1(n11602), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14631 ( .A1(n11317), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11476) );
  INV_X1 U14632 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U14633 ( .A1(n11357), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11478) );
  OAI21_X1 U14634 ( .B1(n11606), .B2(n19845), .A(n11478), .ZN(n14735) );
  NAND2_X1 U14635 ( .A1(n14734), .A2(n14735), .ZN(n14719) );
  NAND2_X1 U14636 ( .A1(n11602), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14637 ( .A1(n11357), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11479) );
  AND2_X1 U14638 ( .A1(n11480), .A2(n11479), .ZN(n14718) );
  NAND2_X1 U14639 ( .A1(n11602), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14640 ( .A1(n11357), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11481) );
  AND2_X1 U14641 ( .A1(n11482), .A2(n11481), .ZN(n11525) );
  INV_X1 U14642 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19851) );
  AOI22_X1 U14643 ( .A1(n11357), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11483) );
  OAI21_X1 U14644 ( .B1(n11606), .B2(n19851), .A(n11483), .ZN(n11485) );
  NOR2_X1 U14645 ( .A1(n11484), .A2(n11485), .ZN(n11486) );
  NAND2_X1 U14646 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15467) );
  INV_X1 U14647 ( .A(n15378), .ZN(n19270) );
  NOR2_X1 U14648 ( .A1(n19255), .A2(n19275), .ZN(n19271) );
  OAI211_X1 U14649 ( .C1(n19270), .C2(n19271), .A(n19269), .B(n15565), .ZN(
        n16342) );
  NOR2_X1 U14650 ( .A1(n11487), .A2(n16342), .ZN(n13794) );
  NAND2_X1 U14651 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n13794), .ZN(
        n15491) );
  NAND2_X1 U14652 ( .A1(n15445), .A2(n11488), .ZN(n15402) );
  NAND2_X1 U14653 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15364), .ZN(
        n11489) );
  NOR2_X1 U14654 ( .A1(n15293), .A2(n11491), .ZN(n11492) );
  NAND2_X1 U14655 ( .A1(n15306), .A2(n11492), .ZN(n15265) );
  OR2_X1 U14656 ( .A1(n15265), .A2(n11493), .ZN(n11524) );
  INV_X1 U14657 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11523) );
  NOR2_X1 U14658 ( .A1(n11524), .A2(n11523), .ZN(n15240) );
  NAND2_X1 U14659 ( .A1(n15240), .A2(n11576), .ZN(n15237) );
  OR2_X1 U14660 ( .A1(n19088), .A2(n19851), .ZN(n11510) );
  OAI211_X1 U14661 ( .C1(n16331), .C2(n14928), .A(n15237), .B(n11510), .ZN(
        n11495) );
  AOI21_X1 U14662 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15236), .A(
        n11495), .ZN(n11496) );
  OAI21_X1 U14663 ( .B1(n14848), .B2(n19257), .A(n11496), .ZN(n11497) );
  INV_X1 U14664 ( .A(n11497), .ZN(n11498) );
  OAI211_X1 U14665 ( .C1(n19264), .C2(n11515), .A(n11499), .B(n11498), .ZN(
        P2_U3018) );
  NAND2_X1 U14666 ( .A1(n15823), .A2(n19905), .ZN(n11500) );
  NAND2_X1 U14667 ( .A1(n11500), .A2(n16370), .ZN(n11501) );
  INV_X1 U14668 ( .A(n12941), .ZN(n11516) );
  INV_X1 U14669 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16384) );
  AOI21_X1 U14670 ( .B1(n19676), .B2(n16384), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n21037) );
  NOR2_X1 U14671 ( .A1(n19676), .A2(n16384), .ZN(n19897) );
  INV_X1 U14672 ( .A(n19897), .ZN(n13073) );
  NAND2_X1 U14673 ( .A1(n21037), .A2(n13073), .ZN(n11502) );
  NAND2_X1 U14674 ( .A1(n16384), .A2(n19678), .ZN(n19866) );
  INV_X1 U14675 ( .A(n19866), .ZN(n19779) );
  OR2_X1 U14676 ( .A1(n19869), .A2(n19779), .ZN(n19892) );
  NAND2_X1 U14677 ( .A1(n19892), .A2(n21039), .ZN(n11504) );
  INV_X1 U14678 ( .A(n13150), .ZN(n11506) );
  INV_X1 U14679 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19467) );
  NAND2_X1 U14680 ( .A1(n19467), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U14681 ( .A1(n11506), .A2(n11505), .ZN(n12993) );
  INV_X1 U14682 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18978) );
  INV_X1 U14683 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15059) );
  INV_X1 U14684 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15038) );
  INV_X1 U14685 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15026) );
  INV_X1 U14686 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14703) );
  NOR2_X1 U14687 ( .A1(n11539), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11508) );
  OR2_X1 U14688 ( .A1(n14645), .A2(n11508), .ZN(n14648) );
  NAND2_X1 U14689 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11509) );
  OAI211_X1 U14690 ( .C1(n16304), .C2(n14648), .A(n11510), .B(n11509), .ZN(
        n11511) );
  INV_X1 U14691 ( .A(n11511), .ZN(n11512) );
  NAND2_X1 U14692 ( .A1(n10072), .A2(n11512), .ZN(n11513) );
  AOI21_X1 U14693 ( .B1(n11514), .B2(n16293), .A(n11513), .ZN(n11520) );
  INV_X1 U14694 ( .A(n11515), .ZN(n11518) );
  NAND2_X1 U14695 ( .A1(n11520), .A2(n11519), .ZN(P2_U2986) );
  NOR2_X1 U14696 ( .A1(n11521), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11537) );
  XNOR2_X1 U14697 ( .A(n11522), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11544) );
  AND2_X1 U14698 ( .A1(n11524), .A2(n11523), .ZN(n11528) );
  AND2_X1 U14699 ( .A1(n9627), .A2(n11525), .ZN(n11526) );
  NOR2_X1 U14700 ( .A1(n11484), .A2(n11526), .ZN(n14706) );
  NAND2_X1 U14701 ( .A1(n14706), .A2(n19261), .ZN(n11527) );
  INV_X1 U14702 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19850) );
  OR2_X1 U14703 ( .A1(n11494), .A2(n19850), .ZN(n11540) );
  OAI211_X1 U14704 ( .C1(n11529), .C2(n11528), .A(n11527), .B(n11540), .ZN(
        n11533) );
  OR2_X1 U14705 ( .A1(n11530), .A2(n11531), .ZN(n11532) );
  OAI21_X1 U14706 ( .B1(n11544), .B2(n19259), .A(n11534), .ZN(n11535) );
  NAND2_X1 U14707 ( .A1(n9573), .A2(n11536), .ZN(P2_U3019) );
  AND2_X1 U14708 ( .A1(n14649), .A2(n14703), .ZN(n11538) );
  NOR2_X1 U14709 ( .A1(n11539), .A2(n11538), .ZN(n14702) );
  NAND2_X1 U14710 ( .A1(n16305), .A2(n14702), .ZN(n11541) );
  OAI211_X1 U14711 ( .C1(n16315), .C2(n14703), .A(n11541), .B(n11540), .ZN(
        n11542) );
  OAI21_X1 U14712 ( .B1(n11544), .B2(n16306), .A(n11543), .ZN(n11545) );
  NAND2_X1 U14713 ( .A1(n9659), .A2(n11546), .ZN(P2_U2987) );
  NAND2_X1 U14714 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14715 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11549) );
  INV_X1 U14716 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U14717 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14718 ( .A1(n9577), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11550) );
  OAI211_X1 U14719 ( .C1(n11258), .C2(n11552), .A(n11551), .B(n11550), .ZN(
        n11553) );
  AOI21_X1 U14720 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11553), .ZN(n14837) );
  INV_X1 U14721 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14722 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11555) );
  NAND2_X1 U14723 ( .A1(n9577), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11554) );
  OAI211_X1 U14724 ( .C1(n11258), .C2(n11556), .A(n11555), .B(n11554), .ZN(
        n11557) );
  AOI21_X1 U14725 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11557), .ZN(n11614) );
  INV_X1 U14726 ( .A(n11614), .ZN(n11558) );
  NAND2_X1 U14727 ( .A1(n14835), .A2(n11558), .ZN(n11566) );
  INV_X1 U14728 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14729 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14730 ( .A1(n9577), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11559) );
  OAI211_X1 U14731 ( .C1(n11258), .C2(n11561), .A(n11560), .B(n11559), .ZN(
        n11563) );
  AOI21_X1 U14732 ( .B1(n11564), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11563), .ZN(n11565) );
  NOR2_X1 U14733 ( .A1(n14130), .A2(n13376), .ZN(n11570) );
  INV_X1 U14734 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11567) );
  NAND2_X1 U14735 ( .A1(n19115), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U14736 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11568) );
  OAI211_X1 U14737 ( .C1(n16304), .C2(n13633), .A(n14124), .B(n11568), .ZN(
        n11569) );
  NOR2_X1 U14738 ( .A1(n11570), .A2(n11569), .ZN(n11601) );
  OAI21_X1 U14739 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n11575), .ZN(n11573) );
  NAND2_X1 U14740 ( .A1(n11574), .A2(n11573), .ZN(n11579) );
  INV_X1 U14741 ( .A(n11575), .ZN(n11577) );
  NAND2_X1 U14742 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  INV_X1 U14743 ( .A(n11580), .ZN(n11581) );
  NAND2_X1 U14744 ( .A1(n11593), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11583) );
  XNOR2_X1 U14745 ( .A(n11584), .B(n11583), .ZN(n11588) );
  INV_X1 U14746 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15239) );
  OAI21_X1 U14747 ( .B1(n11588), .B2(n11587), .A(n15239), .ZN(n15012) );
  NAND2_X1 U14748 ( .A1(n11593), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11585) );
  AOI21_X1 U14749 ( .B1(n11586), .B2(n11596), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11618) );
  INV_X1 U14750 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11613) );
  INV_X1 U14751 ( .A(n11588), .ZN(n16236) );
  NAND3_X1 U14752 ( .A1(n16236), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11596), .ZN(n15011) );
  NOR2_X1 U14753 ( .A1(n11590), .A2(n11589), .ZN(n11591) );
  NOR2_X1 U14754 ( .A1(n11592), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11594) );
  MUX2_X1 U14755 ( .A(n11595), .B(n11594), .S(n11593), .Z(n14676) );
  NAND2_X1 U14756 ( .A1(n14676), .A2(n11596), .ZN(n11597) );
  XOR2_X1 U14757 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11597), .Z(
        n11598) );
  OAI211_X1 U14758 ( .C1(n14132), .C2(n16308), .A(n11601), .B(n11600), .ZN(
        P2_U2983) );
  XNOR2_X1 U14759 ( .A(n15019), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15010) );
  AOI21_X1 U14760 ( .B1(n11610), .B2(n15565), .A(n15236), .ZN(n14127) );
  NAND2_X1 U14761 ( .A1(n11602), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14762 ( .A1(n11357), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11603) );
  AND2_X1 U14763 ( .A1(n11604), .A2(n11603), .ZN(n11608) );
  INV_X1 U14764 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19853) );
  AOI22_X1 U14765 ( .A1(n11357), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11605) );
  OAI21_X1 U14766 ( .B1(n11606), .B2(n19853), .A(n11605), .ZN(n14917) );
  AOI21_X1 U14767 ( .B1(n11608), .B2(n11607), .A(n14123), .ZN(n14686) );
  INV_X1 U14768 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11609) );
  NOR2_X1 U14769 ( .A1(n11494), .A2(n11609), .ZN(n15002) );
  NAND3_X1 U14770 ( .A1(n15240), .A2(n10048), .A3(n11613), .ZN(n11611) );
  OAI211_X1 U14771 ( .C1(n14127), .C2(n11613), .A(n11612), .B(n11611), .ZN(
        n11616) );
  NOR2_X1 U14772 ( .A1(n9575), .A2(n19257), .ZN(n11615) );
  NAND2_X1 U14773 ( .A1(n11617), .A2(n15011), .ZN(n11622) );
  INV_X1 U14774 ( .A(n11618), .ZN(n11620) );
  NAND2_X1 U14775 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  XNOR2_X1 U14776 ( .A(n11622), .B(n11621), .ZN(n15008) );
  NAND2_X1 U14777 ( .A1(n15008), .A2(n16338), .ZN(n11623) );
  AOI22_X1 U14778 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11627) );
  AND2_X2 U14779 ( .A1(n11625), .A2(n11634), .ZN(n12510) );
  AOI22_X1 U14780 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11626) );
  NAND2_X4 U14781 ( .A1(n13476), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11782) );
  INV_X1 U14782 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U14783 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11630) );
  NAND2_X1 U14784 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11629) );
  OAI211_X1 U14785 ( .C1(n11782), .C2(n11631), .A(n11630), .B(n11629), .ZN(
        n11632) );
  INV_X1 U14786 ( .A(n11632), .ZN(n11638) );
  AND2_X2 U14787 ( .A1(n11633), .A2(n11634), .ZN(n11789) );
  AOI22_X1 U14788 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14789 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11636) );
  AND2_X4 U14790 ( .A1(n13476), .A2(n15761), .ZN(n11792) );
  NAND2_X1 U14791 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11635) );
  INV_X1 U14792 ( .A(n11695), .ZN(n13392) );
  INV_X1 U14793 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U14794 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11640) );
  AOI22_X1 U14795 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14796 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11643) );
  NAND2_X1 U14797 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11642) );
  AOI22_X1 U14798 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11648) );
  INV_X2 U14799 ( .A(n12431), .ZN(n11714) );
  AOI22_X1 U14800 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14801 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11646) );
  INV_X1 U14802 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U14803 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11651) );
  NAND2_X1 U14804 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11650) );
  OAI211_X1 U14805 ( .C1(n11782), .C2(n11652), .A(n11651), .B(n11650), .ZN(
        n11653) );
  INV_X1 U14806 ( .A(n11653), .ZN(n11657) );
  AOI22_X1 U14807 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14808 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U14809 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11654) );
  AOI22_X1 U14810 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14811 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11659) );
  INV_X2 U14812 ( .A(n12482), .ZN(n12462) );
  AOI22_X1 U14813 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14814 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U14815 ( .A1(n11663), .A2(n20142), .ZN(n11681) );
  AOI22_X1 U14816 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14817 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14818 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14819 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14820 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14821 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11670) );
  OAI211_X1 U14822 ( .C1(n11782), .C2(n11672), .A(n11671), .B(n11670), .ZN(
        n11673) );
  INV_X1 U14823 ( .A(n11673), .ZN(n11677) );
  AOI22_X1 U14824 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14825 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U14826 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11674) );
  NAND2_X1 U14827 ( .A1(n11681), .A2(n11680), .ZN(n11711) );
  INV_X1 U14828 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U14829 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11683) );
  NAND2_X1 U14830 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11682) );
  OAI211_X1 U14831 ( .C1(n11782), .C2(n12433), .A(n11683), .B(n11682), .ZN(
        n11684) );
  INV_X1 U14832 ( .A(n11684), .ZN(n11688) );
  AOI22_X1 U14833 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14834 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11686) );
  NAND2_X1 U14835 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11685) );
  NAND4_X1 U14836 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11694) );
  AOI22_X1 U14837 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14838 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14839 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14840 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14841 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11693) );
  OR2_X2 U14842 ( .A1(n11694), .A2(n11693), .ZN(n20130) );
  INV_X1 U14843 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11698) );
  NAND2_X1 U14844 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11697) );
  NAND2_X1 U14845 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11696) );
  OAI211_X1 U14846 ( .C1(n11782), .C2(n11698), .A(n11697), .B(n11696), .ZN(
        n11699) );
  INV_X1 U14847 ( .A(n11699), .ZN(n11703) );
  AOI22_X1 U14848 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14849 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11701) );
  NAND2_X1 U14850 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11700) );
  NAND4_X1 U14851 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11709) );
  AOI22_X1 U14852 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14853 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14854 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12545), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14855 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11704) );
  NAND4_X1 U14856 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11708) );
  AND3_X2 U14857 ( .A1(n11711), .A2(n11772), .A3(n11710), .ZN(n13214) );
  AOI22_X1 U14858 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14859 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14860 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9613), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14861 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11665), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11715) );
  INV_X1 U14862 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U14863 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11720) );
  NAND2_X1 U14864 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11719) );
  OAI211_X1 U14865 ( .C1(n11782), .C2(n11721), .A(n11720), .B(n11719), .ZN(
        n11722) );
  INV_X1 U14866 ( .A(n11722), .ZN(n11726) );
  AOI22_X1 U14867 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14868 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11724) );
  NAND2_X1 U14869 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11723) );
  NAND2_X4 U14870 ( .A1(n9650), .A2(n10080), .ZN(n20109) );
  NOR2_X1 U14871 ( .A1(n12835), .A2(n20109), .ZN(n11727) );
  NAND2_X1 U14872 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U14873 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11730) );
  NAND2_X1 U14874 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U14875 ( .A1(n12545), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11728) );
  NAND4_X1 U14876 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n11734) );
  NOR2_X2 U14877 ( .A1(n11734), .A2(n11733), .ZN(n11750) );
  NAND2_X1 U14878 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11738) );
  NAND2_X1 U14879 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U14880 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11736) );
  NAND2_X1 U14881 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11735) );
  NAND2_X1 U14882 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14883 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14884 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U14885 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11739) );
  INV_X1 U14886 ( .A(n11743), .ZN(n11783) );
  NAND2_X1 U14887 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14888 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11744) );
  OAI211_X1 U14889 ( .C1(n11782), .C2(n12386), .A(n11745), .B(n11744), .ZN(
        n11746) );
  INV_X1 U14890 ( .A(n11746), .ZN(n11747) );
  NAND4_X4 U14891 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11757) );
  INV_X2 U14892 ( .A(n11757), .ZN(n13410) );
  NAND2_X1 U14893 ( .A1(n12854), .A2(n13204), .ZN(n13105) );
  NAND2_X1 U14894 ( .A1(n11913), .A2(n20148), .ZN(n11752) );
  NOR2_X2 U14895 ( .A1(n13105), .A2(n11752), .ZN(n12889) );
  NAND2_X1 U14896 ( .A1(n12889), .A2(n13221), .ZN(n11753) );
  AND2_X2 U14897 ( .A1(n12889), .A2(n20109), .ZN(n13411) );
  INV_X1 U14898 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11754) );
  XNOR2_X1 U14899 ( .A(n11754), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12722) );
  NAND3_X1 U14900 ( .A1(n13599), .A2(n13474), .A3(n12585), .ZN(n13215) );
  AOI21_X1 U14901 ( .B1(n13411), .B2(n12722), .A(n13413), .ZN(n11755) );
  NAND2_X1 U14902 ( .A1(n13401), .A2(n11755), .ZN(n11756) );
  INV_X1 U14903 ( .A(n12835), .ZN(n13203) );
  AND2_X2 U14904 ( .A1(n20130), .A2(n11757), .ZN(n12858) );
  NAND2_X1 U14905 ( .A1(n13203), .A2(n12858), .ZN(n11760) );
  NAND2_X1 U14906 ( .A1(n11773), .A2(n20134), .ZN(n11759) );
  NAND2_X1 U14907 ( .A1(n13209), .A2(n11757), .ZN(n13613) );
  NAND2_X1 U14908 ( .A1(n20126), .A2(n20109), .ZN(n11758) );
  NAND4_X1 U14909 ( .A1(n11760), .A2(n11759), .A3(n13613), .A4(n11758), .ZN(
        n11762) );
  NOR2_X1 U14910 ( .A1(n13214), .A2(n20109), .ZN(n11761) );
  NOR2_X2 U14911 ( .A1(n11762), .A2(n11761), .ZN(n11780) );
  NAND2_X1 U14912 ( .A1(n13424), .A2(n13412), .ZN(n11766) );
  NAND2_X1 U14913 ( .A1(n12585), .A2(n20142), .ZN(n11765) );
  AND2_X1 U14914 ( .A1(n20134), .A2(n20148), .ZN(n11767) );
  AOI21_X1 U14915 ( .B1(n13211), .B2(n14623), .A(n13474), .ZN(n11768) );
  NAND2_X1 U14916 ( .A1(n11780), .A2(n11768), .ZN(n12853) );
  NAND2_X1 U14917 ( .A1(n12853), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14918 ( .A1(n11865), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11771) );
  NAND2_X1 U14919 ( .A1(n16214), .A2(n20777), .ZN(n12836) );
  MUX2_X1 U14920 ( .A(n12836), .B(n15781), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11770) );
  NAND2_X1 U14921 ( .A1(n11771), .A2(n11770), .ZN(n11857) );
  INV_X1 U14922 ( .A(n11772), .ZN(n11775) );
  INV_X1 U14923 ( .A(n13599), .ZN(n13102) );
  NAND2_X1 U14924 ( .A1(n13102), .A2(n12624), .ZN(n12997) );
  OAI22_X1 U14925 ( .A1(n11775), .A2(n12997), .B1(n11774), .B2(n13208), .ZN(
        n11777) );
  NAND2_X1 U14926 ( .A1(n13474), .A2(n11913), .ZN(n13405) );
  NAND3_X1 U14927 ( .A1(n13405), .A2(n16214), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11776) );
  NOR2_X1 U14928 ( .A1(n11777), .A2(n11776), .ZN(n11779) );
  NAND3_X1 U14929 ( .A1(n13211), .A2(n11757), .A3(n14623), .ZN(n11778) );
  NAND3_X1 U14930 ( .A1(n11780), .A2(n11779), .A3(n11778), .ZN(n11856) );
  INV_X1 U14931 ( .A(n11856), .ZN(n11781) );
  INV_X1 U14932 ( .A(n11782), .ZN(n11954) );
  INV_X1 U14933 ( .A(n11954), .ZN(n11807) );
  INV_X1 U14934 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11786) );
  INV_X2 U14935 ( .A(n11783), .ZN(n12539) );
  NAND2_X1 U14936 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U14937 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11784) );
  OAI211_X1 U14938 ( .C1(n11807), .C2(n11786), .A(n11785), .B(n11784), .ZN(
        n11787) );
  INV_X1 U14939 ( .A(n11787), .ZN(n11797) );
  AOI22_X1 U14940 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11796) );
  INV_X1 U14941 ( .A(n11790), .ZN(n11791) );
  INV_X2 U14942 ( .A(n11791), .ZN(n11930) );
  AOI22_X1 U14943 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11795) );
  NAND2_X1 U14944 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11794) );
  NAND4_X1 U14945 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11803) );
  AOI22_X1 U14946 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14947 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14948 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14949 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11798) );
  NAND4_X1 U14950 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11802) );
  INV_X1 U14951 ( .A(n12750), .ZN(n11820) );
  INV_X1 U14952 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U14953 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U14954 ( .A1(n9580), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11804) );
  OAI211_X1 U14955 ( .C1(n11807), .C2(n11806), .A(n11805), .B(n11804), .ZN(
        n11808) );
  INV_X1 U14956 ( .A(n11808), .ZN(n11813) );
  AOI22_X1 U14957 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14958 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14959 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11810) );
  NAND4_X1 U14960 ( .A1(n11813), .A2(n11812), .A3(n11811), .A4(n11810), .ZN(
        n11819) );
  AOI22_X1 U14961 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U14962 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14963 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14964 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11814) );
  NAND4_X1 U14965 ( .A1(n11817), .A2(n11816), .A3(n11815), .A4(n11814), .ZN(
        n11818) );
  XNOR2_X1 U14966 ( .A(n11820), .B(n12810), .ZN(n11821) );
  NAND2_X1 U14967 ( .A1(n11860), .A2(n11821), .ZN(n11822) );
  INV_X1 U14968 ( .A(n12810), .ZN(n11825) );
  NAND2_X1 U14969 ( .A1(n12609), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11824) );
  AOI21_X1 U14970 ( .B1(n13209), .B2(n12750), .A(n20777), .ZN(n11823) );
  OAI211_X1 U14971 ( .C1(n11825), .C2(n20134), .A(n11824), .B(n11823), .ZN(
        n11911) );
  NAND2_X1 U14972 ( .A1(n11860), .A2(n12810), .ZN(n11826) );
  INV_X1 U14973 ( .A(n11929), .ZN(n11845) );
  INV_X1 U14974 ( .A(n11954), .ZN(n12354) );
  INV_X1 U14975 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U14976 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U14977 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11829) );
  OAI211_X1 U14978 ( .C1(n12354), .C2(n11831), .A(n11830), .B(n11829), .ZN(
        n11832) );
  INV_X1 U14979 ( .A(n11832), .ZN(n11837) );
  AOI22_X1 U14980 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14981 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U14982 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11834) );
  NAND4_X1 U14983 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11844) );
  AOI22_X1 U14984 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11809), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14985 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U14986 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14987 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11839) );
  NAND4_X1 U14988 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11843) );
  NAND2_X1 U14989 ( .A1(n11845), .A2(n12751), .ZN(n11847) );
  NAND2_X1 U14990 ( .A1(n12609), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11846) );
  OAI211_X1 U14991 ( .C1(n12804), .C2(n12810), .A(n11847), .B(n11846), .ZN(
        n11848) );
  NAND2_X1 U14992 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  NAND2_X1 U14993 ( .A1(n11865), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11853) );
  NAND2_X1 U14994 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11869) );
  OAI21_X1 U14995 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11869), .ZN(n20481) );
  OR2_X1 U14996 ( .A1(n15781), .A2(n20476), .ZN(n11863) );
  OAI21_X1 U14997 ( .B1(n12836), .B2(n20481), .A(n11863), .ZN(n11851) );
  INV_X1 U14998 ( .A(n11851), .ZN(n11852) );
  NAND2_X1 U14999 ( .A1(n11853), .A2(n11852), .ZN(n11855) );
  XNOR2_X2 U15000 ( .A(n11855), .B(n11854), .ZN(n20231) );
  INV_X1 U15001 ( .A(n20231), .ZN(n11858) );
  NAND2_X1 U15002 ( .A1(n11860), .A2(n12751), .ZN(n11861) );
  INV_X1 U15003 ( .A(n11897), .ZN(n11896) );
  AND2_X1 U15004 ( .A1(n11863), .A2(n9998), .ZN(n11864) );
  NOR2_X1 U15005 ( .A1(n15781), .A2(n20560), .ZN(n11867) );
  INV_X1 U15006 ( .A(n12836), .ZN(n11871) );
  INV_X1 U15007 ( .A(n11869), .ZN(n11868) );
  NAND2_X1 U15008 ( .A1(n11868), .A2(n20560), .ZN(n20228) );
  NAND2_X1 U15009 ( .A1(n11869), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U15010 ( .A1(n20228), .A2(n11870), .ZN(n20117) );
  NAND2_X1 U15011 ( .A1(n11871), .A2(n20117), .ZN(n11873) );
  NAND2_X1 U15012 ( .A1(n11875), .A2(n11873), .ZN(n11872) );
  NAND4_X1 U15013 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11877) );
  NAND2_X1 U15014 ( .A1(n13491), .A2(n11877), .ZN(n13458) );
  INV_X1 U15015 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U15016 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11879) );
  NAND2_X1 U15017 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11878) );
  OAI211_X1 U15018 ( .C1(n12354), .C2(n11880), .A(n11879), .B(n11878), .ZN(
        n11881) );
  INV_X1 U15019 ( .A(n11881), .ZN(n11885) );
  AOI22_X1 U15020 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15021 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U15022 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11882) );
  NAND4_X1 U15023 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        n11891) );
  AOI22_X1 U15024 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U15025 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U15026 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U15027 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11886) );
  NAND4_X1 U15028 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11890) );
  NAND2_X1 U15029 ( .A1(n12609), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11892) );
  OAI21_X1 U15030 ( .B1(n12752), .B2(n11929), .A(n11892), .ZN(n11893) );
  XNOR2_X1 U15031 ( .A(n11894), .B(n11893), .ZN(n11898) );
  INV_X1 U15032 ( .A(n11898), .ZN(n11895) );
  NAND2_X1 U15033 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  INV_X1 U15034 ( .A(n13387), .ZN(n12907) );
  NAND2_X1 U15035 ( .A1(n12907), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11973) );
  INV_X1 U15036 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14269) );
  XNOR2_X1 U15037 ( .A(n14269), .B(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19988) );
  NAND2_X1 U15038 ( .A1(n20856), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12098) );
  OAI21_X1 U15039 ( .B1(n19988), .B2(n12559), .A(n12098), .ZN(n11900) );
  AOI21_X1 U15040 ( .B1(n12561), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11900), .ZN(
        n11901) );
  OAI21_X1 U15041 ( .B1(n11902), .B2(n11973), .A(n11901), .ZN(n11903) );
  INV_X1 U15042 ( .A(n11903), .ZN(n11904) );
  NAND2_X1 U15043 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11924) );
  INV_X1 U15044 ( .A(n13357), .ZN(n11923) );
  NAND2_X1 U15045 ( .A1(n13503), .A2(n12192), .ZN(n11910) );
  INV_X1 U15046 ( .A(n11973), .ZN(n11906) );
  NAND2_X1 U15047 ( .A1(n11906), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11908) );
  INV_X2 U15048 ( .A(n9702), .ZN(n12561) );
  AOI22_X1 U15049 ( .A1(n12561), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20856), .ZN(n11907) );
  AND2_X1 U15050 ( .A1(n11908), .A2(n11907), .ZN(n11909) );
  NAND2_X1 U15051 ( .A1(n12741), .A2(n11913), .ZN(n11914) );
  NAND2_X1 U15052 ( .A1(n11914), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13169) );
  NAND2_X1 U15053 ( .A1(n12561), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U15054 ( .A1(n20856), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11917) );
  OAI211_X1 U15055 ( .C1(n11973), .C2(n15761), .A(n11918), .B(n11917), .ZN(
        n11919) );
  AOI21_X1 U15056 ( .B1(n11916), .B2(n12192), .A(n11919), .ZN(n11920) );
  OR2_X1 U15057 ( .A1(n13169), .A2(n11920), .ZN(n13170) );
  INV_X1 U15058 ( .A(n11920), .ZN(n13171) );
  OR2_X1 U15059 ( .A1(n13171), .A2(n12559), .ZN(n11921) );
  NAND2_X1 U15060 ( .A1(n13170), .A2(n11921), .ZN(n13200) );
  NAND2_X1 U15061 ( .A1(n13201), .A2(n13200), .ZN(n13356) );
  NAND2_X1 U15062 ( .A1(n11923), .A2(n11922), .ZN(n13354) );
  NAND2_X1 U15063 ( .A1(n11866), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15064 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10079), .ZN(
        n20408) );
  NAND2_X1 U15065 ( .A1(n20559), .A2(n20408), .ZN(n11925) );
  NOR3_X1 U15066 ( .A1(n20559), .A2(n20560), .A3(n20476), .ZN(n20717) );
  NAND2_X1 U15067 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20717), .ZN(
        n20766) );
  NAND2_X1 U15068 ( .A1(n11925), .A2(n20766), .ZN(n20418) );
  OAI22_X1 U15069 ( .A1(n12836), .A2(n20418), .B1(n15781), .B2(n20559), .ZN(
        n11926) );
  INV_X1 U15070 ( .A(n11926), .ZN(n11927) );
  INV_X1 U15071 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U15072 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U15073 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11931) );
  OAI211_X1 U15074 ( .C1(n12354), .C2(n11933), .A(n11932), .B(n11931), .ZN(
        n11934) );
  INV_X1 U15075 ( .A(n11934), .ZN(n11938) );
  AOI22_X1 U15076 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9585), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15077 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11936) );
  NAND2_X1 U15078 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11935) );
  NAND4_X1 U15079 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11944) );
  AOI22_X1 U15080 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15081 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15082 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15083 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11939) );
  NAND4_X1 U15084 ( .A1(n11942), .A2(n11941), .A3(n11940), .A4(n11939), .ZN(
        n11943) );
  AOI22_X1 U15085 ( .A1(n12583), .A2(n12766), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12609), .ZN(n11945) );
  INV_X1 U15086 ( .A(n13576), .ZN(n13577) );
  NAND2_X1 U15087 ( .A1(n11946), .A2(n13577), .ZN(n11947) );
  INV_X2 U15088 ( .A(n12559), .ZN(n12616) );
  OAI21_X1 U15089 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11949), .A(
        n12002), .ZN(n13618) );
  AOI22_X1 U15090 ( .A1(n12616), .A2(n13618), .B1(n12560), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U15091 ( .A1(n12561), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11950) );
  OAI211_X1 U15092 ( .C1(n11973), .C2(n11948), .A(n11951), .B(n11950), .ZN(
        n11952) );
  INV_X1 U15093 ( .A(n11952), .ZN(n11953) );
  NAND2_X1 U15094 ( .A1(n13511), .A2(n13510), .ZN(n13509) );
  INV_X1 U15095 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U15096 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11956) );
  NAND2_X1 U15097 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11955) );
  OAI211_X1 U15098 ( .C1(n12354), .C2(n11957), .A(n11956), .B(n11955), .ZN(
        n11958) );
  INV_X1 U15099 ( .A(n11958), .ZN(n11962) );
  AOI22_X1 U15100 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9585), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15101 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U15102 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11959) );
  NAND4_X1 U15103 ( .A1(n11962), .A2(n11961), .A3(n11960), .A4(n11959), .ZN(
        n11968) );
  AOI22_X1 U15104 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15105 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15106 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15107 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12511), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11963) );
  NAND4_X1 U15108 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n11967) );
  NAND2_X1 U15109 ( .A1(n12583), .A2(n12777), .ZN(n11970) );
  NAND2_X1 U15110 ( .A1(n12609), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U15111 ( .A1(n11970), .A2(n11969), .ZN(n11978) );
  XNOR2_X1 U15112 ( .A(n11979), .B(n11978), .ZN(n12765) );
  NAND2_X1 U15113 ( .A1(n20856), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U15114 ( .A1(n12561), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11971) );
  OAI211_X1 U15115 ( .C1(n11973), .C2(n16217), .A(n11972), .B(n11971), .ZN(
        n11974) );
  NAND2_X1 U15116 ( .A1(n11974), .A2(n12559), .ZN(n11976) );
  XNOR2_X1 U15117 ( .A(n12002), .B(n14254), .ZN(n14251) );
  NAND2_X1 U15118 ( .A1(n14251), .A2(n12616), .ZN(n11975) );
  NAND2_X1 U15119 ( .A1(n11976), .A2(n11975), .ZN(n11977) );
  AOI21_X1 U15120 ( .B1(n12765), .B2(n12192), .A(n11977), .ZN(n13535) );
  INV_X1 U15121 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U15122 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U15123 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11980) );
  OAI211_X1 U15124 ( .C1(n12354), .C2(n11982), .A(n11981), .B(n11980), .ZN(
        n11983) );
  INV_X1 U15125 ( .A(n11983), .ZN(n11987) );
  AOI22_X1 U15126 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15127 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U15128 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11984) );
  NAND4_X1 U15129 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11993) );
  AOI22_X1 U15130 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15131 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15132 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15133 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11988) );
  NAND4_X1 U15134 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11992) );
  NAND2_X1 U15135 ( .A1(n12583), .A2(n12785), .ZN(n11995) );
  NAND2_X1 U15136 ( .A1(n12609), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11994) );
  NAND2_X1 U15137 ( .A1(n11995), .A2(n11994), .ZN(n11996) );
  OR2_X1 U15138 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  NAND2_X1 U15139 ( .A1(n12028), .A2(n11998), .ZN(n12776) );
  INV_X1 U15140 ( .A(n12776), .ZN(n11999) );
  NAND2_X1 U15141 ( .A1(n11999), .A2(n12192), .ZN(n12008) );
  INV_X1 U15142 ( .A(n12002), .ZN(n12000) );
  AOI21_X1 U15143 ( .B1(n12000), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U15144 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12001) );
  OR2_X1 U15145 ( .A1(n12003), .A2(n12023), .ZN(n16026) );
  NAND2_X1 U15146 ( .A1(n16026), .A2(n12616), .ZN(n12005) );
  NAND2_X1 U15147 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U15148 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  AOI21_X1 U15149 ( .B1(n12561), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12006), .ZN(
        n12007) );
  INV_X1 U15150 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12027) );
  INV_X1 U15151 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U15152 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U15153 ( .A1(n9580), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12009) );
  OAI211_X1 U15154 ( .C1(n12354), .C2(n12011), .A(n12010), .B(n12009), .ZN(
        n12012) );
  INV_X1 U15155 ( .A(n12012), .ZN(n12016) );
  AOI22_X1 U15156 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15157 ( .A1(n11714), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U15158 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12013) );
  NAND4_X1 U15159 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12022) );
  AOI22_X1 U15160 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15161 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15162 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15163 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12017) );
  NAND4_X1 U15164 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n12021) );
  AOI22_X1 U15165 ( .A1(n12583), .A2(n12796), .B1(n12609), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12029) );
  NAND2_X1 U15166 ( .A1(n12028), .A2(n12029), .ZN(n12784) );
  NAND2_X1 U15167 ( .A1(n12784), .A2(n12192), .ZN(n12026) );
  NOR2_X1 U15168 ( .A1(n12023), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12024) );
  OR2_X1 U15169 ( .A1(n12035), .A2(n12024), .ZN(n19975) );
  AOI22_X1 U15170 ( .A1(n19975), .A2(n12616), .B1(n12560), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U15171 ( .C1(n9702), .C2(n12027), .A(n12026), .B(n12025), .ZN(
        n13609) );
  NAND2_X1 U15172 ( .A1(n12583), .A2(n12810), .ZN(n12033) );
  NAND2_X1 U15173 ( .A1(n12609), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12032) );
  NAND2_X1 U15174 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  INV_X1 U15175 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13665) );
  OR2_X1 U15176 ( .A1(n12035), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12036) );
  NAND2_X1 U15177 ( .A1(n12036), .A2(n12059), .ZN(n19967) );
  AOI22_X1 U15178 ( .A1(n19967), .A2(n12616), .B1(n12560), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12037) );
  OAI21_X1 U15179 ( .B1(n9702), .B2(n13665), .A(n12037), .ZN(n12038) );
  AOI21_X1 U15180 ( .B1(n12795), .B2(n12192), .A(n12038), .ZN(n13663) );
  INV_X1 U15181 ( .A(n13663), .ZN(n12039) );
  NAND2_X1 U15182 ( .A1(n12040), .A2(n12039), .ZN(n13662) );
  AOI22_X1 U15183 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15184 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15185 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15186 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12041) );
  NAND4_X1 U15187 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12054) );
  INV_X1 U15188 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U15189 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12046) );
  NAND2_X1 U15190 ( .A1(n9580), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12045) );
  OAI211_X1 U15191 ( .C1(n12354), .C2(n12047), .A(n12046), .B(n12045), .ZN(
        n12048) );
  INV_X1 U15192 ( .A(n12048), .ZN(n12052) );
  AOI22_X1 U15193 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15194 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U15195 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12049) );
  NAND4_X1 U15196 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12053) );
  OAI21_X1 U15197 ( .B1(n12054), .B2(n12053), .A(n12192), .ZN(n12058) );
  NAND2_X1 U15198 ( .A1(n12561), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12057) );
  XNOR2_X1 U15199 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12059), .ZN(
        n19958) );
  OAI22_X1 U15200 ( .A1(n19958), .A2(n12559), .B1(n12098), .B2(n19948), .ZN(
        n12055) );
  INV_X1 U15201 ( .A(n12055), .ZN(n12056) );
  XOR2_X1 U15202 ( .A(n19941), .B(n12090), .Z(n19939) );
  INV_X1 U15203 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U15204 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U15205 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12060) );
  OAI211_X1 U15206 ( .C1(n12354), .C2(n12387), .A(n12061), .B(n12060), .ZN(
        n12062) );
  INV_X1 U15207 ( .A(n12062), .ZN(n12066) );
  AOI22_X1 U15208 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15209 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U15210 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12063) );
  NAND4_X1 U15211 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12072) );
  AOI22_X1 U15212 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11809), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15213 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15214 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15215 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15216 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12071) );
  OR2_X1 U15217 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  AOI22_X1 U15218 ( .A1(n12192), .A2(n12073), .B1(n12560), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12075) );
  NAND2_X1 U15219 ( .A1(n12561), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12074) );
  OAI211_X1 U15220 ( .C1(n19939), .C2(n12559), .A(n12075), .B(n12074), .ZN(
        n13743) );
  INV_X1 U15221 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U15222 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12077) );
  NAND2_X1 U15223 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12076) );
  OAI211_X1 U15224 ( .C1(n12354), .C2(n12078), .A(n12077), .B(n12076), .ZN(
        n12079) );
  INV_X1 U15225 ( .A(n12079), .ZN(n12083) );
  AOI22_X1 U15226 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15227 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U15228 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12080) );
  NAND4_X1 U15229 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12089) );
  AOI22_X1 U15230 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15231 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15232 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15233 ( .A1(n11714), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12084) );
  NAND4_X1 U15234 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12088) );
  NOR2_X1 U15235 ( .A1(n12089), .A2(n12088), .ZN(n12094) );
  XNOR2_X1 U15236 ( .A(n12095), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15934) );
  NAND2_X1 U15237 ( .A1(n15934), .A2(n12616), .ZN(n12092) );
  AOI22_X1 U15238 ( .A1(n12561), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12560), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12091) );
  OAI211_X1 U15239 ( .C1(n12094), .C2(n12093), .A(n12092), .B(n12091), .ZN(
        n13760) );
  INV_X1 U15240 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12099) );
  OAI21_X1 U15241 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12096), .A(
        n12150), .ZN(n16011) );
  NAND2_X1 U15242 ( .A1(n16011), .A2(n12616), .ZN(n12097) );
  OAI21_X1 U15243 ( .B1(n12099), .B2(n12098), .A(n12097), .ZN(n12100) );
  AOI21_X1 U15244 ( .B1(n12561), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12100), .ZN(
        n14236) );
  NAND2_X1 U15245 ( .A1(n9581), .A2(n12101), .ZN(n14235) );
  INV_X1 U15246 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U15247 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U15248 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12102) );
  OAI211_X1 U15249 ( .C1(n12354), .C2(n12104), .A(n12103), .B(n12102), .ZN(
        n12105) );
  INV_X1 U15250 ( .A(n12105), .ZN(n12109) );
  AOI22_X1 U15251 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11809), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15252 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U15253 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12106) );
  NAND4_X1 U15254 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12115) );
  AOI22_X1 U15255 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15256 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15257 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15258 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12110) );
  NAND4_X1 U15259 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12114) );
  OR2_X1 U15260 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  NAND2_X1 U15261 ( .A1(n12192), .A2(n12116), .ZN(n14360) );
  NAND2_X1 U15262 ( .A1(n9581), .A2(n12117), .ZN(n12118) );
  NAND2_X1 U15263 ( .A1(n14235), .A2(n12118), .ZN(n12156) );
  XOR2_X1 U15264 ( .A(n14247), .B(n12157), .Z(n14513) );
  INV_X1 U15265 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12121) );
  NAND2_X1 U15266 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12120) );
  NAND2_X1 U15267 ( .A1(n9580), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12119) );
  OAI211_X1 U15268 ( .C1(n12354), .C2(n12121), .A(n12120), .B(n12119), .ZN(
        n12122) );
  INV_X1 U15269 ( .A(n12122), .ZN(n12126) );
  AOI22_X1 U15270 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15271 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U15272 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12123) );
  NAND4_X1 U15273 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12132) );
  AOI22_X1 U15274 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15275 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15276 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15277 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12127) );
  NAND4_X1 U15278 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12131) );
  OR2_X1 U15279 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  AOI22_X1 U15280 ( .A1(n12192), .A2(n12133), .B1(n12560), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U15281 ( .A1(n12561), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12134) );
  OAI211_X1 U15282 ( .C1(n14513), .C2(n12559), .A(n12135), .B(n12134), .ZN(
        n14240) );
  AOI22_X1 U15283 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9585), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15284 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15285 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15286 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U15287 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12149) );
  INV_X1 U15288 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U15289 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12141) );
  NAND2_X1 U15290 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12140) );
  OAI211_X1 U15291 ( .C1(n12354), .C2(n12142), .A(n12141), .B(n12140), .ZN(
        n12143) );
  INV_X1 U15292 ( .A(n12143), .ZN(n12147) );
  AOI22_X1 U15293 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11809), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15294 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U15295 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12144) );
  NAND4_X1 U15296 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12148) );
  OAI21_X1 U15297 ( .B1(n12149), .B2(n12148), .A(n12192), .ZN(n12154) );
  NAND2_X1 U15298 ( .A1(n12561), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12153) );
  XOR2_X1 U15299 ( .A(n15914), .B(n12150), .Z(n16001) );
  INV_X1 U15300 ( .A(n16001), .ZN(n12151) );
  AOI22_X1 U15301 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12616), .B2(n12151), .ZN(n12152) );
  NAND3_X1 U15302 ( .A1(n12154), .A2(n12153), .A3(n12152), .ZN(n14353) );
  NAND2_X1 U15303 ( .A1(n12156), .A2(n12155), .ZN(n14238) );
  INV_X1 U15304 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12158) );
  XNOR2_X1 U15305 ( .A(n12179), .B(n12158), .ZN(n15911) );
  OR2_X1 U15306 ( .A1(n15911), .A2(n12559), .ZN(n12177) );
  AOI22_X1 U15307 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15308 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11809), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15309 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15310 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12159) );
  NAND4_X1 U15311 ( .A1(n12162), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12172) );
  INV_X1 U15312 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U15313 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12164) );
  NAND2_X1 U15314 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12163) );
  OAI211_X1 U15315 ( .C1(n12354), .C2(n12165), .A(n12164), .B(n12163), .ZN(
        n12166) );
  INV_X1 U15316 ( .A(n12166), .ZN(n12170) );
  AOI22_X1 U15317 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15318 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U15319 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12167) );
  NAND4_X1 U15320 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  OAI21_X1 U15321 ( .B1(n12172), .B2(n12171), .A(n12192), .ZN(n12175) );
  NAND2_X1 U15322 ( .A1(n12561), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12174) );
  NAND2_X1 U15323 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12173) );
  AND3_X1 U15324 ( .A1(n12175), .A2(n12174), .A3(n12173), .ZN(n12176) );
  XOR2_X1 U15325 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12199), .Z(
        n15897) );
  INV_X1 U15326 ( .A(n15897), .ZN(n15994) );
  AOI22_X1 U15327 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15328 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15329 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15330 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12180) );
  NAND4_X1 U15331 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n12194) );
  INV_X1 U15332 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U15333 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12185) );
  NAND2_X1 U15334 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12184) );
  OAI211_X1 U15335 ( .C1(n12354), .C2(n12186), .A(n12185), .B(n12184), .ZN(
        n12187) );
  INV_X1 U15336 ( .A(n12187), .ZN(n12191) );
  AOI22_X1 U15337 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15338 ( .A1(n11714), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12189) );
  NAND2_X1 U15339 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12188) );
  NAND4_X1 U15340 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12193) );
  OAI21_X1 U15341 ( .B1(n12194), .B2(n12193), .A(n12192), .ZN(n12197) );
  NAND2_X1 U15342 ( .A1(n12561), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U15343 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12195) );
  NAND3_X1 U15344 ( .A1(n12197), .A2(n12196), .A3(n12195), .ZN(n12198) );
  AOI21_X1 U15345 ( .B1(n15994), .B2(n12616), .A(n12198), .ZN(n14337) );
  AOI21_X1 U15346 ( .B1(n12200), .B2(n20915), .A(n12257), .ZN(n14495) );
  AOI21_X1 U15347 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20915), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12201) );
  AOI21_X1 U15348 ( .B1(n12561), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12201), .ZN(
        n12217) );
  AOI22_X1 U15349 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15350 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15351 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15352 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U15353 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12215) );
  INV_X1 U15354 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12208) );
  NAND2_X1 U15355 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12207) );
  NAND2_X1 U15356 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12206) );
  OAI211_X1 U15357 ( .C1(n12354), .C2(n12208), .A(n12207), .B(n12206), .ZN(
        n12209) );
  INV_X1 U15358 ( .A(n12209), .ZN(n12213) );
  AOI22_X1 U15359 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15360 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U15361 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12210) );
  NAND4_X1 U15362 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12214) );
  OAI21_X1 U15363 ( .B1(n12215), .B2(n12214), .A(n12520), .ZN(n12216) );
  AOI22_X1 U15364 ( .A1(n14495), .A2(n12616), .B1(n12217), .B2(n12216), .ZN(
        n14223) );
  INV_X1 U15365 ( .A(n14222), .ZN(n12238) );
  INV_X1 U15366 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12220) );
  NAND2_X1 U15367 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12219) );
  NAND2_X1 U15368 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12218) );
  OAI211_X1 U15369 ( .C1(n12354), .C2(n12220), .A(n12219), .B(n12218), .ZN(
        n12221) );
  INV_X1 U15370 ( .A(n12221), .ZN(n12225) );
  AOI22_X1 U15371 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15372 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U15373 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12222) );
  NAND4_X1 U15374 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12231) );
  AOI22_X1 U15375 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15376 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15377 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15378 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12226) );
  NAND4_X1 U15379 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12230) );
  OR2_X1 U15380 ( .A1(n12231), .A2(n12230), .ZN(n12236) );
  INV_X1 U15381 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12234) );
  XOR2_X1 U15382 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12257), .Z(
        n15982) );
  INV_X1 U15383 ( .A(n15982), .ZN(n12232) );
  AOI22_X1 U15384 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12616), .B2(n12232), .ZN(n12233) );
  OAI21_X1 U15385 ( .B1(n9702), .B2(n12234), .A(n12233), .ZN(n12235) );
  AOI21_X1 U15386 ( .B1(n12520), .B2(n12236), .A(n12235), .ZN(n14330) );
  NAND2_X1 U15387 ( .A1(n12238), .A2(n12237), .ZN(n14321) );
  INV_X1 U15388 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U15389 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12240) );
  NAND2_X1 U15390 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12239) );
  OAI211_X1 U15391 ( .C1(n12354), .C2(n12241), .A(n12240), .B(n12239), .ZN(
        n12242) );
  INV_X1 U15392 ( .A(n12242), .ZN(n12247) );
  AOI22_X1 U15393 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15394 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U15395 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12244) );
  NAND4_X1 U15396 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12253) );
  AOI22_X1 U15397 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15398 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15399 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15400 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12248) );
  NAND4_X1 U15401 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12252) );
  NOR2_X1 U15402 ( .A1(n12253), .A2(n12252), .ZN(n12256) );
  OAI21_X1 U15403 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n12277), .A(n12559), 
        .ZN(n12254) );
  AOI21_X1 U15404 ( .B1(n12561), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12254), .ZN(
        n12255) );
  OAI21_X1 U15405 ( .B1(n12556), .B2(n12256), .A(n12255), .ZN(n12259) );
  XNOR2_X1 U15406 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B(n12278), .ZN(
        n15886) );
  NAND2_X1 U15407 ( .A1(n15886), .A2(n12616), .ZN(n12258) );
  NAND2_X1 U15408 ( .A1(n12259), .A2(n12258), .ZN(n14322) );
  NOR2_X2 U15409 ( .A1(n14321), .A2(n14322), .ZN(n14314) );
  AOI22_X1 U15410 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15411 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15412 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15413 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12260) );
  NAND4_X1 U15414 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12273) );
  INV_X1 U15415 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12266) );
  NAND2_X1 U15416 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12265) );
  NAND2_X1 U15417 ( .A1(n9580), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12264) );
  OAI211_X1 U15418 ( .C1(n12354), .C2(n12266), .A(n12265), .B(n12264), .ZN(
        n12267) );
  INV_X1 U15419 ( .A(n12267), .ZN(n12271) );
  AOI22_X1 U15420 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15421 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12269) );
  NAND2_X1 U15422 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12268) );
  NAND4_X1 U15423 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12272) );
  NOR2_X1 U15424 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  OR2_X1 U15425 ( .A1(n12556), .A2(n12274), .ZN(n12282) );
  NAND2_X1 U15426 ( .A1(n20856), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12275) );
  NAND2_X1 U15427 ( .A1(n12559), .A2(n12275), .ZN(n12276) );
  AOI21_X1 U15428 ( .B1(n12561), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12276), .ZN(
        n12281) );
  OAI21_X1 U15429 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12279), .A(
        n12320), .ZN(n15981) );
  NOR2_X1 U15430 ( .A1(n15981), .A2(n12559), .ZN(n12280) );
  AOI21_X1 U15431 ( .B1(n12282), .B2(n12281), .A(n12280), .ZN(n14315) );
  INV_X1 U15432 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U15433 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12284) );
  NAND2_X1 U15434 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12283) );
  OAI211_X1 U15435 ( .C1(n11807), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        n12286) );
  INV_X1 U15436 ( .A(n12286), .ZN(n12290) );
  AOI22_X1 U15437 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11809), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15438 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12243), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U15439 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12287) );
  NAND4_X1 U15440 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12296) );
  AOI22_X1 U15441 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15442 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12511), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15443 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15444 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9585), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12291) );
  NAND4_X1 U15445 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12295) );
  NOR2_X1 U15446 ( .A1(n12296), .A2(n12295), .ZN(n12299) );
  OAI21_X1 U15447 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15867), .A(n12559), 
        .ZN(n12297) );
  AOI21_X1 U15448 ( .B1(n12561), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12297), .ZN(
        n12298) );
  OAI21_X1 U15449 ( .B1(n12556), .B2(n12299), .A(n12298), .ZN(n12301) );
  XNOR2_X1 U15450 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12320), .ZN(
        n15970) );
  NAND2_X1 U15451 ( .A1(n12616), .A2(n15970), .ZN(n12300) );
  NAND2_X1 U15452 ( .A1(n12301), .A2(n12300), .ZN(n14311) );
  AOI22_X1 U15453 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15454 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15455 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15456 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15457 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12315) );
  INV_X1 U15458 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n20888) );
  NAND2_X1 U15459 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12308) );
  NAND2_X1 U15460 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12307) );
  OAI211_X1 U15461 ( .C1(n11807), .C2(n20888), .A(n12308), .B(n12307), .ZN(
        n12309) );
  INV_X1 U15462 ( .A(n12309), .ZN(n12313) );
  AOI22_X1 U15463 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15464 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U15465 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12310) );
  NAND4_X1 U15466 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12314) );
  NOR2_X1 U15467 ( .A1(n12315), .A2(n12314), .ZN(n12319) );
  OAI21_X1 U15468 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20857), .A(
        n20856), .ZN(n12316) );
  INV_X1 U15469 ( .A(n12316), .ZN(n12317) );
  AOI21_X1 U15470 ( .B1(n12561), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12317), .ZN(
        n12318) );
  OAI21_X1 U15471 ( .B1(n12556), .B2(n12319), .A(n12318), .ZN(n12323) );
  OAI21_X1 U15472 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12321), .A(
        n12376), .ZN(n15961) );
  OR2_X1 U15473 ( .A1(n12559), .A2(n15961), .ZN(n12322) );
  NAND2_X1 U15474 ( .A1(n12323), .A2(n12322), .ZN(n14304) );
  NOR2_X1 U15475 ( .A1(n14311), .A2(n14304), .ZN(n12324) );
  INV_X1 U15476 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U15477 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12326) );
  NAND2_X1 U15478 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12325) );
  OAI211_X1 U15479 ( .C1(n12354), .C2(n12327), .A(n12326), .B(n12325), .ZN(
        n12328) );
  INV_X1 U15480 ( .A(n12328), .ZN(n12332) );
  AOI22_X1 U15481 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11809), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15482 ( .A1(n12462), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U15483 ( .A1(n11792), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12329) );
  NAND4_X1 U15484 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12338) );
  AOI22_X1 U15485 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15486 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15487 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9580), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15488 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12333) );
  NAND4_X1 U15489 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12337) );
  NOR2_X1 U15490 ( .A1(n12338), .A2(n12337), .ZN(n12341) );
  INV_X1 U15491 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15840) );
  AOI21_X1 U15492 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15840), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12339) );
  AOI21_X1 U15493 ( .B1(n12561), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12339), .ZN(
        n12340) );
  OAI21_X1 U15494 ( .B1(n12556), .B2(n12341), .A(n12340), .ZN(n12343) );
  XNOR2_X1 U15495 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12376), .ZN(
        n15844) );
  NAND2_X1 U15496 ( .A1(n15844), .A2(n12616), .ZN(n12342) );
  NAND2_X1 U15497 ( .A1(n12343), .A2(n12342), .ZN(n14294) );
  INV_X1 U15498 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12345) );
  INV_X1 U15499 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12344) );
  OAI22_X1 U15500 ( .A1(n9588), .A2(n12345), .B1(n11791), .B2(n12344), .ZN(
        n12349) );
  INV_X1 U15501 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12347) );
  INV_X1 U15502 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12346) );
  OAI22_X1 U15503 ( .A1(n12536), .A2(n12347), .B1(n12534), .B2(n12346), .ZN(
        n12348) );
  AOI211_X1 U15504 ( .C1(n11793), .C2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n12349), .B(n12348), .ZN(n12358) );
  AOI22_X1 U15505 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15506 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15507 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15508 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12350) );
  AND4_X1 U15509 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12357) );
  AOI22_X1 U15510 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U15511 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12355) );
  NAND4_X1 U15512 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12382) );
  INV_X1 U15513 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12360) );
  INV_X1 U15514 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12359) );
  OAI22_X1 U15515 ( .A1(n9588), .A2(n12360), .B1(n11791), .B2(n12359), .ZN(
        n12364) );
  INV_X1 U15516 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12362) );
  INV_X1 U15517 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12361) );
  OAI22_X1 U15518 ( .A1(n12536), .A2(n12362), .B1(n12534), .B2(n12361), .ZN(
        n12363) );
  AOI211_X1 U15519 ( .C1(n11792), .C2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n12364), .B(n12363), .ZN(n12372) );
  AOI22_X1 U15520 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15521 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15522 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15523 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12365) );
  AND4_X1 U15524 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12371) );
  AOI22_X1 U15525 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U15526 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12369) );
  NAND4_X1 U15527 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12383) );
  XOR2_X1 U15528 ( .A(n12382), .B(n12383), .Z(n12373) );
  NAND2_X1 U15529 ( .A1(n12373), .A2(n12520), .ZN(n12380) );
  INV_X1 U15530 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12374) );
  AOI21_X1 U15531 ( .B1(n12374), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12375) );
  AOI21_X1 U15532 ( .B1(n12561), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12375), .ZN(
        n12379) );
  OAI21_X1 U15533 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12377), .A(
        n12381), .ZN(n15959) );
  INV_X1 U15534 ( .A(n15959), .ZN(n12378) );
  AOI22_X1 U15535 ( .A1(n12380), .A2(n12379), .B1(n12616), .B2(n12378), .ZN(
        n14291) );
  XNOR2_X1 U15536 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12422), .ZN(
        n14469) );
  INV_X1 U15537 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15538 ( .A1(n12383), .A2(n12382), .ZN(n12418) );
  INV_X1 U15539 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12392) );
  INV_X1 U15540 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12385) );
  INV_X1 U15541 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12384) );
  OAI22_X1 U15542 ( .A1(n12536), .A2(n12385), .B1(n12534), .B2(n12384), .ZN(
        n12389) );
  OAI22_X1 U15543 ( .A1(n11713), .A2(n12387), .B1(n9579), .B2(n12386), .ZN(
        n12388) );
  AOI211_X1 U15544 ( .C1(n11792), .C2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12389), .B(n12388), .ZN(n12391) );
  AOI22_X1 U15545 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12390) );
  OAI211_X1 U15546 ( .C1(n12354), .C2(n12392), .A(n12391), .B(n12390), .ZN(
        n12398) );
  AOI22_X1 U15547 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15548 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15549 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15550 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12393) );
  NAND4_X1 U15551 ( .A1(n12396), .A2(n12395), .A3(n12394), .A4(n12393), .ZN(
        n12397) );
  NOR2_X1 U15552 ( .A1(n12398), .A2(n12397), .ZN(n12419) );
  XOR2_X1 U15553 ( .A(n12418), .B(n12419), .Z(n12399) );
  NAND2_X1 U15554 ( .A1(n12399), .A2(n12520), .ZN(n12401) );
  AOI21_X1 U15555 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20856), .A(
        n12616), .ZN(n12400) );
  OAI211_X1 U15556 ( .C1(n9702), .C2(n12402), .A(n12401), .B(n12400), .ZN(
        n12403) );
  OAI21_X1 U15557 ( .B1(n14469), .B2(n12559), .A(n12403), .ZN(n14209) );
  NOR2_X2 U15558 ( .A1(n14208), .A2(n14209), .ZN(n14194) );
  INV_X1 U15559 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15560 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12405) );
  NAND2_X1 U15561 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12404) );
  OAI211_X1 U15562 ( .C1(n11807), .C2(n12406), .A(n12405), .B(n12404), .ZN(
        n12407) );
  INV_X1 U15563 ( .A(n12407), .ZN(n12411) );
  AOI22_X1 U15564 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15565 ( .A1(n11809), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U15566 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12408) );
  NAND4_X1 U15567 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12417) );
  AOI22_X1 U15568 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15569 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15570 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15571 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15572 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12416) );
  OR2_X1 U15573 ( .A1(n12417), .A2(n12416), .ZN(n12428) );
  NOR2_X1 U15574 ( .A1(n12419), .A2(n12418), .ZN(n12429) );
  XOR2_X1 U15575 ( .A(n12428), .B(n12429), .Z(n12420) );
  NAND2_X1 U15576 ( .A1(n12420), .A2(n12520), .ZN(n12427) );
  INV_X1 U15577 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14459) );
  NOR2_X1 U15578 ( .A1(n14459), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12421) );
  AOI211_X1 U15579 ( .C1(n12561), .C2(P1_EAX_REG_25__SCAN_IN), .A(n12616), .B(
        n12421), .ZN(n12426) );
  INV_X1 U15580 ( .A(n12423), .ZN(n12424) );
  NAND2_X1 U15581 ( .A1(n12424), .A2(n14459), .ZN(n12425) );
  AND2_X1 U15582 ( .A1(n12471), .A2(n12425), .ZN(n14463) );
  AOI22_X1 U15583 ( .A1(n12427), .A2(n12426), .B1(n12616), .B2(n14463), .ZN(
        n14196) );
  NAND2_X1 U15584 ( .A1(n14194), .A2(n14196), .ZN(n14183) );
  XOR2_X1 U15585 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n12471), .Z(
        n14450) );
  INV_X1 U15586 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U15587 ( .A1(n12429), .A2(n12428), .ZN(n12452) );
  INV_X1 U15588 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12440) );
  INV_X1 U15589 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12432) );
  INV_X1 U15590 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12430) );
  OAI22_X1 U15591 ( .A1(n9588), .A2(n12432), .B1(n12431), .B2(n12430), .ZN(
        n12437) );
  INV_X1 U15592 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12434) );
  OAI22_X1 U15593 ( .A1(n12435), .A2(n12434), .B1(n9579), .B2(n12433), .ZN(
        n12436) );
  AOI211_X1 U15594 ( .C1(n11792), .C2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12437), .B(n12436), .ZN(n12439) );
  AOI22_X1 U15595 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12438) );
  OAI211_X1 U15596 ( .C1(n12354), .C2(n12440), .A(n12439), .B(n12438), .ZN(
        n12446) );
  AOI22_X1 U15597 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15598 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15599 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15600 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12441) );
  NAND4_X1 U15601 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n12445) );
  NOR2_X1 U15602 ( .A1(n12446), .A2(n12445), .ZN(n12453) );
  XOR2_X1 U15603 ( .A(n12452), .B(n12453), .Z(n12447) );
  NAND2_X1 U15604 ( .A1(n12447), .A2(n12520), .ZN(n12449) );
  AOI21_X1 U15605 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20856), .A(
        n12616), .ZN(n12448) );
  OAI211_X1 U15606 ( .C1(n9702), .C2(n12450), .A(n12449), .B(n12448), .ZN(
        n12451) );
  OAI21_X1 U15607 ( .B1(n12559), .B2(n14450), .A(n12451), .ZN(n14185) );
  NOR2_X1 U15608 ( .A1(n12453), .A2(n12452), .ZN(n12478) );
  INV_X1 U15609 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12456) );
  NAND2_X1 U15610 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12455) );
  NAND2_X1 U15611 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12454) );
  OAI211_X1 U15612 ( .C1(n11807), .C2(n12456), .A(n12455), .B(n12454), .ZN(
        n12457) );
  INV_X1 U15613 ( .A(n12457), .ZN(n12461) );
  AOI22_X1 U15614 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9585), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15615 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12459) );
  NAND2_X1 U15616 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12458) );
  NAND4_X1 U15617 ( .A1(n12461), .A2(n12460), .A3(n12459), .A4(n12458), .ZN(
        n12468) );
  AOI22_X1 U15618 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12543), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15619 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12465) );
  INV_X1 U15620 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n20988) );
  AOI22_X1 U15621 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15622 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12511), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12463) );
  NAND4_X1 U15623 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12467) );
  OR2_X1 U15624 ( .A1(n12468), .A2(n12467), .ZN(n12477) );
  XOR2_X1 U15625 ( .A(n12478), .B(n12477), .Z(n12469) );
  NAND2_X1 U15626 ( .A1(n12469), .A2(n12520), .ZN(n12476) );
  INV_X1 U15627 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14439) );
  NOR2_X1 U15628 ( .A1(n14439), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12470) );
  AOI211_X1 U15629 ( .C1(n12561), .C2(P1_EAX_REG_27__SCAN_IN), .A(n12616), .B(
        n12470), .ZN(n12475) );
  INV_X1 U15630 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14186) );
  INV_X1 U15631 ( .A(n12472), .ZN(n12473) );
  NAND2_X1 U15632 ( .A1(n12473), .A2(n14439), .ZN(n12474) );
  AOI22_X1 U15633 ( .A1(n12476), .A2(n12475), .B1(n12616), .B2(n14443), .ZN(
        n14168) );
  NAND2_X1 U15634 ( .A1(n14167), .A2(n14168), .ZN(n14152) );
  INV_X1 U15635 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14158) );
  XNOR2_X1 U15636 ( .A(n12524), .B(n14158), .ZN(n14429) );
  INV_X1 U15637 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12500) );
  NAND2_X1 U15638 ( .A1(n12478), .A2(n12477), .ZN(n12502) );
  INV_X1 U15639 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12490) );
  INV_X1 U15640 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12479) );
  OAI22_X1 U15641 ( .A1(n9579), .A2(n12481), .B1(n12480), .B2(n12479), .ZN(
        n12486) );
  INV_X1 U15642 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12484) );
  INV_X1 U15643 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12483) );
  OAI22_X1 U15644 ( .A1(n12536), .A2(n12484), .B1(n9588), .B2(n12483), .ZN(
        n12485) );
  AOI211_X1 U15645 ( .C1(n11792), .C2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12486), .B(n12485), .ZN(n12489) );
  AOI22_X1 U15646 ( .A1(n12539), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12488) );
  OAI211_X1 U15647 ( .C1(n11807), .C2(n12490), .A(n12489), .B(n12488), .ZN(
        n12496) );
  AOI22_X1 U15648 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15649 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15650 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15651 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U15652 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12495) );
  NOR2_X1 U15653 ( .A1(n12496), .A2(n12495), .ZN(n12503) );
  XOR2_X1 U15654 ( .A(n12502), .B(n12503), .Z(n12497) );
  NAND2_X1 U15655 ( .A1(n12497), .A2(n12520), .ZN(n12499) );
  AOI21_X1 U15656 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20856), .A(
        n12616), .ZN(n12498) );
  OAI211_X1 U15657 ( .C1(n9702), .C2(n12500), .A(n12499), .B(n12498), .ZN(
        n12501) );
  OAI21_X1 U15658 ( .B1(n12559), .B2(n14429), .A(n12501), .ZN(n14153) );
  NOR2_X1 U15659 ( .A1(n12503), .A2(n12502), .ZN(n12522) );
  INV_X1 U15660 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12505) );
  INV_X1 U15661 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12504) );
  OAI22_X1 U15662 ( .A1(n9588), .A2(n12505), .B1(n11791), .B2(n12504), .ZN(
        n12509) );
  INV_X1 U15663 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12507) );
  INV_X1 U15664 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12506) );
  OAI22_X1 U15665 ( .A1(n12536), .A2(n12507), .B1(n12534), .B2(n12506), .ZN(
        n12508) );
  AOI211_X1 U15666 ( .C1(n11793), .C2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12509), .B(n12508), .ZN(n12519) );
  AOI22_X1 U15667 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15668 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15669 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15670 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12512) );
  AND4_X1 U15671 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12518) );
  AOI22_X1 U15672 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U15673 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12516) );
  NAND4_X1 U15674 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12521) );
  NAND2_X1 U15675 ( .A1(n12522), .A2(n12521), .ZN(n12553) );
  OAI211_X1 U15676 ( .C1(n12522), .C2(n12521), .A(n12553), .B(n12520), .ZN(
        n12530) );
  INV_X1 U15677 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12841) );
  NOR2_X1 U15678 ( .A1(n12841), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12523) );
  AOI211_X1 U15679 ( .C1(n12561), .C2(P1_EAX_REG_29__SCAN_IN), .A(n12616), .B(
        n12523), .ZN(n12529) );
  INV_X1 U15680 ( .A(n12524), .ZN(n12525) );
  INV_X1 U15681 ( .A(n12526), .ZN(n12527) );
  NAND2_X1 U15682 ( .A1(n12527), .A2(n12841), .ZN(n12528) );
  AOI22_X1 U15683 ( .A1(n12530), .A2(n12529), .B1(n12616), .B2(n14145), .ZN(
        n12844) );
  XOR2_X1 U15684 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12619), .Z(
        n14417) );
  INV_X1 U15685 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12542) );
  INV_X1 U15686 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12532) );
  INV_X1 U15687 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12531) );
  OAI22_X1 U15688 ( .A1(n9588), .A2(n12532), .B1(n11791), .B2(n12531), .ZN(
        n12538) );
  INV_X1 U15689 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12535) );
  INV_X1 U15690 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12533) );
  OAI22_X1 U15691 ( .A1(n12536), .A2(n12535), .B1(n12534), .B2(n12533), .ZN(
        n12537) );
  AOI211_X1 U15692 ( .C1(n11792), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12538), .B(n12537), .ZN(n12541) );
  AOI22_X1 U15693 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12539), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12540) );
  OAI211_X1 U15694 ( .C1(n11807), .C2(n12542), .A(n12541), .B(n12540), .ZN(
        n12551) );
  AOI22_X1 U15695 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12462), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15696 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15697 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11714), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15698 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9580), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12546) );
  NAND4_X1 U15699 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12550) );
  NOR2_X1 U15700 ( .A1(n12551), .A2(n12550), .ZN(n12552) );
  XNOR2_X1 U15701 ( .A(n12553), .B(n12552), .ZN(n12557) );
  NAND2_X1 U15702 ( .A1(n12561), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12555) );
  OAI21_X1 U15703 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n20856), .ZN(n12554) );
  OAI211_X1 U15704 ( .C1(n12557), .C2(n12556), .A(n12555), .B(n12554), .ZN(
        n12558) );
  OAI21_X1 U15705 ( .B1(n14417), .B2(n12559), .A(n12558), .ZN(n12851) );
  AOI22_X1 U15706 ( .A1(n12561), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12560), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12562) );
  XNOR2_X1 U15707 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12576) );
  NAND2_X1 U15708 ( .A1(n20601), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U15709 ( .A1(n12576), .A2(n12577), .ZN(n12565) );
  NAND2_X1 U15710 ( .A1(n20476), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12564) );
  NAND2_X1 U15711 ( .A1(n12565), .A2(n12564), .ZN(n12579) );
  XNOR2_X1 U15712 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12578) );
  NAND2_X1 U15713 ( .A1(n12579), .A2(n12578), .ZN(n12567) );
  NAND2_X1 U15714 ( .A1(n20560), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12566) );
  NAND2_X1 U15715 ( .A1(n12567), .A2(n12566), .ZN(n12575) );
  XNOR2_X1 U15716 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15717 ( .A1(n12575), .A2(n12574), .ZN(n12569) );
  NAND2_X1 U15718 ( .A1(n20559), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12568) );
  NOR2_X1 U15719 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16217), .ZN(
        n12570) );
  XNOR2_X1 U15720 ( .A(n12575), .B(n12574), .ZN(n12605) );
  XNOR2_X1 U15721 ( .A(n12577), .B(n12576), .ZN(n12592) );
  XNOR2_X1 U15722 ( .A(n12579), .B(n12578), .ZN(n12599) );
  NOR4_X1 U15723 ( .A1(n12608), .A2(n12605), .A3(n12592), .A4(n12599), .ZN(
        n12580) );
  NOR2_X1 U15724 ( .A1(n12581), .A2(n12580), .ZN(n13110) );
  AND2_X1 U15725 ( .A1(n12563), .A2(n13110), .ZN(n13100) );
  NAND2_X1 U15726 ( .A1(n13100), .A2(n13399), .ZN(n12957) );
  NAND2_X1 U15727 ( .A1(n12606), .A2(n12581), .ZN(n12615) );
  NAND2_X1 U15728 ( .A1(n12581), .A2(n12583), .ZN(n12613) );
  INV_X1 U15729 ( .A(n12609), .ZN(n12604) );
  NOR2_X1 U15730 ( .A1(n12592), .A2(n12582), .ZN(n12591) );
  OAI21_X1 U15731 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20601), .A(
        n12584), .ZN(n12587) );
  NOR2_X1 U15732 ( .A1(n12601), .A2(n12587), .ZN(n12590) );
  NAND2_X1 U15733 ( .A1(n12585), .A2(n20109), .ZN(n12586) );
  NAND2_X1 U15734 ( .A1(n12586), .A2(n13410), .ZN(n12600) );
  INV_X1 U15735 ( .A(n12587), .ZN(n12588) );
  OAI211_X1 U15736 ( .C1(n13209), .C2(n12835), .A(n12600), .B(n12588), .ZN(
        n12589) );
  OAI21_X1 U15737 ( .B1(n12606), .B2(n12590), .A(n12589), .ZN(n12593) );
  NAND2_X1 U15738 ( .A1(n12591), .A2(n12593), .ZN(n12598) );
  NAND2_X1 U15739 ( .A1(n12594), .A2(n11757), .ZN(n12611) );
  OAI211_X1 U15740 ( .C1(n12594), .C2(n12593), .A(n12592), .B(n12611), .ZN(
        n12597) );
  NAND2_X1 U15741 ( .A1(n12609), .A2(n12599), .ZN(n12595) );
  OAI211_X1 U15742 ( .C1(n12601), .C2(n12599), .A(n12595), .B(n12600), .ZN(
        n12596) );
  NAND3_X1 U15743 ( .A1(n12598), .A2(n12597), .A3(n12596), .ZN(n12603) );
  INV_X1 U15744 ( .A(n12608), .ZN(n12607) );
  NAND2_X1 U15745 ( .A1(n12609), .A2(n12608), .ZN(n12610) );
  NAND2_X1 U15746 ( .A1(n12613), .A2(n12612), .ZN(n12614) );
  NOR2_X1 U15747 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16227) );
  NAND2_X1 U15748 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16227), .ZN(n16224) );
  OR2_X2 U15749 ( .A1(n12836), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20101) );
  NOR2_X1 U15750 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20776), .ZN(n20859) );
  NAND2_X1 U15751 ( .A1(n12616), .A2(n20859), .ZN(n12617) );
  OAI211_X1 U15752 ( .C1(n16224), .C2(n20777), .A(n20101), .B(n12617), .ZN(
        n12618) );
  INV_X1 U15753 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14133) );
  INV_X1 U15754 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12620) );
  NOR2_X1 U15755 ( .A1(n13601), .A2(n20776), .ZN(n12622) );
  NAND2_X1 U15756 ( .A1(n12896), .A2(n12623), .ZN(n12735) );
  INV_X1 U15757 ( .A(n20130), .ZN(n12625) );
  NAND2_X1 U15758 ( .A1(n12625), .A2(n20109), .ZN(n12642) );
  AOI22_X1 U15759 ( .A1(n12712), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13101), .ZN(n12719) );
  AOI22_X1 U15760 ( .A1(n12712), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13101), .ZN(n12859) );
  AND2_X2 U15761 ( .A1(n13221), .A2(n12858), .ZN(n12706) );
  INV_X1 U15762 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12627) );
  NAND2_X1 U15763 ( .A1(n12706), .A2(n12627), .ZN(n12631) );
  INV_X1 U15764 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12626) );
  NAND2_X1 U15765 ( .A1(n12642), .A2(n12626), .ZN(n12629) );
  NAND2_X1 U15766 ( .A1(n13221), .A2(n12627), .ZN(n12628) );
  NAND3_X1 U15767 ( .A1(n12624), .A2(n12629), .A3(n12628), .ZN(n12630) );
  NAND2_X1 U15768 ( .A1(n12631), .A2(n12630), .ZN(n12633) );
  NAND2_X1 U15769 ( .A1(n12642), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12632) );
  OAI21_X1 U15770 ( .B1(n12858), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12632), .ZN(
        n13167) );
  XNOR2_X1 U15771 ( .A(n12633), .B(n13167), .ZN(n14266) );
  INV_X1 U15772 ( .A(n12633), .ZN(n12634) );
  AOI21_X1 U15773 ( .B1(n14266), .B2(n13221), .A(n12634), .ZN(n13359) );
  INV_X1 U15774 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U15775 ( .A1(n12706), .A2(n12635), .ZN(n12639) );
  INV_X1 U15776 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U15777 ( .A1(n12642), .A2(n13420), .ZN(n12637) );
  NAND2_X1 U15778 ( .A1(n13221), .A2(n12635), .ZN(n12636) );
  NAND3_X1 U15779 ( .A1(n12624), .A2(n12637), .A3(n12636), .ZN(n12638) );
  NAND2_X1 U15780 ( .A1(n12639), .A2(n12638), .ZN(n13358) );
  INV_X1 U15781 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13541) );
  NAND2_X1 U15782 ( .A1(n13205), .A2(n13541), .ZN(n12641) );
  MUX2_X1 U15783 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12640) );
  AND2_X1 U15784 ( .A1(n12641), .A2(n12640), .ZN(n13512) );
  NAND2_X1 U15785 ( .A1(n13513), .A2(n13512), .ZN(n13533) );
  MUX2_X1 U15786 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12646) );
  INV_X1 U15787 ( .A(n12642), .ZN(n12643) );
  NAND2_X1 U15788 ( .A1(n13101), .A2(n12643), .ZN(n12690) );
  NAND2_X1 U15789 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13101), .ZN(
        n12644) );
  AND2_X1 U15790 ( .A1(n12690), .A2(n12644), .ZN(n12645) );
  AND2_X1 U15791 ( .A1(n12646), .A2(n12645), .ZN(n13532) );
  INV_X1 U15792 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16205) );
  INV_X1 U15793 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15794 ( .A1(n13221), .A2(n12647), .ZN(n12648) );
  OAI211_X1 U15795 ( .C1(n12858), .C2(n16205), .A(n12648), .B(n12642), .ZN(
        n12649) );
  OAI21_X1 U15796 ( .B1(n12711), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12649), .ZN(
        n13571) );
  MUX2_X1 U15797 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12652) );
  NAND2_X1 U15798 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13101), .ZN(
        n12650) );
  AND2_X1 U15799 ( .A1(n12690), .A2(n12650), .ZN(n12651) );
  NAND2_X1 U15800 ( .A1(n12652), .A2(n12651), .ZN(n16186) );
  INV_X1 U15801 ( .A(n12711), .ZN(n12653) );
  INV_X1 U15802 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20013) );
  NAND2_X1 U15803 ( .A1(n12653), .A2(n20013), .ZN(n12656) );
  INV_X1 U15804 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16194) );
  NAND2_X1 U15805 ( .A1(n13221), .A2(n20013), .ZN(n12654) );
  OAI211_X1 U15806 ( .C1(n12858), .C2(n16194), .A(n12654), .B(n12642), .ZN(
        n12655) );
  AND2_X1 U15807 ( .A1(n12656), .A2(n12655), .ZN(n16185) );
  NAND2_X1 U15808 ( .A1(n16186), .A2(n16185), .ZN(n12657) );
  MUX2_X1 U15809 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12660) );
  NAND2_X1 U15810 ( .A1(n13101), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12658) );
  AND2_X1 U15811 ( .A1(n12690), .A2(n12658), .ZN(n12659) );
  NAND2_X1 U15812 ( .A1(n12660), .A2(n12659), .ZN(n13700) );
  INV_X1 U15813 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16170) );
  INV_X1 U15814 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20009) );
  NAND2_X1 U15815 ( .A1(n13221), .A2(n20009), .ZN(n12661) );
  OAI211_X1 U15816 ( .C1(n12858), .C2(n16170), .A(n12661), .B(n12642), .ZN(
        n12662) );
  OAI21_X1 U15817 ( .B1(n12711), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12662), .ZN(
        n16163) );
  INV_X1 U15818 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U15819 ( .A1(n12706), .A2(n13764), .ZN(n12666) );
  INV_X1 U15820 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U15821 ( .A1(n12642), .A2(n12823), .ZN(n12664) );
  NAND2_X1 U15822 ( .A1(n13221), .A2(n13764), .ZN(n12663) );
  NAND3_X1 U15823 ( .A1(n12624), .A2(n12664), .A3(n12663), .ZN(n12665) );
  INV_X1 U15824 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16147) );
  NAND2_X1 U15825 ( .A1(n13205), .A2(n16147), .ZN(n12668) );
  MUX2_X1 U15826 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12667) );
  MUX2_X1 U15827 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12671) );
  NAND2_X1 U15828 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13101), .ZN(
        n12669) );
  AND2_X1 U15829 ( .A1(n12690), .A2(n12669), .ZN(n12670) );
  NAND2_X1 U15830 ( .A1(n12671), .A2(n12670), .ZN(n14350) );
  MUX2_X1 U15831 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12672) );
  NAND2_X1 U15832 ( .A1(n12672), .A2(n10077), .ZN(n14245) );
  MUX2_X1 U15833 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12675) );
  NAND2_X1 U15834 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n13101), .ZN(
        n12673) );
  AND2_X1 U15835 ( .A1(n12690), .A2(n12673), .ZN(n12674) );
  INV_X1 U15836 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16115) );
  NAND2_X1 U15837 ( .A1(n13205), .A2(n16115), .ZN(n12677) );
  MUX2_X1 U15838 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12676) );
  AND2_X1 U15839 ( .A1(n12677), .A2(n12676), .ZN(n14339) );
  MUX2_X1 U15840 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12680) );
  NAND2_X1 U15841 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n13101), .ZN(
        n12678) );
  AND2_X1 U15842 ( .A1(n12690), .A2(n12678), .ZN(n12679) );
  MUX2_X1 U15843 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12682) );
  INV_X1 U15844 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U15845 ( .A1(n13205), .A2(n14595), .ZN(n12681) );
  NAND2_X1 U15846 ( .A1(n12682), .A2(n12681), .ZN(n14331) );
  INV_X1 U15847 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15884) );
  NAND2_X1 U15848 ( .A1(n12706), .A2(n15884), .ZN(n12686) );
  INV_X1 U15849 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16101) );
  NAND2_X1 U15850 ( .A1(n12642), .A2(n16101), .ZN(n12684) );
  NAND2_X1 U15851 ( .A1(n13221), .A2(n15884), .ZN(n12683) );
  NAND3_X1 U15852 ( .A1(n12624), .A2(n12684), .A3(n12683), .ZN(n12685) );
  NAND2_X1 U15853 ( .A1(n12686), .A2(n12685), .ZN(n14324) );
  MUX2_X1 U15854 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12688) );
  INV_X1 U15855 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U15856 ( .A1(n13205), .A2(n16091), .ZN(n12687) );
  NAND2_X1 U15857 ( .A1(n12688), .A2(n12687), .ZN(n14319) );
  MUX2_X1 U15858 ( .A(n12717), .B(n12642), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12692) );
  NAND2_X1 U15859 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13101), .ZN(
        n12689) );
  AND2_X1 U15860 ( .A1(n12690), .A2(n12689), .ZN(n12691) );
  MUX2_X1 U15861 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12694) );
  INV_X1 U15862 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U15863 ( .A1(n13205), .A2(n14584), .ZN(n12693) );
  NAND2_X1 U15864 ( .A1(n12694), .A2(n12693), .ZN(n14299) );
  MUX2_X1 U15865 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12695) );
  NAND2_X1 U15866 ( .A1(n12695), .A2(n10074), .ZN(n14286) );
  INV_X1 U15867 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15841) );
  NAND2_X1 U15868 ( .A1(n12706), .A2(n15841), .ZN(n12699) );
  INV_X1 U15869 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U15870 ( .A1(n12642), .A2(n16081), .ZN(n12697) );
  NAND2_X1 U15871 ( .A1(n13221), .A2(n15841), .ZN(n12696) );
  NAND3_X1 U15872 ( .A1(n12624), .A2(n12697), .A3(n12696), .ZN(n12698) );
  AND2_X1 U15873 ( .A1(n12699), .A2(n12698), .ZN(n14285) );
  NOR2_X1 U15874 ( .A1(n14286), .A2(n14285), .ZN(n12700) );
  INV_X1 U15875 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U15876 ( .A1(n12706), .A2(n14281), .ZN(n12704) );
  INV_X1 U15877 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16067) );
  NAND2_X1 U15878 ( .A1(n12642), .A2(n16067), .ZN(n12702) );
  NAND2_X1 U15879 ( .A1(n13221), .A2(n14281), .ZN(n12701) );
  NAND3_X1 U15880 ( .A1(n12624), .A2(n12702), .A3(n12701), .ZN(n12703) );
  NAND2_X1 U15881 ( .A1(n12704), .A2(n12703), .ZN(n14210) );
  MUX2_X1 U15882 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12705) );
  OAI21_X1 U15883 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n12712), .A(
        n12705), .ZN(n14197) );
  INV_X1 U15884 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14278) );
  NAND2_X1 U15885 ( .A1(n12706), .A2(n14278), .ZN(n12710) );
  INV_X1 U15886 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14421) );
  NAND2_X1 U15887 ( .A1(n12642), .A2(n14421), .ZN(n12708) );
  NAND2_X1 U15888 ( .A1(n13221), .A2(n14278), .ZN(n12707) );
  NAND3_X1 U15889 ( .A1(n12624), .A2(n12708), .A3(n12707), .ZN(n12709) );
  AND2_X1 U15890 ( .A1(n12710), .A2(n12709), .ZN(n14180) );
  MUX2_X1 U15891 ( .A(n12711), .B(n12624), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12713) );
  AND2_X1 U15892 ( .A1(n12713), .A2(n10069), .ZN(n14169) );
  INV_X1 U15893 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20953) );
  NAND2_X1 U15894 ( .A1(n12642), .A2(n20953), .ZN(n12715) );
  INV_X1 U15895 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14276) );
  NAND2_X1 U15896 ( .A1(n13221), .A2(n14276), .ZN(n12714) );
  NAND3_X1 U15897 ( .A1(n12624), .A2(n12715), .A3(n12714), .ZN(n12716) );
  OAI21_X1 U15898 ( .B1(n12717), .B2(P1_EBX_REG_28__SCAN_IN), .A(n12716), .ZN(
        n14154) );
  INV_X1 U15899 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14537) );
  NOR2_X1 U15900 ( .A1(n13101), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12718) );
  AOI21_X1 U15901 ( .B1(n13205), .B2(n14537), .A(n12718), .ZN(n12857) );
  MUX2_X1 U15902 ( .A(n12857), .B(n12718), .S(n12858), .Z(n13814) );
  NAND2_X1 U15903 ( .A1(n14156), .A2(n13814), .ZN(n13813) );
  AND2_X1 U15904 ( .A1(n13221), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U15905 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20864) );
  AND2_X1 U15906 ( .A1(n20864), .A2(n20857), .ZN(n15784) );
  INV_X1 U15907 ( .A(n15784), .ZN(n12720) );
  NAND2_X1 U15908 ( .A1(n12727), .A2(n12720), .ZN(n12721) );
  NAND2_X1 U15909 ( .A1(n12722), .A2(n20970), .ZN(n15805) );
  INV_X1 U15910 ( .A(n15805), .ZN(n13336) );
  OR2_X1 U15911 ( .A1(n11757), .A2(n13336), .ZN(n13386) );
  NAND2_X1 U15912 ( .A1(n13386), .A2(n15784), .ZN(n12728) );
  NOR2_X1 U15913 ( .A1(n12728), .A2(n13209), .ZN(n12723) );
  AOI21_X1 U15914 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(P1_REIP_REG_29__SCAN_IN), 
        .A(n19994), .ZN(n12726) );
  INV_X1 U15915 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20818) );
  INV_X1 U15916 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15919) );
  INV_X1 U15917 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15931) );
  INV_X1 U15918 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20799) );
  NAND3_X1 U15919 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14255) );
  NOR2_X1 U15920 ( .A1(n20799), .A2(n14255), .ZN(n14256) );
  NAND3_X1 U15921 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n19952) );
  NOR2_X1 U15922 ( .A1(n13724), .A2(n19952), .ZN(n15918) );
  NAND4_X1 U15923 ( .A1(n14256), .A2(n15918), .A3(P1_REIP_REG_10__SCAN_IN), 
        .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n15925) );
  NOR3_X1 U15924 ( .A1(n15919), .A2(n15931), .A3(n15925), .ZN(n14241) );
  AND3_X1 U15925 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14241), .ZN(n14230) );
  AND4_X1 U15926 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n14230), .ZN(n15873) );
  NAND2_X1 U15927 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15873), .ZN(n15868) );
  NOR2_X1 U15928 ( .A1(n20818), .A2(n15868), .ZN(n15845) );
  INV_X1 U15929 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20823) );
  NAND2_X1 U15930 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15839) );
  NOR2_X1 U15931 ( .A1(n20823), .A2(n15839), .ZN(n15832) );
  NAND3_X1 U15932 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15845), .A3(n15832), 
        .ZN(n14213) );
  NAND2_X1 U15933 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n12724) );
  NOR2_X1 U15934 ( .A1(n14213), .A2(n12724), .ZN(n14187) );
  NAND2_X1 U15935 ( .A1(n14187), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14173) );
  NAND2_X1 U15936 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12725) );
  OR2_X1 U15937 ( .A1(n14173), .A2(n12725), .ZN(n14144) );
  NAND2_X1 U15938 ( .A1(n19962), .A2(n14144), .ZN(n14163) );
  NAND2_X1 U15939 ( .A1(n14163), .A2(n15872), .ZN(n14157) );
  NOR2_X1 U15940 ( .A1(n12726), .A2(n14157), .ZN(n14135) );
  INV_X1 U15941 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20840) );
  INV_X1 U15942 ( .A(n12727), .ZN(n12729) );
  NAND3_X1 U15943 ( .A1(n12729), .A2(n20109), .A3(n12728), .ZN(n12730) );
  INV_X2 U15944 ( .A(n15883), .ZN(n19963) );
  AOI22_X1 U15945 ( .A1(n19963), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19989), .ZN(n12732) );
  INV_X1 U15946 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20836) );
  NOR3_X1 U15947 ( .A1(n19994), .A2(n20836), .A3(n14144), .ZN(n14134) );
  NAND3_X1 U15948 ( .A1(n14134), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n20840), 
        .ZN(n12731) );
  OAI211_X1 U15949 ( .C1(n14135), .C2(n20840), .A(n12732), .B(n12731), .ZN(
        n12733) );
  AOI21_X1 U15950 ( .B1(n14542), .B2(n19977), .A(n12733), .ZN(n12734) );
  NAND2_X1 U15951 ( .A1(n12735), .A2(n12734), .ZN(P1_U2809) );
  XNOR2_X1 U15952 ( .A(n12750), .B(n12751), .ZN(n12737) );
  OAI211_X1 U15953 ( .C1(n13208), .C2(n12737), .A(n13204), .B(n20138), .ZN(
        n12738) );
  INV_X1 U15954 ( .A(n12738), .ZN(n12739) );
  NAND2_X1 U15955 ( .A1(n20107), .A2(n12803), .ZN(n12744) );
  NAND2_X1 U15956 ( .A1(n13209), .A2(n20130), .ZN(n12756) );
  OAI21_X1 U15957 ( .B1(n13208), .B2(n12750), .A(n12756), .ZN(n12742) );
  INV_X1 U15958 ( .A(n12742), .ZN(n12743) );
  NAND2_X1 U15959 ( .A1(n12744), .A2(n12743), .ZN(n20079) );
  NAND2_X1 U15960 ( .A1(n13274), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12748) );
  INV_X1 U15961 ( .A(n12745), .ZN(n12746) );
  OR2_X1 U15962 ( .A1(n20080), .A2(n12746), .ZN(n12747) );
  INV_X1 U15963 ( .A(n12803), .ZN(n12775) );
  NAND2_X1 U15964 ( .A1(n12751), .A2(n12750), .ZN(n12753) );
  AND2_X1 U15965 ( .A1(n12753), .A2(n12752), .ZN(n12767) );
  NOR2_X1 U15966 ( .A1(n12753), .A2(n12752), .ZN(n12754) );
  OAI21_X1 U15967 ( .B1(n12767), .B2(n12754), .A(n11773), .ZN(n12755) );
  NAND2_X1 U15968 ( .A1(n12757), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12758) );
  OR2_X1 U15969 ( .A1(n12759), .A2(n12775), .ZN(n12762) );
  XNOR2_X1 U15970 ( .A(n12767), .B(n12766), .ZN(n12760) );
  NAND2_X1 U15971 ( .A1(n12760), .A2(n11773), .ZN(n12761) );
  NAND2_X1 U15972 ( .A1(n12762), .A2(n12761), .ZN(n13526) );
  NAND2_X1 U15973 ( .A1(n12765), .A2(n12803), .ZN(n12772) );
  INV_X1 U15974 ( .A(n12766), .ZN(n12768) );
  NOR2_X1 U15975 ( .A1(n12768), .A2(n12767), .ZN(n12778) );
  INV_X1 U15976 ( .A(n12778), .ZN(n12769) );
  XNOR2_X1 U15977 ( .A(n12777), .B(n12769), .ZN(n12770) );
  NAND2_X1 U15978 ( .A1(n11773), .A2(n12770), .ZN(n12771) );
  NAND2_X1 U15979 ( .A1(n12772), .A2(n12771), .ZN(n12774) );
  INV_X1 U15980 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12773) );
  XNOR2_X1 U15981 ( .A(n12774), .B(n12773), .ZN(n13548) );
  OR2_X1 U15982 ( .A1(n12776), .A2(n12775), .ZN(n12781) );
  NAND2_X1 U15983 ( .A1(n12778), .A2(n12777), .ZN(n12786) );
  XNOR2_X1 U15984 ( .A(n12785), .B(n12786), .ZN(n12779) );
  NAND2_X1 U15985 ( .A1(n11773), .A2(n12779), .ZN(n12780) );
  NAND2_X1 U15986 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  XNOR2_X1 U15987 ( .A(n12782), .B(n16205), .ZN(n16025) );
  NAND2_X1 U15988 ( .A1(n12782), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12783) );
  NAND3_X1 U15989 ( .A1(n12807), .A2(n12784), .A3(n12803), .ZN(n12791) );
  INV_X1 U15990 ( .A(n12785), .ZN(n12787) );
  NOR2_X1 U15991 ( .A1(n12787), .A2(n12786), .ZN(n12797) );
  INV_X1 U15992 ( .A(n12797), .ZN(n12788) );
  XNOR2_X1 U15993 ( .A(n12796), .B(n12788), .ZN(n12789) );
  NAND2_X1 U15994 ( .A1(n11773), .A2(n12789), .ZN(n12790) );
  AND2_X1 U15995 ( .A1(n12791), .A2(n12790), .ZN(n12792) );
  INV_X1 U15996 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16180) );
  NAND2_X1 U15997 ( .A1(n12792), .A2(n16180), .ZN(n16019) );
  NAND2_X1 U15998 ( .A1(n16017), .A2(n16019), .ZN(n12794) );
  INV_X1 U15999 ( .A(n12792), .ZN(n12793) );
  NAND2_X1 U16000 ( .A1(n12793), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16018) );
  NAND2_X1 U16001 ( .A1(n12795), .A2(n12803), .ZN(n12800) );
  NAND2_X1 U16002 ( .A1(n12797), .A2(n12796), .ZN(n12808) );
  XNOR2_X1 U16003 ( .A(n12810), .B(n12808), .ZN(n12798) );
  NAND2_X1 U16004 ( .A1(n11773), .A2(n12798), .ZN(n12799) );
  NAND2_X1 U16005 ( .A1(n12800), .A2(n12799), .ZN(n16013) );
  OR2_X1 U16006 ( .A1(n16013), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12801) );
  NAND2_X1 U16007 ( .A1(n16013), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12802) );
  NAND2_X1 U16008 ( .A1(n12803), .A2(n12810), .ZN(n12805) );
  NOR2_X1 U16009 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  NAND2_X4 U16010 ( .A1(n12807), .A2(n12806), .ZN(n14579) );
  INV_X1 U16011 ( .A(n12808), .ZN(n12809) );
  NAND3_X1 U16012 ( .A1(n11773), .A2(n12810), .A3(n12809), .ZN(n12811) );
  NAND2_X1 U16013 ( .A1(n14579), .A2(n12811), .ZN(n13722) );
  INV_X1 U16014 ( .A(n13722), .ZN(n12812) );
  INV_X1 U16015 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U16016 ( .A1(n12812), .A2(n16183), .ZN(n12813) );
  INV_X2 U16017 ( .A(n14579), .ZN(n12833) );
  NAND2_X1 U16018 ( .A1(n12833), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12814) );
  NAND2_X1 U16019 ( .A1(n14579), .A2(n16170), .ZN(n12815) );
  NOR2_X1 U16020 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12816) );
  INV_X1 U16021 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16127) );
  NAND2_X1 U16022 ( .A1(n14579), .A2(n16127), .ZN(n14510) );
  NAND2_X1 U16023 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12817) );
  NAND2_X1 U16024 ( .A1(n14579), .A2(n12817), .ZN(n14508) );
  AND2_X1 U16025 ( .A1(n14510), .A2(n14508), .ZN(n12818) );
  INV_X1 U16026 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12819) );
  INV_X1 U16027 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U16028 ( .A1(n12820), .A2(n12819), .ZN(n12821) );
  NAND2_X1 U16029 ( .A1(n12833), .A2(n12821), .ZN(n12825) );
  XNOR2_X1 U16030 ( .A(n14579), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14491) );
  NAND2_X1 U16031 ( .A1(n14579), .A2(n16115), .ZN(n15990) );
  NAND2_X1 U16032 ( .A1(n14491), .A2(n15990), .ZN(n12822) );
  NAND2_X1 U16033 ( .A1(n14589), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12827) );
  NAND2_X1 U16034 ( .A1(n12833), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14509) );
  NAND2_X1 U16035 ( .A1(n16147), .A2(n12823), .ZN(n12824) );
  NAND2_X1 U16036 ( .A1(n12833), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15991) );
  NAND2_X1 U16037 ( .A1(n15987), .A2(n15991), .ZN(n14590) );
  XNOR2_X1 U16038 ( .A(n14579), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14481) );
  AND2_X1 U16039 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U16040 ( .A1(n14546), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12828) );
  OAI21_X2 U16041 ( .B1(n14480), .B2(n12828), .A(n14579), .ZN(n14474) );
  NAND2_X1 U16042 ( .A1(n14474), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12830) );
  INV_X1 U16043 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15816) );
  NAND2_X1 U16044 ( .A1(n14584), .A2(n15816), .ZN(n12829) );
  NAND2_X1 U16045 ( .A1(n12830), .A2(n14473), .ZN(n12831) );
  AND2_X1 U16046 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U16047 ( .A1(n14547), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14534) );
  NAND2_X1 U16048 ( .A1(n12830), .A2(n14579), .ZN(n14454) );
  NOR2_X1 U16049 ( .A1(n12831), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14455) );
  NOR2_X1 U16050 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12832) );
  AOI21_X1 U16051 ( .B1(n14455), .B2(n12832), .A(n14579), .ZN(n14447) );
  AOI21_X2 U16052 ( .B1(n14433), .B2(n14454), .A(n14447), .ZN(n14435) );
  NOR2_X1 U16053 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14574) );
  NAND2_X1 U16054 ( .A1(n14435), .A2(n14574), .ZN(n14413) );
  NAND2_X1 U16055 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14548) );
  NOR2_X2 U16056 ( .A1(n14435), .A2(n14548), .ZN(n12868) );
  AOI21_X2 U16057 ( .B1(n14413), .B2(n12833), .A(n12868), .ZN(n12872) );
  XOR2_X1 U16058 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n14519), .Z(
        n12869) );
  XNOR2_X1 U16059 ( .A(n12872), .B(n12869), .ZN(n14570) );
  NAND2_X1 U16060 ( .A1(n14623), .A2(n13209), .ZN(n12834) );
  NOR2_X1 U16061 ( .A1(n12890), .A2(n12835), .ZN(n13104) );
  NAND2_X1 U16062 ( .A1(n20635), .A2(n12836), .ZN(n20863) );
  AND2_X1 U16063 ( .A1(n20863), .A2(n20777), .ZN(n12837) );
  NAND2_X1 U16064 ( .A1(n20857), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12839) );
  NOR2_X1 U16065 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20856), .ZN(n20858) );
  INV_X1 U16066 ( .A(n20858), .ZN(n12838) );
  NAND2_X1 U16067 ( .A1(n12839), .A2(n12838), .ZN(n20084) );
  NAND2_X1 U16068 ( .A1(n12840), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14561) );
  OAI21_X1 U16069 ( .B1(n16033), .B2(n12841), .A(n14561), .ZN(n12842) );
  AOI21_X1 U16070 ( .B1(n16027), .B2(n14145), .A(n12842), .ZN(n12848) );
  NAND2_X1 U16071 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20859), .ZN(n16221) );
  INV_X1 U16072 ( .A(n16221), .ZN(n12847) );
  NAND3_X1 U16073 ( .A1(n12849), .A2(n12848), .A3(n9662), .ZN(P1_U2970) );
  INV_X1 U16074 ( .A(n14419), .ZN(n14367) );
  NAND2_X1 U16075 ( .A1(n13424), .A2(n11757), .ZN(n12852) );
  NOR2_X1 U16076 ( .A1(n12853), .A2(n12852), .ZN(n13461) );
  NAND2_X1 U16077 ( .A1(n13461), .A2(n13395), .ZN(n13232) );
  NAND4_X1 U16078 ( .A1(n12854), .A2(n13474), .A3(n13810), .A4(n20142), .ZN(
        n12891) );
  OR2_X1 U16079 ( .A1(n12891), .A2(n13101), .ZN(n12855) );
  NAND2_X1 U16080 ( .A1(n13232), .A2(n12855), .ZN(n12856) );
  NAND2_X2 U16081 ( .A1(n20014), .A2(n20148), .ZN(n14364) );
  AOI22_X1 U16082 ( .A1(n13813), .A2(n12858), .B1(n14156), .B2(n12857), .ZN(
        n12860) );
  XNOR2_X1 U16083 ( .A(n12860), .B(n12859), .ZN(n14554) );
  INV_X1 U16084 ( .A(n14554), .ZN(n12864) );
  INV_X1 U16085 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12861) );
  NOR2_X1 U16086 ( .A1(n20101), .A2(n20840), .ZN(n14541) );
  AOI21_X1 U16087 ( .B1(n20085), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14541), .ZN(n12866) );
  OAI21_X1 U16088 ( .B1(n16023), .B2(n13601), .A(n12866), .ZN(n12867) );
  AOI21_X1 U16089 ( .B1(n12896), .B2(n16029), .A(n12867), .ZN(n12875) );
  INV_X1 U16090 ( .A(n12868), .ZN(n14414) );
  NAND2_X1 U16091 ( .A1(n14414), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12871) );
  AOI21_X1 U16092 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14537), .A(
        n12869), .ZN(n12870) );
  OAI211_X1 U16093 ( .C1(n12872), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12871), .B(n12870), .ZN(n12874) );
  INV_X1 U16094 ( .A(n16435), .ZN(n16437) );
  NAND2_X1 U16095 ( .A1(n16434), .A2(n16437), .ZN(n12876) );
  XOR2_X1 U16096 ( .A(n17729), .B(n12876), .Z(n17940) );
  NAND2_X1 U16097 ( .A1(n17581), .A2(n12877), .ZN(n16586) );
  INV_X1 U16098 ( .A(n16586), .ZN(n16585) );
  OAI21_X1 U16099 ( .B1(n16585), .B2(n18771), .A(n17922), .ZN(n12878) );
  AOI21_X1 U16100 ( .B1(n17676), .B2(n12879), .A(n12878), .ZN(n17583) );
  OAI21_X1 U16101 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17702), .A(
        n17583), .ZN(n17571) );
  INV_X1 U16102 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16639) );
  NOR2_X1 U16103 ( .A1(n16639), .A2(n16584), .ZN(n16583) );
  AOI21_X1 U16104 ( .B1(n16639), .B2(n16584), .A(n16583), .ZN(n16638) );
  AOI22_X1 U16105 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17571), .B1(
        n17758), .B2(n16638), .ZN(n12880) );
  NAND2_X1 U16106 ( .A1(n9587), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17938) );
  OAI211_X1 U16107 ( .C1(n17940), .C2(n17807), .A(n12880), .B(n17938), .ZN(
        n12881) );
  INV_X1 U16108 ( .A(n12881), .ZN(n12887) );
  NAND2_X1 U16109 ( .A1(n17582), .A2(n17763), .ZN(n17609) );
  NOR2_X1 U16110 ( .A1(n12882), .A2(n17609), .ZN(n17565) );
  OAI22_X1 U16111 ( .A1(n17926), .A2(n18123), .B1(n17837), .B2(n17792), .ZN(
        n12883) );
  NAND2_X1 U16112 ( .A1(n12884), .A2(n17708), .ZN(n17578) );
  INV_X1 U16113 ( .A(n16407), .ZN(n17932) );
  INV_X1 U16114 ( .A(n16418), .ZN(n17931) );
  OAI22_X1 U16115 ( .A1(n17932), .A2(n17926), .B1(n17931), .B2(n17837), .ZN(
        n17590) );
  NOR2_X1 U16116 ( .A1(n17928), .A2(n17590), .ZN(n17563) );
  INV_X1 U16117 ( .A(n12888), .ZN(n16213) );
  AND2_X1 U16118 ( .A1(n13110), .A2(n20864), .ZN(n13384) );
  NAND2_X1 U16119 ( .A1(n16213), .A2(n13384), .ZN(n13230) );
  NAND2_X1 U16120 ( .A1(n13220), .A2(n20864), .ZN(n13389) );
  INV_X1 U16121 ( .A(n12890), .ZN(n13227) );
  NAND2_X1 U16122 ( .A1(n13227), .A2(n13599), .ZN(n13459) );
  OAI21_X1 U16123 ( .B1(n13389), .B2(n13101), .A(n13459), .ZN(n12893) );
  NOR2_X1 U16124 ( .A1(n12891), .A2(n13102), .ZN(n12892) );
  AOI21_X1 U16125 ( .B1(n12893), .B2(n13390), .A(n12892), .ZN(n12894) );
  NAND2_X1 U16126 ( .A1(n13230), .A2(n12894), .ZN(n12895) );
  INV_X2 U16127 ( .A(n14405), .ZN(n15946) );
  NOR4_X1 U16128 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12900) );
  NOR4_X1 U16129 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12899) );
  NOR4_X1 U16130 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12898) );
  NOR4_X1 U16131 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12897) );
  AND4_X1 U16132 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12905) );
  NOR4_X1 U16133 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12903) );
  NOR4_X1 U16134 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12902) );
  NOR4_X1 U16135 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12901) );
  INV_X1 U16136 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20797) );
  AND4_X1 U16137 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n20797), .ZN(
        n12904) );
  NAND2_X1 U16138 ( .A1(n12905), .A2(n12904), .ZN(n12906) );
  NAND2_X1 U16139 ( .A1(n12907), .A2(n20104), .ZN(n12908) );
  INV_X1 U16140 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16451) );
  NOR2_X1 U16141 ( .A1(n15953), .A2(n16451), .ZN(n12911) );
  NOR3_X4 U16142 ( .A1(n15946), .A2(n20104), .A3(n13387), .ZN(n15949) );
  AOI22_X1 U16143 ( .A1(n15949), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15946), .ZN(n12909) );
  INV_X1 U16144 ( .A(n12909), .ZN(n12910) );
  NOR2_X1 U16145 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  NAND2_X1 U16146 ( .A1(n12913), .A2(n12912), .ZN(P1_U2873) );
  NOR2_X1 U16147 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12915) );
  NOR4_X1 U16148 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12914) );
  NAND4_X1 U16149 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12915), .A4(n12914), .ZN(n12927) );
  INV_X1 U16150 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20855) );
  NOR3_X1 U16151 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20855), .ZN(n12917) );
  NOR4_X1 U16152 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12916) );
  NAND4_X1 U16153 ( .A1(n20104), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12917), .A4(
        n12916), .ZN(U214) );
  NOR4_X1 U16154 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12921) );
  NOR4_X1 U16155 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12920) );
  NOR4_X1 U16156 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12919) );
  NOR4_X1 U16157 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12918) );
  NAND4_X1 U16158 ( .A1(n12921), .A2(n12920), .A3(n12919), .A4(n12918), .ZN(
        n12926) );
  NOR4_X1 U16159 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12924) );
  NOR4_X1 U16160 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12923) );
  NOR4_X1 U16161 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12922) );
  INV_X1 U16162 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19807) );
  NAND4_X1 U16163 ( .A1(n12924), .A2(n12923), .A3(n12922), .A4(n19807), .ZN(
        n12925) );
  NOR2_X1 U16164 ( .A1(n13375), .A2(n12927), .ZN(n16450) );
  NAND2_X1 U16165 ( .A1(n16450), .A2(U214), .ZN(U212) );
  OR2_X1 U16166 ( .A1(n10748), .A2(n16388), .ZN(n13070) );
  NOR2_X1 U16167 ( .A1(n12930), .A2(n13070), .ZN(n13757) );
  INV_X1 U16168 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12933) );
  INV_X1 U16169 ( .A(n12928), .ZN(n12929) );
  NAND2_X1 U16170 ( .A1(n12929), .A2(n19777), .ZN(n12931) );
  INV_X1 U16171 ( .A(n13649), .ZN(n13009) );
  INV_X1 U16172 ( .A(n19869), .ZN(n19722) );
  NOR2_X1 U16173 ( .A1(n19722), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12935) );
  INV_X1 U16174 ( .A(n12935), .ZN(n12932) );
  OAI211_X1 U16175 ( .C1(n13757), .C2(n12933), .A(n13009), .B(n12932), .ZN(
        P2_U2814) );
  INV_X1 U16176 ( .A(n11286), .ZN(n12938) );
  NOR2_X1 U16177 ( .A1(n9594), .A2(n16388), .ZN(n12934) );
  INV_X1 U16178 ( .A(n21033), .ZN(n12937) );
  OAI21_X1 U16179 ( .B1(n12935), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n12937), 
        .ZN(n12936) );
  OAI21_X1 U16180 ( .B1(n12938), .B2(n12937), .A(n12936), .ZN(P2_U3612) );
  NAND2_X1 U16181 ( .A1(n11286), .A2(n21038), .ZN(n12940) );
  NAND4_X1 U16182 ( .A1(n12939), .A2(n16360), .A3(n13639), .A4(n12940), .ZN(
        n16371) );
  NAND2_X1 U16183 ( .A1(n16371), .A2(n19777), .ZN(n19908) );
  INV_X1 U16184 ( .A(n19908), .ZN(n12942) );
  OAI21_X1 U16185 ( .B1(n12950), .B2(n12942), .A(n12941), .ZN(P2_U2819) );
  OR2_X1 U16186 ( .A1(n10748), .A2(n13639), .ZN(n12949) );
  NAND3_X1 U16187 ( .A1(n12943), .A2(n11286), .A3(n12939), .ZN(n12944) );
  OAI21_X1 U16188 ( .B1(n16367), .B2(n13181), .A(n12944), .ZN(n12945) );
  INV_X1 U16189 ( .A(n12945), .ZN(n13123) );
  NAND2_X1 U16190 ( .A1(n16367), .A2(n12946), .ZN(n12982) );
  AND2_X1 U16191 ( .A1(n12982), .A2(n12947), .ZN(n12948) );
  OAI211_X1 U16192 ( .C1(n13071), .C2(n12949), .A(n13123), .B(n12948), .ZN(
        n16376) );
  NOR2_X1 U16193 ( .A1(n21039), .A2(n13073), .ZN(n15824) );
  INV_X1 U16194 ( .A(n15824), .ZN(n16394) );
  OAI22_X1 U16195 ( .A1(n16394), .A2(n12950), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19678), .ZN(n12951) );
  AOI21_X1 U16196 ( .B1(n16376), .B2(n19777), .A(n12951), .ZN(n15599) );
  INV_X1 U16197 ( .A(n15599), .ZN(n12956) );
  INV_X1 U16198 ( .A(n12952), .ZN(n12953) );
  NAND2_X1 U16199 ( .A1(n14062), .A2(n12953), .ZN(n12954) );
  NOR2_X1 U16200 ( .A1(n10748), .A2(n12954), .ZN(n16368) );
  NAND3_X1 U16201 ( .A1(n12956), .A2(n16368), .A3(n19779), .ZN(n12955) );
  OAI21_X1 U16202 ( .B1(n12956), .B2(n16375), .A(n12955), .ZN(P2_U3595) );
  INV_X1 U16203 ( .A(n12957), .ZN(n12958) );
  INV_X1 U16204 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20952) );
  NAND2_X1 U16205 ( .A1(n20716), .A2(n20776), .ZN(n19916) );
  OAI211_X1 U16206 ( .C1(n12958), .C2(n20952), .A(n13287), .B(n19916), .ZN(
        P1_U2801) );
  OAI21_X1 U16207 ( .B1(n13736), .B2(n12960), .A(n12959), .ZN(n12961) );
  XOR2_X1 U16208 ( .A(n12961), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(
        n19260) );
  OAI21_X1 U16209 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n19265) );
  OR2_X1 U16210 ( .A1(n19088), .A2(n19804), .ZN(n19262) );
  INV_X1 U16211 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12965) );
  OR2_X1 U16212 ( .A1(n16315), .A2(n12965), .ZN(n12966) );
  OAI211_X1 U16213 ( .C1(n19265), .C2(n16308), .A(n19262), .B(n12966), .ZN(
        n12969) );
  OAI21_X1 U16214 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13632), .ZN(n13730) );
  INV_X1 U16215 ( .A(n13730), .ZN(n12967) );
  AND2_X1 U16216 ( .A1(n16305), .A2(n12967), .ZN(n12968) );
  NOR2_X1 U16217 ( .A1(n12969), .A2(n12968), .ZN(n12971) );
  NAND2_X1 U16218 ( .A1(n13738), .A2(n16311), .ZN(n12970) );
  OAI211_X1 U16219 ( .C1(n19260), .C2(n16306), .A(n12971), .B(n12970), .ZN(
        P2_U3012) );
  INV_X1 U16220 ( .A(n12972), .ZN(n12973) );
  NAND2_X1 U16221 ( .A1(n13155), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12975) );
  NAND2_X1 U16222 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19375) );
  OAI21_X1 U16223 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n19375), .ZN(n15616) );
  INV_X1 U16224 ( .A(n15616), .ZN(n12974) );
  NAND2_X1 U16225 ( .A1(n12974), .A2(n19869), .ZN(n19581) );
  NAND2_X1 U16226 ( .A1(n12975), .A2(n19581), .ZN(n12976) );
  AOI22_X1 U16227 ( .A1(n13155), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19869), .B2(n19900), .ZN(n12977) );
  NAND2_X1 U16228 ( .A1(n14034), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13061) );
  AOI21_X4 U16229 ( .B1(n12982), .B2(n11295), .A(n16388), .ZN(n19159) );
  NAND2_X1 U16230 ( .A1(n19159), .A2(n13125), .ZN(n19148) );
  MUX2_X1 U16231 ( .A(n12983), .B(n13784), .S(n19159), .Z(n12984) );
  OAI21_X1 U16232 ( .B1(n19278), .B2(n19148), .A(n12984), .ZN(P2_U2886) );
  AOI21_X1 U16233 ( .B1(n13670), .B2(n12986), .A(n12985), .ZN(n13144) );
  NAND2_X1 U16234 ( .A1(n19115), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13140) );
  INV_X1 U16235 ( .A(n13140), .ZN(n12992) );
  INV_X1 U16236 ( .A(n12987), .ZN(n12990) );
  NAND2_X1 U16237 ( .A1(n12988), .A2(n12986), .ZN(n12989) );
  NAND2_X1 U16238 ( .A1(n12990), .A2(n12989), .ZN(n13141) );
  NOR2_X1 U16239 ( .A1(n16308), .A2(n13141), .ZN(n12991) );
  AOI211_X1 U16240 ( .C1(n13144), .C2(n16293), .A(n12992), .B(n12991), .ZN(
        n12995) );
  OAI21_X1 U16241 ( .B1(n16297), .B2(n12993), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12994) );
  OAI211_X1 U16242 ( .C1(n13376), .C2(n15579), .A(n12995), .B(n12994), .ZN(
        P2_U3014) );
  INV_X1 U16243 ( .A(n19916), .ZN(n12996) );
  NOR2_X1 U16244 ( .A1(n12996), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12999)
         );
  NAND2_X1 U16245 ( .A1(n20862), .A2(n12997), .ZN(n12998) );
  OAI21_X1 U16246 ( .B1(n20862), .B2(n12999), .A(n12998), .ZN(P1_U3487) );
  AOI21_X1 U16247 ( .B1(n13776), .B2(n13001), .A(n13000), .ZN(n15570) );
  XOR2_X1 U16248 ( .A(n13002), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n15569) );
  INV_X1 U16249 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n13003) );
  NOR2_X1 U16250 ( .A1(n11494), .A2(n13003), .ZN(n15568) );
  AOI21_X1 U16251 ( .B1(n11517), .B2(n15569), .A(n15568), .ZN(n13006) );
  INV_X1 U16252 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13746) );
  NAND2_X1 U16253 ( .A1(n16305), .A2(n13746), .ZN(n13005) );
  NAND2_X1 U16254 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13004) );
  NAND3_X1 U16255 ( .A1(n13006), .A2(n13005), .A3(n13004), .ZN(n13007) );
  AOI21_X1 U16256 ( .B1(n15570), .B2(n16293), .A(n13007), .ZN(n13008) );
  OAI21_X1 U16257 ( .B1(n13784), .B2(n13376), .A(n13008), .ZN(P2_U3013) );
  NOR3_X1 U16258 ( .A1(n13009), .A2(n14062), .A3(n19786), .ZN(n13010) );
  CLKBUF_X1 U16259 ( .A(n13010), .Z(n13098) );
  OAI22_X1 U16260 ( .A1(n14109), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14110), .ZN(n19303) );
  INV_X1 U16261 ( .A(n19303), .ZN(n16259) );
  NAND2_X1 U16262 ( .A1(n13098), .A2(n16259), .ZN(n13021) );
  OAI21_X1 U16263 ( .B1(n14062), .B2(n21038), .A(n13649), .ZN(n13094) );
  AOI22_X1 U16264 ( .A1(n13078), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13094), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U16265 ( .A1(n13021), .A2(n13011), .ZN(P2_U2958) );
  INV_X1 U16266 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13012) );
  OR2_X1 U16267 ( .A1(n14109), .A2(n13012), .ZN(n13014) );
  NAND2_X1 U16268 ( .A1(n13375), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13013) );
  AND2_X1 U16269 ( .A1(n13014), .A2(n13013), .ZN(n19179) );
  INV_X1 U16270 ( .A(n19179), .ZN(n13015) );
  NAND2_X1 U16271 ( .A1(n13098), .A2(n13015), .ZN(n13042) );
  AOI22_X1 U16272 ( .A1(n13078), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13094), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U16273 ( .A1(n13042), .A2(n13016), .ZN(P2_U2980) );
  AOI22_X1 U16274 ( .A1(n14110), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13375), .ZN(n19223) );
  INV_X1 U16275 ( .A(n19223), .ZN(n14989) );
  NAND2_X1 U16276 ( .A1(n13098), .A2(n14989), .ZN(n13044) );
  INV_X1 U16277 ( .A(n13094), .ZN(n13137) );
  AOI22_X1 U16278 ( .A1(n13078), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U16279 ( .A1(n13044), .A2(n13017), .ZN(P2_U2953) );
  AOI22_X1 U16280 ( .A1(n14110), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13375), .ZN(n19311) );
  INV_X1 U16281 ( .A(n19311), .ZN(n13018) );
  NAND2_X1 U16282 ( .A1(n13098), .A2(n13018), .ZN(n13038) );
  AOI22_X1 U16283 ( .A1(n13078), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16284 ( .A1(n13038), .A2(n13019), .ZN(P2_U2959) );
  AOI22_X1 U16285 ( .A1(n13078), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13020) );
  NAND2_X1 U16286 ( .A1(n13021), .A2(n13020), .ZN(P2_U2973) );
  AOI22_X1 U16287 ( .A1(n14110), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13375), .ZN(n19293) );
  INV_X1 U16288 ( .A(n19293), .ZN(n14980) );
  NAND2_X1 U16289 ( .A1(n13098), .A2(n14980), .ZN(n13029) );
  AOI22_X1 U16290 ( .A1(n13078), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13094), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U16291 ( .A1(n13029), .A2(n13022), .ZN(P2_U2955) );
  INV_X1 U16292 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13023) );
  OR2_X1 U16293 ( .A1(n13375), .A2(n13023), .ZN(n13025) );
  NAND2_X1 U16294 ( .A1(n13375), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13024) );
  AND2_X1 U16295 ( .A1(n13025), .A2(n13024), .ZN(n19184) );
  INV_X1 U16296 ( .A(n19184), .ZN(n13026) );
  NAND2_X1 U16297 ( .A1(n13098), .A2(n13026), .ZN(n13031) );
  AOI22_X1 U16298 ( .A1(n13078), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13094), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U16299 ( .A1(n13031), .A2(n13027), .ZN(P2_U2978) );
  AOI22_X1 U16300 ( .A1(n13078), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U16301 ( .A1(n13029), .A2(n13028), .ZN(P2_U2970) );
  AOI22_X1 U16302 ( .A1(n13078), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U16303 ( .A1(n13031), .A2(n13030), .ZN(P2_U2963) );
  INV_X1 U16304 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n13032) );
  OR2_X1 U16305 ( .A1(n14109), .A2(n13032), .ZN(n13034) );
  NAND2_X1 U16306 ( .A1(n14109), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13033) );
  AND2_X1 U16307 ( .A1(n13034), .A2(n13033), .ZN(n19182) );
  INV_X1 U16308 ( .A(n19182), .ZN(n13035) );
  NAND2_X1 U16309 ( .A1(n13098), .A2(n13035), .ZN(n13040) );
  AOI22_X1 U16310 ( .A1(n13078), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U16311 ( .A1(n13040), .A2(n13036), .ZN(P2_U2964) );
  AOI22_X1 U16312 ( .A1(n13078), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U16313 ( .A1(n13038), .A2(n13037), .ZN(P2_U2974) );
  AOI22_X1 U16314 ( .A1(n13078), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13091), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U16315 ( .A1(n13040), .A2(n13039), .ZN(P2_U2979) );
  AOI22_X1 U16316 ( .A1(n13078), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U16317 ( .A1(n13042), .A2(n13041), .ZN(P2_U2965) );
  AOI22_X1 U16318 ( .A1(n13078), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13043) );
  NAND2_X1 U16319 ( .A1(n13044), .A2(n13043), .ZN(P2_U2968) );
  OAI22_X1 U16320 ( .A1(n14109), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14110), .ZN(n13448) );
  INV_X1 U16321 ( .A(n13448), .ZN(n16271) );
  NAND2_X1 U16322 ( .A1(n13098), .A2(n16271), .ZN(n13047) );
  AOI22_X1 U16323 ( .A1(n13078), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13045) );
  NAND2_X1 U16324 ( .A1(n13047), .A2(n13045), .ZN(P2_U2969) );
  AOI22_X1 U16325 ( .A1(n13078), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13094), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U16326 ( .A1(n13047), .A2(n13046), .ZN(P2_U2954) );
  OAI22_X1 U16327 ( .A1(n14109), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14110), .ZN(n19297) );
  INV_X1 U16328 ( .A(n19297), .ZN(n16265) );
  NAND2_X1 U16329 ( .A1(n13098), .A2(n16265), .ZN(n13050) );
  AOI22_X1 U16330 ( .A1(n13078), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U16331 ( .A1(n13050), .A2(n13048), .ZN(P2_U2971) );
  AOI22_X1 U16332 ( .A1(n13078), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13094), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U16333 ( .A1(n13050), .A2(n13049), .ZN(P2_U2956) );
  MUX2_X1 U16334 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n14109), .Z(n19189) );
  NAND2_X1 U16335 ( .A1(n13098), .A2(n19189), .ZN(n13082) );
  AOI22_X1 U16336 ( .A1(n13078), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13051) );
  NAND2_X1 U16337 ( .A1(n13082), .A2(n13051), .ZN(P2_U2961) );
  NAND2_X1 U16338 ( .A1(n13052), .A2(n13150), .ZN(n13055) );
  NAND2_X1 U16339 ( .A1(n19375), .A2(n19881), .ZN(n13053) );
  NOR2_X1 U16340 ( .A1(n19881), .A2(n19891), .ZN(n19714) );
  AND2_X1 U16341 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19714), .ZN(
        n13152) );
  INV_X1 U16342 ( .A(n13152), .ZN(n13153) );
  AND2_X1 U16343 ( .A1(n13053), .A2(n13153), .ZN(n15617) );
  AOI22_X1 U16344 ( .A1(n13155), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19869), .B2(n15617), .ZN(n13054) );
  NAND2_X1 U16345 ( .A1(n13055), .A2(n13054), .ZN(n13058) );
  NOR2_X1 U16346 ( .A1(n13192), .A2(n13056), .ZN(n13057) );
  NAND2_X1 U16347 ( .A1(n13058), .A2(n13057), .ZN(n13148) );
  NAND2_X1 U16348 ( .A1(n13059), .A2(n13148), .ZN(n13067) );
  NAND2_X1 U16349 ( .A1(n13117), .A2(n13061), .ZN(n13062) );
  NAND2_X1 U16350 ( .A1(n13063), .A2(n13062), .ZN(n13066) );
  NAND2_X1 U16351 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  INV_X1 U16352 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13732) );
  MUX2_X1 U16353 ( .A(n13732), .B(n19258), .S(n19159), .Z(n13069) );
  OAI21_X1 U16354 ( .B1(n19877), .B2(n19148), .A(n13069), .ZN(P2_U2885) );
  INV_X1 U16355 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14929) );
  OAI21_X1 U16356 ( .B1(n13071), .B2(n13070), .A(n13647), .ZN(n13072) );
  NAND2_X1 U16357 ( .A1(n19224), .A2(n10712), .ZN(n13259) );
  NOR2_X4 U16358 ( .A1(n19224), .A2(n21034), .ZN(n19243) );
  AOI22_X1 U16359 ( .A1(n13248), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13074) );
  OAI21_X1 U16360 ( .B1(n14929), .B2(n13259), .A(n13074), .ZN(P2_U2923) );
  INV_X1 U16361 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16362 ( .A1(n13248), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13075) );
  OAI21_X1 U16363 ( .B1(n13088), .B2(n13259), .A(n13075), .ZN(P2_U2925) );
  INV_X1 U16364 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U16365 ( .A1(n13248), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13076) );
  OAI21_X1 U16366 ( .B1(n13097), .B2(n13259), .A(n13076), .ZN(P2_U2927) );
  INV_X1 U16367 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16497) );
  INV_X1 U16368 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18292) );
  OAI22_X1 U16369 ( .A1(n13375), .A2(n16497), .B1(n18292), .B2(n14110), .ZN(
        n19199) );
  NAND2_X1 U16370 ( .A1(n13098), .A2(n19199), .ZN(n13080) );
  AOI22_X1 U16371 ( .A1(n13078), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13091), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13077) );
  NAND2_X1 U16372 ( .A1(n13080), .A2(n13077), .ZN(P2_U2957) );
  AOI22_X1 U16373 ( .A1(n13078), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13091), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13079) );
  NAND2_X1 U16374 ( .A1(n13080), .A2(n13079), .ZN(P2_U2972) );
  INV_X1 U16375 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19237) );
  NAND2_X1 U16376 ( .A1(n13094), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13081) );
  OAI211_X1 U16377 ( .C1(n19237), .C2(n13647), .A(n13082), .B(n13081), .ZN(
        P2_U2976) );
  INV_X1 U16378 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19227) );
  MUX2_X1 U16379 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n14109), .Z(n19176) );
  NAND2_X1 U16380 ( .A1(n13098), .A2(n19176), .ZN(n13090) );
  NAND2_X1 U16381 ( .A1(n13091), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13083) );
  OAI211_X1 U16382 ( .C1(n19227), .C2(n13647), .A(n13090), .B(n13083), .ZN(
        P2_U2981) );
  INV_X1 U16383 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19239) );
  NAND2_X1 U16384 ( .A1(n13375), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13085) );
  INV_X1 U16385 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16491) );
  OR2_X1 U16386 ( .A1(n13375), .A2(n16491), .ZN(n13084) );
  NAND2_X1 U16387 ( .A1(n13085), .A2(n13084), .ZN(n19192) );
  NAND2_X1 U16388 ( .A1(n13098), .A2(n19192), .ZN(n13096) );
  NAND2_X1 U16389 ( .A1(n13094), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13086) );
  OAI211_X1 U16390 ( .C1(n19239), .C2(n13647), .A(n13096), .B(n13086), .ZN(
        P2_U2975) );
  MUX2_X1 U16391 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n14109), .Z(n19186) );
  NAND2_X1 U16392 ( .A1(n13098), .A2(n19186), .ZN(n13093) );
  NAND2_X1 U16393 ( .A1(n13091), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13087) );
  OAI211_X1 U16394 ( .C1(n13088), .C2(n13647), .A(n13093), .B(n13087), .ZN(
        P2_U2962) );
  INV_X1 U16395 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U16396 ( .A1(n13094), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13089) );
  OAI211_X1 U16397 ( .C1(n13247), .C2(n13647), .A(n13090), .B(n13089), .ZN(
        P2_U2966) );
  INV_X1 U16398 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19235) );
  NAND2_X1 U16399 ( .A1(n13091), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13092) );
  OAI211_X1 U16400 ( .C1(n19235), .C2(n13647), .A(n13093), .B(n13092), .ZN(
        P2_U2977) );
  NAND2_X1 U16401 ( .A1(n13094), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13095) );
  OAI211_X1 U16402 ( .C1(n13097), .C2(n13647), .A(n13096), .B(n13095), .ZN(
        P2_U2960) );
  INV_X1 U16403 ( .A(n13098), .ZN(n13136) );
  OAI22_X1 U16404 ( .A1(n13375), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14110), .ZN(n13453) );
  INV_X1 U16405 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13260) );
  INV_X1 U16406 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13099) );
  OAI222_X1 U16407 ( .A1(n13136), .A2(n13453), .B1(n13647), .B2(n13260), .C1(
        n13099), .C2(n13137), .ZN(P2_U2952) );
  OAI22_X1 U16408 ( .A1(n13100), .A2(n13411), .B1(n13599), .B2(n13390), .ZN(
        n19914) );
  NAND3_X1 U16409 ( .A1(n13102), .A2(n13101), .A3(n15805), .ZN(n13103) );
  AND2_X1 U16410 ( .A1(n13103), .A2(n20864), .ZN(n20861) );
  NOR2_X1 U16411 ( .A1(n19914), .A2(n20861), .ZN(n15772) );
  OR2_X1 U16412 ( .A1(n15772), .A2(n19913), .ZN(n13112) );
  INV_X1 U16413 ( .A(n13112), .ZN(n19922) );
  INV_X1 U16414 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13114) );
  INV_X1 U16415 ( .A(n12563), .ZN(n13229) );
  INV_X1 U16416 ( .A(n13104), .ZN(n15775) );
  AND2_X1 U16417 ( .A1(n15775), .A2(n13459), .ZN(n13402) );
  INV_X1 U16418 ( .A(n13402), .ZN(n13107) );
  NOR3_X1 U16419 ( .A1(n13105), .A2(n13209), .A3(n20142), .ZN(n13106) );
  OAI21_X1 U16420 ( .B1(n13107), .B2(n13106), .A(n13395), .ZN(n13109) );
  NAND2_X1 U16421 ( .A1(n13461), .A2(n13390), .ZN(n13108) );
  OAI211_X1 U16422 ( .C1(n13110), .C2(n13229), .A(n13109), .B(n13108), .ZN(
        n13111) );
  NAND2_X1 U16423 ( .A1(n13111), .A2(n20148), .ZN(n15774) );
  OR2_X1 U16424 ( .A1(n15774), .A2(n13112), .ZN(n13113) );
  OAI21_X1 U16425 ( .B1(n19922), .B2(n13114), .A(n13113), .ZN(P1_U3484) );
  NAND2_X1 U16426 ( .A1(n10710), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13115) );
  NAND4_X1 U16427 ( .A1(n10609), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13115), 
        .A4(n19678), .ZN(n13116) );
  NOR2_X1 U16428 ( .A1(n19153), .A2(n15579), .ZN(n13118) );
  AOI21_X1 U16429 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19153), .A(n13118), .ZN(
        n13119) );
  OAI21_X1 U16430 ( .B1(n19148), .B2(n19894), .A(n13119), .ZN(P2_U2887) );
  INV_X1 U16431 ( .A(n13453), .ZN(n19163) );
  NAND2_X1 U16432 ( .A1(n13121), .A2(n13120), .ZN(n13122) );
  NAND2_X1 U16433 ( .A1(n13123), .A2(n13122), .ZN(n13124) );
  AND2_X1 U16434 ( .A1(n13125), .A2(n10743), .ZN(n13126) );
  INV_X1 U16435 ( .A(n13127), .ZN(n13128) );
  OAI21_X1 U16436 ( .B1(n13130), .B2(n13129), .A(n13128), .ZN(n13667) );
  OAI22_X1 U16437 ( .A1(n19173), .A2(n13667), .B1(n19196), .B2(n13135), .ZN(
        n13132) );
  NOR2_X1 U16438 ( .A1(n19894), .A2(n13667), .ZN(n19217) );
  AOI211_X1 U16439 ( .C1(n19894), .C2(n13667), .A(n19218), .B(n19217), .ZN(
        n13131) );
  AOI211_X1 U16440 ( .C1(n19163), .C2(n19198), .A(n13132), .B(n13131), .ZN(
        n13133) );
  INV_X1 U16441 ( .A(n13133), .ZN(P2_U2919) );
  INV_X1 U16442 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13134) );
  OAI222_X1 U16443 ( .A1(n13135), .A2(n13647), .B1(n13134), .B2(n13137), .C1(
        n13136), .C2(n13453), .ZN(P2_U2967) );
  INV_X1 U16444 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13139) );
  INV_X1 U16445 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16446 ( .A1(n14110), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13375), .ZN(n19174) );
  OAI222_X1 U16447 ( .A1(n13647), .A2(n13139), .B1(n13138), .B2(n13137), .C1(
        n13136), .C2(n19174), .ZN(P2_U2982) );
  OAI21_X1 U16448 ( .B1(n19257), .B2(n15579), .A(n13140), .ZN(n13143) );
  OAI22_X1 U16449 ( .A1(n19264), .A2(n13141), .B1(n16331), .B2(n13667), .ZN(
        n13142) );
  AOI211_X1 U16450 ( .C1(n16338), .C2(n13144), .A(n13143), .B(n13142), .ZN(
        n13147) );
  INV_X1 U16451 ( .A(n15567), .ZN(n13145) );
  MUX2_X1 U16452 ( .A(n15382), .B(n13145), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13146) );
  NAND2_X1 U16453 ( .A1(n13147), .A2(n13146), .ZN(P2_U3046) );
  NAND2_X1 U16454 ( .A1(n13152), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19723) );
  NAND2_X1 U16455 ( .A1(n19874), .A2(n13153), .ZN(n13154) );
  AND3_X1 U16456 ( .A1(n19723), .A2(n19869), .A3(n13154), .ZN(n15622) );
  INV_X1 U16457 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13157) );
  NOR2_X1 U16458 ( .A1(n13192), .A2(n13157), .ZN(n13158) );
  NAND2_X1 U16459 ( .A1(n13159), .A2(n13158), .ZN(n13189) );
  NAND2_X1 U16460 ( .A1(n13162), .A2(n13161), .ZN(n13191) );
  INV_X1 U16461 ( .A(n19871), .ZN(n14997) );
  NOR2_X1 U16462 ( .A1(n10798), .A2(n19153), .ZN(n13165) );
  AOI21_X1 U16463 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19153), .A(n13165), .ZN(
        n13166) );
  OAI21_X1 U16464 ( .B1(n14997), .B2(n19148), .A(n13166), .ZN(P2_U2884) );
  INV_X1 U16465 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20082) );
  INV_X1 U16466 ( .A(n13167), .ZN(n13168) );
  AOI21_X1 U16467 ( .B1(n13205), .B2(n20082), .A(n13168), .ZN(n20092) );
  INV_X1 U16468 ( .A(n20092), .ZN(n13174) );
  INV_X1 U16469 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13173) );
  INV_X1 U16470 ( .A(n13169), .ZN(n13172) );
  OAI21_X1 U16471 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(n20091) );
  OAI222_X1 U16472 ( .A1(n13174), .A2(n14358), .B1(n13173), .B2(n20014), .C1(
        n20091), .C2(n14364), .ZN(P1_U2872) );
  NAND2_X1 U16473 ( .A1(n13175), .A2(n11295), .ZN(n15587) );
  INV_X1 U16474 ( .A(n11371), .ZN(n13176) );
  OAI21_X1 U16475 ( .B1(n15584), .B2(n16349), .A(n13176), .ZN(n13180) );
  NOR2_X1 U16476 ( .A1(n10522), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13177) );
  NOR2_X1 U16477 ( .A1(n13178), .A2(n13177), .ZN(n13179) );
  AOI22_X1 U16478 ( .A1(n15587), .A2(n13180), .B1(n13179), .B2(n11275), .ZN(
        n13185) );
  NAND2_X1 U16479 ( .A1(n16366), .A2(n13181), .ZN(n15590) );
  NOR2_X1 U16480 ( .A1(n13182), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15585) );
  XNOR2_X1 U16481 ( .A(n15585), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13183) );
  NAND2_X1 U16482 ( .A1(n15590), .A2(n13183), .ZN(n13184) );
  OAI211_X1 U16483 ( .C1(n10798), .C2(n15593), .A(n13185), .B(n13184), .ZN(
        n16353) );
  AOI22_X1 U16484 ( .A1(n19871), .A2(n15594), .B1(n19779), .B2(n16353), .ZN(
        n13187) );
  NAND2_X1 U16485 ( .A1(n15599), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13186) );
  OAI21_X1 U16486 ( .B1(n13187), .B2(n15599), .A(n13186), .ZN(P2_U3596) );
  NAND2_X1 U16487 ( .A1(n10743), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13188) );
  NOR2_X1 U16488 ( .A1(n13192), .A2(n14015), .ZN(n13681) );
  XOR2_X1 U16489 ( .A(n13280), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13199)
         );
  INV_X1 U16490 ( .A(n13194), .ZN(n13195) );
  AOI21_X1 U16491 ( .B1(n13196), .B2(n13193), .A(n13195), .ZN(n19121) );
  NOR2_X1 U16492 ( .A1(n19159), .A2(n11177), .ZN(n13197) );
  AOI21_X1 U16493 ( .B1(n19121), .B2(n19159), .A(n13197), .ZN(n13198) );
  OAI21_X1 U16494 ( .B1(n13199), .B2(n19148), .A(n13198), .ZN(P2_U2882) );
  OAI21_X1 U16495 ( .B1(n13201), .B2(n13200), .A(n13356), .ZN(n14273) );
  XNOR2_X1 U16496 ( .A(n14266), .B(n13221), .ZN(n13433) );
  AOI22_X1 U16497 ( .A1(n12863), .A2(n13433), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14362), .ZN(n13202) );
  OAI21_X1 U16498 ( .B1(n14273), .B2(n14364), .A(n13202), .ZN(P1_U2871) );
  NOR2_X1 U16499 ( .A1(n13209), .A2(n20126), .ZN(n13213) );
  OAI22_X1 U16500 ( .A1(n13205), .A2(n13204), .B1(n13203), .B2(n13613), .ZN(
        n13206) );
  NOR2_X1 U16501 ( .A1(n13207), .A2(n13206), .ZN(n13212) );
  OAI21_X1 U16502 ( .B1(n13209), .B2(n13424), .A(n13208), .ZN(n13210) );
  NAND2_X1 U16503 ( .A1(n13211), .A2(n13210), .ZN(n13226) );
  OAI211_X1 U16504 ( .C1(n13214), .C2(n13213), .A(n13212), .B(n13226), .ZN(
        n13407) );
  INV_X1 U16505 ( .A(n13215), .ZN(n13216) );
  OR2_X1 U16506 ( .A1(n13220), .A2(n13216), .ZN(n13217) );
  NOR2_X1 U16507 ( .A1(n13407), .A2(n13217), .ZN(n13218) );
  AND2_X1 U16508 ( .A1(n13218), .A2(n12888), .ZN(n13475) );
  INV_X1 U16509 ( .A(n13475), .ZN(n14626) );
  INV_X1 U16510 ( .A(n14623), .ZN(n13394) );
  AOI22_X1 U16511 ( .A1(n11916), .A2(n14626), .B1(n13394), .B2(n15761), .ZN(
        n15759) );
  INV_X1 U16512 ( .A(n16214), .ZN(n14641) );
  AOI22_X1 U16513 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20082), .B1(n15761), 
        .B2(n15785), .ZN(n13219) );
  OAI21_X1 U16514 ( .B1(n15759), .B2(n14641), .A(n13219), .ZN(n13237) );
  NAND2_X1 U16515 ( .A1(n12563), .A2(n11757), .ZN(n15760) );
  OAI21_X1 U16516 ( .B1(n13221), .B2(n13336), .A(n13220), .ZN(n13222) );
  OAI21_X1 U16517 ( .B1(n15760), .B2(n15805), .A(n13222), .ZN(n13223) );
  NAND2_X1 U16518 ( .A1(n13223), .A2(n20864), .ZN(n13224) );
  NAND2_X1 U16519 ( .A1(n13224), .A2(n13459), .ZN(n13225) );
  NAND2_X1 U16520 ( .A1(n13225), .A2(n13390), .ZN(n13234) );
  NAND2_X1 U16521 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  NAND2_X1 U16522 ( .A1(n13229), .A2(n13228), .ZN(n13397) );
  OAI211_X1 U16523 ( .C1(n13613), .C2(n20126), .A(n13230), .B(n13397), .ZN(
        n13231) );
  INV_X1 U16524 ( .A(n13231), .ZN(n13233) );
  INV_X1 U16525 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19921) );
  NOR2_X1 U16526 ( .A1(n20856), .A2(n20776), .ZN(n13498) );
  NAND2_X1 U16527 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13498), .ZN(n16228) );
  OAI22_X1 U16528 ( .A1(n19913), .A2(n13494), .B1(n19921), .B2(n16228), .ZN(
        n13235) );
  INV_X1 U16529 ( .A(n13235), .ZN(n16219) );
  OAI21_X1 U16530 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20566), .A(n16219), 
        .ZN(n16216) );
  OAI21_X1 U16531 ( .B1(n15760), .B2(n14641), .A(n16216), .ZN(n13236) );
  AOI22_X1 U16532 ( .A1(n13237), .A2(n16216), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13236), .ZN(n13238) );
  INV_X1 U16533 ( .A(n13238), .ZN(P1_U3474) );
  INV_X1 U16534 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14938) );
  AOI22_X1 U16535 ( .A1(n13248), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U16536 ( .B1(n14938), .B2(n13259), .A(n13239), .ZN(P2_U2924) );
  INV_X1 U16537 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16538 ( .A1(n13248), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16539 ( .B1(n14972), .B2(n13259), .A(n13240), .ZN(P2_U2930) );
  INV_X1 U16540 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16541 ( .A1(n13248), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13241) );
  OAI21_X1 U16542 ( .B1(n13242), .B2(n13259), .A(n13241), .ZN(P2_U2929) );
  INV_X1 U16543 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U16544 ( .A1(n13248), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13243) );
  OAI21_X1 U16545 ( .B1(n14967), .B2(n13259), .A(n13243), .ZN(P2_U2928) );
  INV_X1 U16546 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U16547 ( .A1(n13248), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13244) );
  OAI21_X1 U16548 ( .B1(n13245), .B2(n13259), .A(n13244), .ZN(P2_U2926) );
  AOI22_X1 U16549 ( .A1(n13248), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13246) );
  OAI21_X1 U16550 ( .B1(n13247), .B2(n13259), .A(n13246), .ZN(P2_U2921) );
  INV_X1 U16551 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U16552 ( .A1(n13248), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U16553 ( .B1(n14922), .B2(n13259), .A(n13249), .ZN(P2_U2922) );
  INV_X1 U16554 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16555 ( .A1(n21034), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13250) );
  OAI21_X1 U16556 ( .B1(n13251), .B2(n13259), .A(n13250), .ZN(P2_U2931) );
  INV_X1 U16557 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13253) );
  AOI22_X1 U16558 ( .A1(n21034), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13252) );
  OAI21_X1 U16559 ( .B1(n13253), .B2(n13259), .A(n13252), .ZN(P2_U2933) );
  INV_X1 U16560 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U16561 ( .A1(n21034), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13254) );
  OAI21_X1 U16562 ( .B1(n13255), .B2(n13259), .A(n13254), .ZN(P2_U2932) );
  INV_X1 U16563 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U16564 ( .A1(n21034), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13256) );
  OAI21_X1 U16565 ( .B1(n13257), .B2(n13259), .A(n13256), .ZN(P2_U2934) );
  AOI22_X1 U16566 ( .A1(n21034), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13258) );
  OAI21_X1 U16567 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(P2_U2935) );
  AOI21_X1 U16568 ( .B1(n13263), .B2(n13262), .A(n13261), .ZN(n14996) );
  XNOR2_X1 U16569 ( .A(n14996), .B(n19877), .ZN(n13270) );
  XNOR2_X1 U16570 ( .A(n13265), .B(n13264), .ZN(n19889) );
  INV_X1 U16571 ( .A(n19889), .ZN(n13266) );
  NAND2_X1 U16572 ( .A1(n19278), .A2(n13266), .ZN(n13267) );
  OAI21_X1 U16573 ( .B1(n19278), .B2(n13266), .A(n13267), .ZN(n19216) );
  NOR2_X1 U16574 ( .A1(n19216), .A2(n19217), .ZN(n19215) );
  INV_X1 U16575 ( .A(n13267), .ZN(n13268) );
  NOR2_X1 U16576 ( .A1(n19215), .A2(n13268), .ZN(n13269) );
  NOR2_X1 U16577 ( .A1(n13269), .A2(n13270), .ZN(n14995) );
  AOI21_X1 U16578 ( .B1(n13270), .B2(n13269), .A(n14995), .ZN(n13273) );
  AOI22_X1 U16579 ( .A1(n19198), .A2(n16271), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19213), .ZN(n13272) );
  INV_X1 U16580 ( .A(n14996), .ZN(n19879) );
  NAND2_X1 U16581 ( .A1(n19879), .A2(n19214), .ZN(n13271) );
  OAI211_X1 U16582 ( .C1(n13273), .C2(n19218), .A(n13272), .B(n13271), .ZN(
        P2_U2917) );
  XNOR2_X1 U16583 ( .A(n13274), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13436) );
  INV_X1 U16584 ( .A(n14273), .ZN(n13277) );
  INV_X1 U16585 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20946) );
  NOR2_X1 U16586 ( .A1(n20101), .A2(n20946), .ZN(n13432) );
  AOI21_X1 U16587 ( .B1(n20085), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13432), .ZN(n13275) );
  OAI21_X1 U16588 ( .B1(n16023), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13275), .ZN(n13276) );
  AOI21_X1 U16589 ( .B1(n13277), .B2(n16029), .A(n13276), .ZN(n13278) );
  OAI21_X1 U16590 ( .B1(n13436), .B2(n19920), .A(n13278), .ZN(P1_U2998) );
  INV_X1 U16591 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13279) );
  NOR2_X1 U16592 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  OAI211_X1 U16593 ( .C1(n13281), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19156), .B(n13518), .ZN(n13285) );
  AND2_X1 U16594 ( .A1(n13194), .A2(n13282), .ZN(n13283) );
  OR2_X1 U16595 ( .A1(n13283), .A2(n13350), .ZN(n16300) );
  INV_X1 U16596 ( .A(n16300), .ZN(n19105) );
  NAND2_X1 U16597 ( .A1(n19105), .A2(n19159), .ZN(n13284) );
  OAI211_X1 U16598 ( .C1(n19159), .C2(n11182), .A(n13285), .B(n13284), .ZN(
        P2_U2881) );
  INV_X2 U16599 ( .A(n13334), .ZN(n20076) );
  NOR2_X1 U16600 ( .A1(n11773), .A2(n20864), .ZN(n13286) );
  INV_X2 U16601 ( .A(n13330), .ZN(n20075) );
  AOI22_X1 U16602 ( .A1(n20076), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20075), .ZN(n13290) );
  INV_X1 U16603 ( .A(n20104), .ZN(n20105) );
  NAND2_X1 U16604 ( .A1(n20105), .A2(DATAI_2_), .ZN(n13289) );
  NAND2_X1 U16605 ( .A1(n20104), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13288) );
  AND2_X1 U16606 ( .A1(n13289), .A2(n13288), .ZN(n20127) );
  INV_X1 U16607 ( .A(n20127), .ZN(n14391) );
  NAND2_X1 U16608 ( .A1(n20061), .A2(n14391), .ZN(n13311) );
  NAND2_X1 U16609 ( .A1(n13290), .A2(n13311), .ZN(P1_U2939) );
  AOI22_X1 U16610 ( .A1(n20076), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20075), .ZN(n13293) );
  NAND2_X1 U16611 ( .A1(n20105), .A2(DATAI_4_), .ZN(n13292) );
  NAND2_X1 U16612 ( .A1(n20104), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13291) );
  AND2_X1 U16613 ( .A1(n13292), .A2(n13291), .ZN(n20135) );
  INV_X1 U16614 ( .A(n20135), .ZN(n15947) );
  NAND2_X1 U16615 ( .A1(n20061), .A2(n15947), .ZN(n13326) );
  NAND2_X1 U16616 ( .A1(n13293), .A2(n13326), .ZN(P1_U2941) );
  AOI22_X1 U16617 ( .A1(n20076), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20075), .ZN(n13296) );
  NAND2_X1 U16618 ( .A1(n20105), .A2(DATAI_5_), .ZN(n13295) );
  NAND2_X1 U16619 ( .A1(n20104), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13294) );
  AND2_X1 U16620 ( .A1(n13295), .A2(n13294), .ZN(n20139) );
  INV_X1 U16621 ( .A(n20139), .ZN(n14385) );
  NAND2_X1 U16622 ( .A1(n20061), .A2(n14385), .ZN(n13309) );
  NAND2_X1 U16623 ( .A1(n13296), .A2(n13309), .ZN(P1_U2942) );
  AOI22_X1 U16624 ( .A1(n20076), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20075), .ZN(n13299) );
  NAND2_X1 U16625 ( .A1(n20105), .A2(DATAI_6_), .ZN(n13298) );
  NAND2_X1 U16626 ( .A1(n20104), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13297) );
  AND2_X1 U16627 ( .A1(n13298), .A2(n13297), .ZN(n20143) );
  INV_X1 U16628 ( .A(n20143), .ZN(n14381) );
  NAND2_X1 U16629 ( .A1(n20061), .A2(n14381), .ZN(n13322) );
  NAND2_X1 U16630 ( .A1(n13299), .A2(n13322), .ZN(P1_U2943) );
  AOI22_X1 U16631 ( .A1(n20076), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20075), .ZN(n13302) );
  NAND2_X1 U16632 ( .A1(n20105), .A2(DATAI_7_), .ZN(n13301) );
  NAND2_X1 U16633 ( .A1(n20104), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13300) );
  AND2_X1 U16634 ( .A1(n13301), .A2(n13300), .ZN(n20151) );
  INV_X1 U16635 ( .A(n20151), .ZN(n15943) );
  NAND2_X1 U16636 ( .A1(n20061), .A2(n15943), .ZN(n13320) );
  NAND2_X1 U16637 ( .A1(n13302), .A2(n13320), .ZN(P1_U2944) );
  AOI22_X1 U16638 ( .A1(n20076), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20075), .ZN(n13305) );
  NAND2_X1 U16639 ( .A1(n20105), .A2(DATAI_3_), .ZN(n13304) );
  NAND2_X1 U16640 ( .A1(n20104), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13303) );
  AND2_X1 U16641 ( .A1(n13304), .A2(n13303), .ZN(n20131) );
  INV_X1 U16642 ( .A(n20131), .ZN(n14388) );
  NAND2_X1 U16643 ( .A1(n20061), .A2(n14388), .ZN(n13313) );
  NAND2_X1 U16644 ( .A1(n13305), .A2(n13313), .ZN(P1_U2940) );
  AOI22_X1 U16645 ( .A1(n20076), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20075), .ZN(n13308) );
  NAND2_X1 U16646 ( .A1(n20105), .A2(DATAI_1_), .ZN(n13307) );
  NAND2_X1 U16647 ( .A1(n20104), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13306) );
  AND2_X1 U16648 ( .A1(n13307), .A2(n13306), .ZN(n20123) );
  INV_X1 U16649 ( .A(n20123), .ZN(n14395) );
  NAND2_X1 U16650 ( .A1(n20061), .A2(n14395), .ZN(n13318) );
  NAND2_X1 U16651 ( .A1(n13308), .A2(n13318), .ZN(P1_U2953) );
  AOI22_X1 U16652 ( .A1(n20076), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20075), .ZN(n13310) );
  NAND2_X1 U16653 ( .A1(n13310), .A2(n13309), .ZN(P1_U2957) );
  AOI22_X1 U16654 ( .A1(n20076), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20075), .ZN(n13312) );
  NAND2_X1 U16655 ( .A1(n13312), .A2(n13311), .ZN(P1_U2954) );
  AOI22_X1 U16656 ( .A1(n20076), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20075), .ZN(n13314) );
  NAND2_X1 U16657 ( .A1(n13314), .A2(n13313), .ZN(P1_U2955) );
  AOI22_X1 U16658 ( .A1(n20076), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20075), .ZN(n13317) );
  NAND2_X1 U16659 ( .A1(n20105), .A2(DATAI_0_), .ZN(n13316) );
  NAND2_X1 U16660 ( .A1(n20104), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13315) );
  AND2_X1 U16661 ( .A1(n13316), .A2(n13315), .ZN(n20115) );
  INV_X1 U16662 ( .A(n20115), .ZN(n14400) );
  NAND2_X1 U16663 ( .A1(n20061), .A2(n14400), .ZN(n13324) );
  NAND2_X1 U16664 ( .A1(n13317), .A2(n13324), .ZN(P1_U2952) );
  AOI22_X1 U16665 ( .A1(n20076), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20075), .ZN(n13319) );
  NAND2_X1 U16666 ( .A1(n13319), .A2(n13318), .ZN(P1_U2938) );
  AOI22_X1 U16667 ( .A1(n20076), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20075), .ZN(n13321) );
  NAND2_X1 U16668 ( .A1(n13321), .A2(n13320), .ZN(P1_U2959) );
  AOI22_X1 U16669 ( .A1(n20076), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20075), .ZN(n13323) );
  NAND2_X1 U16670 ( .A1(n13323), .A2(n13322), .ZN(P1_U2958) );
  AOI22_X1 U16671 ( .A1(n20076), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20075), .ZN(n13325) );
  NAND2_X1 U16672 ( .A1(n13325), .A2(n13324), .ZN(P1_U2937) );
  AOI22_X1 U16673 ( .A1(n20076), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20075), .ZN(n13327) );
  NAND2_X1 U16674 ( .A1(n13327), .A2(n13326), .ZN(P1_U2956) );
  INV_X1 U16675 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13333) );
  INV_X1 U16676 ( .A(n20061), .ZN(n13332) );
  INV_X1 U16677 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13328) );
  NOR2_X1 U16678 ( .A1(n20105), .A2(n13328), .ZN(n13329) );
  AOI21_X1 U16679 ( .B1(DATAI_15_), .B2(n20105), .A(n13329), .ZN(n14403) );
  INV_X1 U16680 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13331) );
  OAI222_X1 U16681 ( .A1(n13334), .A2(n13333), .B1(n13332), .B2(n14403), .C1(
        n13331), .C2(n13330), .ZN(P1_U2967) );
  NAND2_X1 U16682 ( .A1(n13390), .A2(n13399), .ZN(n13335) );
  OAI21_X1 U16683 ( .B1(n15760), .B2(n13335), .A(n13334), .ZN(n13337) );
  NAND2_X1 U16684 ( .A1(n20015), .A2(n20109), .ZN(n13566) );
  INV_X1 U16685 ( .A(n13498), .ZN(n16223) );
  NOR2_X4 U16686 ( .A1(n20015), .A2(n20865), .ZN(n20043) );
  AOI22_X1 U16687 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13338) );
  OAI21_X1 U16688 ( .B1(n12450), .B2(n13566), .A(n13338), .ZN(P1_U2910) );
  INV_X1 U16689 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U16690 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13339) );
  OAI21_X1 U16691 ( .B1(n13340), .B2(n13566), .A(n13339), .ZN(P1_U2909) );
  AOI22_X1 U16692 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13341) );
  OAI21_X1 U16693 ( .B1(n12402), .B2(n13566), .A(n13341), .ZN(P1_U2912) );
  INV_X1 U16694 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U16695 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13342) );
  OAI21_X1 U16696 ( .B1(n13343), .B2(n13566), .A(n13342), .ZN(P1_U2911) );
  INV_X1 U16697 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U16698 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13344) );
  OAI21_X1 U16699 ( .B1(n13345), .B2(n13566), .A(n13344), .ZN(P1_U2906) );
  INV_X1 U16700 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U16701 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13346) );
  OAI21_X1 U16702 ( .B1(n13347), .B2(n13566), .A(n13346), .ZN(P1_U2907) );
  AOI22_X1 U16703 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13348) );
  OAI21_X1 U16704 ( .B1(n12500), .B2(n13566), .A(n13348), .ZN(P1_U2908) );
  XOR2_X1 U16705 ( .A(n13518), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13353)
         );
  OR2_X1 U16706 ( .A1(n13350), .A2(n13349), .ZN(n13351) );
  NAND2_X1 U16707 ( .A1(n13704), .A2(n13351), .ZN(n19091) );
  MUX2_X1 U16708 ( .A(n19091), .B(n11186), .S(n19153), .Z(n13352) );
  OAI21_X1 U16709 ( .B1(n13353), .B2(n19148), .A(n13352), .ZN(P2_U2880) );
  INV_X1 U16710 ( .A(n13354), .ZN(n13355) );
  AOI21_X1 U16711 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n20001) );
  INV_X1 U16712 ( .A(n20001), .ZN(n13426) );
  NOR2_X1 U16713 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  OR2_X1 U16714 ( .A1(n13513), .A2(n13360), .ZN(n20004) );
  INV_X1 U16715 ( .A(n20004), .ZN(n13361) );
  AOI22_X1 U16716 ( .A1(n12863), .A2(n13361), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14362), .ZN(n13362) );
  OAI21_X1 U16717 ( .B1(n13426), .B2(n14364), .A(n13362), .ZN(P1_U2870) );
  XNOR2_X1 U16718 ( .A(n13364), .B(n13363), .ZN(n13423) );
  INV_X1 U16719 ( .A(n19988), .ZN(n13366) );
  AOI22_X1 U16720 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13365) );
  OAI21_X1 U16721 ( .B1(n16023), .B2(n13366), .A(n13365), .ZN(n13367) );
  AOI21_X1 U16722 ( .B1(n20001), .B2(n16029), .A(n13367), .ZN(n13368) );
  OAI21_X1 U16723 ( .B1(n19920), .B2(n13423), .A(n13368), .ZN(P1_U2997) );
  NAND2_X1 U16724 ( .A1(n19871), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19721) );
  NAND3_X1 U16725 ( .A1(n19891), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15614) );
  OAI21_X1 U16726 ( .B1(n19721), .B2(n13377), .A(n15614), .ZN(n13374) );
  NOR2_X1 U16727 ( .A1(n19900), .A2(n15614), .ZN(n19682) );
  INV_X1 U16728 ( .A(n19682), .ZN(n13371) );
  AND2_X1 U16729 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13371), .ZN(n13369) );
  NAND2_X1 U16730 ( .A1(n13370), .A2(n13369), .ZN(n13379) );
  NAND2_X1 U16731 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13371), .ZN(n13372) );
  AND3_X1 U16732 ( .A1(n13379), .A2(n19726), .A3(n13372), .ZN(n13373) );
  NAND2_X1 U16733 ( .A1(n13374), .A2(n13373), .ZN(n19671) );
  INV_X1 U16734 ( .A(n19671), .ZN(n19663) );
  AOI22_X1 U16735 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19306), .ZN(n19692) );
  INV_X1 U16736 ( .A(n19692), .ZN(n19732) );
  AOI22_X1 U16737 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19306), .ZN(n19735) );
  AOI22_X1 U16738 ( .A1(n19670), .A2(n19732), .B1(n19707), .B2(n19689), .ZN(
        n13383) );
  OAI21_X1 U16739 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n15614), .A(n19676), 
        .ZN(n13378) );
  AOI22_X1 U16740 ( .A1(n19669), .A2(n13380), .B1(n13381), .B2(n19682), .ZN(
        n13382) );
  OAI211_X1 U16741 ( .C1(n19663), .C2(n13948), .A(n13383), .B(n13382), .ZN(
        P2_U3153) );
  NAND2_X1 U16742 ( .A1(n11757), .A2(n15805), .ZN(n13385) );
  NAND2_X1 U16743 ( .A1(n13385), .A2(n13384), .ZN(n13393) );
  INV_X1 U16744 ( .A(n13386), .ZN(n13388) );
  OAI211_X1 U16745 ( .C1(n13389), .C2(n13388), .A(n20109), .B(n13387), .ZN(
        n13391) );
  NAND3_X1 U16746 ( .A1(n13395), .A2(n13394), .A3(n11757), .ZN(n13396) );
  NAND3_X1 U16747 ( .A1(n13398), .A2(n13397), .A3(n13396), .ZN(n13400) );
  INV_X1 U16748 ( .A(n13413), .ZN(n13403) );
  OAI211_X1 U16749 ( .C1(n13412), .C2(n13403), .A(n13402), .B(n13401), .ZN(
        n13404) );
  INV_X1 U16750 ( .A(n13405), .ZN(n13406) );
  OR2_X1 U16751 ( .A1(n13407), .A2(n13406), .ZN(n13408) );
  NOR2_X1 U16752 ( .A1(n13420), .A2(n12626), .ZN(n14528) );
  NOR2_X1 U16753 ( .A1(n12840), .A2(n13416), .ZN(n13428) );
  AOI21_X1 U16754 ( .B1(n15810), .B2(n20082), .A(n13428), .ZN(n14610) );
  OAI21_X1 U16755 ( .B1(n14613), .B2(n14528), .A(n14610), .ZN(n16172) );
  INV_X1 U16756 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19993) );
  NOR2_X1 U16757 ( .A1(n20101), .A2(n19993), .ZN(n13419) );
  NOR2_X1 U16758 ( .A1(n20082), .A2(n12626), .ZN(n13409) );
  OAI21_X1 U16759 ( .B1(n20082), .B2(n12626), .A(n13420), .ZN(n14529) );
  INV_X1 U16760 ( .A(n14529), .ZN(n13540) );
  AOI21_X1 U16761 ( .B1(n13409), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13540), .ZN(n13417) );
  NAND2_X1 U16762 ( .A1(n13411), .A2(n13410), .ZN(n15780) );
  NAND2_X1 U16763 ( .A1(n13413), .A2(n13412), .ZN(n13414) );
  NAND2_X1 U16764 ( .A1(n15780), .A2(n13414), .ZN(n13415) );
  OAI22_X1 U16765 ( .A1(n13417), .A2(n15814), .B1(n16159), .B2(n20004), .ZN(
        n13418) );
  AOI211_X1 U16766 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n16172), .A(
        n13419), .B(n13418), .ZN(n13422) );
  NOR2_X1 U16767 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20098), .ZN(
        n13427) );
  NAND3_X1 U16768 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16171), .A3(
        n13420), .ZN(n13421) );
  OAI211_X1 U16769 ( .C1(n16204), .C2(n13423), .A(n13422), .B(n13421), .ZN(
        P1_U3029) );
  NOR2_X1 U16770 ( .A1(n13424), .A2(n13810), .ZN(n13425) );
  OR2_X2 U16771 ( .A1(n15946), .A2(n13425), .ZN(n14411) );
  INV_X1 U16772 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20040) );
  OAI222_X1 U16773 ( .A1(n14411), .A2(n13426), .B1(n14405), .B2(n20040), .C1(
        n14404), .C2(n20127), .ZN(P1_U2902) );
  INV_X1 U16774 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20047) );
  OAI222_X1 U16775 ( .A1(n14411), .A2(n20091), .B1(n14405), .B2(n20047), .C1(
        n14404), .C2(n20115), .ZN(P1_U2904) );
  NOR2_X1 U16776 ( .A1(n14600), .A2(n13427), .ZN(n13430) );
  INV_X1 U16777 ( .A(n15810), .ZN(n14527) );
  NAND2_X1 U16778 ( .A1(n15814), .A2(n14527), .ZN(n20096) );
  AOI21_X1 U16779 ( .B1(n20082), .B2(n20096), .A(n13428), .ZN(n13429) );
  INV_X1 U16780 ( .A(n13429), .ZN(n20097) );
  MUX2_X1 U16781 ( .A(n13430), .B(n20097), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13431) );
  INV_X1 U16782 ( .A(n13431), .ZN(n13435) );
  AOI21_X1 U16783 ( .B1(n20093), .B2(n13433), .A(n13432), .ZN(n13434) );
  OAI211_X1 U16784 ( .C1(n13436), .C2(n16204), .A(n13435), .B(n13434), .ZN(
        P1_U3030) );
  NAND2_X1 U16785 ( .A1(n19881), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19582) );
  INV_X1 U16786 ( .A(n19582), .ZN(n19577) );
  NAND2_X1 U16787 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19577), .ZN(
        n13445) );
  OAI21_X1 U16788 ( .B1(n19721), .B2(n13444), .A(n13445), .ZN(n13443) );
  INV_X1 U16789 ( .A(n19375), .ZN(n13437) );
  NAND2_X1 U16790 ( .A1(n13437), .A2(n19577), .ZN(n13438) );
  INV_X1 U16791 ( .A(n13438), .ZN(n19621) );
  AND2_X1 U16792 ( .A1(n13438), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U16793 ( .A1(n13440), .A2(n13439), .ZN(n13447) );
  OAI211_X1 U16794 ( .C1(n19621), .C2(n19678), .A(n13447), .B(n19726), .ZN(
        n13441) );
  INV_X1 U16795 ( .A(n13441), .ZN(n13442) );
  NAND2_X1 U16796 ( .A1(n13443), .A2(n13442), .ZN(n19617) );
  INV_X1 U16797 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U16798 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19306), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19307), .ZN(n19634) );
  INV_X1 U16799 ( .A(n19651), .ZN(n19637) );
  AOI22_X1 U16800 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19306), .ZN(n19740) );
  INV_X1 U16801 ( .A(n19740), .ZN(n19631) );
  AOI22_X1 U16802 ( .A1(n19623), .A2(n19737), .B1(n19637), .B2(n19631), .ZN(
        n13451) );
  OAI21_X1 U16803 ( .B1(n13445), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19676), 
        .ZN(n13446) );
  AND2_X1 U16804 ( .A1(n13447), .A2(n13446), .ZN(n19622) );
  NOR2_X2 U16805 ( .A1(n10713), .A2(n19308), .ZN(n19736) );
  AOI22_X1 U16806 ( .A1(n19622), .A2(n13449), .B1(n19621), .B2(n19736), .ZN(
        n13450) );
  OAI211_X1 U16807 ( .C1(n19627), .C2(n13452), .A(n13451), .B(n13450), .ZN(
        P2_U3138) );
  INV_X1 U16808 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U16809 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19306), .ZN(n19731) );
  AOI22_X1 U16810 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19306), .ZN(n19507) );
  INV_X1 U16811 ( .A(n19507), .ZN(n19728) );
  AOI22_X1 U16812 ( .A1(n19623), .A2(n19652), .B1(n19637), .B2(n19728), .ZN(
        n13456) );
  NOR2_X2 U16813 ( .A1(n10722), .A2(n19308), .ZN(n19718) );
  AOI22_X1 U16814 ( .A1(n19622), .A2(n13454), .B1(n19718), .B2(n19621), .ZN(
        n13455) );
  OAI211_X1 U16815 ( .C1(n19627), .C2(n13457), .A(n13456), .B(n13455), .ZN(
        P2_U3136) );
  NOR2_X1 U16816 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20776), .ZN(n13496) );
  INV_X1 U16817 ( .A(n20564), .ZN(n20112) );
  XNOR2_X1 U16818 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13465) );
  INV_X1 U16819 ( .A(n13459), .ZN(n13460) );
  OR2_X1 U16820 ( .A1(n13461), .A2(n13460), .ZN(n13471) );
  XNOR2_X1 U16821 ( .A(n14627), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13462) );
  NAND2_X1 U16822 ( .A1(n13471), .A2(n13462), .ZN(n13464) );
  INV_X1 U16823 ( .A(n13462), .ZN(n14634) );
  NAND3_X1 U16824 ( .A1(n13475), .A2(n13474), .A3(n14634), .ZN(n13463) );
  OAI211_X1 U16825 ( .C1(n15760), .C2(n13465), .A(n13464), .B(n13463), .ZN(
        n13466) );
  AOI21_X1 U16826 ( .B1(n20112), .B2(n14626), .A(n13466), .ZN(n14636) );
  INV_X1 U16827 ( .A(n14636), .ZN(n13467) );
  INV_X1 U16828 ( .A(n13494), .ZN(n15763) );
  MUX2_X1 U16829 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13467), .S(
        n15763), .Z(n15769) );
  AOI22_X1 U16830 ( .A1(n13496), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15769), .B2(n20776), .ZN(n13487) );
  MUX2_X1 U16831 ( .A(n11634), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14627), .Z(n13469) );
  NOR2_X1 U16832 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  NAND2_X1 U16833 ( .A1(n13471), .A2(n13470), .ZN(n13482) );
  NAND2_X1 U16834 ( .A1(n14627), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13472) );
  NAND2_X1 U16835 ( .A1(n13472), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13473) );
  NAND2_X1 U16836 ( .A1(n11783), .A2(n13473), .ZN(n14638) );
  NAND3_X1 U16837 ( .A1(n13475), .A2(n13474), .A3(n14638), .ZN(n13481) );
  INV_X1 U16838 ( .A(n13476), .ZN(n13479) );
  NAND2_X1 U16839 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U16840 ( .A1(n11948), .A2(n13477), .ZN(n13478) );
  NAND3_X1 U16841 ( .A1(n9801), .A2(n13479), .A3(n13478), .ZN(n13480) );
  NAND3_X1 U16842 ( .A1(n13482), .A2(n13481), .A3(n13480), .ZN(n13483) );
  AOI21_X1 U16843 ( .B1(n20415), .B2(n14626), .A(n13483), .ZN(n14642) );
  NAND2_X1 U16844 ( .A1(n14642), .A2(n15763), .ZN(n13485) );
  NAND2_X1 U16845 ( .A1(n13494), .A2(n11948), .ZN(n13484) );
  AOI22_X1 U16846 ( .A1(n13496), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20776), .B2(n15758), .ZN(n13486) );
  NOR2_X1 U16847 ( .A1(n13487), .A2(n13486), .ZN(n15778) );
  INV_X1 U16848 ( .A(n13489), .ZN(n13490) );
  NAND2_X1 U16849 ( .A1(n15778), .A2(n13490), .ZN(n13499) );
  INV_X1 U16850 ( .A(n20270), .ZN(n20563) );
  NOR2_X1 U16851 ( .A1(n13491), .A2(n20563), .ZN(n13492) );
  XNOR2_X1 U16852 ( .A(n13492), .B(n16217), .ZN(n16215) );
  AOI21_X1 U16853 ( .B1(n16215), .B2(n16213), .A(n13494), .ZN(n13493) );
  AOI211_X1 U16854 ( .C1(n13494), .C2(n16217), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13493), .ZN(n13495) );
  AOI21_X1 U16855 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13496), .A(
        n13495), .ZN(n15776) );
  AND3_X1 U16856 ( .A1(n13499), .A2(n15776), .A3(n19921), .ZN(n13497) );
  AND3_X1 U16857 ( .A1(n13499), .A2(n15776), .A3(n13498), .ZN(n15788) );
  INV_X1 U16858 ( .A(n11916), .ZN(n13500) );
  AND2_X1 U16859 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20566), .ZN(n14621) );
  OAI22_X1 U16860 ( .A1(n12741), .A2(n20635), .B1(n13500), .B2(n14621), .ZN(
        n13501) );
  OAI21_X1 U16861 ( .B1(n15788), .B2(n13501), .A(n20102), .ZN(n13502) );
  OAI21_X1 U16862 ( .B1(n20102), .B2(n20601), .A(n13502), .ZN(P1_U3478) );
  NOR2_X1 U16863 ( .A1(n20564), .A2(n14621), .ZN(n13507) );
  OR2_X1 U16864 ( .A1(n9615), .A2(n20635), .ZN(n13504) );
  NAND2_X1 U16865 ( .A1(n20377), .A2(n20857), .ZN(n20162) );
  NAND2_X1 U16866 ( .A1(n13504), .A2(n20162), .ZN(n20713) );
  INV_X1 U16867 ( .A(n9615), .ZN(n13578) );
  NOR3_X1 U16868 ( .A1(n13578), .A2(n20857), .A3(n20635), .ZN(n13505) );
  MUX2_X1 U16869 ( .A(n20713), .B(n13505), .S(n12749), .Z(n13506) );
  OAI21_X1 U16870 ( .B1(n13507), .B2(n13506), .A(n20102), .ZN(n13508) );
  OAI21_X1 U16871 ( .B1(n20102), .B2(n20560), .A(n13508), .ZN(P1_U3476) );
  OAI21_X1 U16872 ( .B1(n13511), .B2(n13510), .A(n13509), .ZN(n13625) );
  INV_X1 U16873 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13514) );
  OAI21_X1 U16874 ( .B1(n13513), .B2(n13512), .A(n13533), .ZN(n13542) );
  OAI222_X1 U16875 ( .A1(n13625), .A2(n14364), .B1(n13514), .B2(n20014), .C1(
        n13542), .C2(n14358), .ZN(P1_U2869) );
  NAND2_X1 U16876 ( .A1(n13515), .A2(n13516), .ZN(n13517) );
  NAND2_X1 U16877 ( .A1(n15486), .A2(n13517), .ZN(n19075) );
  NAND2_X1 U16878 ( .A1(n19146), .A2(n13519), .ZN(n13520) );
  INV_X1 U16879 ( .A(n13520), .ZN(n19147) );
  INV_X1 U16880 ( .A(n13521), .ZN(n13522) );
  OAI211_X1 U16881 ( .C1(n19147), .C2(n13522), .A(n19156), .B(n13830), .ZN(
        n13524) );
  NAND2_X1 U16882 ( .A1(n19153), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13523) );
  OAI211_X1 U16883 ( .C1(n19075), .C2(n19153), .A(n13524), .B(n13523), .ZN(
        P2_U2878) );
  XNOR2_X1 U16884 ( .A(n13525), .B(n13526), .ZN(n13546) );
  INV_X1 U16885 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13620) );
  NOR2_X1 U16886 ( .A1(n20101), .A2(n13620), .ZN(n13543) );
  AOI21_X1 U16887 ( .B1(n20085), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13543), .ZN(n13529) );
  INV_X1 U16888 ( .A(n13618), .ZN(n13527) );
  NAND2_X1 U16889 ( .A1(n16027), .A2(n13527), .ZN(n13528) );
  OAI211_X1 U16890 ( .C1(n13625), .C2(n20106), .A(n13529), .B(n13528), .ZN(
        n13530) );
  INV_X1 U16891 ( .A(n13530), .ZN(n13531) );
  OAI21_X1 U16892 ( .B1(n13546), .B2(n19920), .A(n13531), .ZN(P1_U2996) );
  NAND2_X1 U16893 ( .A1(n13533), .A2(n13532), .ZN(n13534) );
  NAND2_X1 U16894 ( .A1(n13572), .A2(n13534), .ZN(n14261) );
  INV_X1 U16895 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13538) );
  AND2_X1 U16896 ( .A1(n13509), .A2(n13535), .ZN(n13537) );
  OR2_X1 U16897 ( .A1(n13537), .A2(n13536), .ZN(n14264) );
  OAI222_X1 U16898 ( .A1(n14261), .A2(n14358), .B1(n20014), .B2(n13538), .C1(
        n14264), .C2(n14364), .ZN(P1_U2868) );
  AOI21_X1 U16899 ( .B1(n16063), .B2(n13540), .A(n16172), .ZN(n13539) );
  INV_X1 U16900 ( .A(n13539), .ZN(n13550) );
  AOI21_X1 U16901 ( .B1(n14528), .B2(n16171), .A(n16063), .ZN(n16125) );
  NOR2_X1 U16902 ( .A1(n13540), .A2(n16125), .ZN(n16201) );
  AOI22_X1 U16903 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13550), .B1(
        n16201), .B2(n13541), .ZN(n13545) );
  INV_X1 U16904 ( .A(n13542), .ZN(n13616) );
  AOI21_X1 U16905 ( .B1(n20093), .B2(n13616), .A(n13543), .ZN(n13544) );
  OAI211_X1 U16906 ( .C1(n16204), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        P1_U3028) );
  XNOR2_X1 U16907 ( .A(n13547), .B(n13548), .ZN(n13598) );
  NOR2_X1 U16908 ( .A1(n20101), .A2(n20799), .ZN(n13592) );
  NOR2_X1 U16909 ( .A1(n16159), .A2(n14261), .ZN(n13549) );
  AOI211_X1 U16910 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13550), .A(
        n13592), .B(n13549), .ZN(n13552) );
  NAND2_X1 U16911 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16174) );
  OAI211_X1 U16912 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n16201), .B(n16174), .ZN(n13551) );
  OAI211_X1 U16913 ( .C1(n13598), .C2(n16204), .A(n13552), .B(n13551), .ZN(
        P1_U3027) );
  INV_X1 U16914 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U16915 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13553) );
  OAI21_X1 U16916 ( .B1(n13554), .B2(n13566), .A(n13553), .ZN(P1_U2920) );
  AOI22_X1 U16917 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16918 ( .B1(n12234), .B2(n13566), .A(n13555), .ZN(P1_U2919) );
  INV_X1 U16919 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13557) );
  AOI22_X1 U16920 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13556) );
  OAI21_X1 U16921 ( .B1(n13557), .B2(n13566), .A(n13556), .ZN(P1_U2918) );
  INV_X1 U16922 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U16923 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13558) );
  OAI21_X1 U16924 ( .B1(n13559), .B2(n13566), .A(n13558), .ZN(P1_U2915) );
  INV_X1 U16925 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U16926 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U16927 ( .B1(n13561), .B2(n13566), .A(n13560), .ZN(P1_U2913) );
  INV_X1 U16928 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U16929 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13562) );
  OAI21_X1 U16930 ( .B1(n13563), .B2(n13566), .A(n13562), .ZN(P1_U2917) );
  INV_X1 U16931 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U16932 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13564) );
  OAI21_X1 U16933 ( .B1(n20873), .B2(n13566), .A(n13564), .ZN(P1_U2914) );
  INV_X1 U16934 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U16935 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13565) );
  OAI21_X1 U16936 ( .B1(n13567), .B2(n13566), .A(n13565), .ZN(P1_U2916) );
  INV_X1 U16937 ( .A(n13568), .ZN(n13570) );
  INV_X1 U16938 ( .A(n13536), .ZN(n13569) );
  AOI21_X1 U16939 ( .B1(n13570), .B2(n13569), .A(n9682), .ZN(n16030) );
  INV_X1 U16940 ( .A(n16030), .ZN(n13607) );
  NAND2_X1 U16941 ( .A1(n13572), .A2(n13571), .ZN(n13573) );
  AND2_X1 U16942 ( .A1(n16184), .A2(n13573), .ZN(n16209) );
  AOI22_X1 U16943 ( .A1(n12863), .A2(n16209), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14362), .ZN(n13574) );
  OAI21_X1 U16944 ( .B1(n13607), .B2(n14364), .A(n13574), .ZN(P1_U2867) );
  MUX2_X1 U16945 ( .A(n20385), .B(n20633), .S(n13578), .Z(n13579) );
  NOR3_X1 U16946 ( .A1(n20528), .A2(n13579), .A3(n20857), .ZN(n13580) );
  AOI211_X1 U16947 ( .C1(n12759), .C2(n20857), .A(n20635), .B(n13580), .ZN(
        n13583) );
  INV_X1 U16948 ( .A(n20415), .ZN(n13581) );
  NOR2_X1 U16949 ( .A1(n13581), .A2(n14621), .ZN(n13582) );
  OAI21_X1 U16950 ( .B1(n13583), .B2(n13582), .A(n20102), .ZN(n13584) );
  OAI21_X1 U16951 ( .B1(n20102), .B2(n20559), .A(n13584), .ZN(P1_U3475) );
  NOR2_X1 U16952 ( .A1(n13830), .A2(n19142), .ZN(n13585) );
  NAND2_X1 U16953 ( .A1(n13585), .A2(n13826), .ZN(n19137) );
  OAI211_X1 U16954 ( .C1(n13585), .C2(n13826), .A(n19137), .B(n19156), .ZN(
        n13590) );
  OR2_X1 U16955 ( .A1(n15485), .A2(n13586), .ZN(n13587) );
  NAND2_X1 U16956 ( .A1(n14820), .A2(n13587), .ZN(n19055) );
  INV_X1 U16957 ( .A(n19055), .ZN(n13588) );
  NAND2_X1 U16958 ( .A1(n13588), .A2(n19159), .ZN(n13589) );
  OAI211_X1 U16959 ( .C1(n19159), .C2(n13591), .A(n13590), .B(n13589), .ZN(
        P2_U2876) );
  AOI21_X1 U16960 ( .B1(n20085), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13592), .ZN(n13595) );
  INV_X1 U16961 ( .A(n14251), .ZN(n13593) );
  NAND2_X1 U16962 ( .A1(n16027), .A2(n13593), .ZN(n13594) );
  OAI211_X1 U16963 ( .C1(n14264), .C2(n20106), .A(n13595), .B(n13594), .ZN(
        n13596) );
  INV_X1 U16964 ( .A(n13596), .ZN(n13597) );
  OAI21_X1 U16965 ( .B1(n13598), .B2(n19920), .A(n13597), .ZN(P1_U2995) );
  INV_X1 U16966 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U16967 ( .A1(n14411), .A2(n14273), .B1(n14405), .B2(n20042), .C1(
        n14404), .C2(n20123), .ZN(P1_U2903) );
  INV_X1 U16968 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20036) );
  OAI222_X1 U16969 ( .A1(n14411), .A2(n14264), .B1(n14405), .B2(n20036), .C1(
        n14404), .C2(n20135), .ZN(P1_U2900) );
  INV_X1 U16970 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20038) );
  OAI222_X1 U16971 ( .A1(n14411), .A2(n13625), .B1(n14405), .B2(n20038), .C1(
        n14404), .C2(n20131), .ZN(P1_U2901) );
  INV_X1 U16972 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20034) );
  OAI222_X1 U16973 ( .A1(n14411), .A2(n13607), .B1(n14405), .B2(n20034), .C1(
        n14404), .C2(n20139), .ZN(P1_U2899) );
  NAND2_X1 U16974 ( .A1(n20862), .A2(n13599), .ZN(n13600) );
  OAI21_X1 U16975 ( .B1(n19994), .B2(n14256), .A(n15872), .ZN(n19961) );
  NAND2_X1 U16976 ( .A1(n19962), .A2(n14256), .ZN(n19981) );
  OAI22_X1 U16977 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19981), .B1(n16026), 
        .B2(n19974), .ZN(n13605) );
  INV_X1 U16978 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16034) );
  AOI22_X1 U16979 ( .A1(n19977), .A2(n16209), .B1(n19963), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13603) );
  OAI211_X1 U16980 ( .C1(n19949), .C2(n16034), .A(n13603), .B(n20101), .ZN(
        n13604) );
  AOI211_X1 U16981 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n19961), .A(n13605), .B(
        n13604), .ZN(n13606) );
  OAI21_X1 U16982 ( .B1(n13607), .B2(n19990), .A(n13606), .ZN(P1_U2835) );
  OR2_X1 U16983 ( .A1(n9682), .A2(n13609), .ZN(n13610) );
  AND2_X1 U16984 ( .A1(n13608), .A2(n13610), .ZN(n19984) );
  INV_X1 U16985 ( .A(n19984), .ZN(n13612) );
  XNOR2_X1 U16986 ( .A(n16184), .B(n16186), .ZN(n19978) );
  AOI22_X1 U16987 ( .A1(n19978), .A2(n12863), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14362), .ZN(n13611) );
  OAI21_X1 U16988 ( .B1(n13612), .B2(n14364), .A(n13611), .ZN(P1_U2866) );
  OAI222_X1 U16989 ( .A1(n14411), .A2(n13612), .B1(n14405), .B2(n12027), .C1(
        n14404), .C2(n20143), .ZN(P1_U2898) );
  NOR2_X1 U16990 ( .A1(n13614), .A2(n13613), .ZN(n19991) );
  INV_X1 U16991 ( .A(n15872), .ZN(n15926) );
  NAND2_X1 U16992 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13615) );
  NAND2_X1 U16993 ( .A1(n19994), .A2(n15872), .ZN(n15924) );
  OAI21_X1 U16994 ( .B1(n15926), .B2(n13615), .A(n15924), .ZN(n19992) );
  AOI22_X1 U16995 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n19989), .B1(
        n19977), .B2(n13616), .ZN(n13617) );
  OAI21_X1 U16996 ( .B1(n19974), .B2(n13618), .A(n13617), .ZN(n13619) );
  AOI21_X1 U16997 ( .B1(n19963), .B2(P1_EBX_REG_3__SCAN_IN), .A(n13619), .ZN(
        n13622) );
  NAND4_X1 U16998 ( .A1(n19962), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n13620), .ZN(n13621) );
  OAI211_X1 U16999 ( .C1(n19992), .C2(n13620), .A(n13622), .B(n13621), .ZN(
        n13623) );
  AOI21_X1 U17000 ( .B1(n20415), .B2(n19991), .A(n13623), .ZN(n13624) );
  OAI21_X1 U17001 ( .B1(n13625), .B2(n19990), .A(n13624), .ZN(P1_U2837) );
  INV_X1 U17002 ( .A(n15924), .ZN(n13629) );
  INV_X1 U17003 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U17004 ( .A1(n19949), .A2(n19974), .ZN(n13626) );
  AOI22_X1 U17005 ( .A1(n19963), .A2(P1_EBX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13626), .ZN(n13628) );
  NAND2_X1 U17006 ( .A1(n19977), .A2(n20092), .ZN(n13627) );
  OAI211_X1 U17007 ( .C1(n13629), .C2(n20847), .A(n13628), .B(n13627), .ZN(
        n13630) );
  AOI21_X1 U17008 ( .B1(n11916), .B2(n19991), .A(n13630), .ZN(n13631) );
  OAI21_X1 U17009 ( .B1(n20091), .B2(n19990), .A(n13631), .ZN(P1_U2840) );
  AOI21_X1 U17010 ( .B1(n13822), .B2(n13632), .A(n13682), .ZN(n13820) );
  OAI22_X1 U17011 ( .A1(n21039), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13777) );
  OAI22_X1 U17012 ( .A1(n21039), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13746), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13754) );
  AND2_X1 U17013 ( .A1(n13777), .A2(n13754), .ZN(n13729) );
  NAND2_X1 U17014 ( .A1(n13729), .A2(n13730), .ZN(n13683) );
  NAND2_X1 U17015 ( .A1(n19118), .A2(n13683), .ZN(n13634) );
  XNOR2_X1 U17016 ( .A(n13820), .B(n13634), .ZN(n13635) );
  NAND4_X1 U17017 ( .A1(n19676), .A2(n21039), .A3(n19467), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19782) );
  INV_X1 U17018 ( .A(n19782), .ZN(n19123) );
  NAND2_X1 U17019 ( .A1(n13635), .A2(n19123), .ZN(n13661) );
  OR2_X1 U17020 ( .A1(n13637), .A2(n13636), .ZN(n13638) );
  NAND2_X1 U17021 ( .A1(n13638), .A2(n13690), .ZN(n19206) );
  NOR2_X1 U17022 ( .A1(n13639), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16380) );
  AND2_X1 U17023 ( .A1(n16380), .A2(n16379), .ZN(n13640) );
  NOR2_X1 U17024 ( .A1(n19678), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19497) );
  INV_X1 U17025 ( .A(n19497), .ZN(n13641) );
  NOR2_X1 U17026 ( .A1(n13642), .A2(n13641), .ZN(n16391) );
  INV_X1 U17027 ( .A(n16391), .ZN(n13643) );
  NAND3_X1 U17028 ( .A1(n13643), .A2(n19088), .A3(n19782), .ZN(n13644) );
  NAND2_X1 U17029 ( .A1(n19096), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19084) );
  INV_X1 U17030 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19806) );
  OAI22_X1 U17031 ( .A1(n13822), .A2(n19084), .B1(n19806), .B2(n19096), .ZN(
        n13654) );
  AND2_X1 U17032 ( .A1(n21033), .A2(n13645), .ZN(n13656) );
  NOR2_X1 U17033 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19786), .ZN(n13655) );
  NOR2_X1 U17034 ( .A1(n13655), .A2(n11561), .ZN(n13646) );
  OR2_X1 U17035 ( .A1(n13647), .A2(n16380), .ZN(n14674) );
  INV_X1 U17036 ( .A(n13655), .ZN(n13648) );
  NAND3_X1 U17037 ( .A1(n13649), .A2(n11561), .A3(n13648), .ZN(n13650) );
  INV_X1 U17038 ( .A(n19110), .ZN(n19097) );
  OAI22_X1 U17039 ( .A1(n19112), .A2(n13652), .B1(n19097), .B2(n13651), .ZN(
        n13653) );
  NOR2_X1 U17040 ( .A1(n13654), .A2(n13653), .ZN(n13658) );
  NAND2_X1 U17041 ( .A1(n13164), .A2(n19122), .ZN(n13657) );
  OAI211_X1 U17042 ( .C1(n19206), .C2(n19127), .A(n13658), .B(n13657), .ZN(
        n13659) );
  AOI21_X1 U17043 ( .B1(n19871), .B2(n13757), .A(n13659), .ZN(n13660) );
  NAND2_X1 U17044 ( .A1(n13661), .A2(n13660), .ZN(P2_U2852) );
  NAND2_X1 U17045 ( .A1(n13608), .A2(n13663), .ZN(n13664) );
  AND2_X1 U17046 ( .A1(n13662), .A2(n13664), .ZN(n20011) );
  INV_X1 U17047 ( .A(n20011), .ZN(n13666) );
  OAI222_X1 U17048 ( .A1(n14411), .A2(n13666), .B1(n14404), .B2(n20151), .C1(
        n13665), .C2(n14405), .ZN(P1_U2897) );
  NOR2_X1 U17049 ( .A1(n19102), .A2(n19782), .ZN(n14795) );
  INV_X1 U17050 ( .A(n14795), .ZN(n13676) );
  NOR2_X1 U17051 ( .A1(n19118), .A2(n19782), .ZN(n13752) );
  OAI21_X1 U17052 ( .B1(n19109), .B2(n13752), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13675) );
  OAI22_X1 U17053 ( .A1(n13667), .A2(n19127), .B1(n19096), .B2(n10738), .ZN(
        n13668) );
  AOI21_X1 U17054 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19110), .A(n13668), .ZN(
        n13669) );
  OAI21_X1 U17055 ( .B1(n13670), .B2(n19112), .A(n13669), .ZN(n13672) );
  INV_X1 U17056 ( .A(n13757), .ZN(n13741) );
  NOR2_X1 U17057 ( .A1(n19894), .A2(n13741), .ZN(n13671) );
  AOI211_X1 U17058 ( .C1(n19122), .C2(n13673), .A(n13672), .B(n13671), .ZN(
        n13674) );
  OAI211_X1 U17059 ( .C1(n13676), .C2(n13777), .A(n13675), .B(n13674), .ZN(
        P2_U2855) );
  AOI21_X1 U17060 ( .B1(n13678), .B2(n13662), .A(n13677), .ZN(n13726) );
  INV_X1 U17061 ( .A(n13726), .ZN(n19955) );
  MUX2_X1 U17062 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20104), .Z(
        n20048) );
  AOI22_X1 U17063 ( .A1(n14409), .A2(n20048), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15946), .ZN(n13679) );
  OAI21_X1 U17064 ( .B1(n19955), .B2(n14411), .A(n13679), .ZN(P1_U2896) );
  OAI21_X1 U17065 ( .B1(n13680), .B2(n13681), .A(n13280), .ZN(n19200) );
  OAI21_X1 U17066 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13682), .A(
        n13706), .ZN(n15230) );
  INV_X1 U17067 ( .A(n15230), .ZN(n13686) );
  NOR2_X1 U17068 ( .A1(n13820), .A2(n13683), .ZN(n13707) );
  NOR2_X1 U17069 ( .A1(n19102), .A2(n13707), .ZN(n13685) );
  AOI21_X1 U17070 ( .B1(n13686), .B2(n13685), .A(n19782), .ZN(n13684) );
  OAI21_X1 U17071 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13699) );
  NAND2_X1 U17072 ( .A1(n13688), .A2(n13687), .ZN(n13689) );
  AND2_X1 U17073 ( .A1(n13193), .A2(n13689), .ZN(n19155) );
  INV_X1 U17074 ( .A(n13690), .ZN(n13691) );
  XNOR2_X1 U17075 ( .A(n13692), .B(n13691), .ZN(n15558) );
  INV_X1 U17076 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19808) );
  AOI22_X1 U17077 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19109), .ZN(n13693) );
  OAI211_X1 U17078 ( .C1(n19096), .C2(n19808), .A(n13693), .B(n11494), .ZN(
        n13694) );
  AOI21_X1 U17079 ( .B1(n14829), .B2(n15558), .A(n13694), .ZN(n13695) );
  OAI21_X1 U17080 ( .B1(n13696), .B2(n19112), .A(n13695), .ZN(n13697) );
  AOI21_X1 U17081 ( .B1(n19155), .B2(n19122), .A(n13697), .ZN(n13698) );
  OAI211_X1 U17082 ( .C1(n19200), .C2(n13741), .A(n13699), .B(n13698), .ZN(
        P2_U2851) );
  INV_X1 U17083 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13703) );
  OR2_X1 U17084 ( .A1(n16188), .A2(n13700), .ZN(n13701) );
  AND2_X1 U17085 ( .A1(n13701), .A2(n16162), .ZN(n19951) );
  INV_X1 U17086 ( .A(n19951), .ZN(n13702) );
  OAI222_X1 U17087 ( .A1(n19955), .A2(n14364), .B1(n20014), .B2(n13703), .C1(
        n13702), .C2(n14358), .ZN(P1_U2864) );
  OAI21_X1 U17088 ( .B1(n11192), .B2(n11191), .A(n13515), .ZN(n19154) );
  AOI21_X1 U17089 ( .B1(n19083), .B2(n13708), .A(n13710), .ZN(n19081) );
  AOI21_X1 U17090 ( .B1(n16314), .B2(n13706), .A(n13709), .ZN(n19120) );
  NAND2_X1 U17091 ( .A1(n13707), .A2(n15230), .ZN(n19117) );
  NOR2_X1 U17092 ( .A1(n19120), .A2(n19117), .ZN(n19101) );
  OAI21_X1 U17093 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13709), .A(
        n13708), .ZN(n19103) );
  NAND2_X1 U17094 ( .A1(n19101), .A2(n19103), .ZN(n19080) );
  NOR2_X1 U17095 ( .A1(n19081), .A2(n19080), .ZN(n14655) );
  NOR2_X1 U17096 ( .A1(n19102), .A2(n14655), .ZN(n13711) );
  OAI21_X1 U17097 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13710), .A(
        n13802), .ZN(n16296) );
  XNOR2_X1 U17098 ( .A(n13711), .B(n16296), .ZN(n13712) );
  NAND2_X1 U17099 ( .A1(n13712), .A2(n19123), .ZN(n13720) );
  INV_X1 U17100 ( .A(n19096), .ZN(n19116) );
  AOI21_X1 U17101 ( .B1(n13713), .B2(n15505), .A(n13795), .ZN(n13714) );
  INV_X1 U17102 ( .A(n13714), .ZN(n19194) );
  AOI22_X1 U17103 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19109), .ZN(n13715) );
  OAI211_X1 U17104 ( .C1(n19127), .C2(n19194), .A(n13715), .B(n11494), .ZN(
        n13718) );
  NOR2_X1 U17105 ( .A1(n13716), .A2(n19112), .ZN(n13717) );
  AOI211_X1 U17106 ( .C1(n19116), .C2(P2_REIP_REG_8__SCAN_IN), .A(n13718), .B(
        n13717), .ZN(n13719) );
  OAI211_X1 U17107 ( .C1(n19090), .C2(n19154), .A(n13720), .B(n13719), .ZN(
        P2_U2847) );
  XNOR2_X1 U17108 ( .A(n13722), .B(n16183), .ZN(n13723) );
  XNOR2_X1 U17109 ( .A(n13721), .B(n13723), .ZN(n16178) );
  INV_X1 U17110 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13724) );
  OAI22_X1 U17111 ( .A1(n16033), .A2(n19948), .B1(n20101), .B2(n13724), .ZN(
        n13725) );
  AOI21_X1 U17112 ( .B1(n16027), .B2(n19958), .A(n13725), .ZN(n13728) );
  NAND2_X1 U17113 ( .A1(n13726), .A2(n16029), .ZN(n13727) );
  OAI211_X1 U17114 ( .C1(n16178), .C2(n19920), .A(n13728), .B(n13727), .ZN(
        P1_U2991) );
  NOR2_X1 U17115 ( .A1(n19102), .A2(n13729), .ZN(n13753) );
  XNOR2_X1 U17116 ( .A(n13753), .B(n13730), .ZN(n13731) );
  NAND2_X1 U17117 ( .A1(n13731), .A2(n19123), .ZN(n13740) );
  OAI22_X1 U17118 ( .A1(n19097), .A2(n13732), .B1(n14996), .B2(n19127), .ZN(
        n13734) );
  NOR2_X1 U17119 ( .A1(n19096), .A2(n19804), .ZN(n13733) );
  AOI211_X1 U17120 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19109), .A(
        n13734), .B(n13733), .ZN(n13735) );
  OAI21_X1 U17121 ( .B1(n13736), .B2(n19112), .A(n13735), .ZN(n13737) );
  AOI21_X1 U17122 ( .B1(n13738), .B2(n19122), .A(n13737), .ZN(n13739) );
  OAI211_X1 U17123 ( .C1(n13741), .C2(n19877), .A(n13740), .B(n13739), .ZN(
        P2_U2853) );
  NOR2_X1 U17124 ( .A1(n13677), .A2(n13743), .ZN(n13744) );
  OR2_X1 U17125 ( .A1(n13742), .A2(n13744), .ZN(n19943) );
  MUX2_X1 U17126 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20104), .Z(
        n20050) );
  AOI22_X1 U17127 ( .A1(n14409), .A2(n20050), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15946), .ZN(n13745) );
  OAI21_X1 U17128 ( .B1(n19943), .B2(n14411), .A(n13745), .ZN(P1_U2895) );
  OAI22_X1 U17129 ( .A1(n19096), .A2(n13003), .B1(n19084), .B2(n13746), .ZN(
        n13749) );
  NOR2_X1 U17130 ( .A1(n19112), .A2(n13747), .ZN(n13748) );
  AOI211_X1 U17131 ( .C1(n19110), .C2(P2_EBX_REG_1__SCAN_IN), .A(n13749), .B(
        n13748), .ZN(n13751) );
  NAND2_X1 U17132 ( .A1(n19889), .A2(n14829), .ZN(n13750) );
  OAI211_X1 U17133 ( .C1(n13784), .C2(n19090), .A(n13751), .B(n13750), .ZN(
        n13756) );
  INV_X1 U17134 ( .A(n13752), .ZN(n19013) );
  OAI21_X1 U17135 ( .B1(n13777), .B2(n13754), .A(n13753), .ZN(n13775) );
  OAI22_X1 U17136 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19013), .B1(
        n13775), .B2(n19782), .ZN(n13755) );
  AOI211_X1 U17137 ( .C1(n13757), .C2(n19887), .A(n13756), .B(n13755), .ZN(
        n13758) );
  INV_X1 U17138 ( .A(n13758), .ZN(P2_U2854) );
  OR2_X1 U17139 ( .A1(n13742), .A2(n13760), .ZN(n13761) );
  AND2_X1 U17140 ( .A1(n13759), .A2(n13761), .ZN(n15938) );
  INV_X1 U17141 ( .A(n14364), .ZN(n20010) );
  NAND2_X1 U17142 ( .A1(n16160), .A2(n13762), .ZN(n13763) );
  NAND2_X1 U17143 ( .A1(n9705), .A2(n13763), .ZN(n16158) );
  OAI22_X1 U17144 ( .A1(n16158), .A2(n14358), .B1(n13764), .B2(n20014), .ZN(
        n13765) );
  AOI21_X1 U17145 ( .B1(n15938), .B2(n20010), .A(n13765), .ZN(n13766) );
  INV_X1 U17146 ( .A(n13766), .ZN(P1_U2862) );
  INV_X1 U17147 ( .A(n15938), .ZN(n13768) );
  MUX2_X1 U17148 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20104), .Z(
        n20052) );
  AOI22_X1 U17149 ( .A1(n14409), .A2(n20052), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15946), .ZN(n13767) );
  OAI21_X1 U17150 ( .B1(n13768), .B2(n14411), .A(n13767), .ZN(P1_U2894) );
  XNOR2_X1 U17151 ( .A(n14579), .B(n16170), .ZN(n13770) );
  XNOR2_X1 U17152 ( .A(n13769), .B(n13770), .ZN(n16165) );
  INV_X1 U17153 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13771) );
  OAI22_X1 U17154 ( .A1(n16033), .A2(n19941), .B1(n20101), .B2(n13771), .ZN(
        n13773) );
  NOR2_X1 U17155 ( .A1(n19943), .A2(n20106), .ZN(n13772) );
  AOI211_X1 U17156 ( .C1(n16027), .C2(n19939), .A(n13773), .B(n13772), .ZN(
        n13774) );
  OAI21_X1 U17157 ( .B1(n19920), .B2(n16165), .A(n13774), .ZN(P1_U2990) );
  OAI21_X1 U17158 ( .B1(n19118), .B2(n13776), .A(n13775), .ZN(n15583) );
  INV_X1 U17159 ( .A(n13777), .ZN(n13778) );
  OAI221_X1 U17160 ( .B1(n13778), .B2(n19102), .C1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19118), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n15597) );
  NAND2_X1 U17161 ( .A1(n13780), .A2(n13779), .ZN(n15575) );
  INV_X1 U17162 ( .A(n13781), .ZN(n13782) );
  AOI22_X1 U17163 ( .A1(n10456), .A2(n11275), .B1(n15575), .B2(n13782), .ZN(
        n13783) );
  OAI22_X1 U17164 ( .A1(n13784), .A2(n15593), .B1(n13182), .B2(n13783), .ZN(
        n16345) );
  AOI22_X1 U17165 ( .A1(n19887), .A2(n15594), .B1(n19779), .B2(n16345), .ZN(
        n13785) );
  OAI21_X1 U17166 ( .B1(n15583), .B2(n15597), .A(n13785), .ZN(n13786) );
  MUX2_X1 U17167 ( .A(n13786), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15599), .Z(P2_U3600) );
  OAI21_X1 U17168 ( .B1(n13788), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n13787), .ZN(n13809) );
  INV_X1 U17169 ( .A(n13789), .ZN(n13792) );
  AOI21_X1 U17170 ( .B1(n13790), .B2(n15479), .A(n9661), .ZN(n13791) );
  AOI21_X1 U17171 ( .B1(n13792), .B2(n15479), .A(n13791), .ZN(n13807) );
  INV_X1 U17172 ( .A(n15459), .ZN(n13793) );
  OAI21_X1 U17173 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n13794), .A(
        n13793), .ZN(n13799) );
  OAI21_X1 U17174 ( .B1(n13796), .B2(n13795), .A(n15489), .ZN(n19191) );
  INV_X1 U17175 ( .A(n19191), .ZN(n13797) );
  AOI22_X1 U17176 ( .A1(n19261), .A2(n13797), .B1(n19115), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n13798) );
  OAI211_X1 U17177 ( .C1(n19257), .C2(n19075), .A(n13799), .B(n13798), .ZN(
        n13800) );
  AOI21_X1 U17178 ( .B1(n13807), .B2(n16338), .A(n13800), .ZN(n13801) );
  OAI21_X1 U17179 ( .B1(n19264), .B2(n13809), .A(n13801), .ZN(P2_U3037) );
  AOI21_X1 U17180 ( .B1(n13803), .B2(n13802), .A(n9680), .ZN(n19071) );
  INV_X1 U17181 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20975) );
  OAI22_X1 U17182 ( .A1(n16315), .A2(n13803), .B1(n20975), .B2(n19088), .ZN(
        n13804) );
  AOI21_X1 U17183 ( .B1(n16305), .B2(n19071), .A(n13804), .ZN(n13805) );
  OAI21_X1 U17184 ( .B1(n19075), .B2(n13376), .A(n13805), .ZN(n13806) );
  AOI21_X1 U17185 ( .B1(n13807), .B2(n16293), .A(n13806), .ZN(n13808) );
  OAI21_X1 U17186 ( .B1(n16308), .B2(n13809), .A(n13808), .ZN(P2_U3005) );
  AOI22_X1 U17187 ( .A1(n15949), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15946), .ZN(n13812) );
  MUX2_X1 U17188 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20104), .Z(
        n20058) );
  AOI22_X1 U17189 ( .A1(n9726), .A2(n20058), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n14399), .ZN(n13811) );
  OAI211_X1 U17190 ( .C1(n14142), .C2(n14411), .A(n13812), .B(n13811), .ZN(
        P1_U2875) );
  INV_X1 U17191 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14147) );
  OAI21_X1 U17192 ( .B1(n14156), .B2(n13814), .A(n13813), .ZN(n14560) );
  OAI222_X1 U17193 ( .A1(n14364), .A2(n14142), .B1(n14147), .B2(n20014), .C1(
        n14560), .C2(n14358), .ZN(P1_U2843) );
  XNOR2_X1 U17194 ( .A(n13815), .B(n13816), .ZN(n16335) );
  XNOR2_X1 U17195 ( .A(n13817), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13818) );
  XNOR2_X1 U17196 ( .A(n13819), .B(n13818), .ZN(n16337) );
  NAND2_X1 U17197 ( .A1(n16337), .A2(n16293), .ZN(n13825) );
  NAND2_X1 U17198 ( .A1(n16305), .A2(n13820), .ZN(n13821) );
  NAND2_X1 U17199 ( .A1(n19115), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16330) );
  OAI211_X1 U17200 ( .C1(n13822), .C2(n16315), .A(n13821), .B(n16330), .ZN(
        n13823) );
  AOI21_X1 U17201 ( .B1(n13164), .B2(n16311), .A(n13823), .ZN(n13824) );
  OAI211_X1 U17202 ( .C1(n16335), .C2(n16308), .A(n13825), .B(n13824), .ZN(
        P2_U3011) );
  OR2_X1 U17203 ( .A1(n14909), .A2(n19138), .ZN(n14910) );
  NOR2_X1 U17204 ( .A1(n14910), .A2(n19133), .ZN(n13827) );
  AOI22_X1 U17205 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13834) );
  AOI22_X1 U17206 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17207 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U17208 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13831) );
  NAND4_X1 U17209 ( .A1(n13834), .A2(n13833), .A3(n13832), .A4(n13831), .ZN(
        n13840) );
  AOI22_X1 U17210 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13838) );
  AOI22_X1 U17211 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13837) );
  AOI22_X1 U17212 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13836) );
  AOI22_X1 U17213 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13835) );
  NAND4_X1 U17214 ( .A1(n13838), .A2(n13837), .A3(n13836), .A4(n13835), .ZN(
        n13839) );
  NAND2_X1 U17215 ( .A1(n14901), .A2(n19128), .ZN(n14895) );
  AOI22_X1 U17216 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10662), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17217 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17218 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17219 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13841) );
  NAND4_X1 U17220 ( .A1(n13844), .A2(n13843), .A3(n13842), .A4(n13841), .ZN(
        n13850) );
  AOI22_X1 U17221 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U17222 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U17223 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17224 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13845) );
  NAND4_X1 U17225 ( .A1(n13848), .A2(n13847), .A3(n13846), .A4(n13845), .ZN(
        n13849) );
  NOR2_X1 U17226 ( .A1(n13850), .A2(n13849), .ZN(n14898) );
  AOI22_X1 U17227 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U17228 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U17229 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13852) );
  AOI22_X1 U17230 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13851) );
  NAND4_X1 U17231 ( .A1(n13854), .A2(n13853), .A3(n13852), .A4(n13851), .ZN(
        n13860) );
  AOI22_X1 U17232 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13858) );
  AOI22_X1 U17233 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U17234 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U17235 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13855) );
  NAND4_X1 U17236 ( .A1(n13858), .A2(n13857), .A3(n13856), .A4(n13855), .ZN(
        n13859) );
  NOR2_X1 U17237 ( .A1(n13860), .A2(n13859), .ZN(n16254) );
  INV_X1 U17238 ( .A(n16254), .ZN(n13861) );
  AOI22_X1 U17239 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10662), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17240 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17241 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13863) );
  AOI22_X1 U17242 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13862) );
  NAND4_X1 U17243 ( .A1(n13865), .A2(n13864), .A3(n13863), .A4(n13862), .ZN(
        n13871) );
  AOI22_X1 U17244 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13869) );
  AOI22_X1 U17245 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U17246 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13867) );
  AOI22_X1 U17247 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13866) );
  NAND4_X1 U17248 ( .A1(n13869), .A2(n13868), .A3(n13867), .A4(n13866), .ZN(
        n13870) );
  OR2_X1 U17249 ( .A1(n13871), .A2(n13870), .ZN(n14885) );
  AOI22_X1 U17250 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U17251 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17252 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17253 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13872) );
  NAND4_X1 U17254 ( .A1(n13875), .A2(n13874), .A3(n13873), .A4(n13872), .ZN(
        n13881) );
  AOI22_X1 U17255 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U17256 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U17257 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U17258 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13876) );
  NAND4_X1 U17259 ( .A1(n13879), .A2(n13878), .A3(n13877), .A4(n13876), .ZN(
        n13880) );
  OR2_X1 U17260 ( .A1(n13881), .A2(n13880), .ZN(n16249) );
  AOI22_X1 U17261 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17262 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U17263 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13883) );
  AOI22_X1 U17264 ( .A1(n13907), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13882) );
  NAND4_X1 U17265 ( .A1(n13885), .A2(n13884), .A3(n13883), .A4(n13882), .ZN(
        n13896) );
  AOI22_X1 U17266 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17267 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13893) );
  INV_X1 U17268 ( .A(n13912), .ZN(n13889) );
  INV_X1 U17269 ( .A(n13886), .ZN(n13888) );
  INV_X1 U17270 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13887) );
  OAI22_X1 U17271 ( .A1(n10879), .A2(n13889), .B1(n13888), .B2(n13887), .ZN(
        n13890) );
  INV_X1 U17272 ( .A(n13890), .ZN(n13892) );
  AOI22_X1 U17273 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13891) );
  NAND4_X1 U17274 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n13891), .ZN(
        n13895) );
  OR2_X1 U17275 ( .A1(n13896), .A2(n13895), .ZN(n14878) );
  AOI22_X1 U17276 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10650), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17277 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U17278 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10906), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U17279 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13907), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13897) );
  NAND4_X1 U17280 ( .A1(n13900), .A2(n13899), .A3(n13898), .A4(n13897), .ZN(
        n13906) );
  AOI22_X1 U17281 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n9625), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17282 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13913), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17283 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17284 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10855), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13901) );
  NAND4_X1 U17285 ( .A1(n13904), .A2(n13903), .A3(n13902), .A4(n13901), .ZN(
        n13905) );
  NOR2_X1 U17286 ( .A1(n13906), .A2(n13905), .ZN(n16246) );
  AOI22_X1 U17287 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10650), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U17288 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U17289 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13907), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17290 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10906), .B1(
        n11371), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13908) );
  NAND4_X1 U17291 ( .A1(n13911), .A2(n13910), .A3(n13909), .A4(n13908), .ZN(
        n13919) );
  AOI22_X1 U17292 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10912), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17293 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13912), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U17294 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n13913), .B1(
        n10855), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U17295 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n9625), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13914) );
  NAND4_X1 U17296 ( .A1(n13917), .A2(n13916), .A3(n13915), .A4(n13914), .ZN(
        n13918) );
  NOR2_X1 U17297 ( .A1(n13919), .A2(n13918), .ZN(n13958) );
  INV_X1 U17298 ( .A(n9628), .ZN(n14079) );
  INV_X1 U17299 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19655) );
  INV_X1 U17300 ( .A(n14099), .ZN(n14074) );
  INV_X1 U17301 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13920) );
  OAI22_X1 U17302 ( .A1(n14079), .A2(n19655), .B1(n14074), .B2(n13920), .ZN(
        n13923) );
  INV_X1 U17303 ( .A(n10621), .ZN(n14076) );
  INV_X1 U17304 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13921) );
  INV_X1 U17305 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19558) );
  OAI22_X1 U17306 ( .A1(n14076), .A2(n13921), .B1(n9620), .B2(n19558), .ZN(
        n13922) );
  NOR2_X1 U17307 ( .A1(n13923), .A2(n13922), .ZN(n13926) );
  AOI22_X1 U17308 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13925) );
  XNOR2_X1 U17309 ( .A(n10459), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14100) );
  AOI22_X1 U17310 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13924) );
  NAND4_X1 U17311 ( .A1(n13926), .A2(n13925), .A3(n14100), .A4(n13924), .ZN(
        n13935) );
  AOI22_X1 U17312 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U17313 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13932) );
  NAND2_X1 U17314 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13930) );
  NAND2_X1 U17315 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13929) );
  NAND2_X1 U17316 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13928) );
  NAND2_X1 U17317 ( .A1(n9621), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13927) );
  AND4_X1 U17318 ( .A1(n13930), .A2(n13929), .A3(n13928), .A4(n13927), .ZN(
        n13931) );
  INV_X1 U17319 ( .A(n14100), .ZN(n14093) );
  NAND4_X1 U17320 ( .A1(n13933), .A2(n13932), .A3(n13931), .A4(n14093), .ZN(
        n13934) );
  NAND2_X1 U17321 ( .A1(n21042), .A2(n13961), .ZN(n13936) );
  XNOR2_X1 U17322 ( .A(n13958), .B(n13936), .ZN(n13964) );
  NAND2_X1 U17323 ( .A1(n14062), .A2(n13961), .ZN(n14966) );
  OAI22_X1 U17325 ( .A1(n14076), .A2(n13940), .B1(n14079), .B2(n10840), .ZN(
        n13944) );
  INV_X1 U17326 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13941) );
  OAI22_X1 U17327 ( .A1(n14074), .A2(n13942), .B1(n9620), .B2(n13941), .ZN(
        n13943) );
  NOR2_X1 U17328 ( .A1(n13944), .A2(n13943), .ZN(n13947) );
  AOI22_X1 U17329 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13946) );
  AOI22_X1 U17330 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13945) );
  NAND4_X1 U17331 ( .A1(n13947), .A2(n13946), .A3(n13945), .A4(n14093), .ZN(
        n13957) );
  OAI22_X1 U17332 ( .A1(n14076), .A2(n13949), .B1(n14079), .B2(n13948), .ZN(
        n13952) );
  OAI22_X1 U17333 ( .A1(n14074), .A2(n13950), .B1(n9620), .B2(n15613), .ZN(
        n13951) );
  NOR2_X1 U17334 ( .A1(n13952), .A2(n13951), .ZN(n13955) );
  AOI22_X1 U17335 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17336 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13953) );
  NAND4_X1 U17337 ( .A1(n13955), .A2(n13954), .A3(n14100), .A4(n13953), .ZN(
        n13956) );
  NAND2_X1 U17338 ( .A1(n13957), .A2(n13956), .ZN(n13966) );
  INV_X1 U17339 ( .A(n13958), .ZN(n13959) );
  NAND2_X1 U17340 ( .A1(n13959), .A2(n13961), .ZN(n13967) );
  XOR2_X1 U17341 ( .A(n13966), .B(n13967), .Z(n13960) );
  NAND2_X1 U17342 ( .A1(n13960), .A2(n14034), .ZN(n14872) );
  INV_X1 U17343 ( .A(n13961), .ZN(n13963) );
  INV_X1 U17344 ( .A(n13966), .ZN(n13962) );
  NAND2_X1 U17345 ( .A1(n14062), .A2(n13962), .ZN(n14874) );
  NOR2_X1 U17346 ( .A1(n13967), .A2(n13966), .ZN(n13984) );
  AOI22_X1 U17347 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17348 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13973) );
  NAND2_X1 U17349 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13971) );
  NAND2_X1 U17350 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13970) );
  NAND2_X1 U17351 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13969) );
  NAND2_X1 U17352 ( .A1(n9621), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13968) );
  AND4_X1 U17353 ( .A1(n13971), .A2(n13970), .A3(n13969), .A4(n13968), .ZN(
        n13972) );
  NAND4_X1 U17354 ( .A1(n13974), .A2(n13973), .A3(n13972), .A4(n14093), .ZN(
        n13983) );
  AOI22_X1 U17355 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13981) );
  AOI22_X1 U17356 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13980) );
  NAND2_X1 U17357 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13978) );
  NAND2_X1 U17358 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13977) );
  NAND2_X1 U17359 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13976) );
  NAND2_X1 U17360 ( .A1(n9621), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13975) );
  AND4_X1 U17361 ( .A1(n13978), .A2(n13977), .A3(n13976), .A4(n13975), .ZN(
        n13979) );
  NAND4_X1 U17362 ( .A1(n13981), .A2(n14100), .A3(n13980), .A4(n13979), .ZN(
        n13982) );
  AND2_X1 U17363 ( .A1(n13983), .A2(n13982), .ZN(n13985) );
  NAND2_X1 U17364 ( .A1(n13984), .A2(n13985), .ZN(n14012) );
  OAI211_X1 U17365 ( .C1(n13984), .C2(n13985), .A(n14034), .B(n14012), .ZN(
        n13987) );
  NAND2_X1 U17366 ( .A1(n14062), .A2(n13985), .ZN(n14866) );
  OR2_X2 U17367 ( .A1(n14862), .A2(n14866), .ZN(n14863) );
  OAI22_X1 U17368 ( .A1(n14076), .A2(n13991), .B1(n14079), .B2(n13990), .ZN(
        n13995) );
  OAI22_X1 U17369 ( .A1(n14074), .A2(n13993), .B1(n9620), .B2(n13992), .ZN(
        n13994) );
  NOR2_X1 U17370 ( .A1(n13995), .A2(n13994), .ZN(n13998) );
  AOI22_X1 U17371 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13997) );
  AOI22_X1 U17372 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13996) );
  NAND4_X1 U17373 ( .A1(n13998), .A2(n13997), .A3(n13996), .A4(n14093), .ZN(
        n14009) );
  OAI22_X1 U17374 ( .A1(n14076), .A2(n14000), .B1(n14079), .B2(n13999), .ZN(
        n14004) );
  OAI22_X1 U17375 ( .A1(n14074), .A2(n14002), .B1(n9620), .B2(n14001), .ZN(
        n14003) );
  NOR2_X1 U17376 ( .A1(n14004), .A2(n14003), .ZN(n14007) );
  AOI22_X1 U17377 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17378 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14005) );
  NAND4_X1 U17379 ( .A1(n14007), .A2(n14006), .A3(n14100), .A4(n14005), .ZN(
        n14008) );
  AND2_X1 U17380 ( .A1(n14009), .A2(n14008), .ZN(n14013) );
  XNOR2_X1 U17381 ( .A(n14012), .B(n14013), .ZN(n14010) );
  NAND2_X1 U17382 ( .A1(n14062), .A2(n14013), .ZN(n14859) );
  INV_X1 U17383 ( .A(n14012), .ZN(n14014) );
  AND2_X1 U17384 ( .A1(n14014), .A2(n14013), .ZN(n14035) );
  OAI22_X1 U17385 ( .A1(n10488), .A2(n14016), .B1(n10573), .B2(n14015), .ZN(
        n14020) );
  INV_X1 U17386 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14018) );
  INV_X1 U17387 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14017) );
  OAI22_X1 U17388 ( .A1(n10620), .A2(n14018), .B1(n10627), .B2(n14017), .ZN(
        n14019) );
  NOR2_X1 U17389 ( .A1(n14020), .A2(n14019), .ZN(n14023) );
  AOI22_X1 U17390 ( .A1(n14099), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9621), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17391 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14021) );
  NAND4_X1 U17392 ( .A1(n14023), .A2(n14022), .A3(n14021), .A4(n14093), .ZN(
        n14033) );
  INV_X1 U17393 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14024) );
  INV_X1 U17394 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n19662) );
  OAI22_X1 U17395 ( .A1(n14076), .A2(n14024), .B1(n14079), .B2(n19662), .ZN(
        n14028) );
  INV_X1 U17396 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14026) );
  INV_X1 U17397 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14025) );
  OAI22_X1 U17398 ( .A1(n14074), .A2(n14026), .B1(n9620), .B2(n14025), .ZN(
        n14027) );
  NOR2_X1 U17399 ( .A1(n14028), .A2(n14027), .ZN(n14031) );
  AOI22_X1 U17400 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17401 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14029) );
  NAND4_X1 U17402 ( .A1(n14031), .A2(n14030), .A3(n14100), .A4(n14029), .ZN(
        n14032) );
  AND2_X1 U17403 ( .A1(n14033), .A2(n14032), .ZN(n14040) );
  NAND2_X1 U17404 ( .A1(n14035), .A2(n14040), .ZN(n14060) );
  OAI211_X1 U17405 ( .C1(n14035), .C2(n14040), .A(n14034), .B(n14060), .ZN(
        n14036) );
  INV_X1 U17406 ( .A(n14845), .ZN(n14039) );
  NAND2_X1 U17407 ( .A1(n14037), .A2(n14036), .ZN(n14038) );
  INV_X1 U17408 ( .A(n14040), .ZN(n14041) );
  OR2_X1 U17409 ( .A1(n10710), .A2(n14041), .ZN(n14853) );
  OAI22_X1 U17410 ( .A1(n14076), .A2(n14043), .B1(n14079), .B2(n14042), .ZN(
        n14047) );
  OAI22_X1 U17411 ( .A1(n14074), .A2(n14045), .B1(n9620), .B2(n14044), .ZN(
        n14046) );
  NOR2_X1 U17412 ( .A1(n14047), .A2(n14046), .ZN(n14050) );
  AOI22_X1 U17413 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U17414 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14048) );
  NAND4_X1 U17415 ( .A1(n14050), .A2(n14049), .A3(n14100), .A4(n14048), .ZN(
        n14059) );
  AOI22_X1 U17416 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17417 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14056) );
  NAND2_X1 U17418 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14054) );
  NAND2_X1 U17419 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14053) );
  NAND2_X1 U17420 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14052) );
  NAND2_X1 U17421 ( .A1(n9621), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n14051) );
  AND4_X1 U17422 ( .A1(n14054), .A2(n14053), .A3(n14052), .A4(n14051), .ZN(
        n14055) );
  NAND4_X1 U17423 ( .A1(n14057), .A2(n14056), .A3(n14055), .A4(n14093), .ZN(
        n14058) );
  AND2_X1 U17424 ( .A1(n14059), .A2(n14058), .ZN(n14061) );
  INV_X1 U17425 ( .A(n14060), .ZN(n14844) );
  INV_X1 U17426 ( .A(n14061), .ZN(n14846) );
  NOR2_X1 U17427 ( .A1(n14062), .A2(n14846), .ZN(n14063) );
  AND2_X1 U17428 ( .A1(n14844), .A2(n14063), .ZN(n14088) );
  OAI22_X1 U17429 ( .A1(n14076), .A2(n14065), .B1(n14079), .B2(n14064), .ZN(
        n14069) );
  OAI22_X1 U17430 ( .A1(n14074), .A2(n14067), .B1(n9620), .B2(n14066), .ZN(
        n14068) );
  NOR2_X1 U17431 ( .A1(n14069), .A2(n14068), .ZN(n14072) );
  AOI22_X1 U17432 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14071) );
  AOI22_X1 U17433 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14070) );
  NAND4_X1 U17434 ( .A1(n14072), .A2(n14071), .A3(n14070), .A4(n14093), .ZN(
        n14086) );
  OAI22_X1 U17435 ( .A1(n14076), .A2(n14075), .B1(n14074), .B2(n14073), .ZN(
        n14081) );
  OAI22_X1 U17436 ( .A1(n14079), .A2(n14078), .B1(n9620), .B2(n14077), .ZN(
        n14080) );
  NOR2_X1 U17437 ( .A1(n14081), .A2(n14080), .ZN(n14084) );
  AOI22_X1 U17438 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17439 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14082) );
  NAND4_X1 U17440 ( .A1(n14084), .A2(n14083), .A3(n14100), .A4(n14082), .ZN(
        n14085) );
  AND2_X1 U17441 ( .A1(n14086), .A2(n14085), .ZN(n14087) );
  NAND2_X1 U17442 ( .A1(n14088), .A2(n14087), .ZN(n14089) );
  OAI21_X1 U17443 ( .B1(n14088), .B2(n14087), .A(n14089), .ZN(n14840) );
  INV_X1 U17444 ( .A(n14089), .ZN(n14090) );
  AOI22_X1 U17445 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17446 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14091) );
  NAND2_X1 U17447 ( .A1(n14092), .A2(n14091), .ZN(n14106) );
  AOI22_X1 U17448 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14099), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17449 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9621), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14094) );
  NAND3_X1 U17450 ( .A1(n14095), .A2(n14094), .A3(n14093), .ZN(n14105) );
  AOI22_X1 U17451 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17452 ( .A1(n15584), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10628), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14097) );
  NAND2_X1 U17453 ( .A1(n14098), .A2(n14097), .ZN(n14104) );
  AOI22_X1 U17454 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9628), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U17455 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9621), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14101) );
  NAND3_X1 U17456 ( .A1(n14102), .A2(n14101), .A3(n14100), .ZN(n14103) );
  OAI22_X1 U17457 ( .A1(n14106), .A2(n14105), .B1(n14104), .B2(n14103), .ZN(
        n14107) );
  XNOR2_X1 U17458 ( .A(n14108), .B(n14107), .ZN(n14119) );
  INV_X1 U17459 ( .A(n19165), .ZN(n14948) );
  INV_X1 U17460 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17461 ( .A1(n19164), .A2(n19176), .B1(n19213), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U17462 ( .A1(n19166), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14112) );
  OAI211_X1 U17463 ( .C1(n14948), .C2(n14114), .A(n14113), .B(n14112), .ZN(
        n14115) );
  AOI21_X1 U17464 ( .B1(n14686), .B2(n19214), .A(n14115), .ZN(n14116) );
  OAI21_X1 U17465 ( .B1(n14119), .B2(n19218), .A(n14116), .ZN(P2_U2889) );
  NOR2_X1 U17466 ( .A1(n9575), .A2(n19153), .ZN(n14117) );
  AOI21_X1 U17467 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19153), .A(n14117), .ZN(
        n14118) );
  OAI21_X1 U17468 ( .B1(n14119), .B2(n19148), .A(n14118), .ZN(P2_U2857) );
  NAND2_X1 U17469 ( .A1(n11602), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17470 ( .A1(n11357), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11318), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U17471 ( .A1(n14121), .A2(n14120), .ZN(n14122) );
  XNOR2_X1 U17472 ( .A(n14123), .B(n14122), .ZN(n14673) );
  NAND4_X1 U17473 ( .A1(n15240), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n10048), .A4(n11548), .ZN(n14125) );
  OAI211_X1 U17474 ( .C1(n14673), .C2(n16331), .A(n14125), .B(n14124), .ZN(
        n14126) );
  OAI21_X1 U17475 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15382), .A(
        n14127), .ZN(n14128) );
  OAI21_X1 U17476 ( .B1(n14130), .B2(n19257), .A(n14129), .ZN(n14131) );
  NAND2_X1 U17477 ( .A1(n14419), .A2(n12623), .ZN(n14141) );
  OAI22_X1 U17478 ( .A1(n14417), .A2(n19974), .B1(n19949), .B2(n14133), .ZN(
        n14139) );
  INV_X1 U17479 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14137) );
  INV_X1 U17480 ( .A(n14134), .ZN(n14136) );
  AOI21_X1 U17481 ( .B1(n14137), .B2(n14136), .A(n14135), .ZN(n14138) );
  AOI211_X1 U17482 ( .C1(n19963), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14139), .B(
        n14138), .ZN(n14140) );
  OAI211_X1 U17483 ( .C1(n20005), .C2(n14554), .A(n14141), .B(n14140), .ZN(
        P1_U2810) );
  NOR3_X1 U17484 ( .A1(n19994), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14144), 
        .ZN(n14149) );
  AOI22_X1 U17485 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19989), .B1(
        n19987), .B2(n14145), .ZN(n14146) );
  OAI21_X1 U17486 ( .B1(n15883), .B2(n14147), .A(n14146), .ZN(n14148) );
  AOI211_X1 U17487 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14157), .A(n14149), 
        .B(n14148), .ZN(n14150) );
  OAI211_X1 U17488 ( .C1(n20005), .C2(n14560), .A(n14151), .B(n14150), .ZN(
        P1_U2811) );
  AOI21_X1 U17489 ( .B1(n14153), .B2(n14152), .A(n12843), .ZN(n14431) );
  INV_X1 U17490 ( .A(n14431), .ZN(n14370) );
  NOR2_X1 U17491 ( .A1(n14171), .A2(n14154), .ZN(n14155) );
  OR2_X1 U17492 ( .A1(n14156), .A2(n14155), .ZN(n14571) );
  INV_X1 U17493 ( .A(n14571), .ZN(n14165) );
  INV_X1 U17494 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14438) );
  OR2_X1 U17495 ( .A1(n14173), .A2(n14438), .ZN(n14162) );
  NAND2_X1 U17496 ( .A1(n14157), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14161) );
  OAI22_X1 U17497 ( .A1(n14158), .A2(n19949), .B1(n19974), .B2(n14429), .ZN(
        n14159) );
  AOI21_X1 U17498 ( .B1(n19963), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14159), .ZN(
        n14160) );
  OAI211_X1 U17499 ( .C1(n14163), .C2(n14162), .A(n14161), .B(n14160), .ZN(
        n14164) );
  AOI21_X1 U17500 ( .B1(n14165), .B2(n19977), .A(n14164), .ZN(n14166) );
  OAI21_X1 U17501 ( .B1(n14370), .B2(n19954), .A(n14166), .ZN(P1_U2812) );
  NOR2_X1 U17502 ( .A1(n14181), .A2(n14169), .ZN(n14170) );
  OR2_X1 U17503 ( .A1(n14171), .A2(n14170), .ZN(n16041) );
  INV_X1 U17504 ( .A(n16041), .ZN(n14178) );
  AOI21_X1 U17505 ( .B1(n19962), .B2(n14173), .A(n15926), .ZN(n14189) );
  INV_X1 U17506 ( .A(n14443), .ZN(n14172) );
  OAI22_X1 U17507 ( .A1(n14439), .A2(n19949), .B1(n19974), .B2(n14172), .ZN(
        n14175) );
  NOR3_X1 U17508 ( .A1(n19994), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14173), 
        .ZN(n14174) );
  AOI211_X1 U17509 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n19963), .A(n14175), .B(
        n14174), .ZN(n14176) );
  OAI21_X1 U17510 ( .B1(n14189), .B2(n14438), .A(n14176), .ZN(n14177) );
  AOI21_X1 U17511 ( .B1(n14178), .B2(n19977), .A(n14177), .ZN(n14179) );
  OAI21_X1 U17512 ( .B1(n14440), .B2(n19954), .A(n14179), .ZN(P1_U2813) );
  AND2_X1 U17513 ( .A1(n9694), .A2(n14180), .ZN(n14182) );
  OR2_X1 U17514 ( .A1(n14182), .A2(n14181), .ZN(n16050) );
  AOI21_X1 U17515 ( .B1(n14185), .B2(n14183), .A(n14184), .ZN(n14452) );
  NAND2_X1 U17516 ( .A1(n14452), .A2(n12623), .ZN(n14193) );
  OAI22_X1 U17517 ( .A1(n14186), .A2(n19949), .B1(n19974), .B2(n14450), .ZN(
        n14191) );
  AOI21_X1 U17518 ( .B1(n19962), .B2(n14187), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14188) );
  NOR2_X1 U17519 ( .A1(n14189), .A2(n14188), .ZN(n14190) );
  AOI211_X1 U17520 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n19963), .A(n14191), .B(
        n14190), .ZN(n14192) );
  OAI211_X1 U17521 ( .C1(n16050), .C2(n20005), .A(n14193), .B(n14192), .ZN(
        P1_U2814) );
  OAI21_X1 U17522 ( .B1(n14195), .B2(n14196), .A(n14183), .ZN(n14460) );
  NAND2_X1 U17523 ( .A1(n14212), .A2(n14197), .ZN(n14198) );
  NAND2_X1 U17524 ( .A1(n9694), .A2(n14198), .ZN(n14279) );
  INV_X1 U17525 ( .A(n14279), .ZN(n16053) );
  INV_X1 U17526 ( .A(n14213), .ZN(n14199) );
  NAND2_X1 U17527 ( .A1(n15872), .A2(n14199), .ZN(n14200) );
  NAND2_X1 U17528 ( .A1(n15924), .A2(n14200), .ZN(n15833) );
  INV_X1 U17529 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14458) );
  INV_X1 U17530 ( .A(n14463), .ZN(n14201) );
  OAI22_X1 U17531 ( .A1(n14459), .A2(n19949), .B1(n19974), .B2(n14201), .ZN(
        n14202) );
  AOI21_X1 U17532 ( .B1(n19963), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14202), .ZN(
        n14205) );
  OAI21_X1 U17533 ( .B1(n14213), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14203) );
  OAI211_X1 U17534 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(P1_REIP_REG_24__SCAN_IN), .A(n19962), .B(n14203), .ZN(n14204) );
  OAI211_X1 U17535 ( .C1(n15833), .C2(n14458), .A(n14205), .B(n14204), .ZN(
        n14206) );
  AOI21_X1 U17536 ( .B1(n16053), .B2(n19977), .A(n14206), .ZN(n14207) );
  OAI21_X1 U17537 ( .B1(n14460), .B2(n19954), .A(n14207), .ZN(P1_U2815) );
  AOI21_X1 U17538 ( .B1(n14209), .B2(n14208), .A(n14195), .ZN(n14471) );
  INV_X1 U17539 ( .A(n14471), .ZN(n14380) );
  OR2_X1 U17540 ( .A1(n14289), .A2(n14210), .ZN(n14211) );
  NAND2_X1 U17541 ( .A1(n14212), .A2(n14211), .ZN(n14282) );
  INV_X1 U17542 ( .A(n14282), .ZN(n16060) );
  INV_X1 U17543 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20825) );
  NOR2_X1 U17544 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14213), .ZN(n14216) );
  INV_X1 U17545 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14214) );
  OAI22_X1 U17546 ( .A1(n14469), .A2(n19974), .B1(n19949), .B2(n14214), .ZN(
        n14215) );
  AOI21_X1 U17547 ( .B1(n19962), .B2(n14216), .A(n14215), .ZN(n14218) );
  NAND2_X1 U17548 ( .A1(n19963), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14217) );
  OAI211_X1 U17549 ( .C1(n15833), .C2(n20825), .A(n14218), .B(n14217), .ZN(
        n14219) );
  AOI21_X1 U17550 ( .B1(n16060), .B2(n19977), .A(n14219), .ZN(n14220) );
  OAI21_X1 U17551 ( .B1(n14380), .B2(n19954), .A(n14220), .ZN(P1_U2816) );
  OAI21_X1 U17552 ( .B1(n14221), .B2(n14223), .A(n14222), .ZN(n14492) );
  NAND2_X1 U17553 ( .A1(n9712), .A2(n14224), .ZN(n14225) );
  NAND2_X1 U17554 ( .A1(n9695), .A2(n14225), .ZN(n16113) );
  AOI22_X1 U17555 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n19963), .B1(n14495), 
        .B2(n19987), .ZN(n14226) );
  OAI21_X1 U17556 ( .B1(n20005), .B2(n16113), .A(n14226), .ZN(n14227) );
  AOI211_X1 U17557 ( .C1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19989), .A(
        n14227), .B(n12840), .ZN(n14234) );
  INV_X1 U17558 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20812) );
  INV_X1 U17559 ( .A(n14241), .ZN(n14228) );
  NOR2_X1 U17560 ( .A1(n19994), .A2(n14228), .ZN(n15904) );
  NAND3_X1 U17561 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n15904), .ZN(n14229) );
  NOR2_X1 U17562 ( .A1(n20812), .A2(n14229), .ZN(n15892) );
  NOR2_X1 U17563 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14229), .ZN(n15898) );
  INV_X1 U17564 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14231) );
  OAI21_X1 U17565 ( .B1(n19994), .B2(n14230), .A(n15872), .ZN(n15910) );
  OR3_X1 U17566 ( .A1(n15898), .A2(n14231), .A3(n15910), .ZN(n14232) );
  OAI21_X1 U17567 ( .B1(n15892), .B2(P1_REIP_REG_16__SCAN_IN), .A(n14232), 
        .ZN(n14233) );
  OAI211_X1 U17568 ( .C1(n14492), .C2(n19954), .A(n14234), .B(n14233), .ZN(
        P1_U2824) );
  NAND2_X1 U17569 ( .A1(n13759), .A2(n14236), .ZN(n14237) );
  NAND2_X1 U17570 ( .A1(n14235), .A2(n14237), .ZN(n14359) );
  OAI21_X1 U17571 ( .B1(n14359), .B2(n14360), .A(n14235), .ZN(n14354) );
  AND2_X1 U17572 ( .A1(n14354), .A2(n14353), .ZN(n14356) );
  OAI21_X1 U17573 ( .B1(n14356), .B2(n14240), .A(n14239), .ZN(n14516) );
  OAI21_X1 U17574 ( .B1(n19994), .B2(n14241), .A(n15872), .ZN(n15921) );
  INV_X1 U17575 ( .A(n14513), .ZN(n14243) );
  INV_X1 U17576 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20810) );
  NAND2_X1 U17577 ( .A1(n15904), .A2(n20810), .ZN(n14242) );
  OAI211_X1 U17578 ( .C1(n14243), .C2(n19974), .A(n14242), .B(n20101), .ZN(
        n14249) );
  INV_X1 U17579 ( .A(n14343), .ZN(n14244) );
  AOI21_X1 U17580 ( .B1(n14245), .B2(n14352), .A(n14244), .ZN(n16136) );
  AOI22_X1 U17581 ( .A1(n16136), .A2(n19977), .B1(n19963), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14246) );
  OAI21_X1 U17582 ( .B1(n14247), .B2(n19949), .A(n14246), .ZN(n14248) );
  AOI211_X1 U17583 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n15921), .A(n14249), 
        .B(n14248), .ZN(n14250) );
  OAI21_X1 U17584 ( .B1(n14516), .B2(n19954), .A(n14250), .ZN(P1_U2827) );
  INV_X1 U17585 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14254) );
  NOR2_X1 U17586 ( .A1(n14251), .A2(n19974), .ZN(n14252) );
  NOR2_X1 U17587 ( .A1(n12840), .A2(n14252), .ZN(n14253) );
  OAI21_X1 U17588 ( .B1(n14254), .B2(n19949), .A(n14253), .ZN(n14258) );
  NOR3_X1 U17589 ( .A1(n19994), .A2(n14256), .A3(n14255), .ZN(n14257) );
  AOI211_X1 U17590 ( .C1(n19963), .C2(P1_EBX_REG_4__SCAN_IN), .A(n14258), .B(
        n14257), .ZN(n14260) );
  NAND2_X1 U17591 ( .A1(n19961), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n14259) );
  OAI211_X1 U17592 ( .C1(n14261), .C2(n20005), .A(n14260), .B(n14259), .ZN(
        n14262) );
  AOI21_X1 U17593 ( .B1(n19991), .B2(n16215), .A(n14262), .ZN(n14263) );
  OAI21_X1 U17594 ( .B1(n14264), .B2(n19990), .A(n14263), .ZN(P1_U2836) );
  INV_X1 U17595 ( .A(n14265), .ZN(n20646) );
  NAND2_X1 U17596 ( .A1(n19977), .A2(n14266), .ZN(n14268) );
  AOI22_X1 U17597 ( .A1(n19987), .A2(n14269), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n15926), .ZN(n14267) );
  OAI211_X1 U17598 ( .C1(n19949), .C2(n14269), .A(n14268), .B(n14267), .ZN(
        n14271) );
  OAI22_X1 U17599 ( .A1(n15883), .A2(n12627), .B1(n19994), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14270) );
  AOI211_X1 U17600 ( .C1(n20646), .C2(n19991), .A(n14271), .B(n14270), .ZN(
        n14272) );
  OAI21_X1 U17601 ( .B1(n14273), .B2(n19990), .A(n14272), .ZN(P1_U2839) );
  INV_X1 U17602 ( .A(n14542), .ZN(n14275) );
  INV_X1 U17603 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14274) );
  OAI22_X1 U17604 ( .A1(n14275), .A2(n14358), .B1(n20014), .B2(n14274), .ZN(
        P1_U2841) );
  OAI222_X1 U17605 ( .A1(n14364), .A2(n14370), .B1(n14276), .B2(n20014), .C1(
        n14571), .C2(n14358), .ZN(P1_U2844) );
  INV_X1 U17606 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14277) );
  OAI222_X1 U17607 ( .A1(n16041), .A2(n14358), .B1(n14277), .B2(n20014), .C1(
        n14440), .C2(n14364), .ZN(P1_U2845) );
  INV_X1 U17608 ( .A(n14452), .ZN(n14375) );
  OAI222_X1 U17609 ( .A1(n16050), .A2(n14358), .B1(n14278), .B2(n20014), .C1(
        n14375), .C2(n14364), .ZN(P1_U2846) );
  INV_X1 U17610 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14280) );
  OAI222_X1 U17611 ( .A1(n14364), .A2(n14460), .B1(n14280), .B2(n20014), .C1(
        n14279), .C2(n14358), .ZN(P1_U2847) );
  OAI22_X1 U17612 ( .A1(n14282), .A2(n14358), .B1(n14281), .B2(n20014), .ZN(
        n14283) );
  AOI21_X1 U17613 ( .B1(n14471), .B2(n20010), .A(n14283), .ZN(n14284) );
  INV_X1 U17614 ( .A(n14284), .ZN(P1_U2848) );
  INV_X1 U17615 ( .A(n14285), .ZN(n14296) );
  INV_X1 U17616 ( .A(n14286), .ZN(n14287) );
  AOI21_X1 U17617 ( .B1(n14300), .B2(n14296), .A(n14287), .ZN(n14288) );
  OR2_X1 U17618 ( .A1(n14289), .A2(n14288), .ZN(n16078) );
  INV_X1 U17619 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14292) );
  OAI21_X1 U17620 ( .B1(n14290), .B2(n14291), .A(n14208), .ZN(n15830) );
  OAI222_X1 U17621 ( .A1(n16078), .A2(n14358), .B1(n14292), .B2(n20014), .C1(
        n15830), .C2(n14364), .ZN(P1_U2849) );
  AND2_X1 U17622 ( .A1(n14293), .A2(n14294), .ZN(n14295) );
  OR2_X1 U17623 ( .A1(n14290), .A2(n14295), .ZN(n14384) );
  XNOR2_X1 U17624 ( .A(n14300), .B(n14296), .ZN(n16082) );
  OAI22_X1 U17625 ( .A1(n16082), .A2(n14358), .B1(n15841), .B2(n20014), .ZN(
        n14297) );
  AOI21_X1 U17626 ( .B1(n15848), .B2(n20010), .A(n14297), .ZN(n14298) );
  INV_X1 U17627 ( .A(n14298), .ZN(P1_U2850) );
  AND2_X1 U17628 ( .A1(n14310), .A2(n14299), .ZN(n14301) );
  OR2_X1 U17629 ( .A1(n14301), .A2(n14300), .ZN(n15856) );
  INV_X1 U17630 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14307) );
  INV_X1 U17631 ( .A(n14311), .ZN(n14303) );
  NAND2_X1 U17632 ( .A1(n14302), .A2(n14303), .ZN(n14305) );
  NAND2_X1 U17633 ( .A1(n14305), .A2(n14304), .ZN(n14306) );
  NAND2_X1 U17634 ( .A1(n14306), .A2(n14293), .ZN(n15965) );
  OAI222_X1 U17635 ( .A1(n14358), .A2(n15856), .B1(n14307), .B2(n20014), .C1(
        n15965), .C2(n14364), .ZN(P1_U2851) );
  NAND2_X1 U17636 ( .A1(n14317), .A2(n14308), .ZN(n14309) );
  NAND2_X1 U17637 ( .A1(n14310), .A2(n14309), .ZN(n15861) );
  INV_X1 U17638 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14313) );
  XNOR2_X1 U17639 ( .A(n14302), .B(n14311), .ZN(n15971) );
  INV_X1 U17640 ( .A(n15971), .ZN(n14312) );
  OAI222_X1 U17641 ( .A1(n15861), .A2(n14358), .B1(n14313), .B2(n20014), .C1(
        n14312), .C2(n14364), .ZN(P1_U2852) );
  NOR2_X1 U17642 ( .A1(n14314), .A2(n14315), .ZN(n14316) );
  OR2_X1 U17643 ( .A1(n14302), .A2(n14316), .ZN(n15871) );
  INV_X1 U17644 ( .A(n14317), .ZN(n14318) );
  AOI21_X1 U17645 ( .B1(n14319), .B2(n14326), .A(n14318), .ZN(n16089) );
  AOI22_X1 U17646 ( .A1(n16089), .A2(n12863), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14362), .ZN(n14320) );
  OAI21_X1 U17647 ( .B1(n15871), .B2(n14364), .A(n14320), .ZN(P1_U2853) );
  AND2_X1 U17648 ( .A1(n14321), .A2(n14322), .ZN(n14323) );
  OR2_X1 U17649 ( .A1(n14323), .A2(n14314), .ZN(n14394) );
  OR2_X1 U17650 ( .A1(n14333), .A2(n14324), .ZN(n14325) );
  NAND2_X1 U17651 ( .A1(n14326), .A2(n14325), .ZN(n16096) );
  OAI22_X1 U17652 ( .A1(n16096), .A2(n14358), .B1(n15884), .B2(n20014), .ZN(
        n14327) );
  AOI21_X1 U17653 ( .B1(n15887), .B2(n20010), .A(n14327), .ZN(n14328) );
  INV_X1 U17654 ( .A(n14328), .ZN(P1_U2854) );
  INV_X1 U17655 ( .A(n14321), .ZN(n14329) );
  AOI21_X1 U17656 ( .B1(n14330), .B2(n14222), .A(n14329), .ZN(n15983) );
  INV_X1 U17657 ( .A(n15983), .ZN(n14398) );
  AND2_X1 U17658 ( .A1(n9695), .A2(n14331), .ZN(n14332) );
  NOR2_X1 U17659 ( .A1(n14333), .A2(n14332), .ZN(n15890) );
  AOI22_X1 U17660 ( .A1(n15890), .A2(n12863), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14362), .ZN(n14334) );
  OAI21_X1 U17661 ( .B1(n14398), .B2(n14364), .A(n14334), .ZN(P1_U2855) );
  INV_X1 U17662 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14335) );
  OAI222_X1 U17663 ( .A1(n16113), .A2(n14358), .B1(n20014), .B2(n14335), .C1(
        n14492), .C2(n14364), .ZN(P1_U2856) );
  AND2_X1 U17664 ( .A1(n14336), .A2(n14337), .ZN(n14338) );
  OR2_X1 U17665 ( .A1(n14338), .A2(n14221), .ZN(n15995) );
  OR2_X1 U17666 ( .A1(n14344), .A2(n14339), .ZN(n14340) );
  AND2_X1 U17667 ( .A1(n9712), .A2(n14340), .ZN(n16119) );
  AOI22_X1 U17668 ( .A1(n16119), .A2(n12863), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14362), .ZN(n14341) );
  OAI21_X1 U17669 ( .B1(n15995), .B2(n14364), .A(n14341), .ZN(P1_U2857) );
  AND2_X1 U17670 ( .A1(n14343), .A2(n14342), .ZN(n14345) );
  OR2_X1 U17671 ( .A1(n14345), .A2(n14344), .ZN(n16133) );
  INV_X1 U17672 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14348) );
  INV_X1 U17673 ( .A(n14336), .ZN(n14346) );
  AOI21_X1 U17674 ( .B1(n14347), .B2(n14239), .A(n14346), .ZN(n14505) );
  INV_X1 U17675 ( .A(n14505), .ZN(n15907) );
  OAI222_X1 U17676 ( .A1(n16133), .A2(n14358), .B1(n20014), .B2(n14348), .C1(
        n15907), .C2(n14364), .ZN(P1_U2858) );
  AOI22_X1 U17677 ( .A1(n16136), .A2(n12863), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14362), .ZN(n14349) );
  OAI21_X1 U17678 ( .B1(n14516), .B2(n14364), .A(n14349), .ZN(P1_U2859) );
  OR2_X1 U17679 ( .A1(n14361), .A2(n14350), .ZN(n14351) );
  NAND2_X1 U17680 ( .A1(n14352), .A2(n14351), .ZN(n15915) );
  INV_X1 U17681 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14357) );
  NOR2_X1 U17682 ( .A1(n14354), .A2(n14353), .ZN(n14355) );
  OAI222_X1 U17683 ( .A1(n15915), .A2(n14358), .B1(n20014), .B2(n14357), .C1(
        n15999), .C2(n14364), .ZN(P1_U2860) );
  XOR2_X1 U17684 ( .A(n14360), .B(n14359), .Z(n16008) );
  INV_X1 U17685 ( .A(n16008), .ZN(n14412) );
  AOI21_X1 U17686 ( .B1(n9721), .B2(n9705), .A(n14361), .ZN(n16142) );
  AOI22_X1 U17687 ( .A1(n16142), .A2(n12863), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14362), .ZN(n14363) );
  OAI21_X1 U17688 ( .B1(n14412), .B2(n14364), .A(n14363), .ZN(P1_U2861) );
  AOI22_X1 U17689 ( .A1(n15949), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15946), .ZN(n14366) );
  MUX2_X1 U17690 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20104), .Z(
        n20060) );
  AOI22_X1 U17691 ( .A1(n9726), .A2(n20060), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n14399), .ZN(n14365) );
  OAI211_X1 U17692 ( .C1(n14367), .C2(n14411), .A(n14366), .B(n14365), .ZN(
        P1_U2874) );
  AOI22_X1 U17693 ( .A1(n15949), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n15946), .ZN(n14369) );
  MUX2_X1 U17694 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20104), .Z(
        n20056) );
  AOI22_X1 U17695 ( .A1(n9726), .A2(n20056), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n14399), .ZN(n14368) );
  OAI211_X1 U17696 ( .C1(n14370), .C2(n14411), .A(n14369), .B(n14368), .ZN(
        P1_U2876) );
  AOI22_X1 U17697 ( .A1(n15949), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15946), .ZN(n14372) );
  MUX2_X1 U17698 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20104), .Z(
        n20054) );
  AOI22_X1 U17699 ( .A1(n9726), .A2(n20054), .B1(BUF1_REG_27__SCAN_IN), .B2(
        n14399), .ZN(n14371) );
  OAI211_X1 U17700 ( .C1(n14440), .C2(n14411), .A(n14372), .B(n14371), .ZN(
        P1_U2877) );
  AOI22_X1 U17701 ( .A1(n15949), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15946), .ZN(n14374) );
  AOI22_X1 U17702 ( .A1(n9726), .A2(n20052), .B1(BUF1_REG_26__SCAN_IN), .B2(
        n14399), .ZN(n14373) );
  OAI211_X1 U17703 ( .C1(n14375), .C2(n14411), .A(n14374), .B(n14373), .ZN(
        P1_U2878) );
  AOI22_X1 U17704 ( .A1(n15949), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n15946), .ZN(n14377) );
  AOI22_X1 U17705 ( .A1(n9726), .A2(n20050), .B1(BUF1_REG_25__SCAN_IN), .B2(
        n14399), .ZN(n14376) );
  OAI211_X1 U17706 ( .C1(n14460), .C2(n14411), .A(n14377), .B(n14376), .ZN(
        P1_U2879) );
  AOI22_X1 U17707 ( .A1(n15949), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15946), .ZN(n14379) );
  AOI22_X1 U17708 ( .A1(n9726), .A2(n20048), .B1(n14399), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14378) );
  OAI211_X1 U17709 ( .C1(n14380), .C2(n14411), .A(n14379), .B(n14378), .ZN(
        P1_U2880) );
  AOI22_X1 U17710 ( .A1(n15949), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15946), .ZN(n14383) );
  AOI22_X1 U17711 ( .A1(n9726), .A2(n14381), .B1(n14399), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14382) );
  OAI211_X1 U17712 ( .C1(n14384), .C2(n14411), .A(n14383), .B(n14382), .ZN(
        P1_U2882) );
  AOI22_X1 U17713 ( .A1(n15949), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15946), .ZN(n14387) );
  AOI22_X1 U17714 ( .A1(n9726), .A2(n14385), .B1(n14399), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14386) );
  OAI211_X1 U17715 ( .C1(n15965), .C2(n14411), .A(n14387), .B(n14386), .ZN(
        P1_U2883) );
  AOI22_X1 U17716 ( .A1(n15949), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15946), .ZN(n14390) );
  AOI22_X1 U17717 ( .A1(n9726), .A2(n14388), .B1(n14399), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14389) );
  OAI211_X1 U17718 ( .C1(n15871), .C2(n14411), .A(n14390), .B(n14389), .ZN(
        P1_U2885) );
  AOI22_X1 U17719 ( .A1(n15949), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15946), .ZN(n14393) );
  AOI22_X1 U17720 ( .A1(n9726), .A2(n14391), .B1(n14399), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14392) );
  OAI211_X1 U17721 ( .C1(n14394), .C2(n14411), .A(n14393), .B(n14392), .ZN(
        P1_U2886) );
  AOI22_X1 U17722 ( .A1(n15949), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15946), .ZN(n14397) );
  AOI22_X1 U17723 ( .A1(n9726), .A2(n14395), .B1(n14399), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14396) );
  OAI211_X1 U17724 ( .C1(n14398), .C2(n14411), .A(n14397), .B(n14396), .ZN(
        P1_U2887) );
  AOI22_X1 U17725 ( .A1(n15949), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15946), .ZN(n14402) );
  AOI22_X1 U17726 ( .A1(n9726), .A2(n14400), .B1(n14399), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14401) );
  OAI211_X1 U17727 ( .C1(n14492), .C2(n14411), .A(n14402), .B(n14401), .ZN(
        P1_U2888) );
  OAI222_X1 U17728 ( .A1(n14411), .A2(n15995), .B1(n14405), .B2(n13333), .C1(
        n14404), .C2(n14403), .ZN(P1_U2889) );
  AOI22_X1 U17729 ( .A1(n14409), .A2(n20060), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15946), .ZN(n14406) );
  OAI21_X1 U17730 ( .B1(n15907), .B2(n14411), .A(n14406), .ZN(P1_U2890) );
  AOI22_X1 U17731 ( .A1(n14409), .A2(n20058), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15946), .ZN(n14407) );
  OAI21_X1 U17732 ( .B1(n14516), .B2(n14411), .A(n14407), .ZN(P1_U2891) );
  AOI22_X1 U17733 ( .A1(n14409), .A2(n20056), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15946), .ZN(n14408) );
  OAI21_X1 U17734 ( .B1(n15999), .B2(n14411), .A(n14408), .ZN(P1_U2892) );
  AOI22_X1 U17735 ( .A1(n14409), .A2(n20054), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15946), .ZN(n14410) );
  OAI21_X1 U17736 ( .B1(n14412), .B2(n14411), .A(n14410), .ZN(P1_U2893) );
  NOR2_X1 U17737 ( .A1(n14413), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14415) );
  NAND2_X1 U17738 ( .A1(n12840), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14553) );
  NAND2_X1 U17739 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14416) );
  OAI211_X1 U17740 ( .C1(n16023), .C2(n14417), .A(n14553), .B(n14416), .ZN(
        n14418) );
  AOI21_X1 U17741 ( .B1(n14419), .B2(n16029), .A(n14418), .ZN(n14420) );
  NOR3_X1 U17742 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14422) );
  NAND4_X1 U17743 ( .A1(n12833), .A2(n14422), .A3(n14421), .A4(n16067), .ZN(
        n14426) );
  NAND3_X1 U17744 ( .A1(n14519), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14425) );
  INV_X1 U17745 ( .A(n15955), .ZN(n14423) );
  AOI21_X1 U17746 ( .B1(n14519), .B2(n14534), .A(n14423), .ZN(n14424) );
  MUX2_X1 U17747 ( .A(n14426), .B(n14425), .S(n14424), .Z(n14427) );
  XNOR2_X1 U17748 ( .A(n14427), .B(n20953), .ZN(n14578) );
  INV_X1 U17749 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20831) );
  NOR2_X1 U17750 ( .A1(n20101), .A2(n20831), .ZN(n14573) );
  AOI21_X1 U17751 ( .B1(n20085), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14573), .ZN(n14428) );
  OAI21_X1 U17752 ( .B1(n16023), .B2(n14429), .A(n14428), .ZN(n14430) );
  AOI21_X1 U17753 ( .B1(n14431), .B2(n16029), .A(n14430), .ZN(n14432) );
  OAI21_X1 U17754 ( .B1(n14578), .B2(n19920), .A(n14432), .ZN(P1_U2971) );
  INV_X1 U17755 ( .A(n14433), .ZN(n14434) );
  NOR2_X1 U17756 ( .A1(n14434), .A2(n12830), .ZN(n14436) );
  MUX2_X1 U17757 ( .A(n14436), .B(n14435), .S(n12833), .Z(n14437) );
  OAI22_X1 U17758 ( .A1(n16033), .A2(n14439), .B1(n20101), .B2(n14438), .ZN(
        n14442) );
  NOR2_X1 U17759 ( .A1(n14440), .A2(n20106), .ZN(n14441) );
  OAI21_X1 U17760 ( .B1(n19920), .B2(n16038), .A(n14444), .ZN(P1_U2972) );
  INV_X1 U17761 ( .A(n14534), .ZN(n14445) );
  AOI21_X1 U17762 ( .B1(n15955), .B2(n14445), .A(n12833), .ZN(n14446) );
  NOR2_X1 U17763 ( .A1(n14447), .A2(n14446), .ZN(n14448) );
  XNOR2_X1 U17764 ( .A(n14448), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16042) );
  INV_X1 U17765 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20829) );
  NOR2_X1 U17766 ( .A1(n20101), .A2(n20829), .ZN(n16043) );
  AOI21_X1 U17767 ( .B1(n20085), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16043), .ZN(n14449) );
  OAI21_X1 U17768 ( .B1(n16023), .B2(n14450), .A(n14449), .ZN(n14451) );
  AOI21_X1 U17769 ( .B1(n14452), .B2(n16029), .A(n14451), .ZN(n14453) );
  OAI21_X1 U17770 ( .B1(n19920), .B2(n16042), .A(n14453), .ZN(P1_U2973) );
  MUX2_X1 U17771 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14455), .S(
        n15975), .Z(n14456) );
  OAI21_X1 U17772 ( .B1(n14466), .B2(n16067), .A(n14456), .ZN(n14457) );
  XOR2_X1 U17773 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n14457), .Z(
        n16052) );
  OAI22_X1 U17774 ( .A1(n16033), .A2(n14459), .B1(n20101), .B2(n14458), .ZN(
        n14462) );
  NOR2_X1 U17775 ( .A1(n14460), .A2(n20106), .ZN(n14461) );
  AOI211_X1 U17776 ( .C1(n16027), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n14464) );
  OAI21_X1 U17777 ( .B1(n19920), .B2(n16052), .A(n14464), .ZN(P1_U2974) );
  NOR2_X1 U17778 ( .A1(n14466), .A2(n15955), .ZN(n14465) );
  MUX2_X1 U17779 ( .A(n14466), .B(n14465), .S(n15975), .Z(n14467) );
  XNOR2_X1 U17780 ( .A(n14467), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16059) );
  AOI22_X1 U17781 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n14468) );
  OAI21_X1 U17782 ( .B1(n16023), .B2(n14469), .A(n14468), .ZN(n14470) );
  AOI21_X1 U17783 ( .B1(n14471), .B2(n16029), .A(n14470), .ZN(n14472) );
  OAI21_X1 U17784 ( .B1(n19920), .B2(n16059), .A(n14472), .ZN(P1_U2975) );
  NAND2_X1 U17785 ( .A1(n14473), .A2(n14474), .ZN(n14475) );
  XNOR2_X1 U17786 ( .A(n14475), .B(n16081), .ZN(n16083) );
  INV_X1 U17787 ( .A(n15844), .ZN(n14477) );
  AOI22_X1 U17788 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14476) );
  OAI21_X1 U17789 ( .B1(n16023), .B2(n14477), .A(n14476), .ZN(n14478) );
  AOI21_X1 U17790 ( .B1(n15848), .B2(n16029), .A(n14478), .ZN(n14479) );
  OAI21_X1 U17791 ( .B1(n19920), .B2(n16083), .A(n14479), .ZN(P1_U2977) );
  OR2_X1 U17792 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U17793 ( .A1(n14480), .A2(n14483), .ZN(n16097) );
  INV_X1 U17794 ( .A(n15886), .ZN(n14485) );
  AOI22_X1 U17795 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14484) );
  OAI21_X1 U17796 ( .B1(n16023), .B2(n14485), .A(n14484), .ZN(n14486) );
  AOI21_X1 U17797 ( .B1(n15887), .B2(n16029), .A(n14486), .ZN(n14487) );
  OAI21_X1 U17798 ( .B1(n19920), .B2(n16097), .A(n14487), .ZN(P1_U2981) );
  NOR2_X1 U17799 ( .A1(n14488), .A2(n14489), .ZN(n15989) );
  OAI21_X1 U17800 ( .B1(n15989), .B2(n14590), .A(n15990), .ZN(n14490) );
  XOR2_X1 U17801 ( .A(n14491), .B(n14490), .Z(n16105) );
  OAI22_X1 U17802 ( .A1(n16033), .A2(n20915), .B1(n20101), .B2(n14231), .ZN(
        n14494) );
  NOR2_X1 U17803 ( .A1(n14492), .A2(n20106), .ZN(n14493) );
  AOI211_X1 U17804 ( .C1(n16027), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        n14496) );
  OAI21_X1 U17805 ( .B1(n19920), .B2(n16105), .A(n14496), .ZN(P1_U2983) );
  MUX2_X1 U17806 ( .A(n12819), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n14519), .Z(n14501) );
  AOI21_X1 U17807 ( .B1(n14488), .B2(n14498), .A(n14497), .ZN(n14499) );
  AOI21_X1 U17808 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n12833), .A(
        n14499), .ZN(n14500) );
  XOR2_X1 U17809 ( .A(n14501), .B(n14500), .Z(n16122) );
  INV_X1 U17810 ( .A(n15911), .ZN(n14503) );
  AOI22_X1 U17811 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14502) );
  OAI21_X1 U17812 ( .B1(n16023), .B2(n14503), .A(n14502), .ZN(n14504) );
  AOI21_X1 U17813 ( .B1(n14505), .B2(n16029), .A(n14504), .ZN(n14506) );
  OAI21_X1 U17814 ( .B1(n16122), .B2(n19920), .A(n14506), .ZN(P1_U2985) );
  INV_X1 U17815 ( .A(n14488), .ZN(n14591) );
  AOI21_X1 U17816 ( .B1(n14591), .B2(n14508), .A(n14507), .ZN(n14606) );
  AND2_X1 U17817 ( .A1(n14509), .A2(n14510), .ZN(n14605) );
  NAND2_X1 U17818 ( .A1(n14606), .A2(n14605), .ZN(n14604) );
  NAND2_X1 U17819 ( .A1(n14604), .A2(n14510), .ZN(n14512) );
  XNOR2_X1 U17820 ( .A(n14512), .B(n14511), .ZN(n16138) );
  AOI22_X1 U17821 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14515) );
  NAND2_X1 U17822 ( .A1(n16027), .A2(n14513), .ZN(n14514) );
  OAI211_X1 U17823 ( .C1(n14516), .C2(n20106), .A(n14515), .B(n14514), .ZN(
        n14517) );
  AOI21_X1 U17824 ( .B1(n16138), .B2(n20087), .A(n14517), .ZN(n14518) );
  INV_X1 U17825 ( .A(n14518), .ZN(P1_U2986) );
  AND2_X1 U17826 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14521) );
  XNOR2_X1 U17827 ( .A(n14488), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14520) );
  MUX2_X1 U17828 ( .A(n14521), .B(n14520), .S(n14519), .Z(n14523) );
  NOR3_X1 U17829 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14579), .ZN(n16005) );
  NOR2_X1 U17830 ( .A1(n14523), .A2(n16005), .ZN(n16149) );
  AOI22_X1 U17831 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14524) );
  OAI21_X1 U17832 ( .B1(n16023), .B2(n15934), .A(n14524), .ZN(n14525) );
  AOI21_X1 U17833 ( .B1(n15938), .B2(n16029), .A(n14525), .ZN(n14526) );
  OAI21_X1 U17834 ( .B1(n16149), .B2(n19920), .A(n14526), .ZN(P1_U2989) );
  AOI21_X1 U17835 ( .B1(n15814), .B2(n14527), .A(n14547), .ZN(n14533) );
  NOR2_X1 U17836 ( .A1(n14584), .A2(n16081), .ZN(n14543) );
  INV_X1 U17837 ( .A(n14546), .ZN(n16062) );
  INV_X1 U17838 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16107) );
  NOR4_X1 U17839 ( .A1(n12819), .A2(n16115), .A3(n16107), .A4(n14595), .ZN(
        n16102) );
  NAND2_X1 U17840 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16102), .ZN(
        n14545) );
  NAND3_X1 U17841 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U17842 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16152) );
  NOR2_X1 U17843 ( .A1(n16123), .A2(n16152), .ZN(n14612) );
  NAND2_X1 U17844 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14612), .ZN(
        n14615) );
  NOR2_X1 U17845 ( .A1(n16127), .A2(n14615), .ZN(n14530) );
  NOR2_X1 U17846 ( .A1(n16205), .A2(n16174), .ZN(n14608) );
  AND2_X1 U17847 ( .A1(n14608), .A2(n14528), .ZN(n14611) );
  NAND2_X1 U17848 ( .A1(n14530), .A2(n14611), .ZN(n15812) );
  INV_X1 U17849 ( .A(n15812), .ZN(n16135) );
  NAND2_X1 U17850 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16135), .ZN(
        n14599) );
  NOR2_X1 U17851 ( .A1(n14545), .A2(n14599), .ZN(n14532) );
  NAND2_X1 U17852 ( .A1(n14529), .A2(n14608), .ZN(n16124) );
  INV_X1 U17853 ( .A(n16124), .ZN(n14609) );
  NAND2_X1 U17854 ( .A1(n14609), .A2(n14530), .ZN(n15813) );
  NOR2_X1 U17855 ( .A1(n12820), .A2(n15813), .ZN(n14597) );
  INV_X1 U17856 ( .A(n14597), .ZN(n14544) );
  OAI21_X1 U17857 ( .B1(n14544), .B2(n14545), .A(n16063), .ZN(n14531) );
  OAI211_X1 U17858 ( .C1(n14613), .C2(n14532), .A(n14610), .B(n14531), .ZN(
        n16093) );
  NAND2_X1 U17859 ( .A1(n14600), .A2(n14610), .ZN(n16150) );
  OAI21_X1 U17860 ( .B1(n16062), .B2(n16093), .A(n16150), .ZN(n16080) );
  OAI21_X1 U17861 ( .B1(n14600), .B2(n14543), .A(n16080), .ZN(n16074) );
  AOI211_X1 U17862 ( .C1(n20098), .C2(n14534), .A(n14533), .B(n16074), .ZN(
        n16058) );
  NAND2_X1 U17863 ( .A1(n16058), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16046) );
  INV_X1 U17864 ( .A(n16046), .ZN(n14536) );
  INV_X1 U17865 ( .A(n16058), .ZN(n14535) );
  INV_X1 U17866 ( .A(n14600), .ZN(n16177) );
  NOR2_X1 U17867 ( .A1(n14535), .A2(n16177), .ZN(n14565) );
  AOI21_X1 U17868 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14536), .A(
        n14565), .ZN(n16039) );
  NOR2_X1 U17869 ( .A1(n16039), .A2(n14537), .ZN(n14564) );
  INV_X1 U17870 ( .A(n14548), .ZN(n14575) );
  NAND2_X1 U17871 ( .A1(n14564), .A2(n14575), .ZN(n14539) );
  INV_X1 U17872 ( .A(n14565), .ZN(n14538) );
  INV_X1 U17873 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14552) );
  AOI21_X1 U17874 ( .B1(n14539), .B2(n14538), .A(n14552), .ZN(n14550) );
  NOR3_X1 U17875 ( .A1(n14550), .A2(n14565), .A3(n12873), .ZN(n14540) );
  INV_X1 U17876 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16057) );
  INV_X1 U17877 ( .A(n14543), .ZN(n16079) );
  OAI22_X1 U17878 ( .A1(n15814), .A2(n14544), .B1(n14599), .B2(n16176), .ZN(
        n16100) );
  NAND2_X1 U17879 ( .A1(n14547), .A2(n16068), .ZN(n16045) );
  INV_X1 U17880 ( .A(n14550), .ZN(n14557) );
  NAND2_X1 U17881 ( .A1(n14552), .A2(n14551), .ZN(n14556) );
  OAI21_X1 U17882 ( .B1(n14554), .B2(n16159), .A(n14553), .ZN(n14555) );
  AOI21_X1 U17883 ( .B1(n14557), .B2(n14556), .A(n14555), .ZN(n14558) );
  OAI21_X1 U17884 ( .B1(n14559), .B2(n16204), .A(n14558), .ZN(P1_U3001) );
  INV_X1 U17885 ( .A(n14560), .ZN(n14563) );
  INV_X1 U17886 ( .A(n14561), .ZN(n14562) );
  AOI21_X1 U17887 ( .B1(n14563), .B2(n20093), .A(n14562), .ZN(n14569) );
  OAI21_X1 U17888 ( .B1(n14575), .B2(n14565), .A(n14564), .ZN(n14566) );
  OAI21_X1 U17889 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14567), .A(
        n14566), .ZN(n14568) );
  OAI211_X1 U17890 ( .C1(n14570), .C2(n16204), .A(n14569), .B(n14568), .ZN(
        P1_U3002) );
  NOR2_X1 U17891 ( .A1(n14571), .A2(n16159), .ZN(n14572) );
  AOI211_X1 U17892 ( .C1(n16039), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14573), .B(n14572), .ZN(n14577) );
  OR3_X1 U17893 ( .A1(n16035), .A2(n14575), .A3(n14574), .ZN(n14576) );
  OAI211_X1 U17894 ( .C1(n14578), .C2(n16204), .A(n14577), .B(n14576), .ZN(
        P1_U3003) );
  NAND2_X1 U17895 ( .A1(n14579), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14580) );
  OR2_X1 U17896 ( .A1(n14480), .A2(n14580), .ZN(n14582) );
  OAI21_X1 U17897 ( .B1(n14581), .B2(n14579), .A(n14582), .ZN(n15808) );
  NAND2_X1 U17898 ( .A1(n15808), .A2(n15816), .ZN(n15807) );
  OAI22_X1 U17899 ( .A1(n15807), .A2(n14579), .B1(n15816), .B2(n14582), .ZN(
        n14583) );
  XNOR2_X1 U17900 ( .A(n14583), .B(n14584), .ZN(n15960) );
  INV_X1 U17901 ( .A(n15960), .ZN(n14588) );
  INV_X1 U17902 ( .A(n15856), .ZN(n14586) );
  NAND2_X1 U17903 ( .A1(n12840), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15967) );
  OAI221_X1 U17904 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n16088), 
        .C1(n14584), .C2(n16080), .A(n15967), .ZN(n14585) );
  AOI21_X1 U17905 ( .B1(n14586), .B2(n20093), .A(n14585), .ZN(n14587) );
  OAI21_X1 U17906 ( .B1(n14588), .B2(n16204), .A(n14587), .ZN(P1_U3010) );
  OAI21_X1 U17907 ( .B1(n14591), .B2(n14590), .A(n14589), .ZN(n14593) );
  NAND2_X1 U17908 ( .A1(n14593), .A2(n16107), .ZN(n14592) );
  MUX2_X1 U17909 ( .A(n14593), .B(n14592), .S(n15975), .Z(n14594) );
  XNOR2_X1 U17910 ( .A(n14594), .B(n14595), .ZN(n15986) );
  AOI22_X1 U17911 ( .A1(n15890), .A2(n20093), .B1(n12840), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14603) );
  NAND2_X1 U17912 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U17913 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16100), .ZN(
        n16106) );
  OAI21_X1 U17914 ( .B1(n14596), .B2(n16106), .A(n14595), .ZN(n14601) );
  INV_X1 U17915 ( .A(n14613), .ZN(n16175) );
  OAI21_X1 U17916 ( .B1(n14597), .B2(n15814), .A(n14610), .ZN(n14598) );
  AOI21_X1 U17917 ( .B1(n16175), .B2(n14599), .A(n14598), .ZN(n16128) );
  OAI21_X1 U17918 ( .B1(n14600), .B2(n16102), .A(n16128), .ZN(n16099) );
  NAND2_X1 U17919 ( .A1(n14601), .A2(n16099), .ZN(n14602) );
  OAI211_X1 U17920 ( .C1(n15986), .C2(n16204), .A(n14603), .B(n14602), .ZN(
        P1_U3014) );
  OAI21_X1 U17921 ( .B1(n14606), .B2(n14605), .A(n14604), .ZN(n14607) );
  INV_X1 U17922 ( .A(n14607), .ZN(n16004) );
  NAND2_X1 U17923 ( .A1(n14608), .A2(n16201), .ZN(n16200) );
  NOR2_X1 U17924 ( .A1(n14615), .A2(n16200), .ZN(n14618) );
  NOR2_X1 U17925 ( .A1(n14609), .A2(n15814), .ZN(n16173) );
  OAI221_X1 U17926 ( .B1(n14613), .B2(n14612), .C1(n14613), .C2(n14611), .A(
        n14610), .ZN(n14614) );
  AOI211_X1 U17927 ( .C1(n16063), .C2(n14615), .A(n16173), .B(n14614), .ZN(
        n16148) );
  OAI21_X1 U17928 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16176), .A(
        n16148), .ZN(n14617) );
  OAI22_X1 U17929 ( .A1(n20101), .A2(n15919), .B1(n16159), .B2(n15915), .ZN(
        n14616) );
  AOI221_X1 U17930 ( .B1(n14618), .B2(n16127), .C1(n14617), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n14616), .ZN(n14619) );
  OAI21_X1 U17931 ( .B1(n16004), .B2(n16204), .A(n14619), .ZN(P1_U3019) );
  OAI21_X1 U17932 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9615), .A(n20713), 
        .ZN(n14620) );
  OAI21_X1 U17933 ( .B1(n14265), .B2(n14621), .A(n14620), .ZN(n14622) );
  MUX2_X1 U17934 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14622), .S(
        n20102), .Z(P1_U3477) );
  NOR2_X1 U17935 ( .A1(n15760), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14625) );
  NOR3_X1 U17936 ( .A1(n14623), .A2(n13489), .A3(n14627), .ZN(n14624) );
  AOI211_X1 U17937 ( .C1(n20646), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        n15762) );
  OAI22_X1 U17938 ( .A1(n12873), .A2(n12626), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14631) );
  NOR2_X1 U17939 ( .A1(n20776), .A2(n20082), .ZN(n14633) );
  NOR3_X1 U17940 ( .A1(n13489), .A2(n14627), .A3(n14639), .ZN(n14628) );
  AOI21_X1 U17941 ( .B1(n14631), .B2(n14633), .A(n14628), .ZN(n14629) );
  OAI21_X1 U17942 ( .B1(n15762), .B2(n14641), .A(n14629), .ZN(n14630) );
  MUX2_X1 U17943 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14630), .S(
        n16216), .Z(P1_U3473) );
  INV_X1 U17944 ( .A(n14631), .ZN(n14632) );
  AOI22_X1 U17945 ( .A1(n14634), .A2(n15785), .B1(n14633), .B2(n14632), .ZN(
        n14635) );
  OAI21_X1 U17946 ( .B1(n14636), .B2(n14641), .A(n14635), .ZN(n14637) );
  MUX2_X1 U17947 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14637), .S(
        n16216), .Z(P1_U3472) );
  INV_X1 U17948 ( .A(n14638), .ZN(n14640) );
  OAI22_X1 U17949 ( .A1(n14642), .A2(n14641), .B1(n14640), .B2(n14639), .ZN(
        n14643) );
  MUX2_X1 U17950 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14643), .S(
        n16216), .Z(P1_U3469) );
  INV_X1 U17951 ( .A(n14130), .ZN(n14644) );
  NAND2_X1 U17952 ( .A1(n14644), .A2(n19122), .ZN(n14680) );
  XOR2_X1 U17953 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n14647), .Z(
        n15003) );
  NOR2_X1 U17954 ( .A1(n14645), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14646) );
  OR2_X1 U17955 ( .A1(n14647), .A2(n14646), .ZN(n15016) );
  INV_X1 U17956 ( .A(n15016), .ZN(n16232) );
  INV_X1 U17957 ( .A(n14648), .ZN(n14691) );
  INV_X1 U17958 ( .A(n14649), .ZN(n14650) );
  AOI21_X1 U17959 ( .B1(n15026), .B2(n14651), .A(n14650), .ZN(n15029) );
  INV_X1 U17960 ( .A(n14651), .ZN(n14652) );
  AOI21_X1 U17961 ( .B1(n15038), .B2(n14671), .A(n14652), .ZN(n15040) );
  AOI21_X1 U17962 ( .B1(n15059), .B2(n14668), .A(n9683), .ZN(n15061) );
  INV_X1 U17963 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15099) );
  AOI21_X1 U17964 ( .B1(n14667), .B2(n15099), .A(n14669), .ZN(n15097) );
  AOI21_X1 U17965 ( .B1(n18978), .B2(n14665), .A(n9679), .ZN(n18977) );
  NOR2_X1 U17966 ( .A1(n14662), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14653) );
  OR2_X1 U17967 ( .A1(n14666), .A2(n14653), .ZN(n19014) );
  INV_X1 U17968 ( .A(n19014), .ZN(n14664) );
  AOI21_X1 U17969 ( .B1(n15166), .B2(n9638), .A(n9849), .ZN(n19020) );
  AOI21_X1 U17970 ( .B1(n14657), .B2(n15194), .A(n14659), .ZN(n19043) );
  AOI21_X1 U17971 ( .B1(n14654), .B2(n14656), .A(n14658), .ZN(n19050) );
  NAND2_X1 U17972 ( .A1(n14655), .A2(n16296), .ZN(n19070) );
  NOR2_X1 U17973 ( .A1(n19071), .A2(n19070), .ZN(n19063) );
  OAI21_X1 U17974 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9680), .A(
        n14656), .ZN(n19064) );
  NAND2_X1 U17975 ( .A1(n19063), .A2(n19064), .ZN(n19049) );
  NOR2_X1 U17976 ( .A1(n19050), .A2(n19049), .ZN(n14816) );
  OAI21_X1 U17977 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n14658), .A(
        n14657), .ZN(n15202) );
  NAND2_X1 U17978 ( .A1(n14816), .A2(n15202), .ZN(n19042) );
  NOR2_X1 U17979 ( .A1(n19043), .A2(n19042), .ZN(n19026) );
  OR2_X1 U17980 ( .A1(n14659), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14660) );
  NAND2_X1 U17981 ( .A1(n9638), .A2(n14660), .ZN(n19027) );
  NAND2_X1 U17982 ( .A1(n19026), .A2(n19027), .ZN(n19019) );
  NOR2_X1 U17983 ( .A1(n19020), .A2(n19019), .ZN(n14804) );
  AND2_X1 U17984 ( .A1(n14661), .A2(n15155), .ZN(n14663) );
  OR2_X1 U17985 ( .A1(n14663), .A2(n14662), .ZN(n15152) );
  NAND2_X1 U17986 ( .A1(n14804), .A2(n15152), .ZN(n19001) );
  NOR2_X1 U17987 ( .A1(n14664), .A2(n19001), .ZN(n18988) );
  OAI21_X1 U17988 ( .B1(n14666), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14665), .ZN(n18989) );
  NAND2_X1 U17989 ( .A1(n18988), .A2(n18989), .ZN(n18975) );
  NOR2_X1 U17990 ( .A1(n18977), .A2(n18975), .ZN(n18961) );
  OAI21_X1 U17991 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9679), .A(
        n14667), .ZN(n18962) );
  NAND2_X1 U17992 ( .A1(n18961), .A2(n18962), .ZN(n14794) );
  NOR2_X1 U17993 ( .A1(n15097), .A2(n14794), .ZN(n14776) );
  OAI21_X1 U17994 ( .B1(n14669), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14668), .ZN(n15072) );
  NAND2_X1 U17995 ( .A1(n14776), .A2(n15072), .ZN(n14762) );
  NOR2_X1 U17996 ( .A1(n15061), .A2(n14762), .ZN(n14743) );
  OR2_X1 U17997 ( .A1(n9683), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14670) );
  AND2_X1 U17998 ( .A1(n14671), .A2(n14670), .ZN(n14746) );
  INV_X1 U17999 ( .A(n14746), .ZN(n15051) );
  NAND2_X1 U18000 ( .A1(n14743), .A2(n15051), .ZN(n14729) );
  OAI21_X1 U18001 ( .B1(n15040), .B2(n14729), .A(n19118), .ZN(n14672) );
  NOR2_X1 U18002 ( .A1(n19102), .A2(n14700), .ZN(n14690) );
  NOR2_X1 U18003 ( .A1(n14691), .A2(n14690), .ZN(n14689) );
  NOR2_X1 U18004 ( .A1(n19102), .A2(n14689), .ZN(n16231) );
  NOR2_X1 U18005 ( .A1(n16232), .A2(n16231), .ZN(n16230) );
  NOR2_X1 U18006 ( .A1(n19102), .A2(n16230), .ZN(n14682) );
  NOR2_X1 U18007 ( .A1(n15003), .A2(n14682), .ZN(n14681) );
  AOI22_X1 U18008 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19109), .B1(
        n14795), .B2(n14681), .ZN(n14679) );
  INV_X1 U18009 ( .A(n14673), .ZN(n19160) );
  INV_X1 U18010 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20991) );
  OAI22_X1 U18011 ( .A1(n11561), .A2(n14674), .B1(n19096), .B2(n20991), .ZN(
        n14675) );
  AOI21_X1 U18012 ( .B1(n19160), .B2(n14829), .A(n14675), .ZN(n14678) );
  NAND2_X1 U18013 ( .A1(n14676), .A2(n19086), .ZN(n14677) );
  NAND4_X1 U18014 ( .A1(n14680), .A2(n14679), .A3(n14678), .A4(n14677), .ZN(
        P2_U2824) );
  AOI211_X1 U18015 ( .C1(n15003), .C2(n14682), .A(n14681), .B(n19782), .ZN(
        n14685) );
  AOI22_X1 U18016 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19109), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19116), .ZN(n14683) );
  INV_X1 U18017 ( .A(n14683), .ZN(n14684) );
  AOI211_X1 U18018 ( .C1(P2_EBX_REG_30__SCAN_IN), .C2(n19110), .A(n14685), .B(
        n14684), .ZN(n14688) );
  AOI22_X1 U18019 ( .A1(n11586), .A2(n19086), .B1(n14686), .B2(n14829), .ZN(
        n14687) );
  OAI211_X1 U18020 ( .C1(n9575), .C2(n19090), .A(n14688), .B(n14687), .ZN(
        P2_U2825) );
  AOI211_X1 U18021 ( .C1(n14691), .C2(n14690), .A(n14689), .B(n19782), .ZN(
        n14694) );
  AOI22_X1 U18022 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19109), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19116), .ZN(n14692) );
  INV_X1 U18023 ( .A(n14692), .ZN(n14693) );
  AOI211_X1 U18024 ( .C1(P2_EBX_REG_28__SCAN_IN), .C2(n19110), .A(n14694), .B(
        n14693), .ZN(n14698) );
  OAI22_X1 U18025 ( .A1(n14695), .A2(n19112), .B1(n14928), .B2(n19127), .ZN(
        n14696) );
  INV_X1 U18026 ( .A(n14696), .ZN(n14697) );
  OAI211_X1 U18027 ( .C1(n14848), .C2(n19090), .A(n14698), .B(n14697), .ZN(
        P2_U2827) );
  AOI211_X1 U18028 ( .C1(n14702), .C2(n14701), .A(n14700), .B(n19782), .ZN(
        n14705) );
  OAI22_X1 U18029 ( .A1(n14703), .A2(n19084), .B1(n19850), .B2(n19096), .ZN(
        n14704) );
  AOI211_X1 U18030 ( .C1(P2_EBX_REG_27__SCAN_IN), .C2(n19110), .A(n14705), .B(
        n14704), .ZN(n14710) );
  INV_X1 U18031 ( .A(n14706), .ZN(n14943) );
  OAI22_X1 U18032 ( .A1(n14707), .A2(n19112), .B1(n14943), .B2(n19127), .ZN(
        n14708) );
  INV_X1 U18033 ( .A(n14708), .ZN(n14709) );
  OAI211_X1 U18034 ( .C1(n14856), .C2(n19090), .A(n14710), .B(n14709), .ZN(
        P2_U2828) );
  NOR2_X1 U18035 ( .A1(n14728), .A2(n14711), .ZN(n14712) );
  AOI211_X1 U18036 ( .C1(n15029), .C2(n14714), .A(n14713), .B(n19782), .ZN(
        n14717) );
  INV_X1 U18037 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19847) );
  OAI22_X1 U18038 ( .A1(n19097), .A2(n14715), .B1(n19847), .B2(n19096), .ZN(
        n14716) );
  AOI211_X1 U18039 ( .C1(n19109), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14717), .B(n14716), .ZN(n14722) );
  NAND2_X1 U18040 ( .A1(n14719), .A2(n14718), .ZN(n14720) );
  AND2_X1 U18041 ( .A1(n9627), .A2(n14720), .ZN(n15254) );
  NAND2_X1 U18042 ( .A1(n15254), .A2(n14829), .ZN(n14721) );
  NAND2_X1 U18043 ( .A1(n14722), .A2(n14721), .ZN(n14723) );
  AOI21_X1 U18044 ( .B1(n14724), .B2(n19086), .A(n14723), .ZN(n14725) );
  OAI21_X1 U18045 ( .B1(n15250), .B2(n19090), .A(n14725), .ZN(P2_U2829) );
  NOR2_X1 U18046 ( .A1(n14741), .A2(n14726), .ZN(n14727) );
  OR2_X1 U18047 ( .A1(n14728), .A2(n14727), .ZN(n15274) );
  AND2_X1 U18048 ( .A1(n19118), .A2(n14729), .ZN(n14731) );
  OAI21_X1 U18049 ( .B1(n15040), .B2(n14731), .A(n19123), .ZN(n14730) );
  AOI21_X1 U18050 ( .B1(n15040), .B2(n14731), .A(n14730), .ZN(n14733) );
  OAI22_X1 U18051 ( .A1(n15038), .A2(n19084), .B1(n19845), .B2(n19096), .ZN(
        n14732) );
  AOI211_X1 U18052 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n19110), .A(n14733), .B(
        n14732), .ZN(n14739) );
  XNOR2_X1 U18053 ( .A(n14734), .B(n14735), .ZN(n15267) );
  INV_X1 U18054 ( .A(n15267), .ZN(n14736) );
  AOI22_X1 U18055 ( .A1(n14737), .A2(n19086), .B1(n14829), .B2(n14736), .ZN(
        n14738) );
  OAI211_X1 U18056 ( .C1(n15274), .C2(n19090), .A(n14739), .B(n14738), .ZN(
        P2_U2830) );
  AND2_X1 U18057 ( .A1(n14761), .A2(n14740), .ZN(n14742) );
  OR2_X1 U18058 ( .A1(n14742), .A2(n14741), .ZN(n15279) );
  NOR2_X1 U18059 ( .A1(n19102), .A2(n14743), .ZN(n14745) );
  OAI21_X1 U18060 ( .B1(n14746), .B2(n14745), .A(n19123), .ZN(n14744) );
  AOI21_X1 U18061 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n14749) );
  INV_X1 U18062 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19843) );
  OAI22_X1 U18063 ( .A1(n19097), .A2(n14747), .B1(n19843), .B2(n19096), .ZN(
        n14748) );
  AOI211_X1 U18064 ( .C1(n19109), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14749), .B(n14748), .ZN(n14757) );
  INV_X1 U18065 ( .A(n14750), .ZN(n14755) );
  INV_X1 U18066 ( .A(n14734), .ZN(n14753) );
  NAND2_X1 U18067 ( .A1(n14766), .A2(n14751), .ZN(n14752) );
  NAND2_X1 U18068 ( .A1(n14753), .A2(n14752), .ZN(n15285) );
  INV_X1 U18069 ( .A(n15285), .ZN(n14754) );
  AOI22_X1 U18070 ( .A1(n14755), .A2(n19086), .B1(n14829), .B2(n14754), .ZN(
        n14756) );
  OAI211_X1 U18071 ( .C1(n15279), .C2(n19090), .A(n14757), .B(n14756), .ZN(
        P2_U2831) );
  NAND2_X1 U18072 ( .A1(n14758), .A2(n14759), .ZN(n14760) );
  NAND2_X1 U18073 ( .A1(n14761), .A2(n14760), .ZN(n16241) );
  NAND2_X1 U18074 ( .A1(n19118), .A2(n14762), .ZN(n14763) );
  XNOR2_X1 U18075 ( .A(n15061), .B(n14763), .ZN(n14764) );
  AOI22_X1 U18076 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19110), .B1(n19123), 
        .B2(n14764), .ZN(n14774) );
  INV_X1 U18077 ( .A(n14766), .ZN(n14767) );
  AOI21_X1 U18078 ( .B1(n14768), .B2(n14765), .A(n14767), .ZN(n15292) );
  INV_X1 U18079 ( .A(n15292), .ZN(n14770) );
  AOI22_X1 U18080 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19109), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19116), .ZN(n14769) );
  OAI21_X1 U18081 ( .B1(n14770), .B2(n19127), .A(n14769), .ZN(n14771) );
  AOI21_X1 U18082 ( .B1(n14772), .B2(n19086), .A(n14771), .ZN(n14773) );
  OAI211_X1 U18083 ( .C1(n16241), .C2(n19090), .A(n14774), .B(n14773), .ZN(
        P2_U2832) );
  OAI21_X1 U18084 ( .B1(n14786), .B2(n14775), .A(n14758), .ZN(n16248) );
  NOR2_X1 U18085 ( .A1(n19102), .A2(n14776), .ZN(n14777) );
  XOR2_X1 U18086 ( .A(n15072), .B(n14777), .Z(n14779) );
  AOI22_X1 U18087 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19109), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19116), .ZN(n14778) );
  OAI21_X1 U18088 ( .B1(n19782), .B2(n14779), .A(n14778), .ZN(n14780) );
  AOI21_X1 U18089 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n19110), .A(n14780), .ZN(
        n14785) );
  OR2_X1 U18090 ( .A1(n14789), .A2(n14781), .ZN(n14782) );
  NAND2_X1 U18091 ( .A1(n14765), .A2(n14782), .ZN(n15304) );
  INV_X1 U18092 ( .A(n15304), .ZN(n16260) );
  AOI22_X1 U18093 ( .A1(n14783), .A2(n19086), .B1(n16260), .B2(n14829), .ZN(
        n14784) );
  OAI211_X1 U18094 ( .C1(n16248), .C2(n19090), .A(n14785), .B(n14784), .ZN(
        P2_U2833) );
  AOI21_X1 U18095 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n15324) );
  INV_X1 U18096 ( .A(n15324), .ZN(n14800) );
  AOI21_X1 U18097 ( .B1(n19118), .B2(n14794), .A(n19782), .ZN(n14798) );
  AOI21_X1 U18098 ( .B1(n14790), .B2(n15332), .A(n14789), .ZN(n15316) );
  INV_X1 U18099 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19837) );
  OAI22_X1 U18100 ( .A1(n15099), .A2(n19084), .B1(n19837), .B2(n19096), .ZN(
        n14791) );
  AOI21_X1 U18101 ( .B1(n15316), .B2(n14829), .A(n14791), .ZN(n14792) );
  OAI21_X1 U18102 ( .B1(n14793), .B2(n19112), .A(n14792), .ZN(n14797) );
  NAND2_X1 U18103 ( .A1(n14795), .A2(n14794), .ZN(n18964) );
  OAI22_X1 U18104 ( .A1(n15097), .A2(n18964), .B1(n19097), .B2(n14879), .ZN(
        n14796) );
  AOI211_X1 U18105 ( .C1(n15097), .C2(n14798), .A(n14797), .B(n14796), .ZN(
        n14799) );
  OAI21_X1 U18106 ( .B1(n14800), .B2(n19090), .A(n14799), .ZN(P2_U2834) );
  INV_X1 U18107 ( .A(n14801), .ZN(n14906) );
  AND2_X1 U18108 ( .A1(n14906), .A2(n14802), .ZN(n14803) );
  OR2_X1 U18109 ( .A1(n14803), .A2(n14893), .ZN(n19131) );
  NOR2_X1 U18110 ( .A1(n19102), .A2(n14804), .ZN(n14805) );
  XNOR2_X1 U18111 ( .A(n14805), .B(n15152), .ZN(n14814) );
  AND2_X1 U18112 ( .A1(n15397), .A2(n14807), .ZN(n14808) );
  NOR2_X1 U18113 ( .A1(n14806), .A2(n14808), .ZN(n19167) );
  INV_X1 U18114 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U18115 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19109), .ZN(n14809) );
  OAI211_X1 U18116 ( .C1(n19096), .C2(n15153), .A(n14809), .B(n11494), .ZN(
        n14810) );
  AOI21_X1 U18117 ( .B1(n19167), .B2(n14829), .A(n14810), .ZN(n14811) );
  OAI21_X1 U18118 ( .B1(n14812), .B2(n19112), .A(n14811), .ZN(n14813) );
  AOI21_X1 U18119 ( .B1(n14814), .B2(n19123), .A(n14813), .ZN(n14815) );
  OAI21_X1 U18120 ( .B1(n19131), .B2(n19090), .A(n14815), .ZN(P2_U2839) );
  NOR2_X1 U18121 ( .A1(n19102), .A2(n14816), .ZN(n14817) );
  XNOR2_X1 U18122 ( .A(n14817), .B(n15202), .ZN(n14833) );
  NAND2_X1 U18123 ( .A1(n14820), .A2(n14819), .ZN(n14821) );
  NAND2_X1 U18124 ( .A1(n14818), .A2(n14821), .ZN(n19141) );
  INV_X1 U18125 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U18126 ( .A1(n14822), .A2(n19086), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19110), .ZN(n14823) );
  OAI211_X1 U18127 ( .C1(n19823), .C2(n19096), .A(n14823), .B(n19088), .ZN(
        n14824) );
  AOI21_X1 U18128 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19109), .A(
        n14824), .ZN(n14831) );
  NOR2_X1 U18129 ( .A1(n14826), .A2(n14827), .ZN(n14828) );
  NOR2_X1 U18130 ( .A1(n14825), .A2(n14828), .ZN(n19181) );
  NAND2_X1 U18131 ( .A1(n14829), .A2(n19181), .ZN(n14830) );
  OAI211_X1 U18132 ( .C1(n19090), .C2(n19141), .A(n14831), .B(n14830), .ZN(
        n14832) );
  AOI21_X1 U18133 ( .B1(n14833), .B2(n19123), .A(n14832), .ZN(n14834) );
  INV_X1 U18134 ( .A(n14834), .ZN(P2_U2843) );
  AOI21_X1 U18135 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n16237) );
  INV_X1 U18136 ( .A(n16237), .ZN(n14843) );
  INV_X1 U18137 ( .A(n14838), .ZN(n14921) );
  NAND2_X1 U18138 ( .A1(n14839), .A2(n14840), .ZN(n14920) );
  NAND3_X1 U18139 ( .A1(n14921), .A2(n19156), .A3(n14920), .ZN(n14842) );
  NAND2_X1 U18140 ( .A1(n19153), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14841) );
  OAI211_X1 U18141 ( .C1(n19153), .C2(n14843), .A(n14842), .B(n14841), .ZN(
        P2_U2858) );
  NOR2_X1 U18142 ( .A1(n14845), .A2(n14844), .ZN(n14847) );
  XNOR2_X1 U18143 ( .A(n14847), .B(n14846), .ZN(n14936) );
  NOR2_X1 U18144 ( .A1(n14848), .A2(n19153), .ZN(n14849) );
  AOI21_X1 U18145 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19153), .A(n14849), .ZN(
        n14850) );
  OAI21_X1 U18146 ( .B1(n14936), .B2(n19148), .A(n14850), .ZN(P2_U2859) );
  NAND2_X1 U18147 ( .A1(n14937), .A2(n19156), .ZN(n14855) );
  NAND2_X1 U18148 ( .A1(n19153), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14854) );
  OAI211_X1 U18149 ( .C1(n14856), .C2(n19153), .A(n14855), .B(n14854), .ZN(
        P2_U2860) );
  AOI21_X1 U18150 ( .B1(n14857), .B2(n14859), .A(n14858), .ZN(n14944) );
  NAND2_X1 U18151 ( .A1(n14944), .A2(n19156), .ZN(n14861) );
  NAND2_X1 U18152 ( .A1(n19153), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14860) );
  OAI211_X1 U18153 ( .C1(n15250), .C2(n19153), .A(n14861), .B(n14860), .ZN(
        P2_U2861) );
  INV_X1 U18154 ( .A(n14864), .ZN(n14865) );
  AOI21_X1 U18155 ( .B1(n14862), .B2(n14866), .A(n14865), .ZN(n14952) );
  NAND2_X1 U18156 ( .A1(n14952), .A2(n19156), .ZN(n14868) );
  NAND2_X1 U18157 ( .A1(n19153), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14867) );
  OAI211_X1 U18158 ( .C1(n15274), .C2(n19153), .A(n14868), .B(n14867), .ZN(
        P2_U2862) );
  AOI21_X1 U18159 ( .B1(n14870), .B2(n14872), .A(n14871), .ZN(n14873) );
  XOR2_X1 U18160 ( .A(n14874), .B(n14873), .Z(n14963) );
  MUX2_X1 U18161 ( .A(n15279), .B(n14747), .S(n19153), .Z(n14875) );
  OAI21_X1 U18162 ( .B1(n14963), .B2(n19148), .A(n14875), .ZN(P2_U2863) );
  OAI21_X1 U18163 ( .B1(n14876), .B2(n14878), .A(n14877), .ZN(n14977) );
  NOR2_X1 U18164 ( .A1(n19159), .A2(n14879), .ZN(n14880) );
  AOI21_X1 U18165 ( .B1(n15324), .B2(n19159), .A(n14880), .ZN(n14881) );
  OAI21_X1 U18166 ( .B1(n14977), .B2(n19148), .A(n14881), .ZN(P2_U2866) );
  INV_X1 U18167 ( .A(n14883), .ZN(n14884) );
  OAI21_X1 U18168 ( .B1(n14882), .B2(n14885), .A(n14884), .ZN(n14985) );
  NAND2_X1 U18169 ( .A1(n14886), .A2(n14887), .ZN(n14888) );
  NAND2_X1 U18170 ( .A1(n15110), .A2(n14888), .ZN(n18983) );
  NOR2_X1 U18171 ( .A1(n18983), .A2(n19153), .ZN(n14889) );
  AOI21_X1 U18172 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19153), .A(n14889), .ZN(
        n14890) );
  OAI21_X1 U18173 ( .B1(n14985), .B2(n19148), .A(n14890), .ZN(P2_U2868) );
  NOR2_X1 U18174 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  OR2_X1 U18175 ( .A1(n14891), .A2(n14894), .ZN(n19009) );
  INV_X1 U18176 ( .A(n14896), .ZN(n14897) );
  AOI21_X1 U18177 ( .B1(n14898), .B2(n14895), .A(n14896), .ZN(n14993) );
  NAND2_X1 U18178 ( .A1(n14993), .A2(n19156), .ZN(n14900) );
  NAND2_X1 U18179 ( .A1(n19153), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14899) );
  OAI211_X1 U18180 ( .C1(n19009), .C2(n19153), .A(n14900), .B(n14899), .ZN(
        P2_U2870) );
  INV_X1 U18181 ( .A(n14901), .ZN(n14902) );
  OAI211_X1 U18182 ( .C1(n9713), .C2(n14903), .A(n14902), .B(n19156), .ZN(
        n14908) );
  NAND2_X1 U18183 ( .A1(n15181), .A2(n14904), .ZN(n14905) );
  NAND2_X1 U18184 ( .A1(n14906), .A2(n14905), .ZN(n15169) );
  INV_X1 U18185 ( .A(n15169), .ZN(n19022) );
  NAND2_X1 U18186 ( .A1(n19022), .A2(n19159), .ZN(n14907) );
  OAI211_X1 U18187 ( .C1(n19159), .C2(n19015), .A(n14908), .B(n14907), .ZN(
        P2_U2872) );
  NOR2_X1 U18188 ( .A1(n19137), .A2(n19138), .ZN(n14912) );
  INV_X1 U18189 ( .A(n14909), .ZN(n14911) );
  OR2_X1 U18190 ( .A1(n19137), .A2(n14910), .ZN(n19132) );
  OAI211_X1 U18191 ( .C1(n14912), .C2(n14911), .A(n19156), .B(n19132), .ZN(
        n14916) );
  AND2_X1 U18192 ( .A1(n14818), .A2(n14913), .ZN(n14914) );
  OR2_X1 U18193 ( .A1(n14914), .A2(n15179), .ZN(n15430) );
  INV_X1 U18194 ( .A(n15430), .ZN(n19045) );
  NAND2_X1 U18195 ( .A1(n19045), .A2(n19159), .ZN(n14915) );
  OAI211_X1 U18196 ( .C1(n19159), .C2(n11215), .A(n14916), .B(n14915), .ZN(
        P2_U2874) );
  OR2_X1 U18197 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  NAND2_X1 U18198 ( .A1(n11607), .A2(n14919), .ZN(n16240) );
  INV_X1 U18199 ( .A(n19218), .ZN(n19168) );
  NAND3_X1 U18200 ( .A1(n14921), .A2(n19168), .A3(n14920), .ZN(n14927) );
  INV_X1 U18201 ( .A(n19164), .ZN(n14973) );
  OAI22_X1 U18202 ( .A1(n14973), .A2(n19179), .B1(n19196), .B2(n14922), .ZN(
        n14925) );
  INV_X1 U18203 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n14923) );
  NOR2_X1 U18204 ( .A1(n14948), .A2(n14923), .ZN(n14924) );
  AOI211_X1 U18205 ( .C1(n19166), .C2(BUF1_REG_29__SCAN_IN), .A(n14925), .B(
        n14924), .ZN(n14926) );
  OAI211_X1 U18206 ( .C1(n19173), .C2(n16240), .A(n14927), .B(n14926), .ZN(
        P2_U2890) );
  INV_X1 U18207 ( .A(n14928), .ZN(n14934) );
  INV_X1 U18208 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n14932) );
  OAI22_X1 U18209 ( .A1(n14973), .A2(n19182), .B1(n19196), .B2(n14929), .ZN(
        n14930) );
  AOI21_X1 U18210 ( .B1(n19166), .B2(BUF1_REG_28__SCAN_IN), .A(n14930), .ZN(
        n14931) );
  OAI21_X1 U18211 ( .B1(n14948), .B2(n14932), .A(n14931), .ZN(n14933) );
  AOI21_X1 U18212 ( .B1(n14934), .B2(n19214), .A(n14933), .ZN(n14935) );
  OAI21_X1 U18213 ( .B1(n14936), .B2(n19218), .A(n14935), .ZN(P2_U2891) );
  NAND2_X1 U18214 ( .A1(n14937), .A2(n19168), .ZN(n14942) );
  OAI22_X1 U18215 ( .A1(n14973), .A2(n19184), .B1(n19196), .B2(n14938), .ZN(
        n14940) );
  INV_X1 U18216 ( .A(n19166), .ZN(n14955) );
  INV_X1 U18217 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16459) );
  NOR2_X1 U18218 ( .A1(n14955), .A2(n16459), .ZN(n14939) );
  AOI211_X1 U18219 ( .C1(BUF2_REG_27__SCAN_IN), .C2(n19165), .A(n14940), .B(
        n14939), .ZN(n14941) );
  OAI211_X1 U18220 ( .C1(n14943), .C2(n19173), .A(n14942), .B(n14941), .ZN(
        P2_U2892) );
  INV_X1 U18221 ( .A(n14944), .ZN(n14951) );
  INV_X1 U18222 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n14947) );
  AOI22_X1 U18223 ( .A1(n19164), .A2(n19186), .B1(n19213), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n14946) );
  NAND2_X1 U18224 ( .A1(n19166), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14945) );
  OAI211_X1 U18225 ( .C1(n14948), .C2(n14947), .A(n14946), .B(n14945), .ZN(
        n14949) );
  AOI21_X1 U18226 ( .B1(n15254), .B2(n19214), .A(n14949), .ZN(n14950) );
  OAI21_X1 U18227 ( .B1(n14951), .B2(n19218), .A(n14950), .ZN(P2_U2893) );
  NAND2_X1 U18228 ( .A1(n14952), .A2(n19168), .ZN(n14958) );
  INV_X1 U18229 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U18230 ( .A1(n19164), .A2(n19189), .B1(n19213), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n14953) );
  OAI21_X1 U18231 ( .B1(n14955), .B2(n14954), .A(n14953), .ZN(n14956) );
  AOI21_X1 U18232 ( .B1(n19165), .B2(BUF2_REG_25__SCAN_IN), .A(n14956), .ZN(
        n14957) );
  OAI211_X1 U18233 ( .C1(n15267), .C2(n19173), .A(n14958), .B(n14957), .ZN(
        P2_U2894) );
  AOI22_X1 U18234 ( .A1(n19164), .A2(n19192), .B1(n19213), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U18235 ( .A1(n19165), .A2(BUF2_REG_24__SCAN_IN), .B1(n19166), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14959) );
  OAI211_X1 U18236 ( .C1(n15285), .C2(n19173), .A(n14960), .B(n14959), .ZN(
        n14961) );
  INV_X1 U18237 ( .A(n14961), .ZN(n14962) );
  OAI21_X1 U18238 ( .B1(n14963), .B2(n19218), .A(n14962), .ZN(P2_U2895) );
  AOI21_X1 U18239 ( .B1(n14964), .B2(n14966), .A(n14965), .ZN(n16243) );
  INV_X1 U18240 ( .A(n16243), .ZN(n14971) );
  OAI22_X1 U18241 ( .A1(n14973), .A2(n19311), .B1(n19196), .B2(n14967), .ZN(
        n14968) );
  AOI21_X1 U18242 ( .B1(n15292), .B2(n19214), .A(n14968), .ZN(n14970) );
  AOI22_X1 U18243 ( .A1(n19165), .A2(BUF2_REG_23__SCAN_IN), .B1(n19166), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14969) );
  OAI211_X1 U18244 ( .C1(n14971), .C2(n19218), .A(n14970), .B(n14969), .ZN(
        P2_U2896) );
  INV_X1 U18245 ( .A(n19199), .ZN(n19300) );
  OAI22_X1 U18246 ( .A1(n14973), .A2(n19300), .B1(n19196), .B2(n14972), .ZN(
        n14974) );
  AOI21_X1 U18247 ( .B1(n15316), .B2(n19214), .A(n14974), .ZN(n14976) );
  AOI22_X1 U18248 ( .A1(n19165), .A2(BUF2_REG_21__SCAN_IN), .B1(n19166), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14975) );
  OAI211_X1 U18249 ( .C1(n14977), .C2(n19218), .A(n14976), .B(n14975), .ZN(
        P2_U2898) );
  NAND2_X1 U18250 ( .A1(n15358), .A2(n14978), .ZN(n14979) );
  NAND2_X1 U18251 ( .A1(n15330), .A2(n14979), .ZN(n18982) );
  AOI22_X1 U18252 ( .A1(n19165), .A2(BUF2_REG_19__SCAN_IN), .B1(n19166), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U18253 ( .A1(n19164), .A2(n14980), .B1(n19213), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14981) );
  OAI211_X1 U18254 ( .C1(n19173), .C2(n18982), .A(n14982), .B(n14981), .ZN(
        n14983) );
  INV_X1 U18255 ( .A(n14983), .ZN(n14984) );
  OAI21_X1 U18256 ( .B1(n14985), .B2(n19218), .A(n14984), .ZN(P2_U2900) );
  NOR2_X1 U18257 ( .A1(n14806), .A2(n14987), .ZN(n14988) );
  OR2_X1 U18258 ( .A1(n14986), .A2(n14988), .ZN(n19008) );
  AOI22_X1 U18259 ( .A1(n19165), .A2(BUF2_REG_17__SCAN_IN), .B1(n19166), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U18260 ( .A1(n19164), .A2(n14989), .B1(n19213), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14990) );
  OAI211_X1 U18261 ( .C1(n19173), .C2(n19008), .A(n14991), .B(n14990), .ZN(
        n14992) );
  AOI21_X1 U18262 ( .B1(n14993), .B2(n19168), .A(n14992), .ZN(n14994) );
  INV_X1 U18263 ( .A(n14994), .ZN(P2_U2902) );
  AOI21_X1 U18264 ( .B1(n14996), .B2(n19877), .A(n14995), .ZN(n19209) );
  XOR2_X1 U18265 ( .A(n19206), .B(n19871), .Z(n19208) );
  NOR2_X1 U18266 ( .A1(n19209), .A2(n19208), .ZN(n19207) );
  AOI21_X1 U18267 ( .B1(n19206), .B2(n14997), .A(n19207), .ZN(n14998) );
  NOR2_X1 U18268 ( .A1(n14998), .A2(n15558), .ZN(n19201) );
  XNOR2_X1 U18269 ( .A(n19201), .B(n19200), .ZN(n15001) );
  AOI22_X1 U18270 ( .A1(n19214), .A2(n15558), .B1(n19213), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n15000) );
  NAND2_X1 U18271 ( .A1(n19198), .A2(n16265), .ZN(n14999) );
  OAI211_X1 U18272 ( .C1(n15001), .C2(n19218), .A(n15000), .B(n14999), .ZN(
        P2_U2915) );
  AOI21_X1 U18273 ( .B1(n16297), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15002), .ZN(n15005) );
  NAND2_X1 U18274 ( .A1(n16305), .A2(n15003), .ZN(n15004) );
  OAI211_X1 U18275 ( .C1(n9575), .C2(n13376), .A(n15005), .B(n15004), .ZN(
        n15007) );
  AOI21_X1 U18276 ( .B1(n15008), .B2(n16293), .A(n15007), .ZN(n15009) );
  OAI21_X1 U18277 ( .B1(n16308), .B2(n15010), .A(n15009), .ZN(P2_U2984) );
  NAND2_X1 U18278 ( .A1(n15012), .A2(n15011), .ZN(n15014) );
  XOR2_X1 U18279 ( .A(n15014), .B(n15013), .Z(n15249) );
  NOR2_X1 U18280 ( .A1(n11494), .A2(n19853), .ZN(n15241) );
  AOI21_X1 U18281 ( .B1(n16297), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15241), .ZN(n15015) );
  OAI21_X1 U18282 ( .B1(n16304), .B2(n15016), .A(n15015), .ZN(n15017) );
  AOI21_X1 U18283 ( .B1(n16237), .B2(n16311), .A(n15017), .ZN(n15022) );
  AOI21_X1 U18284 ( .B1(n15018), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15020) );
  NOR2_X2 U18285 ( .A1(n15020), .A2(n15019), .ZN(n15246) );
  NAND2_X1 U18286 ( .A1(n15246), .A2(n11517), .ZN(n15021) );
  OAI211_X1 U18287 ( .C1(n15249), .C2(n16306), .A(n15022), .B(n15021), .ZN(
        P2_U2985) );
  AOI21_X1 U18288 ( .B1(n15023), .B2(n15034), .A(n15036), .ZN(n15024) );
  XOR2_X1 U18289 ( .A(n15025), .B(n15024), .Z(n15264) );
  NAND2_X1 U18290 ( .A1(n19115), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15256) );
  OAI21_X1 U18291 ( .B1(n16315), .B2(n15026), .A(n15256), .ZN(n15028) );
  NOR2_X1 U18292 ( .A1(n15250), .A2(n13376), .ZN(n15027) );
  AOI211_X1 U18293 ( .C1(n16305), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        n15032) );
  AOI21_X1 U18294 ( .B1(n15251), .B2(n15030), .A(n11521), .ZN(n15261) );
  NAND2_X1 U18295 ( .A1(n15261), .A2(n11517), .ZN(n15031) );
  OAI211_X1 U18296 ( .C1(n15264), .C2(n16306), .A(n15032), .B(n15031), .ZN(
        P2_U2988) );
  OAI21_X1 U18297 ( .B1(n15033), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15030), .ZN(n15278) );
  INV_X1 U18298 ( .A(n15034), .ZN(n15035) );
  NOR2_X1 U18299 ( .A1(n15036), .A2(n15035), .ZN(n15037) );
  XNOR2_X1 U18300 ( .A(n15023), .B(n15037), .ZN(n15276) );
  NAND2_X1 U18301 ( .A1(n19115), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15266) );
  OAI21_X1 U18302 ( .B1(n16315), .B2(n15038), .A(n15266), .ZN(n15039) );
  AOI21_X1 U18303 ( .B1(n16305), .B2(n15040), .A(n15039), .ZN(n15041) );
  OAI21_X1 U18304 ( .B1(n15274), .B2(n13376), .A(n15041), .ZN(n15042) );
  AOI21_X1 U18305 ( .B1(n15276), .B2(n16293), .A(n15042), .ZN(n15043) );
  OAI21_X1 U18306 ( .B1(n16308), .B2(n15278), .A(n15043), .ZN(P2_U2989) );
  INV_X1 U18307 ( .A(n15056), .ZN(n15046) );
  INV_X1 U18308 ( .A(n15033), .ZN(n15045) );
  OAI21_X1 U18309 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15046), .A(
        n15045), .ZN(n15290) );
  XOR2_X1 U18310 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15047), .Z(
        n15048) );
  XNOR2_X1 U18311 ( .A(n15049), .B(n15048), .ZN(n15288) );
  NOR2_X1 U18312 ( .A1(n15279), .A2(n13376), .ZN(n15053) );
  NAND2_X1 U18313 ( .A1(n19115), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15283) );
  NAND2_X1 U18314 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15050) );
  OAI211_X1 U18315 ( .C1(n16304), .C2(n15051), .A(n15283), .B(n15050), .ZN(
        n15052) );
  AOI211_X1 U18316 ( .C1(n15288), .C2(n16293), .A(n15053), .B(n15052), .ZN(
        n15054) );
  OAI21_X1 U18317 ( .B1(n16308), .B2(n15290), .A(n15054), .ZN(P2_U2990) );
  INV_X1 U18318 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15308) );
  NOR2_X1 U18319 ( .A1(n15055), .A2(n15308), .ZN(n15070) );
  OAI21_X1 U18320 ( .B1(n15070), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15056), .ZN(n15301) );
  XOR2_X1 U18321 ( .A(n15058), .B(n15057), .Z(n15299) );
  INV_X1 U18322 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19841) );
  NOR2_X1 U18323 ( .A1(n11494), .A2(n19841), .ZN(n15291) );
  NOR2_X1 U18324 ( .A1(n16315), .A2(n15059), .ZN(n15060) );
  AOI211_X1 U18325 ( .C1(n15061), .C2(n16305), .A(n15291), .B(n15060), .ZN(
        n15062) );
  OAI21_X1 U18326 ( .B1(n16241), .B2(n13376), .A(n15062), .ZN(n15063) );
  AOI21_X1 U18327 ( .B1(n15299), .B2(n16293), .A(n15063), .ZN(n15064) );
  OAI21_X1 U18328 ( .B1(n16308), .B2(n15301), .A(n15064), .ZN(P2_U2991) );
  INV_X1 U18329 ( .A(n15066), .ZN(n15068) );
  NAND2_X1 U18330 ( .A1(n15068), .A2(n15067), .ZN(n15069) );
  XNOR2_X1 U18331 ( .A(n15065), .B(n15069), .ZN(n15313) );
  AOI21_X1 U18332 ( .B1(n15308), .B2(n15055), .A(n15070), .ZN(n15302) );
  NAND2_X1 U18333 ( .A1(n15302), .A2(n11517), .ZN(n15075) );
  INV_X1 U18334 ( .A(n16248), .ZN(n15310) );
  NAND2_X1 U18335 ( .A1(n19115), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15303) );
  NAND2_X1 U18336 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15071) );
  OAI211_X1 U18337 ( .C1(n16304), .C2(n15072), .A(n15303), .B(n15071), .ZN(
        n15073) );
  AOI21_X1 U18338 ( .B1(n15310), .B2(n16311), .A(n15073), .ZN(n15074) );
  OAI211_X1 U18339 ( .C1(n15313), .C2(n16306), .A(n15075), .B(n15074), .ZN(
        P2_U2992) );
  XNOR2_X1 U18340 ( .A(n15078), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15200) );
  INV_X1 U18341 ( .A(n15079), .ZN(n15080) );
  INV_X1 U18342 ( .A(n15189), .ZN(n15081) );
  INV_X1 U18343 ( .A(n15172), .ZN(n15082) );
  INV_X1 U18344 ( .A(n15083), .ZN(n15147) );
  INV_X1 U18345 ( .A(n15086), .ZN(n15087) );
  NAND2_X1 U18346 ( .A1(n15129), .A2(n15127), .ZN(n15115) );
  INV_X1 U18347 ( .A(n15116), .ZN(n15090) );
  INV_X1 U18348 ( .A(n15088), .ZN(n15089) );
  OAI21_X1 U18349 ( .B1(n15115), .B2(n15090), .A(n15089), .ZN(n15106) );
  INV_X1 U18350 ( .A(n15093), .ZN(n15092) );
  NAND2_X1 U18351 ( .A1(n15092), .A2(n15091), .ZN(n15105) );
  NOR2_X1 U18352 ( .A1(n15107), .A2(n15093), .ZN(n15096) );
  NAND2_X1 U18353 ( .A1(n9655), .A2(n15094), .ZN(n15095) );
  XNOR2_X1 U18354 ( .A(n15096), .B(n15095), .ZN(n15326) );
  NAND2_X1 U18355 ( .A1(n16305), .A2(n15097), .ZN(n15098) );
  NAND2_X1 U18356 ( .A1(n19115), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15314) );
  OAI211_X1 U18357 ( .C1(n16315), .C2(n15099), .A(n15098), .B(n15314), .ZN(
        n15101) );
  OAI21_X1 U18358 ( .B1(n9674), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15055), .ZN(n15321) );
  NOR2_X1 U18359 ( .A1(n15321), .A2(n16308), .ZN(n15100) );
  AOI211_X1 U18360 ( .C1(n16311), .C2(n15324), .A(n15101), .B(n15100), .ZN(
        n15102) );
  OAI21_X1 U18361 ( .B1(n15326), .B2(n16306), .A(n15102), .ZN(P2_U2993) );
  INV_X1 U18362 ( .A(n9674), .ZN(n15104) );
  OAI21_X1 U18363 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15103), .A(
        n15104), .ZN(n15343) );
  AND2_X1 U18364 ( .A1(n15106), .A2(n15105), .ZN(n15108) );
  NOR2_X1 U18365 ( .A1(n15108), .A2(n15107), .ZN(n15327) );
  NAND2_X1 U18366 ( .A1(n15327), .A2(n16293), .ZN(n15114) );
  XNOR2_X1 U18367 ( .A(n15110), .B(n9942), .ZN(n18972) );
  INV_X1 U18368 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19835) );
  NOR2_X1 U18369 ( .A1(n11494), .A2(n19835), .ZN(n15336) );
  AOI21_X1 U18370 ( .B1(n16297), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15336), .ZN(n15111) );
  OAI21_X1 U18371 ( .B1(n16304), .B2(n18962), .A(n15111), .ZN(n15112) );
  AOI21_X1 U18372 ( .B1(n18972), .B2(n16311), .A(n15112), .ZN(n15113) );
  OAI211_X1 U18373 ( .C1(n16308), .C2(n15343), .A(n15114), .B(n15113), .ZN(
        P2_U2994) );
  NAND2_X1 U18374 ( .A1(n15115), .A2(n15126), .ZN(n15119) );
  NAND2_X1 U18375 ( .A1(n15117), .A2(n15116), .ZN(n15118) );
  XNOR2_X1 U18376 ( .A(n15119), .B(n15118), .ZN(n15354) );
  INV_X1 U18377 ( .A(n15120), .ZN(n15121) );
  AOI21_X1 U18378 ( .B1(n15348), .B2(n15121), .A(n15103), .ZN(n15352) );
  INV_X1 U18379 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19833) );
  NOR2_X1 U18380 ( .A1(n19088), .A2(n19833), .ZN(n15344) );
  NOR2_X1 U18381 ( .A1(n16315), .A2(n18978), .ZN(n15122) );
  AOI211_X1 U18382 ( .C1(n18977), .C2(n16305), .A(n15344), .B(n15122), .ZN(
        n15123) );
  OAI21_X1 U18383 ( .B1(n18983), .B2(n13376), .A(n15123), .ZN(n15124) );
  AOI21_X1 U18384 ( .B1(n15352), .B2(n11517), .A(n15124), .ZN(n15125) );
  OAI21_X1 U18385 ( .B1(n15354), .B2(n16306), .A(n15125), .ZN(P2_U2995) );
  NAND2_X1 U18386 ( .A1(n15127), .A2(n15126), .ZN(n15128) );
  XNOR2_X1 U18387 ( .A(n15129), .B(n15128), .ZN(n15371) );
  INV_X1 U18388 ( .A(n15130), .ZN(n15131) );
  AOI21_X1 U18389 ( .B1(n15131), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U18390 ( .A1(n15132), .A2(n15120), .ZN(n15369) );
  OR2_X1 U18391 ( .A1(n14891), .A2(n15133), .ZN(n15134) );
  NAND2_X1 U18392 ( .A1(n14886), .A2(n15134), .ZN(n18995) );
  INV_X1 U18393 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U18394 ( .A1(n11494), .A2(n15135), .ZN(n15359) );
  NOR2_X1 U18395 ( .A1(n18989), .A2(n16304), .ZN(n15136) );
  AOI211_X1 U18396 ( .C1(n16297), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15359), .B(n15136), .ZN(n15137) );
  OAI21_X1 U18397 ( .B1(n18995), .B2(n13376), .A(n15137), .ZN(n15138) );
  AOI21_X1 U18398 ( .B1(n15369), .B2(n11517), .A(n15138), .ZN(n15139) );
  OAI21_X1 U18399 ( .B1(n15371), .B2(n16306), .A(n15139), .ZN(P2_U2996) );
  XNOR2_X1 U18400 ( .A(n15141), .B(n15140), .ZN(n15386) );
  XNOR2_X1 U18401 ( .A(n15130), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15145) );
  NOR2_X1 U18402 ( .A1(n19009), .A2(n13376), .ZN(n15144) );
  OR2_X1 U18403 ( .A1(n19088), .A2(n19830), .ZN(n15373) );
  NAND2_X1 U18404 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15142) );
  OAI211_X1 U18405 ( .C1(n16304), .C2(n19014), .A(n15373), .B(n15142), .ZN(
        n15143) );
  AOI211_X1 U18406 ( .C1(n15145), .C2(n11517), .A(n15144), .B(n15143), .ZN(
        n15146) );
  OAI21_X1 U18407 ( .B1(n15386), .B2(n16306), .A(n15146), .ZN(P2_U2997) );
  XNOR2_X1 U18408 ( .A(n15148), .B(n15147), .ZN(n15396) );
  INV_X1 U18409 ( .A(n15149), .ZN(n15150) );
  OAI21_X1 U18410 ( .B1(n15150), .B2(n15403), .A(n15388), .ZN(n15151) );
  NAND3_X1 U18411 ( .A1(n15130), .A2(n15151), .A3(n11517), .ZN(n15159) );
  INV_X1 U18412 ( .A(n15152), .ZN(n15157) );
  NOR2_X1 U18413 ( .A1(n11494), .A2(n15153), .ZN(n15390) );
  INV_X1 U18414 ( .A(n15390), .ZN(n15154) );
  OAI21_X1 U18415 ( .B1(n16315), .B2(n15155), .A(n15154), .ZN(n15156) );
  AOI21_X1 U18416 ( .B1(n16305), .B2(n15157), .A(n15156), .ZN(n15158) );
  OAI211_X1 U18417 ( .C1(n13376), .C2(n19131), .A(n15159), .B(n15158), .ZN(
        n15160) );
  INV_X1 U18418 ( .A(n15160), .ZN(n15161) );
  OAI21_X1 U18419 ( .B1(n15396), .B2(n16306), .A(n15161), .ZN(P2_U2998) );
  NAND2_X1 U18420 ( .A1(n15163), .A2(n15162), .ZN(n15165) );
  XOR2_X1 U18421 ( .A(n15165), .B(n15164), .Z(n15410) );
  XNOR2_X1 U18422 ( .A(n15150), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15407) );
  NOR2_X1 U18423 ( .A1(n19088), .A2(n19827), .ZN(n15399) );
  NOR2_X1 U18424 ( .A1(n16315), .A2(n15166), .ZN(n15167) );
  AOI211_X1 U18425 ( .C1(n19020), .C2(n16305), .A(n15399), .B(n15167), .ZN(
        n15168) );
  OAI21_X1 U18426 ( .B1(n15169), .B2(n13376), .A(n15168), .ZN(n15170) );
  AOI21_X1 U18427 ( .B1(n15407), .B2(n11517), .A(n15170), .ZN(n15171) );
  OAI21_X1 U18428 ( .B1(n15410), .B2(n16306), .A(n15171), .ZN(P2_U2999) );
  NAND2_X1 U18429 ( .A1(n15173), .A2(n15172), .ZN(n15174) );
  XNOR2_X1 U18430 ( .A(n15175), .B(n15174), .ZN(n15428) );
  INV_X1 U18431 ( .A(n15176), .ZN(n15177) );
  INV_X1 U18432 ( .A(n15436), .ZN(n15415) );
  NAND2_X1 U18433 ( .A1(n15177), .A2(n15415), .ZN(n15188) );
  AOI21_X1 U18434 ( .B1(n15414), .B2(n15188), .A(n15149), .ZN(n15426) );
  OR2_X1 U18435 ( .A1(n15179), .A2(n15178), .ZN(n15180) );
  NAND2_X1 U18436 ( .A1(n15181), .A2(n15180), .ZN(n19136) );
  INV_X1 U18437 ( .A(n19027), .ZN(n15184) );
  INV_X1 U18438 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n15182) );
  OR2_X1 U18439 ( .A1(n19088), .A2(n15182), .ZN(n15422) );
  OAI21_X1 U18440 ( .B1(n16315), .B2(n9852), .A(n15422), .ZN(n15183) );
  AOI21_X1 U18441 ( .B1(n16305), .B2(n15184), .A(n15183), .ZN(n15185) );
  OAI21_X1 U18442 ( .B1(n19136), .B2(n13376), .A(n15185), .ZN(n15186) );
  AOI21_X1 U18443 ( .B1(n15426), .B2(n11517), .A(n15186), .ZN(n15187) );
  OAI21_X1 U18444 ( .B1(n15428), .B2(n16306), .A(n15187), .ZN(P2_U3000) );
  NOR2_X1 U18445 ( .A1(n15176), .A2(n15447), .ZN(n15204) );
  OAI21_X1 U18446 ( .B1(n15204), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15188), .ZN(n15444) );
  NAND2_X1 U18447 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  XNOR2_X1 U18448 ( .A(n15192), .B(n15191), .ZN(n15429) );
  INV_X1 U18449 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15193) );
  OR2_X1 U18450 ( .A1(n19088), .A2(n15193), .ZN(n15437) );
  OAI21_X1 U18451 ( .B1(n16315), .B2(n15194), .A(n15437), .ZN(n15195) );
  AOI21_X1 U18452 ( .B1(n16305), .B2(n19043), .A(n15195), .ZN(n15196) );
  OAI21_X1 U18453 ( .B1(n15430), .B2(n13376), .A(n15196), .ZN(n15197) );
  AOI21_X1 U18454 ( .B1(n15429), .B2(n16293), .A(n15197), .ZN(n15198) );
  OAI21_X1 U18455 ( .B1(n16308), .B2(n15444), .A(n15198), .ZN(P2_U3001) );
  XOR2_X1 U18456 ( .A(n15200), .B(n15199), .Z(n15458) );
  INV_X1 U18457 ( .A(n19141), .ZN(n15453) );
  NOR2_X1 U18458 ( .A1(n11494), .A2(n19823), .ZN(n15449) );
  AOI21_X1 U18459 ( .B1(n16297), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15449), .ZN(n15201) );
  OAI21_X1 U18460 ( .B1(n16304), .B2(n15202), .A(n15201), .ZN(n15203) );
  AOI21_X1 U18461 ( .B1(n15453), .B2(n16311), .A(n15203), .ZN(n15206) );
  INV_X1 U18462 ( .A(n15204), .ZN(n15455) );
  NAND2_X1 U18463 ( .A1(n15176), .A2(n15447), .ZN(n15454) );
  NAND3_X1 U18464 ( .A1(n15455), .A2(n11517), .A3(n15454), .ZN(n15205) );
  OAI211_X1 U18465 ( .C1(n15458), .C2(n16306), .A(n15206), .B(n15205), .ZN(
        P2_U3002) );
  OAI21_X1 U18466 ( .B1(n9677), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15176), .ZN(n15477) );
  XNOR2_X1 U18467 ( .A(n15207), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15208) );
  XNOR2_X1 U18468 ( .A(n15209), .B(n15208), .ZN(n15475) );
  AOI22_X1 U18469 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16305), .B2(n19050), .ZN(n15210) );
  NAND2_X1 U18470 ( .A1(n19115), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n15466) );
  OAI211_X1 U18471 ( .C1(n19055), .C2(n13376), .A(n15210), .B(n15466), .ZN(
        n15211) );
  AOI21_X1 U18472 ( .B1(n15475), .B2(n16293), .A(n15211), .ZN(n15212) );
  OAI21_X1 U18473 ( .B1(n16308), .B2(n15477), .A(n15212), .ZN(P2_U3003) );
  NOR2_X1 U18474 ( .A1(n15213), .A2(n15214), .ZN(n16283) );
  INV_X1 U18475 ( .A(n16283), .ZN(n15216) );
  OAI21_X1 U18476 ( .B1(n16282), .B2(n15214), .A(n15213), .ZN(n15215) );
  OAI21_X1 U18477 ( .B1(n15216), .B2(n16282), .A(n15215), .ZN(n15514) );
  INV_X1 U18478 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19814) );
  OAI22_X1 U18479 ( .A1(n16315), .A2(n19083), .B1(n19814), .B2(n19088), .ZN(
        n15218) );
  NOR2_X1 U18480 ( .A1(n19091), .A2(n13376), .ZN(n15217) );
  AOI211_X1 U18481 ( .C1(n16305), .C2(n19081), .A(n15218), .B(n15217), .ZN(
        n15225) );
  AND2_X1 U18482 ( .A1(n15220), .A2(n15219), .ZN(n15221) );
  XNOR2_X1 U18483 ( .A(n15222), .B(n16325), .ZN(n15223) );
  XNOR2_X1 U18484 ( .A(n15221), .B(n15223), .ZN(n15511) );
  NAND2_X1 U18485 ( .A1(n15511), .A2(n11517), .ZN(n15224) );
  OAI211_X1 U18486 ( .C1(n15514), .C2(n16306), .A(n15225), .B(n15224), .ZN(
        P2_U3007) );
  XNOR2_X1 U18487 ( .A(n15227), .B(n15226), .ZN(n15564) );
  OAI21_X1 U18488 ( .B1(n15228), .B2(n15555), .A(n15539), .ZN(n15562) );
  INV_X1 U18489 ( .A(n19155), .ZN(n15233) );
  OAI22_X1 U18490 ( .A1(n19808), .A2(n19088), .B1(n16304), .B2(n15230), .ZN(
        n15231) );
  AOI21_X1 U18491 ( .B1(n16297), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n15231), .ZN(n15232) );
  OAI21_X1 U18492 ( .B1(n13376), .B2(n15233), .A(n15232), .ZN(n15234) );
  AOI21_X1 U18493 ( .B1(n15562), .B2(n11517), .A(n15234), .ZN(n15235) );
  OAI21_X1 U18494 ( .B1(n15564), .B2(n16306), .A(n15235), .ZN(P2_U3010) );
  INV_X1 U18495 ( .A(n15236), .ZN(n15238) );
  AOI21_X1 U18496 ( .B1(n15238), .B2(n15237), .A(n15239), .ZN(n15245) );
  NAND3_X1 U18497 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n15240), .A3(
        n15239), .ZN(n15243) );
  INV_X1 U18498 ( .A(n15241), .ZN(n15242) );
  OAI211_X1 U18499 ( .C1(n16240), .C2(n16331), .A(n15243), .B(n15242), .ZN(
        n15244) );
  AOI211_X1 U18500 ( .C1(n16237), .C2(n16333), .A(n15245), .B(n15244), .ZN(
        n15248) );
  NAND2_X1 U18501 ( .A1(n15246), .A2(n16319), .ZN(n15247) );
  OAI211_X1 U18502 ( .C1(n15249), .C2(n19259), .A(n15248), .B(n15247), .ZN(
        P2_U3017) );
  INV_X1 U18503 ( .A(n15250), .ZN(n15260) );
  INV_X1 U18504 ( .A(n15281), .ZN(n15252) );
  NOR3_X1 U18505 ( .A1(n15253), .A2(n15252), .A3(n15251), .ZN(n15259) );
  XNOR2_X1 U18506 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15257) );
  NAND2_X1 U18507 ( .A1(n15254), .A2(n19261), .ZN(n15255) );
  OAI211_X1 U18508 ( .C1(n15265), .C2(n15257), .A(n15256), .B(n15255), .ZN(
        n15258) );
  AOI211_X1 U18509 ( .C1(n15260), .C2(n16333), .A(n15259), .B(n15258), .ZN(
        n15263) );
  NAND2_X1 U18510 ( .A1(n15261), .A2(n16319), .ZN(n15262) );
  OAI211_X1 U18511 ( .C1(n15264), .C2(n19259), .A(n15263), .B(n15262), .ZN(
        P2_U3020) );
  INV_X1 U18512 ( .A(n15265), .ZN(n15270) );
  OAI21_X1 U18513 ( .B1(n15267), .B2(n16331), .A(n15266), .ZN(n15268) );
  AOI21_X1 U18514 ( .B1(n15270), .B2(n15269), .A(n15268), .ZN(n15273) );
  NAND3_X1 U18515 ( .A1(n15271), .A2(n15281), .A3(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15272) );
  OAI211_X1 U18516 ( .C1(n15274), .C2(n19257), .A(n15273), .B(n15272), .ZN(
        n15275) );
  AOI21_X1 U18517 ( .B1(n15276), .B2(n16338), .A(n15275), .ZN(n15277) );
  OAI21_X1 U18518 ( .B1(n19264), .B2(n15278), .A(n15277), .ZN(P2_U3021) );
  NOR2_X1 U18519 ( .A1(n15279), .A2(n19257), .ZN(n15287) );
  INV_X1 U18520 ( .A(n15306), .ZN(n15280) );
  NOR2_X1 U18521 ( .A1(n15280), .A2(n15293), .ZN(n15282) );
  OAI21_X1 U18522 ( .B1(n15282), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15281), .ZN(n15284) );
  OAI211_X1 U18523 ( .C1(n16331), .C2(n15285), .A(n15284), .B(n15283), .ZN(
        n15286) );
  AOI211_X1 U18524 ( .C1(n15288), .C2(n16338), .A(n15287), .B(n15286), .ZN(
        n15289) );
  OAI21_X1 U18525 ( .B1(n19264), .B2(n15290), .A(n15289), .ZN(P2_U3022) );
  NOR2_X1 U18526 ( .A1(n16241), .A2(n19257), .ZN(n15298) );
  AOI21_X1 U18527 ( .B1(n15292), .B2(n19261), .A(n15291), .ZN(n15295) );
  OAI211_X1 U18528 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15306), .B(n15293), .ZN(
        n15294) );
  OAI211_X1 U18529 ( .C1(n15320), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        n15297) );
  AOI211_X1 U18530 ( .C1(n15299), .C2(n16338), .A(n15298), .B(n15297), .ZN(
        n15300) );
  OAI21_X1 U18531 ( .B1(n19264), .B2(n15301), .A(n15300), .ZN(P2_U3023) );
  NAND2_X1 U18532 ( .A1(n15302), .A2(n16319), .ZN(n15312) );
  OAI21_X1 U18533 ( .B1(n15304), .B2(n16331), .A(n15303), .ZN(n15305) );
  AOI21_X1 U18534 ( .B1(n15306), .B2(n15308), .A(n15305), .ZN(n15307) );
  OAI21_X1 U18535 ( .B1(n15320), .B2(n15308), .A(n15307), .ZN(n15309) );
  AOI21_X1 U18536 ( .B1(n15310), .B2(n16333), .A(n15309), .ZN(n15311) );
  OAI211_X1 U18537 ( .C1(n15313), .C2(n19259), .A(n15312), .B(n15311), .ZN(
        P2_U3024) );
  INV_X1 U18538 ( .A(n15314), .ZN(n15315) );
  AOI21_X1 U18539 ( .B1(n15316), .B2(n19261), .A(n15315), .ZN(n15318) );
  INV_X1 U18540 ( .A(n15333), .ZN(n15346) );
  NAND3_X1 U18541 ( .A1(n15346), .A2(n15334), .A3(n15319), .ZN(n15317) );
  OAI211_X1 U18542 ( .C1(n15320), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        n15323) );
  NOR2_X1 U18543 ( .A1(n15321), .A2(n19264), .ZN(n15322) );
  OAI21_X1 U18544 ( .B1(n15326), .B2(n19259), .A(n15325), .ZN(P2_U3025) );
  NAND2_X1 U18545 ( .A1(n15327), .A2(n16338), .ZN(n15342) );
  NAND2_X1 U18546 ( .A1(n15411), .A2(n15328), .ZN(n15349) );
  NAND2_X1 U18547 ( .A1(n15330), .A2(n15329), .ZN(n15331) );
  NAND2_X1 U18548 ( .A1(n15332), .A2(n15331), .ZN(n18970) );
  INV_X1 U18549 ( .A(n18970), .ZN(n15337) );
  AOI211_X1 U18550 ( .C1(n15339), .C2(n15348), .A(n15334), .B(n15333), .ZN(
        n15335) );
  AOI211_X1 U18551 ( .C1(n19261), .C2(n15337), .A(n15336), .B(n15335), .ZN(
        n15338) );
  OAI21_X1 U18552 ( .B1(n15349), .B2(n15339), .A(n15338), .ZN(n15340) );
  AOI21_X1 U18553 ( .B1(n16333), .B2(n18972), .A(n15340), .ZN(n15341) );
  OAI211_X1 U18554 ( .C1(n15343), .C2(n19264), .A(n15342), .B(n15341), .ZN(
        P2_U3026) );
  NOR2_X1 U18555 ( .A1(n18983), .A2(n19257), .ZN(n15351) );
  NOR2_X1 U18556 ( .A1(n18982), .A2(n16331), .ZN(n15345) );
  AOI211_X1 U18557 ( .C1(n15346), .C2(n15348), .A(n15345), .B(n15344), .ZN(
        n15347) );
  OAI21_X1 U18558 ( .B1(n15349), .B2(n15348), .A(n15347), .ZN(n15350) );
  AOI211_X1 U18559 ( .C1(n15352), .C2(n16319), .A(n15351), .B(n15350), .ZN(
        n15353) );
  OAI21_X1 U18560 ( .B1(n15354), .B2(n19259), .A(n15353), .ZN(P2_U3027) );
  NAND2_X1 U18561 ( .A1(n15355), .A2(n15364), .ZN(n15361) );
  OR2_X1 U18562 ( .A1(n14986), .A2(n15356), .ZN(n15357) );
  AND2_X1 U18563 ( .A1(n15358), .A2(n15357), .ZN(n16272) );
  AOI21_X1 U18564 ( .B1(n19261), .B2(n16272), .A(n15359), .ZN(n15360) );
  OAI21_X1 U18565 ( .B1(n15402), .B2(n15361), .A(n15360), .ZN(n15362) );
  INV_X1 U18566 ( .A(n15362), .ZN(n15367) );
  INV_X1 U18567 ( .A(n15411), .ZN(n15521) );
  OR2_X1 U18568 ( .A1(n15363), .A2(n15521), .ZN(n15404) );
  OAI21_X1 U18569 ( .B1(n15382), .B2(n15364), .A(n15404), .ZN(n15365) );
  NAND2_X1 U18570 ( .A1(n15365), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15366) );
  OAI211_X1 U18571 ( .C1(n18995), .C2(n19257), .A(n15367), .B(n15366), .ZN(
        n15368) );
  AOI21_X1 U18572 ( .B1(n15369), .B2(n16319), .A(n15368), .ZN(n15370) );
  OAI21_X1 U18573 ( .B1(n15371), .B2(n19259), .A(n15370), .ZN(P2_U3028) );
  OAI22_X1 U18574 ( .A1(n15130), .A2(n19264), .B1(n15372), .B2(n15402), .ZN(
        n15377) );
  NOR2_X1 U18575 ( .A1(n19009), .A2(n19257), .ZN(n15375) );
  OAI21_X1 U18576 ( .B1(n16331), .B2(n19008), .A(n15373), .ZN(n15374) );
  AOI211_X1 U18577 ( .C1(n15377), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15385) );
  NAND2_X1 U18578 ( .A1(n15378), .A2(n19264), .ZN(n15381) );
  OAI21_X1 U18579 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15379), .A(
        n15404), .ZN(n15380) );
  AOI21_X1 U18580 ( .B1(n15130), .B2(n15381), .A(n15380), .ZN(n15387) );
  OAI21_X1 U18581 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15382), .A(
        n15387), .ZN(n15383) );
  NAND2_X1 U18582 ( .A1(n15383), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15384) );
  OAI211_X1 U18583 ( .C1(n15386), .C2(n19259), .A(n15385), .B(n15384), .ZN(
        P2_U3029) );
  INV_X1 U18584 ( .A(n15387), .ZN(n15394) );
  OAI21_X1 U18585 ( .B1(n15150), .B2(n19264), .A(n15402), .ZN(n15389) );
  NAND3_X1 U18586 ( .A1(n15389), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15388), .ZN(n15392) );
  AOI21_X1 U18587 ( .B1(n19261), .B2(n19167), .A(n15390), .ZN(n15391) );
  OAI211_X1 U18588 ( .C1(n19131), .C2(n19257), .A(n15392), .B(n15391), .ZN(
        n15393) );
  AOI21_X1 U18589 ( .B1(n15394), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15393), .ZN(n15395) );
  OAI21_X1 U18590 ( .B1(n15396), .B2(n19259), .A(n15395), .ZN(P2_U3030) );
  OAI21_X1 U18591 ( .B1(n15419), .B2(n15398), .A(n15397), .ZN(n19175) );
  INV_X1 U18592 ( .A(n19175), .ZN(n15400) );
  AOI21_X1 U18593 ( .B1(n19261), .B2(n15400), .A(n15399), .ZN(n15401) );
  OAI21_X1 U18594 ( .B1(n15402), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15401), .ZN(n15406) );
  NOR2_X1 U18595 ( .A1(n15404), .A2(n15403), .ZN(n15405) );
  AOI211_X1 U18596 ( .C1(n19022), .C2(n16333), .A(n15406), .B(n15405), .ZN(
        n15409) );
  NAND2_X1 U18597 ( .A1(n15407), .A2(n16319), .ZN(n15408) );
  OAI211_X1 U18598 ( .C1(n15410), .C2(n19259), .A(n15409), .B(n15408), .ZN(
        P2_U3031) );
  NOR2_X1 U18599 ( .A1(n19136), .A2(n19257), .ZN(n15425) );
  NAND2_X1 U18600 ( .A1(n15412), .A2(n15411), .ZN(n15446) );
  NAND2_X1 U18601 ( .A1(n15445), .A2(n15436), .ZN(n15413) );
  NAND2_X1 U18602 ( .A1(n15446), .A2(n15413), .ZN(n15441) );
  NAND2_X1 U18603 ( .A1(n15441), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15423) );
  NAND3_X1 U18604 ( .A1(n15445), .A2(n15415), .A3(n15414), .ZN(n15421) );
  NOR2_X1 U18605 ( .A1(n15416), .A2(n15417), .ZN(n15418) );
  NOR2_X1 U18606 ( .A1(n15419), .A2(n15418), .ZN(n19033) );
  NAND2_X1 U18607 ( .A1(n19261), .A2(n19033), .ZN(n15420) );
  NAND4_X1 U18608 ( .A1(n15423), .A2(n15422), .A3(n15421), .A4(n15420), .ZN(
        n15424) );
  AOI211_X1 U18609 ( .C1(n15426), .C2(n16319), .A(n15425), .B(n15424), .ZN(
        n15427) );
  OAI21_X1 U18610 ( .B1(n15428), .B2(n19259), .A(n15427), .ZN(P2_U3032) );
  NAND2_X1 U18611 ( .A1(n15429), .A2(n16338), .ZN(n15443) );
  NOR2_X1 U18612 ( .A1(n15430), .A2(n19257), .ZN(n15440) );
  INV_X1 U18613 ( .A(n15416), .ZN(n15435) );
  INV_X1 U18614 ( .A(n14825), .ZN(n15433) );
  INV_X1 U18615 ( .A(n15431), .ZN(n15432) );
  NAND2_X1 U18616 ( .A1(n15433), .A2(n15432), .ZN(n15434) );
  NAND2_X1 U18617 ( .A1(n15435), .A2(n15434), .ZN(n19180) );
  NAND3_X1 U18618 ( .A1(n15445), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n15436), .ZN(n15438) );
  OAI211_X1 U18619 ( .C1(n16331), .C2(n19180), .A(n15438), .B(n15437), .ZN(
        n15439) );
  AOI211_X1 U18620 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15441), .A(
        n15440), .B(n15439), .ZN(n15442) );
  OAI211_X1 U18621 ( .C1(n15444), .C2(n19264), .A(n15443), .B(n15442), .ZN(
        P2_U3033) );
  INV_X1 U18622 ( .A(n15445), .ZN(n15451) );
  NOR2_X1 U18623 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  AOI211_X1 U18624 ( .C1(n19261), .C2(n19181), .A(n15449), .B(n15448), .ZN(
        n15450) );
  OAI21_X1 U18625 ( .B1(n15451), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15450), .ZN(n15452) );
  AOI21_X1 U18626 ( .B1(n16333), .B2(n15453), .A(n15452), .ZN(n15457) );
  NAND3_X1 U18627 ( .A1(n15455), .A2(n16319), .A3(n15454), .ZN(n15456) );
  OAI211_X1 U18628 ( .C1(n15458), .C2(n19259), .A(n15457), .B(n15456), .ZN(
        P2_U3034) );
  NOR2_X1 U18629 ( .A1(n15521), .A2(n15459), .ZN(n15488) );
  NAND2_X1 U18630 ( .A1(n15488), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15473) );
  INV_X1 U18631 ( .A(n14826), .ZN(n15465) );
  INV_X1 U18632 ( .A(n15460), .ZN(n15463) );
  INV_X1 U18633 ( .A(n15461), .ZN(n15462) );
  NAND2_X1 U18634 ( .A1(n15463), .A2(n15462), .ZN(n15464) );
  NAND2_X1 U18635 ( .A1(n15465), .A2(n15464), .ZN(n19185) );
  INV_X1 U18636 ( .A(n19185), .ZN(n15471) );
  INV_X1 U18637 ( .A(n15466), .ZN(n15470) );
  OAI21_X1 U18638 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15467), .ZN(n15468) );
  NOR2_X1 U18639 ( .A1(n15468), .A2(n15491), .ZN(n15469) );
  AOI211_X1 U18640 ( .C1(n19261), .C2(n15471), .A(n15470), .B(n15469), .ZN(
        n15472) );
  OAI211_X1 U18641 ( .C1(n19055), .C2(n19257), .A(n15473), .B(n15472), .ZN(
        n15474) );
  AOI21_X1 U18642 ( .B1(n15475), .B2(n16338), .A(n15474), .ZN(n15476) );
  OAI21_X1 U18643 ( .B1(n19264), .B2(n15477), .A(n15476), .ZN(P2_U3035) );
  AOI21_X1 U18644 ( .B1(n15478), .B2(n13787), .A(n9677), .ZN(n16278) );
  INV_X1 U18645 ( .A(n16278), .ZN(n15499) );
  NAND2_X1 U18646 ( .A1(n13789), .A2(n15479), .ZN(n15484) );
  INV_X1 U18647 ( .A(n15480), .ZN(n15482) );
  NAND2_X1 U18648 ( .A1(n15482), .A2(n15481), .ZN(n15483) );
  XNOR2_X1 U18649 ( .A(n15484), .B(n15483), .ZN(n16279) );
  AOI21_X1 U18650 ( .B1(n15487), .B2(n15486), .A(n15485), .ZN(n19066) );
  INV_X1 U18651 ( .A(n19066), .ZN(n19145) );
  NAND2_X1 U18652 ( .A1(n15488), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15496) );
  XNOR2_X1 U18653 ( .A(n15490), .B(n15489), .ZN(n19188) );
  INV_X1 U18654 ( .A(n19188), .ZN(n15494) );
  INV_X1 U18655 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19819) );
  NOR2_X1 U18656 ( .A1(n19819), .A2(n11494), .ZN(n15493) );
  NOR2_X1 U18657 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15491), .ZN(
        n15492) );
  AOI211_X1 U18658 ( .C1(n19261), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15495) );
  OAI211_X1 U18659 ( .C1(n19145), .C2(n19257), .A(n15496), .B(n15495), .ZN(
        n15497) );
  AOI21_X1 U18660 ( .B1(n16279), .B2(n16338), .A(n15497), .ZN(n15498) );
  OAI21_X1 U18661 ( .B1(n15499), .B2(n19264), .A(n15498), .ZN(P2_U3036) );
  INV_X1 U18662 ( .A(n15500), .ZN(n15501) );
  NOR2_X1 U18663 ( .A1(n15501), .A2(n16342), .ZN(n16323) );
  AND2_X1 U18664 ( .A1(n15565), .A2(n15501), .ZN(n15502) );
  NOR2_X1 U18665 ( .A1(n15520), .A2(n15502), .ZN(n16316) );
  INV_X1 U18666 ( .A(n19091), .ZN(n15508) );
  OR2_X1 U18667 ( .A1(n15504), .A2(n15503), .ZN(n15506) );
  NAND2_X1 U18668 ( .A1(n15506), .A2(n15505), .ZN(n19195) );
  OAI22_X1 U18669 ( .A1(n16331), .A2(n19195), .B1(n19814), .B2(n11494), .ZN(
        n15507) );
  AOI21_X1 U18670 ( .B1(n15508), .B2(n16333), .A(n15507), .ZN(n15509) );
  OAI21_X1 U18671 ( .B1(n16316), .B2(n16325), .A(n15509), .ZN(n15510) );
  AOI21_X1 U18672 ( .B1(n16323), .B2(n16325), .A(n15510), .ZN(n15513) );
  NAND2_X1 U18673 ( .A1(n15511), .A2(n16319), .ZN(n15512) );
  OAI211_X1 U18674 ( .C1(n15514), .C2(n19259), .A(n15513), .B(n15512), .ZN(
        P2_U3039) );
  OR2_X1 U18675 ( .A1(n15537), .A2(n15515), .ZN(n15516) );
  NAND2_X1 U18676 ( .A1(n15517), .A2(n15516), .ZN(n15519) );
  NAND2_X1 U18677 ( .A1(n15519), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15518) );
  OAI21_X1 U18678 ( .B1(n15519), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15518), .ZN(n16299) );
  NAND2_X1 U18679 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15545) );
  INV_X1 U18680 ( .A(n15520), .ZN(n16340) );
  AOI21_X1 U18681 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16340), .A(
        n15521), .ZN(n15557) );
  AOI21_X1 U18682 ( .B1(n15565), .B2(n15545), .A(n15557), .ZN(n15527) );
  XNOR2_X1 U18683 ( .A(n15522), .B(n15523), .ZN(n19197) );
  INV_X1 U18684 ( .A(n19197), .ZN(n15524) );
  AOI22_X1 U18685 ( .A1(n19261), .A2(n15524), .B1(P2_REIP_REG_6__SCAN_IN), 
        .B2(n16322), .ZN(n15525) );
  OAI21_X1 U18686 ( .B1(n15527), .B2(n15526), .A(n15525), .ZN(n15530) );
  NOR3_X1 U18687 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15528), .A3(
        n16342), .ZN(n15529) );
  AOI211_X1 U18688 ( .C1(n19105), .C2(n16333), .A(n15530), .B(n15529), .ZN(
        n15534) );
  XNOR2_X1 U18689 ( .A(n15532), .B(n9607), .ZN(n16298) );
  OR2_X1 U18690 ( .A1(n16298), .A2(n19259), .ZN(n15533) );
  OAI211_X1 U18691 ( .C1(n16299), .C2(n19264), .A(n15534), .B(n15533), .ZN(
        P2_U3040) );
  XNOR2_X1 U18692 ( .A(n15536), .B(n15535), .ZN(n16307) );
  INV_X1 U18693 ( .A(n15537), .ZN(n15543) );
  NAND2_X1 U18694 ( .A1(n15539), .A2(n15538), .ZN(n15540) );
  OAI21_X1 U18695 ( .B1(n15543), .B2(n15541), .A(n15540), .ZN(n15542) );
  OAI21_X1 U18696 ( .B1(n9602), .B2(n15543), .A(n15542), .ZN(n16309) );
  NOR2_X1 U18697 ( .A1(n16341), .A2(n16342), .ZN(n15556) );
  OAI211_X1 U18698 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15556), .B(n15545), .ZN(n15551) );
  XNOR2_X1 U18699 ( .A(n15547), .B(n15546), .ZN(n19204) );
  AOI22_X1 U18700 ( .A1(n19115), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15557), .ZN(n15548) );
  OAI21_X1 U18701 ( .B1(n16331), .B2(n19204), .A(n15548), .ZN(n15549) );
  AOI21_X1 U18702 ( .B1(n19121), .B2(n16333), .A(n15549), .ZN(n15550) );
  OAI211_X1 U18703 ( .C1(n16309), .C2(n19264), .A(n15551), .B(n15550), .ZN(
        n15552) );
  INV_X1 U18704 ( .A(n15552), .ZN(n15553) );
  OAI21_X1 U18705 ( .B1(n19259), .B2(n16307), .A(n15553), .ZN(P2_U3041) );
  NOR2_X1 U18706 ( .A1(n19808), .A2(n11494), .ZN(n15554) );
  AOI221_X1 U18707 ( .B1(n15557), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n15556), .C2(n15555), .A(n15554), .ZN(n15560) );
  AOI22_X1 U18708 ( .A1(n19155), .A2(n16333), .B1(n19261), .B2(n15558), .ZN(
        n15559) );
  NAND2_X1 U18709 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  AOI21_X1 U18710 ( .B1(n16319), .B2(n15562), .A(n15561), .ZN(n15563) );
  OAI21_X1 U18711 ( .B1(n15564), .B2(n19259), .A(n15563), .ZN(P2_U3042) );
  OAI211_X1 U18712 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15565), .B(n19275), .ZN(n15574) );
  AOI22_X1 U18713 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15567), .B1(
        n16333), .B2(n15566), .ZN(n15573) );
  AOI21_X1 U18714 ( .B1(n16319), .B2(n15569), .A(n15568), .ZN(n15572) );
  AOI22_X1 U18715 ( .A1(n19261), .A2(n19889), .B1(n15570), .B2(n16338), .ZN(
        n15571) );
  NAND4_X1 U18716 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        P2_U3045) );
  INV_X1 U18717 ( .A(n15575), .ZN(n15577) );
  INV_X1 U18718 ( .A(n11275), .ZN(n15576) );
  MUX2_X1 U18719 ( .A(n15577), .B(n15576), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15578) );
  OAI21_X1 U18720 ( .B1(n15579), .B2(n15593), .A(n15578), .ZN(n16344) );
  INV_X1 U18721 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19678) );
  AOI21_X1 U18722 ( .B1(n16344), .B2(n19678), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n15581) );
  INV_X1 U18723 ( .A(n15597), .ZN(n15580) );
  INV_X1 U18724 ( .A(n15594), .ZN(n16387) );
  OAI22_X1 U18725 ( .A1(n15581), .A2(n15580), .B1(n13060), .B2(n16387), .ZN(
        n15582) );
  MUX2_X1 U18726 ( .A(n15582), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15599), .Z(P2_U3601) );
  INV_X1 U18727 ( .A(n15583), .ZN(n15598) );
  INV_X1 U18728 ( .A(n19877), .ZN(n15595) );
  NOR2_X1 U18729 ( .A1(n15585), .A2(n15584), .ZN(n15588) );
  XNOR2_X1 U18730 ( .A(n10459), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15586) );
  AOI22_X1 U18731 ( .A1(n15587), .A2(n15588), .B1(n15586), .B2(n11275), .ZN(
        n15592) );
  INV_X1 U18732 ( .A(n15588), .ZN(n15589) );
  NAND2_X1 U18733 ( .A1(n15590), .A2(n15589), .ZN(n15591) );
  OAI211_X1 U18734 ( .C1(n19258), .C2(n15593), .A(n15592), .B(n15591), .ZN(
        n16343) );
  AOI22_X1 U18735 ( .A1(n15595), .A2(n15594), .B1(n19779), .B2(n16343), .ZN(
        n15596) );
  OAI21_X1 U18736 ( .B1(n15598), .B2(n15597), .A(n15596), .ZN(n15600) );
  MUX2_X1 U18737 ( .A(n15600), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15599), .Z(P2_U3599) );
  OAI21_X1 U18738 ( .B1(n19721), .B2(n15609), .A(n19869), .ZN(n15608) );
  NAND2_X1 U18739 ( .A1(n19577), .A2(n19891), .ZN(n19525) );
  INV_X1 U18740 ( .A(n19525), .ZN(n15601) );
  OR2_X1 U18741 ( .A1(n15608), .A2(n15601), .ZN(n15605) );
  OR2_X1 U18742 ( .A1(n10896), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15603) );
  NAND2_X1 U18743 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19891), .ZN(
        n19316) );
  NOR2_X1 U18744 ( .A1(n19316), .A2(n19582), .ZN(n19583) );
  NOR2_X1 U18745 ( .A1(n19583), .A2(n19869), .ZN(n15602) );
  AOI21_X1 U18746 ( .B1(n15603), .B2(n15602), .A(n19680), .ZN(n15604) );
  NAND2_X1 U18747 ( .A1(n15605), .A2(n15604), .ZN(n19574) );
  INV_X1 U18748 ( .A(n19574), .ZN(n19559) );
  INV_X1 U18749 ( .A(n10896), .ZN(n15606) );
  OAI21_X1 U18750 ( .B1(n15606), .B2(n19583), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15607) );
  OAI21_X1 U18751 ( .B1(n15608), .B2(n19525), .A(n15607), .ZN(n19573) );
  INV_X1 U18752 ( .A(n19572), .ZN(n19567) );
  AOI22_X1 U18753 ( .A1(n19689), .A2(n19584), .B1(n13381), .B2(n19583), .ZN(
        n15610) );
  OAI21_X1 U18754 ( .B1(n19567), .B2(n19692), .A(n15610), .ZN(n15611) );
  AOI21_X1 U18755 ( .B1(n13380), .B2(n19573), .A(n15611), .ZN(n15612) );
  OAI21_X1 U18756 ( .B1(n19559), .B2(n15613), .A(n15612), .ZN(P2_U3121) );
  NOR2_X1 U18757 ( .A1(n15614), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19646) );
  INV_X1 U18758 ( .A(n19646), .ZN(n15621) );
  INV_X1 U18759 ( .A(n15615), .ZN(n15623) );
  OAI21_X1 U18760 ( .B1(n15623), .B2(n19676), .A(n19678), .ZN(n15620) );
  AND2_X1 U18761 ( .A1(n15617), .A2(n15616), .ZN(n19406) );
  AOI21_X1 U18762 ( .B1(n19668), .B2(n19651), .A(n19467), .ZN(n15618) );
  AOI21_X1 U18763 ( .B1(n19406), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n15618), .ZN(n15619) );
  AOI211_X1 U18764 ( .C1(n15621), .C2(n15620), .A(n19680), .B(n15619), .ZN(
        n19628) );
  INV_X1 U18765 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U18766 ( .A1(n19637), .A2(n19652), .B1(n19670), .B2(n19728), .ZN(
        n15628) );
  INV_X1 U18767 ( .A(n15622), .ZN(n15626) );
  INV_X1 U18768 ( .A(n19406), .ZN(n15625) );
  OAI21_X1 U18769 ( .B1(n15623), .B2(n19646), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15624) );
  OAI21_X1 U18770 ( .B1(n15626), .B2(n15625), .A(n15624), .ZN(n19647) );
  AOI22_X1 U18771 ( .A1(n19647), .A2(n13454), .B1(n19718), .B2(n19646), .ZN(
        n15627) );
  OAI211_X1 U18772 ( .C1(n19628), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        P2_U3144) );
  INV_X1 U18773 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17061) );
  INV_X1 U18774 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20919) );
  INV_X1 U18775 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17121) );
  INV_X1 U18776 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17205) );
  INV_X1 U18777 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17267) );
  NOR3_X1 U18778 ( .A1(n18299), .A2(n18287), .A3(n15630), .ZN(n15631) );
  INV_X1 U18779 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16931) );
  NAND2_X1 U18780 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17285) );
  NOR2_X1 U18781 ( .A1(n16931), .A2(n17285), .ZN(n17276) );
  NAND3_X1 U18782 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17276), .ZN(n17278) );
  INV_X1 U18783 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17262) );
  INV_X1 U18784 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16801) );
  INV_X1 U18785 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16787) );
  NAND3_X1 U18786 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .ZN(n15634) );
  INV_X1 U18787 ( .A(n17016), .ZN(n17019) );
  NAND2_X1 U18788 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17019), .ZN(n15712) );
  INV_X1 U18789 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16969) );
  INV_X1 U18790 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16968) );
  NOR2_X1 U18791 ( .A1(n17295), .A2(n17009), .ZN(n17010) );
  AOI22_X1 U18792 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15635) );
  OAI21_X1 U18793 ( .B1(n17148), .B2(n17079), .A(n15635), .ZN(n15644) );
  AOI22_X1 U18794 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15642) );
  OAI22_X1 U18795 ( .A1(n10131), .A2(n17087), .B1(n9616), .B2(n18605), .ZN(
        n15640) );
  AOI22_X1 U18796 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15638) );
  AOI22_X1 U18797 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U18798 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17258), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15636) );
  NAND3_X1 U18799 ( .A1(n15638), .A2(n15637), .A3(n15636), .ZN(n15639) );
  AOI211_X1 U18800 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n15640), .B(n15639), .ZN(n15641) );
  OAI211_X1 U18801 ( .C1(n9651), .C2(n17282), .A(n15642), .B(n15641), .ZN(
        n15643) );
  AOI211_X1 U18802 ( .C1(n9576), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15644), .B(n15643), .ZN(n17017) );
  AOI22_X1 U18803 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9586), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10178), .ZN(n15645) );
  OAI21_X1 U18804 ( .B1(n9652), .B2(n17106), .A(n15645), .ZN(n15654) );
  AOI22_X1 U18805 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17251), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17244), .ZN(n15652) );
  OAI22_X1 U18806 ( .A1(n17107), .A2(n17156), .B1(n18597), .B2(n9616), .ZN(
        n15650) );
  AOI22_X1 U18807 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15648) );
  AOI22_X1 U18808 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17243), .ZN(n15647) );
  AOI22_X1 U18809 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10247), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17258), .ZN(n15646) );
  NAND3_X1 U18810 ( .A1(n15648), .A2(n15647), .A3(n15646), .ZN(n15649) );
  AOI211_X1 U18811 ( .C1(n10142), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n15650), .B(n15649), .ZN(n15651) );
  OAI211_X1 U18812 ( .C1(n9651), .C2(n17290), .A(n15652), .B(n15651), .ZN(
        n15653) );
  AOI211_X1 U18813 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n15654), .B(n15653), .ZN(n17025) );
  AOI22_X1 U18814 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10247), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U18815 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18816 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15655) );
  OAI211_X1 U18817 ( .C1(n9616), .C2(n18593), .A(n15656), .B(n15655), .ZN(
        n15662) );
  AOI22_X1 U18818 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18819 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15659) );
  AOI22_X1 U18820 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15658) );
  NAND2_X1 U18821 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15657) );
  NAND4_X1 U18822 ( .A1(n15660), .A2(n15659), .A3(n15658), .A4(n15657), .ZN(
        n15661) );
  AOI211_X1 U18823 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n15662), .B(n15661), .ZN(n15663) );
  OAI211_X1 U18824 ( .C1(n9651), .C2(n20925), .A(n15664), .B(n15663), .ZN(
        n17029) );
  AOI22_X1 U18825 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15675) );
  INV_X1 U18826 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U18827 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18828 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15665) );
  OAI211_X1 U18829 ( .C1(n9616), .C2(n15667), .A(n15666), .B(n15665), .ZN(
        n15673) );
  AOI22_X1 U18830 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U18831 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U18832 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15669) );
  NAND2_X1 U18833 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15668) );
  NAND4_X1 U18834 ( .A1(n15671), .A2(n15670), .A3(n15669), .A4(n15668), .ZN(
        n15672) );
  AOI211_X1 U18835 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15673), .B(n15672), .ZN(n15674) );
  OAI211_X1 U18836 ( .C1(n17224), .C2(n17264), .A(n15675), .B(n15674), .ZN(
        n17030) );
  NAND2_X1 U18837 ( .A1(n17029), .A2(n17030), .ZN(n17028) );
  NOR2_X1 U18838 ( .A1(n17025), .A2(n17028), .ZN(n17022) );
  AOI22_X1 U18839 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18840 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18841 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15676) );
  OAI211_X1 U18842 ( .C1(n17142), .C2(n15678), .A(n15677), .B(n15676), .ZN(
        n15684) );
  AOI22_X1 U18843 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18844 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15681) );
  AOI22_X1 U18845 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15680) );
  NAND2_X1 U18846 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n15679) );
  NAND4_X1 U18847 ( .A1(n15682), .A2(n15681), .A3(n15680), .A4(n15679), .ZN(
        n15683) );
  AOI211_X1 U18848 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n15684), .B(n15683), .ZN(n15685) );
  OAI211_X1 U18849 ( .C1(n15688), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        n17021) );
  NAND2_X1 U18850 ( .A1(n17022), .A2(n17021), .ZN(n17020) );
  NOR2_X1 U18851 ( .A1(n17017), .A2(n17020), .ZN(n17014) );
  AOI22_X1 U18852 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15698) );
  AOI22_X1 U18853 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15697) );
  AOI22_X1 U18854 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15696) );
  OAI22_X1 U18855 ( .A1(n10131), .A2(n17182), .B1(n17199), .B2(n17173), .ZN(
        n15694) );
  AOI22_X1 U18856 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15692) );
  AOI22_X1 U18857 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15691) );
  AOI22_X1 U18858 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15690) );
  NAND2_X1 U18859 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n15689) );
  NAND4_X1 U18860 ( .A1(n15692), .A2(n15691), .A3(n15690), .A4(n15689), .ZN(
        n15693) );
  NAND4_X1 U18861 ( .A1(n15698), .A2(n15697), .A3(n15696), .A4(n15695), .ZN(
        n17013) );
  NAND2_X1 U18862 ( .A1(n17014), .A2(n17013), .ZN(n17012) );
  INV_X1 U18863 ( .A(n17012), .ZN(n17004) );
  AOI22_X1 U18864 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U18865 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U18866 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17258), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15708) );
  OAI22_X1 U18867 ( .A1(n17199), .A2(n15700), .B1(n9722), .B2(n15699), .ZN(
        n15706) );
  AOI22_X1 U18868 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U18869 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18870 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15702) );
  NAND2_X1 U18871 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n15701) );
  NAND4_X1 U18872 ( .A1(n15704), .A2(n15703), .A3(n15702), .A4(n15701), .ZN(
        n15705) );
  AOI211_X1 U18873 ( .C1(n10178), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n15706), .B(n15705), .ZN(n15707) );
  NAND4_X1 U18874 ( .A1(n15710), .A2(n15709), .A3(n15708), .A4(n15707), .ZN(
        n17005) );
  XOR2_X1 U18875 ( .A(n17004), .B(n17005), .Z(n17317) );
  AOI22_X1 U18876 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17010), .B1(n17295), 
        .B2(n17317), .ZN(n15711) );
  OAI21_X1 U18877 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15712), .A(n15711), .ZN(
        P3_U2675) );
  AOI22_X1 U18878 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15713) );
  OAI21_X1 U18879 ( .B1(n9722), .B2(n17050), .A(n15713), .ZN(n15724) );
  INV_X1 U18880 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15722) );
  AOI22_X1 U18881 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15721) );
  AOI22_X1 U18882 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15714) );
  OAI21_X1 U18883 ( .B1(n9612), .B2(n17275), .A(n15714), .ZN(n15719) );
  INV_X1 U18884 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15717) );
  AOI22_X1 U18885 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15716) );
  AOI22_X1 U18886 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15715) );
  OAI211_X1 U18887 ( .C1(n9649), .C2(n15717), .A(n15716), .B(n15715), .ZN(
        n15718) );
  AOI211_X1 U18888 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15719), .B(n15718), .ZN(n15720) );
  OAI211_X1 U18889 ( .C1(n17199), .C2(n15722), .A(n15721), .B(n15720), .ZN(
        n15723) );
  AOI211_X1 U18890 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n15724), .B(n15723), .ZN(n17394) );
  NOR2_X1 U18891 ( .A1(n18299), .A2(n17202), .ZN(n17185) );
  NAND2_X1 U18892 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17185), .ZN(n15725) );
  NOR2_X1 U18893 ( .A1(n16801), .A2(n15725), .ZN(n17153) );
  INV_X1 U18894 ( .A(n15725), .ZN(n17187) );
  AOI21_X1 U18895 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n9582), .A(n17187), .ZN(
        n15726) );
  OAI22_X1 U18896 ( .A1(n17394), .A2(n9582), .B1(n17153), .B2(n15726), .ZN(
        P3_U2690) );
  INV_X1 U18897 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18273) );
  NAND2_X1 U18898 ( .A1(n18273), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18307) );
  NAND3_X1 U18899 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18861)
         );
  INV_X1 U18900 ( .A(n18732), .ZN(n18715) );
  AOI211_X1 U18901 ( .C1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n18715), .A(
        n17244), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18258) );
  INV_X1 U18902 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16558) );
  OR2_X1 U18903 ( .A1(n16558), .A2(n18861), .ZN(n15739) );
  OAI211_X1 U18904 ( .C1(n18861), .C2(n18258), .A(n18372), .B(n15739), .ZN(
        n18265) );
  NAND2_X1 U18905 ( .A1(n18307), .A2(n18265), .ZN(n15729) );
  INV_X1 U18906 ( .A(n15729), .ZN(n15728) );
  OAI22_X1 U18907 ( .A1(n18909), .A2(n17676), .B1(n18273), .B2(n18862), .ZN(
        n15731) );
  NAND3_X1 U18908 ( .A1(n18397), .A2(n18265), .A3(n15731), .ZN(n15727) );
  OAI221_X1 U18909 ( .B1(n18397), .B2(n15728), .C1(n18397), .C2(n18513), .A(
        n15727), .ZN(P3_U2864) );
  NAND2_X1 U18910 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18490) );
  NOR2_X1 U18911 ( .A1(n18909), .A2(n17676), .ZN(n15730) );
  AOI221_X1 U18912 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18490), .C1(n15730), 
        .C2(n18490), .A(n15729), .ZN(n18264) );
  INV_X1 U18913 ( .A(n18513), .ZN(n18621) );
  OAI221_X1 U18914 ( .B1(n18621), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18621), .C2(n15731), .A(n18265), .ZN(n18262) );
  AOI22_X1 U18915 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18264), .B1(
        n18262), .B2(n18271), .ZN(P3_U2865) );
  INV_X1 U18916 ( .A(n18918), .ZN(n18912) );
  INV_X1 U18917 ( .A(n16555), .ZN(n18702) );
  NAND2_X1 U18918 ( .A1(n18702), .A2(n18918), .ZN(n15735) );
  INV_X1 U18919 ( .A(n18915), .ZN(n16577) );
  OAI21_X1 U18920 ( .B1(n15735), .B2(n17457), .A(n15734), .ZN(n15736) );
  NAND2_X1 U18921 ( .A1(n18859), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18267) );
  INV_X1 U18922 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16901) );
  INV_X1 U18923 ( .A(n18928), .ZN(n18889) );
  AOI21_X1 U18924 ( .B1(n18715), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15742) );
  NAND2_X1 U18925 ( .A1(n16575), .A2(n15740), .ZN(n15741) );
  NOR2_X1 U18926 ( .A1(n15742), .A2(n15741), .ZN(n18709) );
  NAND3_X1 U18927 ( .A1(n18891), .A2(n18889), .A3(n18709), .ZN(n15743) );
  OAI21_X1 U18928 ( .B1(n18891), .B2(n16901), .A(n15743), .ZN(P3_U3284) );
  INV_X1 U18929 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15754) );
  AOI21_X1 U18930 ( .B1(n16433), .B2(n15745), .A(n15744), .ZN(n15746) );
  XNOR2_X1 U18931 ( .A(n15754), .B(n15746), .ZN(n16424) );
  INV_X1 U18932 ( .A(n18057), .ZN(n18136) );
  AOI21_X1 U18933 ( .B1(n18136), .B2(n17928), .A(n15747), .ZN(n16441) );
  OAI22_X1 U18934 ( .A1(n16420), .A2(n18172), .B1(n16406), .B2(n18210), .ZN(
        n15748) );
  NOR2_X1 U18935 ( .A1(n18211), .A2(n15748), .ZN(n15801) );
  OR2_X1 U18936 ( .A1(n18240), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15749) );
  OAI211_X1 U18937 ( .C1(n16441), .C2(n18254), .A(n15801), .B(n15749), .ZN(
        n15750) );
  AOI22_X1 U18938 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15750), .B1(
        n9587), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U18939 ( .A1(n17932), .A2(n18250), .B1(n17931), .B2(n15751), .ZN(
        n15753) );
  NAND2_X1 U18940 ( .A1(n15753), .A2(n15752), .ZN(n15803) );
  NAND3_X1 U18941 ( .A1(n15755), .A2(n15754), .A3(n15803), .ZN(n15756) );
  OAI211_X1 U18942 ( .C1(n16424), .C2(n18144), .A(n15757), .B(n15756), .ZN(
        P3_U2833) );
  INV_X1 U18943 ( .A(n15758), .ZN(n15771) );
  OAI211_X1 U18944 ( .C1(n15761), .C2(n15760), .A(n15759), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15765) );
  INV_X1 U18945 ( .A(n15762), .ZN(n15764) );
  OAI211_X1 U18946 ( .C1(n20476), .C2(n15765), .A(n15764), .B(n15763), .ZN(
        n15767) );
  NAND2_X1 U18947 ( .A1(n15765), .A2(n20476), .ZN(n15766) );
  NAND2_X1 U18948 ( .A1(n15767), .A2(n15766), .ZN(n15768) );
  AOI222_X1 U18949 ( .A1(n15769), .A2(n15768), .B1(n15769), .B2(n20560), .C1(
        n15768), .C2(n20560), .ZN(n15770) );
  AOI222_X1 U18950 ( .A1(n15771), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n15771), .B2(n15770), .C1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n15770), .ZN(n15779) );
  OAI21_X1 U18951 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15772), .ZN(n15773) );
  NAND4_X1 U18952 ( .A1(n15776), .A2(n15775), .A3(n15774), .A4(n15773), .ZN(
        n15777) );
  AOI211_X1 U18953 ( .C1(n20103), .C2(n15779), .A(n15778), .B(n15777), .ZN(
        n15793) );
  NOR2_X1 U18954 ( .A1(n15780), .A2(n15805), .ZN(n15783) );
  INV_X1 U18955 ( .A(n20864), .ZN(n20781) );
  AOI21_X1 U18956 ( .B1(n20858), .B2(n20781), .A(n15781), .ZN(n15782) );
  AOI21_X1 U18957 ( .B1(n15784), .B2(n15783), .A(n15782), .ZN(n16222) );
  OAI221_X1 U18958 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15793), 
        .A(n16222), .ZN(n16229) );
  AND2_X1 U18959 ( .A1(n16227), .A2(n15785), .ZN(n15786) );
  NOR2_X1 U18960 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15786), .ZN(n15791) );
  INV_X1 U18961 ( .A(n16224), .ZN(n15787) );
  AOI211_X1 U18962 ( .C1(n20781), .C2(n20856), .A(n15788), .B(n15787), .ZN(
        n15789) );
  NAND2_X1 U18963 ( .A1(n16229), .A2(n15789), .ZN(n15790) );
  AOI22_X1 U18964 ( .A1(n16229), .A2(n15791), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15790), .ZN(n15792) );
  OAI21_X1 U18965 ( .B1(n15793), .B2(n19913), .A(n15792), .ZN(P1_U3161) );
  INV_X1 U18966 ( .A(n15794), .ZN(n15796) );
  NOR2_X1 U18967 ( .A1(n15796), .A2(n15795), .ZN(n15797) );
  XOR2_X1 U18968 ( .A(n15797), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16405) );
  NOR2_X1 U18969 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15798), .ZN(
        n16400) );
  AOI21_X1 U18970 ( .B1(n15801), .B2(n15800), .A(n15799), .ZN(n15802) );
  AOI21_X1 U18971 ( .B1(n16400), .B2(n15803), .A(n15802), .ZN(n15804) );
  NAND2_X1 U18972 ( .A1(n9587), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16396) );
  OAI211_X1 U18973 ( .C1(n16405), .C2(n18144), .A(n15804), .B(n16396), .ZN(
        P3_U2832) );
  INV_X1 U18974 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20790) );
  NOR2_X1 U18975 ( .A1(n20970), .A2(n20790), .ZN(n20786) );
  INV_X1 U18976 ( .A(HOLD), .ZN(n20782) );
  INV_X1 U18977 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20794) );
  OAI222_X1 U18978 ( .A1(n20786), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n20786), 
        .B2(HOLD), .C1(n20782), .C2(n20794), .ZN(n15806) );
  OAI211_X1 U18979 ( .C1(n20864), .C2(n11754), .A(n15806), .B(n15805), .ZN(
        P1_U3195) );
  AND2_X1 U18980 ( .A1(n20043), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AND3_X1 U18981 ( .A1(n15816), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16092), .ZN(n15819) );
  OAI21_X1 U18982 ( .B1(n15808), .B2(n15816), .A(n15807), .ZN(n15809) );
  INV_X1 U18983 ( .A(n15809), .ZN(n15974) );
  NAND2_X1 U18984 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15810), .ZN(
        n15811) );
  OAI22_X1 U18985 ( .A1(n15814), .A2(n15813), .B1(n15812), .B2(n15811), .ZN(
        n16134) );
  OR2_X1 U18986 ( .A1(n16134), .A2(n20098), .ZN(n15815) );
  AOI21_X1 U18987 ( .B1(n16091), .B2(n15815), .A(n16093), .ZN(n15817) );
  OAI22_X1 U18988 ( .A1(n15974), .A2(n16204), .B1(n15817), .B2(n15816), .ZN(
        n15818) );
  AOI211_X1 U18989 ( .C1(P1_REIP_REG_20__SCAN_IN), .C2(n12840), .A(n15819), 
        .B(n15818), .ZN(n15820) );
  OAI21_X1 U18990 ( .B1(n16159), .B2(n15861), .A(n15820), .ZN(P1_U3011) );
  NOR2_X1 U18991 ( .A1(n19786), .A2(n21039), .ZN(n19778) );
  NAND2_X1 U18992 ( .A1(n19778), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15822) );
  AND2_X1 U18993 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19883) );
  AOI21_X1 U18994 ( .B1(n19883), .B2(n21039), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15821) );
  AOI21_X1 U18995 ( .B1(n15822), .B2(n15821), .A(n15824), .ZN(P2_U3178) );
  INV_X1 U18996 ( .A(n15823), .ZN(n19904) );
  AOI221_X1 U18997 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15824), .C1(n19904), .C2(
        n15824), .A(n19726), .ZN(n19901) );
  AND2_X1 U18998 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19901), .ZN(
        P2_U3047) );
  NOR3_X1 U18999 ( .A1(n15825), .A2(n18269), .A3(n18277), .ZN(n15826) );
  INV_X1 U19000 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17527) );
  NOR2_X2 U19001 ( .A1(n15828), .A2(n17527), .ZN(n17454) );
  OR2_X1 U19002 ( .A1(n18299), .A2(n15828), .ZN(n17304) );
  AOI22_X1 U19003 ( .A1(n17451), .A2(BUF2_REG_0__SCAN_IN), .B1(n17450), .B2(
        n17921), .ZN(n15829) );
  OAI221_X1 U19004 ( .B1(n17454), .B2(n17527), .C1(n17454), .C2(n17304), .A(
        n15829), .ZN(P3_U2735) );
  AOI22_X1 U19005 ( .A1(n19963), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19989), .ZN(n15837) );
  INV_X1 U19006 ( .A(n15830), .ZN(n15956) );
  INV_X1 U19007 ( .A(n15845), .ZN(n15831) );
  NOR2_X1 U19008 ( .A1(n19994), .A2(n15831), .ZN(n15860) );
  AOI21_X1 U19009 ( .B1(n15832), .B2(n15860), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15834) );
  OAI22_X1 U19010 ( .A1(n16078), .A2(n20005), .B1(n15834), .B2(n15833), .ZN(
        n15835) );
  AOI21_X1 U19011 ( .B1(n15956), .B2(n12623), .A(n15835), .ZN(n15836) );
  OAI211_X1 U19012 ( .C1(n15959), .C2(n19974), .A(n15837), .B(n15836), .ZN(
        P1_U2817) );
  INV_X1 U19013 ( .A(n15860), .ZN(n15838) );
  NOR3_X1 U19014 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15839), .A3(n15838), 
        .ZN(n15843) );
  OAI22_X1 U19015 ( .A1(n15883), .A2(n15841), .B1(n15840), .B2(n19949), .ZN(
        n15842) );
  AOI211_X1 U19016 ( .C1(n19987), .C2(n15844), .A(n15843), .B(n15842), .ZN(
        n15850) );
  AND2_X1 U19017 ( .A1(n15845), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15852) );
  NAND2_X1 U19018 ( .A1(n15872), .A2(n15852), .ZN(n15846) );
  NAND2_X1 U19019 ( .A1(n15924), .A2(n15846), .ZN(n15862) );
  OAI21_X1 U19020 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19994), .A(n15862), 
        .ZN(n15847) );
  AOI22_X1 U19021 ( .A1(n15848), .A2(n12623), .B1(P1_REIP_REG_22__SCAN_IN), 
        .B2(n15847), .ZN(n15849) );
  OAI211_X1 U19022 ( .C1(n20005), .C2(n16082), .A(n15850), .B(n15849), .ZN(
        P1_U2818) );
  INV_X1 U19023 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20820) );
  INV_X1 U19024 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15969) );
  OAI22_X1 U19025 ( .A1(n15969), .A2(n19949), .B1(n19974), .B2(n15961), .ZN(
        n15851) );
  AOI21_X1 U19026 ( .B1(n19963), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15851), .ZN(
        n15854) );
  NAND3_X1 U19027 ( .A1(n19962), .A2(n20820), .A3(n15852), .ZN(n15853) );
  OAI211_X1 U19028 ( .C1(n15862), .C2(n20820), .A(n15854), .B(n15853), .ZN(
        n15855) );
  INV_X1 U19029 ( .A(n15855), .ZN(n15859) );
  OAI22_X1 U19030 ( .A1(n15965), .A2(n19954), .B1(n15856), .B2(n20005), .ZN(
        n15857) );
  INV_X1 U19031 ( .A(n15857), .ZN(n15858) );
  NAND2_X1 U19032 ( .A1(n15859), .A2(n15858), .ZN(P1_U2819) );
  AOI22_X1 U19033 ( .A1(n19963), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n19987), 
        .B2(n15970), .ZN(n15866) );
  NOR2_X1 U19034 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15860), .ZN(n15863) );
  OAI22_X1 U19035 ( .A1(n15863), .A2(n15862), .B1(n15861), .B2(n20005), .ZN(
        n15864) );
  AOI21_X1 U19036 ( .B1(n15971), .B2(n12623), .A(n15864), .ZN(n15865) );
  OAI211_X1 U19037 ( .C1(n15867), .C2(n19949), .A(n15866), .B(n15865), .ZN(
        P1_U2820) );
  NOR3_X1 U19038 ( .A1(n19994), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15868), 
        .ZN(n15869) );
  AOI211_X1 U19039 ( .C1(n19989), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15869), .B(n12840), .ZN(n15879) );
  INV_X1 U19040 ( .A(n15981), .ZN(n15870) );
  AOI22_X1 U19041 ( .A1(n19963), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n15870), 
        .B2(n19987), .ZN(n15878) );
  INV_X1 U19042 ( .A(n15871), .ZN(n15978) );
  AOI22_X1 U19043 ( .A1(n15978), .A2(n12623), .B1(n16089), .B2(n19977), .ZN(
        n15877) );
  OAI21_X1 U19044 ( .B1(n19994), .B2(n15873), .A(n15872), .ZN(n15891) );
  INV_X1 U19045 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15874) );
  NAND2_X1 U19046 ( .A1(n15874), .A2(n15873), .ZN(n15875) );
  NOR2_X1 U19047 ( .A1(n19994), .A2(n15875), .ZN(n15880) );
  OAI21_X1 U19048 ( .B1(n15891), .B2(n15880), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15876) );
  NAND4_X1 U19049 ( .A1(n15879), .A2(n15878), .A3(n15877), .A4(n15876), .ZN(
        P1_U2821) );
  INV_X1 U19050 ( .A(n15880), .ZN(n15882) );
  AOI21_X1 U19051 ( .B1(n19989), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12840), .ZN(n15881) );
  OAI211_X1 U19052 ( .C1(n15884), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15885) );
  AOI21_X1 U19053 ( .B1(n15886), .B2(n19987), .A(n15885), .ZN(n15889) );
  AOI22_X1 U19054 ( .A1(n15887), .A2(n12623), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n15891), .ZN(n15888) );
  OAI211_X1 U19055 ( .C1(n20005), .C2(n16096), .A(n15889), .B(n15888), .ZN(
        P1_U2822) );
  AOI22_X1 U19056 ( .A1(n19963), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19989), .ZN(n15896) );
  AOI21_X1 U19057 ( .B1(n19987), .B2(n15982), .A(n12840), .ZN(n15895) );
  AOI22_X1 U19058 ( .A1(n15983), .A2(n12623), .B1(n19977), .B2(n15890), .ZN(
        n15894) );
  OAI221_X1 U19059 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n15892), .A(n15891), .ZN(n15893) );
  NAND4_X1 U19060 ( .A1(n15896), .A2(n15895), .A3(n15894), .A4(n15893), .ZN(
        P1_U2823) );
  AOI22_X1 U19061 ( .A1(n15897), .A2(n19987), .B1(n19977), .B2(n16119), .ZN(
        n15903) );
  AOI22_X1 U19062 ( .A1(n15910), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n19963), 
        .B2(P1_EBX_REG_15__SCAN_IN), .ZN(n15902) );
  AOI21_X1 U19063 ( .B1(n19989), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n12840), .ZN(n15901) );
  INV_X1 U19064 ( .A(n15995), .ZN(n15899) );
  AOI21_X1 U19065 ( .B1(n15899), .B2(n12623), .A(n15898), .ZN(n15900) );
  NAND4_X1 U19066 ( .A1(n15903), .A2(n15902), .A3(n15901), .A4(n15900), .ZN(
        P1_U2825) );
  AND2_X1 U19067 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15904), .ZN(n15909) );
  AOI21_X1 U19068 ( .B1(n19989), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n12840), .ZN(n15906) );
  NAND2_X1 U19069 ( .A1(n19963), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n15905) );
  OAI211_X1 U19070 ( .C1(n15907), .C2(n19954), .A(n15906), .B(n15905), .ZN(
        n15908) );
  AOI221_X1 U19071 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15910), .C1(n15909), 
        .C2(n15910), .A(n15908), .ZN(n15913) );
  NAND2_X1 U19072 ( .A1(n15911), .A2(n19987), .ZN(n15912) );
  OAI211_X1 U19073 ( .C1(n16133), .C2(n20005), .A(n15913), .B(n15912), .ZN(
        P1_U2826) );
  OAI21_X1 U19074 ( .B1(n19949), .B2(n15914), .A(n20101), .ZN(n15917) );
  NOR2_X1 U19075 ( .A1(n15915), .A2(n20005), .ZN(n15916) );
  AOI211_X1 U19076 ( .C1(n19963), .C2(P1_EBX_REG_12__SCAN_IN), .A(n15917), .B(
        n15916), .ZN(n15923) );
  INV_X1 U19077 ( .A(n15918), .ZN(n19938) );
  NOR2_X1 U19078 ( .A1(n19981), .A2(n19938), .ZN(n19944) );
  NAND3_X1 U19079 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n19944), .ZN(n15932) );
  OAI21_X1 U19080 ( .B1(n15931), .B2(n15932), .A(n15919), .ZN(n15920) );
  AOI22_X1 U19081 ( .A1(n16001), .A2(n19987), .B1(n15921), .B2(n15920), .ZN(
        n15922) );
  OAI211_X1 U19082 ( .C1(n19954), .C2(n15999), .A(n15923), .B(n15922), .ZN(
        P1_U2828) );
  OAI21_X1 U19083 ( .B1(n15926), .B2(n15925), .A(n15924), .ZN(n15940) );
  AOI21_X1 U19084 ( .B1(n19989), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n12840), .ZN(n15928) );
  AOI22_X1 U19085 ( .A1(n16142), .A2(n19977), .B1(n19963), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15927) );
  OAI211_X1 U19086 ( .C1(n16011), .C2(n19974), .A(n15928), .B(n15927), .ZN(
        n15929) );
  AOI21_X1 U19087 ( .B1(n12623), .B2(n16008), .A(n15929), .ZN(n15930) );
  OAI221_X1 U19088 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15932), .C1(n15931), 
        .C2(n15940), .A(n15930), .ZN(P1_U2829) );
  NAND2_X1 U19089 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19944), .ZN(n15942) );
  INV_X1 U19090 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15941) );
  AOI21_X1 U19091 ( .B1(n19989), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n12840), .ZN(n15933) );
  OAI21_X1 U19092 ( .B1(n19974), .B2(n15934), .A(n15933), .ZN(n15935) );
  AOI21_X1 U19093 ( .B1(n19963), .B2(P1_EBX_REG_10__SCAN_IN), .A(n15935), .ZN(
        n15936) );
  OAI21_X1 U19094 ( .B1(n16158), .B2(n20005), .A(n15936), .ZN(n15937) );
  AOI21_X1 U19095 ( .B1(n15938), .B2(n12623), .A(n15937), .ZN(n15939) );
  OAI221_X1 U19096 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15942), .C1(n15941), 
        .C2(n15940), .A(n15939), .ZN(P1_U2830) );
  INV_X1 U19097 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19098 ( .A1(n9726), .A2(n15943), .B1(P1_EAX_REG_23__SCAN_IN), .B2(
        n15946), .ZN(n15945) );
  AOI22_X1 U19099 ( .A1(n15956), .A2(n15950), .B1(n15949), .B2(DATAI_23_), 
        .ZN(n15944) );
  OAI211_X1 U19100 ( .C1(n15953), .C2(n16465), .A(n15945), .B(n15944), .ZN(
        P1_U2881) );
  INV_X1 U19101 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U19102 ( .A1(n9726), .A2(n15947), .B1(P1_EAX_REG_20__SCAN_IN), .B2(
        n15946), .ZN(n15952) );
  AOI22_X1 U19103 ( .A1(n15971), .A2(n15950), .B1(n15949), .B2(DATAI_20_), 
        .ZN(n15951) );
  OAI211_X1 U19104 ( .C1(n15953), .C2(n16471), .A(n15952), .B(n15951), .ZN(
        P1_U2884) );
  AOI22_X1 U19105 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15958) );
  XNOR2_X1 U19106 ( .A(n12833), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15954) );
  XNOR2_X1 U19107 ( .A(n15955), .B(n15954), .ZN(n16075) );
  AOI22_X1 U19108 ( .A1(n15956), .A2(n16029), .B1(n20087), .B2(n16075), .ZN(
        n15957) );
  OAI211_X1 U19109 ( .C1(n16023), .C2(n15959), .A(n15958), .B(n15957), .ZN(
        P1_U2976) );
  NAND2_X1 U19110 ( .A1(n15960), .A2(n20087), .ZN(n15964) );
  INV_X1 U19111 ( .A(n15961), .ZN(n15962) );
  NAND2_X1 U19112 ( .A1(n16027), .A2(n15962), .ZN(n15963) );
  OAI211_X1 U19113 ( .C1(n20106), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        n15966) );
  INV_X1 U19114 ( .A(n15966), .ZN(n15968) );
  OAI211_X1 U19115 ( .C1(n15969), .C2(n16033), .A(n15968), .B(n15967), .ZN(
        P1_U2978) );
  AOI22_X1 U19116 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15973) );
  AOI22_X1 U19117 ( .A1(n15971), .A2(n16029), .B1(n16027), .B2(n15970), .ZN(
        n15972) );
  OAI211_X1 U19118 ( .C1(n15974), .C2(n19920), .A(n15973), .B(n15972), .ZN(
        P1_U2979) );
  AOI22_X1 U19119 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15980) );
  NAND2_X1 U19120 ( .A1(n14480), .A2(n16101), .ZN(n15976) );
  MUX2_X1 U19121 ( .A(n14480), .B(n15976), .S(n15975), .Z(n15977) );
  XNOR2_X1 U19122 ( .A(n15977), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16090) );
  AOI22_X1 U19123 ( .A1(n15978), .A2(n16029), .B1(n20087), .B2(n16090), .ZN(
        n15979) );
  OAI211_X1 U19124 ( .C1(n16023), .C2(n15981), .A(n15980), .B(n15979), .ZN(
        P1_U2980) );
  AOI22_X1 U19125 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15985) );
  AOI22_X1 U19126 ( .A1(n15983), .A2(n16029), .B1(n15982), .B2(n16027), .ZN(
        n15984) );
  OAI211_X1 U19127 ( .C1(n19920), .C2(n15986), .A(n15985), .B(n15984), .ZN(
        P1_U2982) );
  INV_X1 U19128 ( .A(n15987), .ZN(n15988) );
  NOR2_X1 U19129 ( .A1(n15989), .A2(n15988), .ZN(n15993) );
  NAND2_X1 U19130 ( .A1(n15991), .A2(n15990), .ZN(n15992) );
  XNOR2_X1 U19131 ( .A(n15993), .B(n15992), .ZN(n16116) );
  AOI22_X1 U19132 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15998) );
  OAI22_X1 U19133 ( .A1(n15995), .A2(n20106), .B1(n15994), .B2(n16023), .ZN(
        n15996) );
  INV_X1 U19134 ( .A(n15996), .ZN(n15997) );
  OAI211_X1 U19135 ( .C1(n16116), .C2(n19920), .A(n15998), .B(n15997), .ZN(
        P1_U2984) );
  AOI22_X1 U19136 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16003) );
  INV_X1 U19137 ( .A(n15999), .ZN(n16000) );
  AOI22_X1 U19138 ( .A1(n16027), .A2(n16001), .B1(n16029), .B2(n16000), .ZN(
        n16002) );
  OAI211_X1 U19139 ( .C1(n16004), .C2(n19920), .A(n16003), .B(n16002), .ZN(
        P1_U2987) );
  AOI22_X1 U19140 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16010) );
  NOR3_X1 U19141 ( .A1(n14488), .A2(n12833), .A3(n12823), .ZN(n16006) );
  NOR2_X1 U19142 ( .A1(n16006), .A2(n16005), .ZN(n16007) );
  XNOR2_X1 U19143 ( .A(n16007), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16144) );
  AOI22_X1 U19144 ( .A1(n20087), .A2(n16144), .B1(n16029), .B2(n16008), .ZN(
        n16009) );
  OAI211_X1 U19145 ( .C1(n16023), .C2(n16011), .A(n16010), .B(n16009), .ZN(
        P1_U2988) );
  AOI22_X1 U19146 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16016) );
  XNOR2_X1 U19147 ( .A(n16013), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16014) );
  XNOR2_X1 U19148 ( .A(n16012), .B(n16014), .ZN(n16191) );
  AOI22_X1 U19149 ( .A1(n16191), .A2(n20087), .B1(n16029), .B2(n20011), .ZN(
        n16015) );
  OAI211_X1 U19150 ( .C1(n16023), .C2(n19967), .A(n16016), .B(n16015), .ZN(
        P1_U2992) );
  AOI22_X1 U19151 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12840), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16022) );
  NAND2_X1 U19152 ( .A1(n16019), .A2(n16018), .ZN(n16020) );
  XNOR2_X1 U19153 ( .A(n16017), .B(n16020), .ZN(n16197) );
  AOI22_X1 U19154 ( .A1(n16197), .A2(n20087), .B1(n16029), .B2(n19984), .ZN(
        n16021) );
  OAI211_X1 U19155 ( .C1(n16023), .C2(n19975), .A(n16022), .B(n16021), .ZN(
        P1_U2993) );
  XNOR2_X1 U19156 ( .A(n16024), .B(n16025), .ZN(n16203) );
  INV_X1 U19157 ( .A(n16203), .ZN(n16031) );
  INV_X1 U19158 ( .A(n16026), .ZN(n16028) );
  AOI222_X1 U19159 ( .A1(n16031), .A2(n20087), .B1(n16030), .B2(n16029), .C1(
        n16028), .C2(n16027), .ZN(n16032) );
  NAND2_X1 U19160 ( .A1(n12840), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16202) );
  OAI211_X1 U19161 ( .C1(n16034), .C2(n16033), .A(n16032), .B(n16202), .ZN(
        P1_U2994) );
  INV_X1 U19162 ( .A(n16035), .ZN(n16037) );
  INV_X1 U19163 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U19164 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n12840), .B1(n16037), 
        .B2(n16036), .ZN(n16040) );
  INV_X1 U19165 ( .A(n16042), .ZN(n16044) );
  AOI21_X1 U19166 ( .B1(n16044), .B2(n20094), .A(n16043), .ZN(n16049) );
  NOR2_X1 U19167 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16045), .ZN(
        n16051) );
  OAI22_X1 U19168 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16047), .B1(
        n16051), .B2(n16046), .ZN(n16048) );
  OAI211_X1 U19169 ( .C1(n16159), .C2(n16050), .A(n16049), .B(n16048), .ZN(
        P1_U3005) );
  AOI21_X1 U19170 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n12840), .A(n16051), 
        .ZN(n16056) );
  INV_X1 U19171 ( .A(n16052), .ZN(n16054) );
  AOI22_X1 U19172 ( .A1(n16054), .A2(n20094), .B1(n20093), .B2(n16053), .ZN(
        n16055) );
  OAI211_X1 U19173 ( .C1(n16058), .C2(n16057), .A(n16056), .B(n16055), .ZN(
        P1_U3006) );
  INV_X1 U19174 ( .A(n16059), .ZN(n16061) );
  AOI22_X1 U19175 ( .A1(n16061), .A2(n20094), .B1(n20093), .B2(n16060), .ZN(
        n16072) );
  NAND2_X1 U19176 ( .A1(n12840), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16071) );
  INV_X1 U19177 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16064) );
  NOR3_X1 U19178 ( .A1(n16062), .A2(n16079), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16073) );
  AOI22_X1 U19179 ( .A1(n16064), .A2(n16063), .B1(n16073), .B2(n16171), .ZN(
        n16065) );
  INV_X1 U19180 ( .A(n16065), .ZN(n16066) );
  OAI21_X1 U19181 ( .B1(n16074), .B2(n16066), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16070) );
  NAND3_X1 U19182 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16068), .A3(
        n16067), .ZN(n16069) );
  NAND4_X1 U19183 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        P1_U3007) );
  AOI22_X1 U19184 ( .A1(n12840), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n16092), 
        .B2(n16073), .ZN(n16077) );
  AOI22_X1 U19185 ( .A1(n16075), .A2(n20094), .B1(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16074), .ZN(n16076) );
  OAI211_X1 U19186 ( .C1(n16159), .C2(n16078), .A(n16077), .B(n16076), .ZN(
        P1_U3008) );
  OAI21_X1 U19187 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16079), .ZN(n16087) );
  OAI222_X1 U19188 ( .A1(n16083), .A2(n16204), .B1(n16159), .B2(n16082), .C1(
        n16081), .C2(n16080), .ZN(n16084) );
  INV_X1 U19189 ( .A(n16084), .ZN(n16086) );
  NAND2_X1 U19190 ( .A1(n12840), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16085) );
  OAI211_X1 U19191 ( .C1(n16088), .C2(n16087), .A(n16086), .B(n16085), .ZN(
        P1_U3009) );
  AOI22_X1 U19192 ( .A1(n16090), .A2(n20094), .B1(n20093), .B2(n16089), .ZN(
        n16095) );
  AOI22_X1 U19193 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16093), .B1(
        n16092), .B2(n16091), .ZN(n16094) );
  OAI211_X1 U19194 ( .C1(n20818), .C2(n20101), .A(n16095), .B(n16094), .ZN(
        P1_U3012) );
  OAI22_X1 U19195 ( .A1(n16097), .A2(n16204), .B1(n16159), .B2(n16096), .ZN(
        n16098) );
  AOI21_X1 U19196 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16099), .A(
        n16098), .ZN(n16104) );
  NAND3_X1 U19197 ( .A1(n16102), .A2(n16101), .A3(n16100), .ZN(n16103) );
  OAI211_X1 U19198 ( .C1(n15874), .C2(n20101), .A(n16104), .B(n16103), .ZN(
        P1_U3013) );
  INV_X1 U19199 ( .A(n16105), .ZN(n16110) );
  NOR3_X1 U19200 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16115), .A3(
        n16106), .ZN(n16109) );
  INV_X1 U19201 ( .A(n16128), .ZN(n16137) );
  AOI21_X1 U19202 ( .B1(n12819), .B2(n16177), .A(n16137), .ZN(n16114) );
  OR2_X1 U19203 ( .A1(n16106), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16120) );
  AOI21_X1 U19204 ( .B1(n16114), .B2(n16120), .A(n16107), .ZN(n16108) );
  AOI211_X1 U19205 ( .C1(n16110), .C2(n20094), .A(n16109), .B(n16108), .ZN(
        n16112) );
  NAND2_X1 U19206 ( .A1(n12840), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16111) );
  OAI211_X1 U19207 ( .C1(n16159), .C2(n16113), .A(n16112), .B(n16111), .ZN(
        P1_U3015) );
  NOR2_X1 U19208 ( .A1(n20101), .A2(n20812), .ZN(n16118) );
  OAI22_X1 U19209 ( .A1(n16116), .A2(n16204), .B1(n16115), .B2(n16114), .ZN(
        n16117) );
  AOI211_X1 U19210 ( .C1(n20093), .C2(n16119), .A(n16118), .B(n16117), .ZN(
        n16121) );
  NAND2_X1 U19211 ( .A1(n16121), .A2(n16120), .ZN(P1_U3016) );
  INV_X1 U19212 ( .A(n16122), .ZN(n16130) );
  OR2_X1 U19213 ( .A1(n16124), .A2(n16123), .ZN(n16151) );
  OR2_X1 U19214 ( .A1(n16151), .A2(n16125), .ZN(n16164) );
  NOR2_X1 U19215 ( .A1(n16152), .A2(n16164), .ZN(n16143) );
  NAND4_X1 U19216 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n16143), .A4(n12819), .ZN(
        n16126) );
  OAI22_X1 U19217 ( .A1(n16128), .A2(n12819), .B1(n16127), .B2(n16126), .ZN(
        n16129) );
  AOI21_X1 U19218 ( .B1(n16130), .B2(n20094), .A(n16129), .ZN(n16132) );
  NAND2_X1 U19219 ( .A1(n12840), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16131) );
  OAI211_X1 U19220 ( .C1(n16159), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        P1_U3017) );
  AOI21_X1 U19221 ( .B1(n20098), .B2(n16135), .A(n16134), .ZN(n16141) );
  AOI22_X1 U19222 ( .A1(n12840), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n20093), 
        .B2(n16136), .ZN(n16140) );
  AOI22_X1 U19223 ( .A1(n16138), .A2(n20094), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16137), .ZN(n16139) );
  OAI211_X1 U19224 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16141), .A(
        n16140), .B(n16139), .ZN(P1_U3018) );
  AOI22_X1 U19225 ( .A1(n12840), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20093), 
        .B2(n16142), .ZN(n16146) );
  AOI22_X1 U19226 ( .A1(n16144), .A2(n20094), .B1(n16147), .B2(n16143), .ZN(
        n16145) );
  OAI211_X1 U19227 ( .C1(n16148), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P1_U3020) );
  INV_X1 U19228 ( .A(n16149), .ZN(n16155) );
  OAI21_X1 U19229 ( .B1(n16151), .B2(n16172), .A(n16150), .ZN(n16169) );
  OAI21_X1 U19230 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16152), .ZN(n16153) );
  OAI22_X1 U19231 ( .A1(n12823), .A2(n16169), .B1(n16164), .B2(n16153), .ZN(
        n16154) );
  AOI21_X1 U19232 ( .B1(n16155), .B2(n20094), .A(n16154), .ZN(n16157) );
  NAND2_X1 U19233 ( .A1(n12840), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16156) );
  OAI211_X1 U19234 ( .C1(n16159), .C2(n16158), .A(n16157), .B(n16156), .ZN(
        P1_U3021) );
  INV_X1 U19235 ( .A(n16160), .ZN(n16161) );
  AOI21_X1 U19236 ( .B1(n16163), .B2(n16162), .A(n16161), .ZN(n20006) );
  NOR2_X1 U19237 ( .A1(n20101), .A2(n13771), .ZN(n16167) );
  OAI22_X1 U19238 ( .A1(n16165), .A2(n16204), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16164), .ZN(n16166) );
  AOI211_X1 U19239 ( .C1(n20093), .C2(n20006), .A(n16167), .B(n16166), .ZN(
        n16168) );
  OAI21_X1 U19240 ( .B1(n16170), .B2(n16169), .A(n16168), .ZN(P1_U3022) );
  INV_X1 U19241 ( .A(n16171), .ZN(n16176) );
  OR2_X1 U19242 ( .A1(n16174), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16211) );
  AOI211_X1 U19243 ( .C1(n16175), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        n16206) );
  OAI21_X1 U19244 ( .B1(n16176), .B2(n16211), .A(n16206), .ZN(n16196) );
  AOI21_X1 U19245 ( .B1(n16180), .B2(n16177), .A(n16196), .ZN(n16195) );
  INV_X1 U19246 ( .A(n16178), .ZN(n16179) );
  AOI222_X1 U19247 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n12840), .B1(n20093), 
        .B2(n19951), .C1(n20094), .C2(n16179), .ZN(n16182) );
  NOR2_X1 U19248 ( .A1(n16180), .A2(n16200), .ZN(n16190) );
  OAI221_X1 U19249 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16183), .C2(n16194), .A(
        n16190), .ZN(n16181) );
  OAI211_X1 U19250 ( .C1(n16195), .C2(n16183), .A(n16182), .B(n16181), .ZN(
        P1_U3023) );
  INV_X1 U19251 ( .A(n16184), .ZN(n16187) );
  AOI21_X1 U19252 ( .B1(n16187), .B2(n16186), .A(n16185), .ZN(n16189) );
  AOI22_X1 U19253 ( .A1(n12840), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20093), 
        .B2(n9704), .ZN(n16193) );
  AOI22_X1 U19254 ( .A1(n16191), .A2(n20094), .B1(n16194), .B2(n16190), .ZN(
        n16192) );
  OAI211_X1 U19255 ( .C1(n16195), .C2(n16194), .A(n16193), .B(n16192), .ZN(
        P1_U3024) );
  AOI22_X1 U19256 ( .A1(n12840), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20093), 
        .B2(n19978), .ZN(n16199) );
  AOI22_X1 U19257 ( .A1(n16197), .A2(n20094), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16196), .ZN(n16198) );
  OAI211_X1 U19258 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16200), .A(
        n16199), .B(n16198), .ZN(P1_U3025) );
  INV_X1 U19259 ( .A(n16201), .ZN(n16212) );
  INV_X1 U19260 ( .A(n16202), .ZN(n16208) );
  OAI22_X1 U19261 ( .A1(n16206), .A2(n16205), .B1(n16204), .B2(n16203), .ZN(
        n16207) );
  AOI211_X1 U19262 ( .C1(n20093), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        n16210) );
  OAI21_X1 U19263 ( .B1(n16212), .B2(n16211), .A(n16210), .ZN(P1_U3026) );
  NAND3_X1 U19264 ( .A1(n16215), .A2(n16214), .A3(n16213), .ZN(n16218) );
  OAI22_X1 U19265 ( .A1(n16219), .A2(n16218), .B1(n16217), .B2(n16216), .ZN(
        P1_U3468) );
  NAND4_X1 U19266 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20856), .A4(n20864), .ZN(n16220) );
  AND2_X1 U19267 ( .A1(n16221), .A2(n16220), .ZN(n20778) );
  AOI21_X1 U19268 ( .B1(n20778), .B2(n16223), .A(n16222), .ZN(n16226) );
  OAI221_X1 U19269 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16229), 
        .A(n16224), .ZN(n16225) );
  AOI211_X1 U19270 ( .C1(n16227), .C2(n20781), .A(n16226), .B(n16225), .ZN(
        P1_U3162) );
  OAI221_X1 U19271 ( .B1(n20566), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20566), 
        .C2(n16229), .A(n16228), .ZN(P1_U3466) );
  AOI211_X1 U19272 ( .C1(n16232), .C2(n16231), .A(n16230), .B(n19782), .ZN(
        n16235) );
  INV_X1 U19273 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16233) );
  OAI22_X1 U19274 ( .A1(n16233), .A2(n19084), .B1(n19853), .B2(n19096), .ZN(
        n16234) );
  AOI211_X1 U19275 ( .C1(P2_EBX_REG_29__SCAN_IN), .C2(n19110), .A(n16235), .B(
        n16234), .ZN(n16239) );
  AOI22_X1 U19276 ( .A1(n16237), .A2(n19122), .B1(n19086), .B2(n16236), .ZN(
        n16238) );
  OAI211_X1 U19277 ( .C1(n16240), .C2(n19127), .A(n16239), .B(n16238), .ZN(
        P2_U2826) );
  AOI22_X1 U19278 ( .A1(n19159), .A2(n14130), .B1(n11561), .B2(n19153), .ZN(
        P2_U2856) );
  INV_X1 U19279 ( .A(n16241), .ZN(n16242) );
  AOI22_X1 U19280 ( .A1(n16243), .A2(n19156), .B1(n19159), .B2(n16242), .ZN(
        n16244) );
  OAI21_X1 U19281 ( .B1(n19159), .B2(n11250), .A(n16244), .ZN(P2_U2864) );
  AOI21_X1 U19282 ( .B1(n16246), .B2(n14877), .A(n16245), .ZN(n16261) );
  AOI22_X1 U19283 ( .A1(n16261), .A2(n19156), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19153), .ZN(n16247) );
  OAI21_X1 U19284 ( .B1(n19153), .B2(n16248), .A(n16247), .ZN(P2_U2865) );
  NOR2_X1 U19285 ( .A1(n14883), .A2(n16249), .ZN(n16250) );
  OR2_X1 U19286 ( .A1(n14876), .A2(n16250), .ZN(n16266) );
  INV_X1 U19287 ( .A(n18972), .ZN(n16251) );
  OAI22_X1 U19288 ( .A1(n16266), .A2(n19148), .B1(n16251), .B2(n19153), .ZN(
        n16252) );
  INV_X1 U19289 ( .A(n16252), .ZN(n16253) );
  OAI21_X1 U19290 ( .B1(n19159), .B2(n11240), .A(n16253), .ZN(P2_U2867) );
  AND2_X1 U19291 ( .A1(n14897), .A2(n16254), .ZN(n16255) );
  OR2_X1 U19292 ( .A1(n16255), .A2(n14882), .ZN(n16273) );
  OAI22_X1 U19293 ( .A1(n16273), .A2(n19148), .B1(n19159), .B2(n16256), .ZN(
        n16257) );
  INV_X1 U19294 ( .A(n16257), .ZN(n16258) );
  OAI21_X1 U19295 ( .B1(n19153), .B2(n18995), .A(n16258), .ZN(P2_U2869) );
  AOI22_X1 U19296 ( .A1(n19164), .A2(n16259), .B1(n19213), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16264) );
  AOI22_X1 U19297 ( .A1(n19166), .A2(BUF1_REG_22__SCAN_IN), .B1(n19165), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16263) );
  AOI22_X1 U19298 ( .A1(n16261), .A2(n19168), .B1(n19214), .B2(n16260), .ZN(
        n16262) );
  NAND3_X1 U19299 ( .A1(n16264), .A2(n16263), .A3(n16262), .ZN(P2_U2897) );
  AOI22_X1 U19300 ( .A1(n19164), .A2(n16265), .B1(n19213), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16270) );
  AOI22_X1 U19301 ( .A1(n19166), .A2(BUF1_REG_20__SCAN_IN), .B1(n19165), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16269) );
  OAI22_X1 U19302 ( .A1(n16266), .A2(n19218), .B1(n19173), .B2(n18970), .ZN(
        n16267) );
  INV_X1 U19303 ( .A(n16267), .ZN(n16268) );
  NAND3_X1 U19304 ( .A1(n16270), .A2(n16269), .A3(n16268), .ZN(P2_U2899) );
  AOI22_X1 U19305 ( .A1(n19164), .A2(n16271), .B1(n19213), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16277) );
  AOI22_X1 U19306 ( .A1(n19166), .A2(BUF1_REG_18__SCAN_IN), .B1(n19165), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16276) );
  INV_X1 U19307 ( .A(n16272), .ZN(n18994) );
  OAI22_X1 U19308 ( .A1(n16273), .A2(n19218), .B1(n19173), .B2(n18994), .ZN(
        n16274) );
  INV_X1 U19309 ( .A(n16274), .ZN(n16275) );
  NAND3_X1 U19310 ( .A1(n16277), .A2(n16276), .A3(n16275), .ZN(P2_U2901) );
  AOI22_X1 U19311 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19115), .ZN(n16281) );
  AOI222_X1 U19312 ( .A1(n16279), .A2(n16293), .B1(n16311), .B2(n19066), .C1(
        n11517), .C2(n16278), .ZN(n16280) );
  OAI211_X1 U19313 ( .C1(n16304), .C2(n19064), .A(n16281), .B(n16280), .ZN(
        P2_U3004) );
  AOI22_X1 U19314 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19115), .ZN(n16295) );
  NOR2_X1 U19315 ( .A1(n16283), .A2(n16282), .ZN(n16287) );
  NOR2_X1 U19316 ( .A1(n16285), .A2(n16284), .ZN(n16286) );
  XNOR2_X1 U19317 ( .A(n16287), .B(n16286), .ZN(n16321) );
  INV_X1 U19318 ( .A(n19154), .ZN(n16320) );
  NAND2_X1 U19319 ( .A1(n16288), .A2(n16325), .ZN(n16289) );
  NAND2_X1 U19320 ( .A1(n16290), .A2(n16289), .ZN(n16291) );
  XOR2_X1 U19321 ( .A(n16292), .B(n16291), .Z(n16318) );
  AOI222_X1 U19322 ( .A1(n16321), .A2(n16293), .B1(n16311), .B2(n16320), .C1(
        n11517), .C2(n16318), .ZN(n16294) );
  OAI211_X1 U19323 ( .C1(n16304), .C2(n16296), .A(n16295), .B(n16294), .ZN(
        P2_U3006) );
  AOI22_X1 U19324 ( .A1(n16297), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19115), .ZN(n16303) );
  OAI222_X1 U19325 ( .A1(n16300), .A2(n13376), .B1(n16299), .B2(n16308), .C1(
        n16306), .C2(n16298), .ZN(n16301) );
  INV_X1 U19326 ( .A(n16301), .ZN(n16302) );
  OAI211_X1 U19327 ( .C1(n16304), .C2(n19103), .A(n16303), .B(n16302), .ZN(
        P2_U3008) );
  AOI22_X1 U19328 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19115), .B1(n16305), 
        .B2(n19120), .ZN(n16313) );
  OAI22_X1 U19329 ( .A1(n16309), .A2(n16308), .B1(n16307), .B2(n16306), .ZN(
        n16310) );
  AOI21_X1 U19330 ( .B1(n16311), .B2(n19121), .A(n16310), .ZN(n16312) );
  OAI211_X1 U19331 ( .C1(n16315), .C2(n16314), .A(n16313), .B(n16312), .ZN(
        P2_U3009) );
  OAI22_X1 U19332 ( .A1(n16316), .A2(n16324), .B1(n16331), .B2(n19194), .ZN(
        n16317) );
  INV_X1 U19333 ( .A(n16317), .ZN(n16329) );
  AOI222_X1 U19334 ( .A1(n16321), .A2(n16338), .B1(n16333), .B2(n16320), .C1(
        n16319), .C2(n16318), .ZN(n16328) );
  NAND2_X1 U19335 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16322), .ZN(n16327) );
  OAI221_X1 U19336 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n16325), .C2(n16324), .A(
        n16323), .ZN(n16326) );
  NAND4_X1 U19337 ( .A1(n16329), .A2(n16328), .A3(n16327), .A4(n16326), .ZN(
        P2_U3038) );
  OAI21_X1 U19338 ( .B1(n19206), .B2(n16331), .A(n16330), .ZN(n16332) );
  AOI21_X1 U19339 ( .B1(n13164), .B2(n16333), .A(n16332), .ZN(n16334) );
  OAI21_X1 U19340 ( .B1(n16335), .B2(n19264), .A(n16334), .ZN(n16336) );
  AOI21_X1 U19341 ( .B1(n16338), .B2(n16337), .A(n16336), .ZN(n16339) );
  OAI221_X1 U19342 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16342), .C1(
        n16341), .C2(n16340), .A(n16339), .ZN(P2_U3043) );
  INV_X1 U19343 ( .A(n16343), .ZN(n16348) );
  OAI21_X1 U19344 ( .B1(n16345), .B2(n19891), .A(n16376), .ZN(n16347) );
  AOI211_X1 U19345 ( .C1(n16345), .C2(n19891), .A(n19900), .B(n16344), .ZN(
        n16346) );
  AOI211_X1 U19346 ( .C1(n16348), .C2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16347), .B(n16346), .ZN(n16354) );
  MUX2_X1 U19347 ( .A(n10430), .B(n16348), .S(n16376), .Z(n16355) );
  INV_X1 U19348 ( .A(n16376), .ZN(n16351) );
  NAND2_X1 U19349 ( .A1(n16351), .A2(n16349), .ZN(n16350) );
  OAI21_X1 U19350 ( .B1(n16353), .B2(n16351), .A(n16350), .ZN(n16356) );
  OAI21_X1 U19351 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16355), .A(
        n16356), .ZN(n16352) );
  AOI222_X1 U19352 ( .A1(n16354), .A2(n19874), .B1(n16354), .B2(n16353), .C1(
        n19874), .C2(n16352), .ZN(n16357) );
  OAI22_X1 U19353 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16357), .B1(
        n16356), .B2(n16355), .ZN(n16378) );
  NAND2_X1 U19354 ( .A1(n16367), .A2(n16358), .ZN(n16365) );
  INV_X1 U19355 ( .A(n16359), .ZN(n16361) );
  OAI22_X1 U19356 ( .A1(n16362), .A2(n16361), .B1(n9594), .B2(n16360), .ZN(
        n16363) );
  INV_X1 U19357 ( .A(n16363), .ZN(n16364) );
  OAI211_X1 U19358 ( .C1(n16367), .C2(n16366), .A(n16365), .B(n16364), .ZN(
        n19903) );
  NOR2_X1 U19359 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16372) );
  NOR2_X1 U19360 ( .A1(n16368), .A2(n19905), .ZN(n16369) );
  OAI211_X1 U19361 ( .C1(n16372), .C2(n16371), .A(n16370), .B(n16369), .ZN(
        n16373) );
  NOR2_X1 U19362 ( .A1(n19903), .A2(n16373), .ZN(n16374) );
  OAI21_X1 U19363 ( .B1(n16376), .B2(n16375), .A(n16374), .ZN(n16377) );
  NOR2_X1 U19364 ( .A1(n16378), .A2(n16377), .ZN(n16389) );
  AOI21_X1 U19365 ( .B1(n16389), .B2(n16384), .A(n21039), .ZN(n16383) );
  NAND3_X1 U19366 ( .A1(n16380), .A2(n10747), .A3(n16379), .ZN(n16382) );
  NOR2_X1 U19367 ( .A1(n16381), .A2(n19676), .ZN(n21036) );
  NAND2_X1 U19368 ( .A1(n16382), .A2(n21036), .ZN(n16385) );
  NOR2_X1 U19369 ( .A1(n16383), .A2(n16385), .ZN(n19784) );
  NOR2_X1 U19370 ( .A1(n19784), .A2(n21039), .ZN(n16395) );
  NAND2_X1 U19371 ( .A1(n19676), .A2(n16384), .ZN(n16386) );
  OAI22_X1 U19372 ( .A1(n16387), .A2(n16386), .B1(n21038), .B2(n16385), .ZN(
        n16393) );
  NAND2_X1 U19373 ( .A1(n19676), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18936) );
  INV_X1 U19374 ( .A(n18936), .ZN(n19780) );
  OAI22_X1 U19375 ( .A1(n16389), .A2(n16388), .B1(n19904), .B2(n16394), .ZN(
        n16390) );
  AOI211_X1 U19376 ( .C1(n19786), .C2(n19780), .A(n16391), .B(n16390), .ZN(
        n16392) );
  OAI221_X1 U19377 ( .B1(n16395), .B2(n21039), .C1(n16395), .C2(n16393), .A(
        n16392), .ZN(P2_U3176) );
  OAI21_X1 U19378 ( .B1(n16395), .B2(n19678), .A(n16394), .ZN(P2_U3593) );
  INV_X1 U19379 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16607) );
  XNOR2_X1 U19380 ( .A(n16607), .B(n16410), .ZN(n16606) );
  OAI221_X1 U19381 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16398), .C1(
        n16607), .C2(n16397), .A(n16396), .ZN(n16399) );
  AOI21_X1 U19382 ( .B1(n17758), .B2(n16606), .A(n16399), .ZN(n16404) );
  OAI22_X1 U19383 ( .A1(n16406), .A2(n17926), .B1(n16420), .B2(n17837), .ZN(
        n16402) );
  INV_X1 U19384 ( .A(n17578), .ZN(n16401) );
  AOI22_X1 U19385 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16402), .B1(
        n16401), .B2(n16400), .ZN(n16403) );
  OAI211_X1 U19386 ( .C1(n16405), .C2(n17807), .A(n16404), .B(n16403), .ZN(
        P3_U2800) );
  NOR2_X1 U19387 ( .A1(n16406), .A2(n17926), .ZN(n16417) );
  NOR2_X1 U19388 ( .A1(n16407), .A2(n16419), .ZN(n16442) );
  AOI22_X1 U19389 ( .A1(n9587), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16408), .ZN(n16413) );
  INV_X1 U19390 ( .A(n16409), .ZN(n16582) );
  AOI21_X1 U19391 ( .B1(n16617), .B2(n16582), .A(n16410), .ZN(n16616) );
  OAI21_X1 U19392 ( .B1(n16411), .B2(n17758), .A(n16616), .ZN(n16412) );
  OAI211_X1 U19393 ( .C1(n16415), .C2(n16414), .A(n16413), .B(n16412), .ZN(
        n16416) );
  AOI221_X1 U19394 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16417), 
        .C1(n16442), .C2(n16417), .A(n16416), .ZN(n16423) );
  NOR2_X1 U19395 ( .A1(n16419), .A2(n16418), .ZN(n16440) );
  NOR2_X1 U19396 ( .A1(n16420), .A2(n17837), .ZN(n16421) );
  OAI21_X1 U19397 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16440), .A(
        n16421), .ZN(n16422) );
  OAI211_X1 U19398 ( .C1(n16424), .C2(n17807), .A(n16423), .B(n16422), .ZN(
        P3_U2801) );
  NAND2_X1 U19399 ( .A1(n9587), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17566) );
  NOR2_X1 U19400 ( .A1(n18700), .A2(n16439), .ZN(n18101) );
  OAI22_X1 U19401 ( .A1(n18123), .A2(n18104), .B1(n17792), .B2(n18125), .ZN(
        n18031) );
  INV_X1 U19402 ( .A(n18052), .ZN(n16425) );
  OAI22_X1 U19403 ( .A1(n18736), .A2(n16425), .B1(n18097), .B2(n18220), .ZN(
        n16426) );
  OAI21_X1 U19404 ( .B1(n18031), .B2(n16426), .A(n17691), .ZN(n18000) );
  NOR2_X1 U19405 ( .A1(n16427), .A2(n18000), .ZN(n17978) );
  NAND2_X1 U19406 ( .A1(n16428), .A2(n17978), .ZN(n17927) );
  INV_X1 U19407 ( .A(n17927), .ZN(n16431) );
  INV_X1 U19408 ( .A(n18252), .ZN(n18246) );
  NOR3_X1 U19409 ( .A1(n17729), .A2(n16429), .A3(n18246), .ZN(n16430) );
  OAI211_X1 U19410 ( .C1(n16431), .C2(n16430), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17562), .ZN(n16447) );
  NOR2_X1 U19411 ( .A1(n16433), .A2(n16432), .ZN(n17574) );
  OR3_X1 U19412 ( .A1(n18144), .A2(n16434), .A3(n17574), .ZN(n16446) );
  OAI21_X1 U19413 ( .B1(n16435), .B2(n17729), .A(n16434), .ZN(n17573) );
  OAI21_X1 U19414 ( .B1(n16437), .B2(n16436), .A(n17572), .ZN(n16438) );
  AOI221_X1 U19415 ( .B1(n17427), .B2(n16440), .C1(n16439), .C2(n16438), .A(
        n18700), .ZN(n16444) );
  OAI211_X1 U19416 ( .C1(n16442), .C2(n18104), .A(n16441), .B(n18239), .ZN(
        n16443) );
  OAI211_X1 U19417 ( .C1(n16444), .C2(n16443), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18253), .ZN(n16445) );
  NAND4_X1 U19418 ( .A1(n17566), .A2(n16447), .A3(n16446), .A4(n16445), .ZN(
        P3_U2834) );
  NOR3_X1 U19419 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16449) );
  NOR4_X1 U19420 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16448) );
  NAND4_X1 U19421 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16449), .A3(n16448), .A4(
        U215), .ZN(U213) );
  INV_X1 U19422 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16543) );
  INV_X2 U19423 ( .A(U214), .ZN(n16507) );
  NOR2_X1 U19424 ( .A1(n16507), .A2(n16450), .ZN(n16494) );
  INV_X1 U19425 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16544) );
  OAI222_X1 U19426 ( .A1(U212), .A2(n16543), .B1(n16509), .B2(n16451), .C1(
        U214), .C2(n16544), .ZN(U216) );
  INV_X1 U19427 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16453) );
  INV_X2 U19428 ( .A(U212), .ZN(n16500) );
  AOI22_X1 U19429 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16500), .ZN(n16452) );
  OAI21_X1 U19430 ( .B1(n16453), .B2(n16509), .A(n16452), .ZN(U217) );
  INV_X1 U19431 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U19432 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16500), .ZN(n16454) );
  OAI21_X1 U19433 ( .B1(n16455), .B2(n16509), .A(n16454), .ZN(U218) );
  INV_X1 U19434 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16457) );
  AOI22_X1 U19435 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16500), .ZN(n16456) );
  OAI21_X1 U19436 ( .B1(n16457), .B2(n16509), .A(n16456), .ZN(U219) );
  AOI22_X1 U19437 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16500), .ZN(n16458) );
  OAI21_X1 U19438 ( .B1(n16459), .B2(n16509), .A(n16458), .ZN(U220) );
  AOI222_X1 U19439 ( .A1(n16500), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(n16494), 
        .B2(BUF1_REG_26__SCAN_IN), .C1(n16507), .C2(P1_DATAO_REG_26__SCAN_IN), 
        .ZN(n16460) );
  INV_X1 U19440 ( .A(n16460), .ZN(U221) );
  AOI22_X1 U19441 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16500), .ZN(n16461) );
  OAI21_X1 U19442 ( .B1(n14954), .B2(n16509), .A(n16461), .ZN(U222) );
  INV_X1 U19443 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16463) );
  AOI22_X1 U19444 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16500), .ZN(n16462) );
  OAI21_X1 U19445 ( .B1(n16463), .B2(n16509), .A(n16462), .ZN(U223) );
  AOI22_X1 U19446 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16500), .ZN(n16464) );
  OAI21_X1 U19447 ( .B1(n16465), .B2(n16509), .A(n16464), .ZN(U224) );
  INV_X1 U19448 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19449 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16500), .ZN(n16466) );
  OAI21_X1 U19450 ( .B1(n16467), .B2(n16509), .A(n16466), .ZN(U225) );
  INV_X1 U19451 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19452 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16500), .ZN(n16468) );
  OAI21_X1 U19453 ( .B1(n16469), .B2(n16509), .A(n16468), .ZN(U226) );
  AOI22_X1 U19454 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16500), .ZN(n16470) );
  OAI21_X1 U19455 ( .B1(n16471), .B2(n16509), .A(n16470), .ZN(U227) );
  INV_X1 U19456 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16473) );
  AOI22_X1 U19457 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16500), .ZN(n16472) );
  OAI21_X1 U19458 ( .B1(n16473), .B2(n16509), .A(n16472), .ZN(U228) );
  INV_X1 U19459 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19460 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16500), .ZN(n16474) );
  OAI21_X1 U19461 ( .B1(n16475), .B2(n16509), .A(n16474), .ZN(U229) );
  INV_X1 U19462 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16477) );
  AOI22_X1 U19463 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16500), .ZN(n16476) );
  OAI21_X1 U19464 ( .B1(n16477), .B2(n16509), .A(n16476), .ZN(U230) );
  INV_X1 U19465 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U19466 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16500), .ZN(n16478) );
  OAI21_X1 U19467 ( .B1(n16479), .B2(n16509), .A(n16478), .ZN(U231) );
  AOI22_X1 U19468 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16500), .ZN(n16480) );
  OAI21_X1 U19469 ( .B1(n13328), .B2(n16509), .A(n16480), .ZN(U232) );
  INV_X1 U19470 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19471 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16500), .ZN(n16481) );
  OAI21_X1 U19472 ( .B1(n16482), .B2(n16509), .A(n16481), .ZN(U233) );
  AOI22_X1 U19473 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16500), .ZN(n16483) );
  OAI21_X1 U19474 ( .B1(n13012), .B2(n16509), .A(n16483), .ZN(U234) );
  AOI22_X1 U19475 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16500), .ZN(n16484) );
  OAI21_X1 U19476 ( .B1(n13032), .B2(n16509), .A(n16484), .ZN(U235) );
  AOI22_X1 U19477 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16500), .ZN(n16485) );
  OAI21_X1 U19478 ( .B1(n13023), .B2(n16509), .A(n16485), .ZN(U236) );
  INV_X1 U19479 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16487) );
  AOI22_X1 U19480 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16500), .ZN(n16486) );
  OAI21_X1 U19481 ( .B1(n16487), .B2(n16509), .A(n16486), .ZN(U237) );
  INV_X1 U19482 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19483 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16500), .ZN(n16488) );
  OAI21_X1 U19484 ( .B1(n16489), .B2(n16509), .A(n16488), .ZN(U238) );
  AOI22_X1 U19485 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16500), .ZN(n16490) );
  OAI21_X1 U19486 ( .B1(n16491), .B2(n16509), .A(n16490), .ZN(U239) );
  INV_X1 U19487 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16493) );
  AOI22_X1 U19488 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16500), .ZN(n16492) );
  OAI21_X1 U19489 ( .B1(n16493), .B2(n16509), .A(n16492), .ZN(U240) );
  AOI222_X1 U19490 ( .A1(n16500), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n16494), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n16507), .C2(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n16495) );
  INV_X1 U19491 ( .A(n16495), .ZN(U241) );
  AOI22_X1 U19492 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16500), .ZN(n16496) );
  OAI21_X1 U19493 ( .B1(n16497), .B2(n16509), .A(n16496), .ZN(U242) );
  INV_X1 U19494 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16499) );
  AOI22_X1 U19495 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16500), .ZN(n16498) );
  OAI21_X1 U19496 ( .B1(n16499), .B2(n16509), .A(n16498), .ZN(U243) );
  INV_X1 U19497 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16502) );
  AOI22_X1 U19498 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16500), .ZN(n16501) );
  OAI21_X1 U19499 ( .B1(n16502), .B2(n16509), .A(n16501), .ZN(U244) );
  INV_X1 U19500 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19501 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16500), .ZN(n16503) );
  OAI21_X1 U19502 ( .B1(n16504), .B2(n16509), .A(n16503), .ZN(U245) );
  INV_X1 U19503 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16506) );
  AOI22_X1 U19504 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16500), .ZN(n16505) );
  OAI21_X1 U19505 ( .B1(n16506), .B2(n16509), .A(n16505), .ZN(U246) );
  INV_X1 U19506 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16510) );
  AOI22_X1 U19507 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16507), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16500), .ZN(n16508) );
  OAI21_X1 U19508 ( .B1(n16510), .B2(n16509), .A(n16508), .ZN(U247) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16541), .ZN(n16511) );
  INV_X1 U19510 ( .A(n16511), .ZN(U251) );
  OAI22_X1 U19511 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16541), .ZN(n16512) );
  INV_X1 U19512 ( .A(n16512), .ZN(U252) );
  OAI22_X1 U19513 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16541), .ZN(n16513) );
  INV_X1 U19514 ( .A(n16513), .ZN(U253) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16541), .ZN(n16514) );
  INV_X1 U19516 ( .A(n16514), .ZN(U254) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16541), .ZN(n16515) );
  INV_X1 U19518 ( .A(n16515), .ZN(U255) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16541), .ZN(n16516) );
  INV_X1 U19520 ( .A(n16516), .ZN(U256) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n20934) );
  INV_X1 U19522 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U19523 ( .A1(n16541), .A2(n20934), .B1(n18296), .B2(U215), .ZN(U257) );
  OAI22_X1 U19524 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16541), .ZN(n16517) );
  INV_X1 U19525 ( .A(n16517), .ZN(U258) );
  OAI22_X1 U19526 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16541), .ZN(n16518) );
  INV_X1 U19527 ( .A(n16518), .ZN(U259) );
  OAI22_X1 U19528 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16541), .ZN(n16519) );
  INV_X1 U19529 ( .A(n16519), .ZN(U260) );
  OAI22_X1 U19530 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16533), .ZN(n16520) );
  INV_X1 U19531 ( .A(n16520), .ZN(U261) );
  OAI22_X1 U19532 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16533), .ZN(n16521) );
  INV_X1 U19533 ( .A(n16521), .ZN(U262) );
  OAI22_X1 U19534 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16541), .ZN(n16522) );
  INV_X1 U19535 ( .A(n16522), .ZN(U263) );
  OAI22_X1 U19536 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16533), .ZN(n16523) );
  INV_X1 U19537 ( .A(n16523), .ZN(U264) );
  OAI22_X1 U19538 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16541), .ZN(n16524) );
  INV_X1 U19539 ( .A(n16524), .ZN(U265) );
  OAI22_X1 U19540 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16541), .ZN(n16525) );
  INV_X1 U19541 ( .A(n16525), .ZN(U266) );
  OAI22_X1 U19542 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16533), .ZN(n16526) );
  INV_X1 U19543 ( .A(n16526), .ZN(U267) );
  OAI22_X1 U19544 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16533), .ZN(n16527) );
  INV_X1 U19545 ( .A(n16527), .ZN(U268) );
  OAI22_X1 U19546 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16533), .ZN(n16528) );
  INV_X1 U19547 ( .A(n16528), .ZN(U269) );
  OAI22_X1 U19548 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16533), .ZN(n16529) );
  INV_X1 U19549 ( .A(n16529), .ZN(U270) );
  OAI22_X1 U19550 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16533), .ZN(n16530) );
  INV_X1 U19551 ( .A(n16530), .ZN(U271) );
  OAI22_X1 U19552 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16533), .ZN(n16531) );
  INV_X1 U19553 ( .A(n16531), .ZN(U272) );
  OAI22_X1 U19554 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16541), .ZN(n16532) );
  INV_X1 U19555 ( .A(n16532), .ZN(U273) );
  OAI22_X1 U19556 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16533), .ZN(n16534) );
  INV_X1 U19557 ( .A(n16534), .ZN(U274) );
  OAI22_X1 U19558 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16541), .ZN(n16535) );
  INV_X1 U19559 ( .A(n16535), .ZN(U275) );
  OAI22_X1 U19560 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16541), .ZN(n16536) );
  INV_X1 U19561 ( .A(n16536), .ZN(U276) );
  INV_X1 U19562 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U19563 ( .A1(n16541), .A2(n20967), .B1(n14947), .B2(U215), .ZN(U277) );
  OAI22_X1 U19564 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16541), .ZN(n16537) );
  INV_X1 U19565 ( .A(n16537), .ZN(U278) );
  OAI22_X1 U19566 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16541), .ZN(n16538) );
  INV_X1 U19567 ( .A(n16538), .ZN(U279) );
  OAI22_X1 U19568 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16541), .ZN(n16539) );
  INV_X1 U19569 ( .A(n16539), .ZN(U280) );
  OAI22_X1 U19570 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16541), .ZN(n16540) );
  INV_X1 U19571 ( .A(n16540), .ZN(U281) );
  INV_X1 U19572 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U19573 ( .A1(n16541), .A2(n16543), .B1(n18303), .B2(U215), .ZN(U282) );
  INV_X1 U19574 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16542) );
  AOI222_X1 U19575 ( .A1(n16544), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16543), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16542), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16545) );
  INV_X2 U19576 ( .A(n16547), .ZN(n16546) );
  INV_X1 U19577 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18808) );
  INV_X1 U19578 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19820) );
  AOI22_X1 U19579 ( .A1(n16546), .A2(n18808), .B1(n19820), .B2(n16547), .ZN(
        U347) );
  INV_X1 U19580 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18806) );
  INV_X1 U19581 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U19582 ( .A1(n16546), .A2(n18806), .B1(n19818), .B2(n16547), .ZN(
        U348) );
  INV_X1 U19583 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18803) );
  INV_X1 U19584 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19817) );
  AOI22_X1 U19585 ( .A1(n16546), .A2(n18803), .B1(n19817), .B2(n16547), .ZN(
        U349) );
  INV_X1 U19586 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18802) );
  INV_X1 U19587 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U19588 ( .A1(n16546), .A2(n18802), .B1(n19815), .B2(n16547), .ZN(
        U350) );
  INV_X1 U19589 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18800) );
  INV_X1 U19590 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19813) );
  AOI22_X1 U19591 ( .A1(n16546), .A2(n18800), .B1(n19813), .B2(n16547), .ZN(
        U351) );
  INV_X1 U19592 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18798) );
  INV_X1 U19593 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U19594 ( .A1(n16546), .A2(n18798), .B1(n19811), .B2(n16547), .ZN(
        U352) );
  INV_X1 U19595 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18796) );
  INV_X1 U19596 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19597 ( .A1(n16546), .A2(n18796), .B1(n19809), .B2(n16547), .ZN(
        U353) );
  INV_X1 U19598 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18794) );
  AOI22_X1 U19599 ( .A1(n16546), .A2(n18794), .B1(n19807), .B2(n16547), .ZN(
        U354) );
  INV_X1 U19600 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18848) );
  INV_X1 U19601 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19856) );
  AOI22_X1 U19602 ( .A1(n16546), .A2(n18848), .B1(n19856), .B2(n16547), .ZN(
        U355) );
  INV_X1 U19603 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18845) );
  INV_X1 U19604 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U19605 ( .A1(n16546), .A2(n18845), .B1(n19854), .B2(n16547), .ZN(
        U356) );
  INV_X1 U19606 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18842) );
  INV_X1 U19607 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U19608 ( .A1(n16546), .A2(n18842), .B1(n19852), .B2(n16547), .ZN(
        U357) );
  INV_X1 U19609 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18841) );
  INV_X1 U19610 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U19611 ( .A1(n16546), .A2(n18841), .B1(n19849), .B2(n16547), .ZN(
        U358) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18839) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19848) );
  AOI22_X1 U19614 ( .A1(n16546), .A2(n18839), .B1(n19848), .B2(n16547), .ZN(
        U359) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18837) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U19617 ( .A1(n16546), .A2(n18837), .B1(n19846), .B2(n16547), .ZN(
        U360) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18835) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U19620 ( .A1(n16546), .A2(n18835), .B1(n19844), .B2(n16547), .ZN(
        U361) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18832) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19842) );
  AOI22_X1 U19623 ( .A1(n16546), .A2(n18832), .B1(n19842), .B2(n16547), .ZN(
        U362) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18831) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19840) );
  AOI22_X1 U19626 ( .A1(n16546), .A2(n18831), .B1(n19840), .B2(n16547), .ZN(
        U363) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18828) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19838) );
  AOI22_X1 U19629 ( .A1(n16546), .A2(n18828), .B1(n19838), .B2(n16547), .ZN(
        U364) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18792) );
  INV_X1 U19631 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19805) );
  AOI22_X1 U19632 ( .A1(n16546), .A2(n18792), .B1(n19805), .B2(n16547), .ZN(
        U365) );
  INV_X1 U19633 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18827) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19836) );
  AOI22_X1 U19635 ( .A1(n16546), .A2(n18827), .B1(n19836), .B2(n16547), .ZN(
        U366) );
  INV_X1 U19636 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18824) );
  INV_X1 U19637 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19834) );
  AOI22_X1 U19638 ( .A1(n16546), .A2(n18824), .B1(n19834), .B2(n16547), .ZN(
        U367) );
  INV_X1 U19639 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18823) );
  INV_X1 U19640 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19832) );
  AOI22_X1 U19641 ( .A1(n16546), .A2(n18823), .B1(n19832), .B2(n16547), .ZN(
        U368) );
  INV_X1 U19642 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18821) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U19644 ( .A1(n16546), .A2(n18821), .B1(n19831), .B2(n16547), .ZN(
        U369) );
  INV_X1 U19645 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18820) );
  INV_X1 U19646 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U19647 ( .A1(n16546), .A2(n18820), .B1(n19829), .B2(n16547), .ZN(
        U370) );
  INV_X1 U19648 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18818) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19828) );
  AOI22_X1 U19650 ( .A1(n16546), .A2(n18818), .B1(n19828), .B2(n16547), .ZN(
        U371) );
  INV_X1 U19651 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18815) );
  INV_X1 U19652 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U19653 ( .A1(n16546), .A2(n18815), .B1(n19826), .B2(n16547), .ZN(
        U372) );
  INV_X1 U19654 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18814) );
  INV_X1 U19655 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U19656 ( .A1(n16546), .A2(n18814), .B1(n19825), .B2(n16547), .ZN(
        U373) );
  INV_X1 U19657 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18811) );
  INV_X1 U19658 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19824) );
  AOI22_X1 U19659 ( .A1(n16546), .A2(n18811), .B1(n19824), .B2(n16547), .ZN(
        U374) );
  INV_X1 U19660 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18810) );
  INV_X1 U19661 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19822) );
  AOI22_X1 U19662 ( .A1(n16546), .A2(n18810), .B1(n19822), .B2(n16547), .ZN(
        U375) );
  INV_X1 U19663 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18790) );
  INV_X1 U19664 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19803) );
  AOI22_X1 U19665 ( .A1(n16546), .A2(n18790), .B1(n19803), .B2(n16547), .ZN(
        U376) );
  INV_X1 U19666 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18789) );
  NAND2_X1 U19667 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18789), .ZN(n18776) );
  AOI22_X1 U19668 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18776), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18787), .ZN(n18858) );
  AOI21_X1 U19669 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18858), .ZN(n16548) );
  INV_X1 U19670 ( .A(n16548), .ZN(P3_U2633) );
  INV_X1 U19671 ( .A(n18763), .ZN(n18754) );
  OAI21_X1 U19672 ( .B1(n16556), .B2(n17458), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16549) );
  OAI21_X1 U19673 ( .B1(n16550), .B2(n18754), .A(n16549), .ZN(P3_U2634) );
  AOI21_X1 U19674 ( .B1(n18787), .B2(n18789), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16551) );
  AOI22_X1 U19675 ( .A1(n18925), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16551), 
        .B2(n18926), .ZN(P3_U2635) );
  NOR2_X1 U19676 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16552) );
  OAI21_X1 U19677 ( .B1(n16552), .B2(BS16), .A(n18858), .ZN(n18856) );
  OAI21_X1 U19678 ( .B1(n18858), .B2(n18916), .A(n18856), .ZN(P3_U2636) );
  INV_X1 U19679 ( .A(n16553), .ZN(n16554) );
  NOR3_X1 U19680 ( .A1(n16556), .A2(n16555), .A3(n16554), .ZN(n18746) );
  NOR2_X1 U19681 ( .A1(n18746), .A2(n18750), .ZN(n18905) );
  OAI21_X1 U19682 ( .B1(n18905), .B2(n16558), .A(n16557), .ZN(P3_U2637) );
  NOR4_X1 U19683 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16562) );
  NOR4_X1 U19684 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16561) );
  NOR4_X1 U19685 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16560) );
  NOR4_X1 U19686 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16559) );
  NAND4_X1 U19687 ( .A1(n16562), .A2(n16561), .A3(n16560), .A4(n16559), .ZN(
        n16568) );
  NOR4_X1 U19688 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16566) );
  AOI211_X1 U19689 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_11__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16565) );
  NOR4_X1 U19690 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16564) );
  NOR4_X1 U19691 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16563) );
  NAND4_X1 U19692 ( .A1(n16566), .A2(n16565), .A3(n16564), .A4(n16563), .ZN(
        n16567) );
  NOR2_X1 U19693 ( .A1(n16568), .A2(n16567), .ZN(n18899) );
  INV_X1 U19694 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16570) );
  NOR3_X1 U19695 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16571) );
  OAI21_X1 U19696 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16571), .A(n18899), .ZN(
        n16569) );
  OAI21_X1 U19697 ( .B1(n18899), .B2(n16570), .A(n16569), .ZN(P3_U2638) );
  INV_X1 U19698 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18895) );
  INV_X1 U19699 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18857) );
  AOI21_X1 U19700 ( .B1(n18895), .B2(n18857), .A(n16571), .ZN(n16573) );
  INV_X1 U19701 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16572) );
  INV_X1 U19702 ( .A(n18899), .ZN(n18902) );
  AOI22_X1 U19703 ( .A1(n18899), .A2(n16573), .B1(n16572), .B2(n18902), .ZN(
        P3_U2639) );
  NAND4_X1 U19704 ( .A1(n18753), .A2(n18859), .A3(n18916), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18767) );
  NAND2_X1 U19705 ( .A1(n18253), .A2(n18767), .ZN(n16758) );
  NOR3_X1 U19706 ( .A1(n16576), .A2(n16575), .A3(n16574), .ZN(n18703) );
  AOI211_X4 U19707 ( .C1(n18763), .C2(n18589), .A(n16758), .B(n18914), .ZN(
        n16961) );
  OAI211_X1 U19708 ( .C1(n18277), .C2(n16577), .A(n18918), .B(n18916), .ZN(
        n16578) );
  INV_X1 U19709 ( .A(n16578), .ZN(n18752) );
  AOI211_X4 U19710 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18277), .A(n18752), .B(
        n16581), .ZN(n16965) );
  INV_X1 U19711 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18849) );
  INV_X1 U19712 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18836) );
  INV_X1 U19713 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18833) );
  INV_X1 U19714 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18829) );
  INV_X1 U19715 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18825) );
  INV_X1 U19716 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20986) );
  INV_X1 U19717 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18812) );
  INV_X1 U19718 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18804) );
  INV_X1 U19719 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18799) );
  INV_X1 U19720 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18795) );
  NAND3_X1 U19721 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16909) );
  NOR2_X1 U19722 ( .A1(n18795), .A2(n16909), .ZN(n16888) );
  NAND2_X1 U19723 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16888), .ZN(n16864) );
  NOR2_X1 U19724 ( .A1(n18799), .A2(n16864), .ZN(n16867) );
  NAND2_X1 U19725 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16867), .ZN(n16853) );
  NOR2_X1 U19726 ( .A1(n18804), .A2(n16853), .ZN(n16816) );
  NAND4_X1 U19727 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16816), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16811) );
  NOR2_X1 U19728 ( .A1(n18812), .A2(n16811), .ZN(n16782) );
  NAND3_X1 U19729 ( .A1(n16782), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .ZN(n16781) );
  NAND2_X1 U19730 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16765) );
  NOR3_X1 U19731 ( .A1(n20986), .A2(n16781), .A3(n16765), .ZN(n16726) );
  NAND2_X1 U19732 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16726), .ZN(n16725) );
  NOR2_X1 U19733 ( .A1(n18825), .A2(n16725), .ZN(n16717) );
  NAND2_X1 U19734 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16717), .ZN(n16701) );
  NOR2_X1 U19735 ( .A1(n18829), .A2(n16701), .ZN(n16697) );
  NAND2_X1 U19736 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16697), .ZN(n16684) );
  NOR2_X1 U19737 ( .A1(n18833), .A2(n16684), .ZN(n16682) );
  NAND2_X1 U19738 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16682), .ZN(n16662) );
  NOR2_X1 U19739 ( .A1(n18836), .A2(n16662), .ZN(n16648) );
  NAND2_X1 U19740 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16648), .ZN(n16596) );
  NOR2_X1 U19741 ( .A1(n16959), .A2(n16596), .ZN(n16642) );
  NAND4_X1 U19742 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16642), .ZN(n16598) );
  NOR3_X1 U19743 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18849), .A3(n16598), 
        .ZN(n16579) );
  AOI21_X1 U19744 ( .B1(n16965), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16579), .ZN(
        n16602) );
  NAND2_X1 U19745 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18277), .ZN(n16580) );
  AOI211_X4 U19746 ( .C1(n18916), .C2(n18918), .A(n16581), .B(n16580), .ZN(
        n16964) );
  NOR3_X1 U19747 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16934) );
  INV_X1 U19748 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16928) );
  NAND2_X1 U19749 ( .A1(n16934), .A2(n16928), .ZN(n16925) );
  NOR2_X1 U19750 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16925), .ZN(n16910) );
  INV_X1 U19751 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16893) );
  NAND2_X1 U19752 ( .A1(n16910), .A2(n16893), .ZN(n16892) );
  INV_X1 U19753 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16873) );
  NAND2_X1 U19754 ( .A1(n16876), .A2(n16873), .ZN(n16872) );
  INV_X1 U19755 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16843) );
  NAND2_X1 U19756 ( .A1(n16850), .A2(n16843), .ZN(n16842) );
  INV_X1 U19757 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16822) );
  NAND2_X1 U19758 ( .A1(n16827), .A2(n16822), .ZN(n16821) );
  NAND2_X1 U19759 ( .A1(n16809), .A2(n16801), .ZN(n16800) );
  INV_X1 U19760 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16773) );
  NAND2_X1 U19761 ( .A1(n16783), .A2(n16773), .ZN(n16772) );
  INV_X1 U19762 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16756) );
  NAND2_X1 U19763 ( .A1(n16757), .A2(n16756), .ZN(n16749) );
  INV_X1 U19764 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16735) );
  NAND2_X1 U19765 ( .A1(n16736), .A2(n16735), .ZN(n16727) );
  NAND2_X1 U19766 ( .A1(n16714), .A2(n17061), .ZN(n16704) );
  INV_X1 U19767 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20891) );
  NAND2_X1 U19768 ( .A1(n16691), .A2(n20891), .ZN(n16687) );
  INV_X1 U19769 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16666) );
  NAND2_X1 U19770 ( .A1(n16678), .A2(n16666), .ZN(n16665) );
  NOR2_X1 U19771 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16665), .ZN(n16649) );
  NAND2_X1 U19772 ( .A1(n16649), .A2(n16968), .ZN(n16643) );
  NOR2_X1 U19773 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16643), .ZN(n16626) );
  INV_X1 U19774 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17008) );
  NAND2_X1 U19775 ( .A1(n16626), .A2(n17008), .ZN(n16604) );
  NOR2_X1 U19776 ( .A1(n16952), .A2(n16604), .ZN(n16611) );
  INV_X1 U19777 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16976) );
  OAI21_X1 U19778 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16583), .A(
        n16582), .ZN(n17568) );
  INV_X1 U19779 ( .A(n17568), .ZN(n16629) );
  OAI21_X1 U19780 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16585), .A(
        n16584), .ZN(n17586) );
  INV_X1 U19781 ( .A(n17586), .ZN(n16652) );
  INV_X1 U19782 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16588) );
  NOR2_X1 U19783 ( .A1(n16588), .A2(n16589), .ZN(n16587) );
  OAI21_X1 U19784 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16587), .A(
        n16586), .ZN(n17598) );
  INV_X1 U19785 ( .A(n17598), .ZN(n16660) );
  AOI21_X1 U19786 ( .B1(n16588), .B2(n16589), .A(n16587), .ZN(n17607) );
  AND2_X1 U19787 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17622), .ZN(
        n17623) );
  OAI21_X1 U19788 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17623), .A(
        n16589), .ZN(n16590) );
  INV_X1 U19789 ( .A(n16590), .ZN(n17625) );
  INV_X1 U19790 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17636) );
  NOR2_X1 U19791 ( .A1(n17918), .A2(n17679), .ZN(n16593) );
  INV_X1 U19792 ( .A(n16593), .ZN(n16745) );
  NOR2_X1 U19793 ( .A1(n16591), .A2(n16745), .ZN(n16594) );
  NAND2_X1 U19794 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16594), .ZN(
        n16592) );
  AOI21_X1 U19795 ( .B1(n17636), .B2(n16592), .A(n17623), .ZN(n17638) );
  INV_X1 U19796 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17637) );
  XOR2_X1 U19797 ( .A(n17637), .B(n16594), .Z(n17653) );
  INV_X1 U19798 ( .A(n17653), .ZN(n16703) );
  INV_X1 U19799 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16595) );
  NAND2_X1 U19800 ( .A1(n17664), .A2(n16593), .ZN(n17634) );
  AOI21_X1 U19801 ( .B1(n16595), .B2(n17634), .A(n16594), .ZN(n17669) );
  NOR3_X1 U19802 ( .A1(n17918), .A2(n17679), .A3(n17678), .ZN(n17677) );
  NAND2_X1 U19803 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17677), .ZN(
        n16738) );
  NOR2_X1 U19804 ( .A1(n17918), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16937) );
  INV_X1 U19805 ( .A(n16937), .ZN(n16908) );
  NOR3_X1 U19806 ( .A1(n17742), .A2(n17741), .A3(n16908), .ZN(n16769) );
  NAND2_X1 U19807 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16769), .ZN(
        n16759) );
  OAI21_X1 U19808 ( .B1(n16738), .B2(n16759), .A(n16949), .ZN(n16723) );
  NOR2_X1 U19809 ( .A1(n16702), .A2(n16918), .ZN(n16693) );
  NOR2_X1 U19810 ( .A1(n17607), .A2(n16673), .ZN(n16672) );
  NOR2_X1 U19811 ( .A1(n16672), .A2(n16918), .ZN(n16659) );
  NOR2_X1 U19812 ( .A1(n16638), .A2(n16637), .ZN(n16636) );
  NOR2_X1 U19813 ( .A1(n16636), .A2(n16918), .ZN(n16628) );
  NOR2_X1 U19814 ( .A1(n16629), .A2(n16628), .ZN(n16627) );
  NOR2_X1 U19815 ( .A1(n16627), .A2(n16918), .ZN(n16615) );
  NAND3_X1 U19816 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16597) );
  AND2_X1 U19817 ( .A1(n16920), .A2(n16596), .ZN(n16647) );
  NOR2_X1 U19818 ( .A1(n16961), .A2(n16647), .ZN(n16646) );
  INV_X1 U19819 ( .A(n16646), .ZN(n16655) );
  AOI21_X1 U19820 ( .B1(n16920), .B2(n16597), .A(n16655), .ZN(n16625) );
  NOR2_X1 U19821 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16598), .ZN(n16609) );
  INV_X1 U19822 ( .A(n16609), .ZN(n16599) );
  AOI21_X1 U19823 ( .B1(n16625), .B2(n16599), .A(n18847), .ZN(n16600) );
  OAI211_X1 U19824 ( .C1(n16603), .C2(n16947), .A(n16602), .B(n16601), .ZN(
        P3_U2640) );
  NAND2_X1 U19825 ( .A1(n16964), .A2(n16604), .ZN(n16621) );
  XOR2_X1 U19826 ( .A(n16606), .B(n16605), .Z(n16610) );
  INV_X1 U19827 ( .A(n18767), .ZN(n16946) );
  OAI22_X1 U19828 ( .A1(n16625), .A2(n18849), .B1(n16607), .B2(n16947), .ZN(
        n16608) );
  AOI211_X1 U19829 ( .C1(n16610), .C2(n16946), .A(n16609), .B(n16608), .ZN(
        n16613) );
  OAI21_X1 U19830 ( .B1(n16965), .B2(n16611), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16612) );
  OAI211_X1 U19831 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16621), .A(n16613), .B(
        n16612), .ZN(P3_U2641) );
  INV_X1 U19832 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18844) );
  AOI211_X1 U19833 ( .C1(n16616), .C2(n16615), .A(n16614), .B(n18767), .ZN(
        n16620) );
  NAND3_X1 U19834 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16642), .ZN(n16618) );
  OAI22_X1 U19835 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16618), .B1(n16617), 
        .B2(n16947), .ZN(n16619) );
  AOI211_X1 U19836 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16965), .A(n16620), .B(
        n16619), .ZN(n16624) );
  INV_X1 U19837 ( .A(n16621), .ZN(n16622) );
  OAI21_X1 U19838 ( .B1(n16626), .B2(n17008), .A(n16622), .ZN(n16623) );
  OAI211_X1 U19839 ( .C1(n16625), .C2(n18844), .A(n16624), .B(n16623), .ZN(
        P3_U2642) );
  AOI22_X1 U19840 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16900), .B1(
        n16965), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16635) );
  AOI211_X1 U19841 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16643), .A(n16626), .B(
        n16952), .ZN(n16631) );
  AOI211_X1 U19842 ( .C1(n16629), .C2(n16628), .A(n16627), .B(n18767), .ZN(
        n16630) );
  AOI211_X1 U19843 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16655), .A(n16631), 
        .B(n16630), .ZN(n16634) );
  NAND2_X1 U19844 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16632) );
  OAI211_X1 U19845 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16642), .B(n16632), .ZN(n16633) );
  NAND3_X1 U19846 ( .A1(n16635), .A2(n16634), .A3(n16633), .ZN(P3_U2643) );
  INV_X1 U19847 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18840) );
  AOI211_X1 U19848 ( .C1(n16638), .C2(n16637), .A(n16636), .B(n18767), .ZN(
        n16641) );
  OAI22_X1 U19849 ( .A1(n16639), .A2(n16947), .B1(n16953), .B2(n16968), .ZN(
        n16640) );
  AOI211_X1 U19850 ( .C1(n16642), .C2(n18840), .A(n16641), .B(n16640), .ZN(
        n16645) );
  OAI211_X1 U19851 ( .C1(n16649), .C2(n16968), .A(n16964), .B(n16643), .ZN(
        n16644) );
  OAI211_X1 U19852 ( .C1(n16646), .C2(n18840), .A(n16645), .B(n16644), .ZN(
        P3_U2644) );
  INV_X1 U19853 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17585) );
  AOI22_X1 U19854 ( .A1(n16965), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16648), 
        .B2(n16647), .ZN(n16657) );
  AOI211_X1 U19855 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16665), .A(n16649), .B(
        n16952), .ZN(n16654) );
  AOI211_X1 U19856 ( .C1(n16652), .C2(n16651), .A(n16650), .B(n18767), .ZN(
        n16653) );
  AOI211_X1 U19857 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16655), .A(n16654), 
        .B(n16653), .ZN(n16656) );
  OAI211_X1 U19858 ( .C1(n17585), .C2(n16947), .A(n16657), .B(n16656), .ZN(
        P3_U2645) );
  INV_X1 U19859 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18834) );
  INV_X1 U19860 ( .A(n16961), .ZN(n16932) );
  OAI21_X1 U19861 ( .B1(n16682), .B2(n16959), .A(n16932), .ZN(n16679) );
  AOI21_X1 U19862 ( .B1(n16920), .B2(n18834), .A(n16679), .ZN(n16669) );
  AOI211_X1 U19863 ( .C1(n16660), .C2(n16659), .A(n16658), .B(n18767), .ZN(
        n16664) );
  NAND2_X1 U19864 ( .A1(n16920), .A2(n18836), .ZN(n16661) );
  OAI22_X1 U19865 ( .A1(n16953), .A2(n16666), .B1(n16662), .B2(n16661), .ZN(
        n16663) );
  AOI211_X1 U19866 ( .C1(n16900), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16664), .B(n16663), .ZN(n16668) );
  OAI211_X1 U19867 ( .C1(n16678), .C2(n16666), .A(n16964), .B(n16665), .ZN(
        n16667) );
  OAI211_X1 U19868 ( .C1(n16669), .C2(n18836), .A(n16668), .B(n16667), .ZN(
        P3_U2646) );
  AOI21_X1 U19869 ( .B1(n16687), .B2(P3_EBX_REG_24__SCAN_IN), .A(n16952), .ZN(
        n16670) );
  AOI21_X1 U19870 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16965), .A(n16670), .ZN(
        n16677) );
  NOR2_X1 U19871 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16959), .ZN(n16671) );
  AOI22_X1 U19872 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16900), .B1(
        n16682), .B2(n16671), .ZN(n16676) );
  AOI211_X1 U19873 ( .C1(n17607), .C2(n16673), .A(n16672), .B(n18767), .ZN(
        n16674) );
  AOI21_X1 U19874 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16679), .A(n16674), 
        .ZN(n16675) );
  OAI211_X1 U19875 ( .C1(n16678), .C2(n16677), .A(n16676), .B(n16675), .ZN(
        P3_U2647) );
  INV_X1 U19876 ( .A(n16679), .ZN(n16690) );
  AOI211_X1 U19877 ( .C1(n17625), .C2(n16681), .A(n16680), .B(n18767), .ZN(
        n16686) );
  OR2_X1 U19878 ( .A1(n16959), .A2(n16682), .ZN(n16683) );
  OAI22_X1 U19879 ( .A1(n16953), .A2(n20891), .B1(n16684), .B2(n16683), .ZN(
        n16685) );
  AOI211_X1 U19880 ( .C1(n16900), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16686), .B(n16685), .ZN(n16689) );
  OAI211_X1 U19881 ( .C1(n16691), .C2(n20891), .A(n16964), .B(n16687), .ZN(
        n16688) );
  OAI211_X1 U19882 ( .C1(n16690), .C2(n18833), .A(n16689), .B(n16688), .ZN(
        P3_U2648) );
  AOI221_X1 U19883 ( .B1(n18829), .B2(n16920), .C1(n16701), .C2(n16920), .A(
        n16961), .ZN(n16700) );
  INV_X1 U19884 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18830) );
  AOI22_X1 U19885 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16900), .B1(
        n16965), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16699) );
  NOR2_X1 U19886 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16959), .ZN(n16696) );
  AOI211_X1 U19887 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16704), .A(n16691), .B(
        n16952), .ZN(n16695) );
  AOI211_X1 U19888 ( .C1(n17638), .C2(n16693), .A(n16692), .B(n18767), .ZN(
        n16694) );
  AOI211_X1 U19889 ( .C1(n16697), .C2(n16696), .A(n16695), .B(n16694), .ZN(
        n16698) );
  OAI211_X1 U19890 ( .C1(n16700), .C2(n18830), .A(n16699), .B(n16698), .ZN(
        P3_U2649) );
  INV_X1 U19891 ( .A(n16701), .ZN(n16708) );
  NOR2_X1 U19892 ( .A1(n16959), .A2(n16708), .ZN(n16716) );
  OR2_X1 U19893 ( .A1(n16961), .A2(n16716), .ZN(n16718) );
  AOI211_X1 U19894 ( .C1(n16703), .C2(n9716), .A(n16702), .B(n18767), .ZN(
        n16707) );
  OAI211_X1 U19895 ( .C1(n16714), .C2(n17061), .A(n16964), .B(n16704), .ZN(
        n16705) );
  OAI21_X1 U19896 ( .B1(n16947), .B2(n17637), .A(n16705), .ZN(n16706) );
  AOI211_X1 U19897 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16718), .A(n16707), 
        .B(n16706), .ZN(n16710) );
  NAND3_X1 U19898 ( .A1(n16920), .A2(n16708), .A3(n18829), .ZN(n16709) );
  OAI211_X1 U19899 ( .C1(n17061), .C2(n16953), .A(n16710), .B(n16709), .ZN(
        P3_U2650) );
  AOI211_X1 U19900 ( .C1(n17669), .C2(n16712), .A(n16711), .B(n18767), .ZN(
        n16713) );
  AOI21_X1 U19901 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16965), .A(n16713), .ZN(
        n16721) );
  AOI211_X1 U19902 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16727), .A(n16714), .B(
        n16952), .ZN(n16715) );
  AOI21_X1 U19903 ( .B1(n16900), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16715), .ZN(n16720) );
  AOI22_X1 U19904 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16718), .B1(n16717), 
        .B2(n16716), .ZN(n16719) );
  NAND3_X1 U19905 ( .A1(n16721), .A2(n16720), .A3(n16719), .ZN(P3_U2651) );
  INV_X1 U19906 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16730) );
  INV_X1 U19907 ( .A(n17634), .ZN(n16722) );
  AOI21_X1 U19908 ( .B1(n16730), .B2(n16738), .A(n16722), .ZN(n16724) );
  INV_X1 U19909 ( .A(n16724), .ZN(n17683) );
  OAI221_X1 U19910 ( .B1(n16724), .B2(n16723), .C1(n17683), .C2(n9890), .A(
        n18253), .ZN(n16733) );
  NOR3_X1 U19911 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16959), .A3(n16725), 
        .ZN(n16732) );
  OAI21_X1 U19912 ( .B1(n16726), .B2(n16959), .A(n16932), .ZN(n16754) );
  INV_X1 U19913 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18822) );
  AND3_X1 U19914 ( .A1(n18822), .A2(n16920), .A3(n16726), .ZN(n16740) );
  OAI21_X1 U19915 ( .B1(n16754), .B2(n16740), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16729) );
  OAI211_X1 U19916 ( .C1(n16736), .C2(n16735), .A(n16964), .B(n16727), .ZN(
        n16728) );
  OAI211_X1 U19917 ( .C1(n16947), .C2(n16730), .A(n16729), .B(n16728), .ZN(
        n16731) );
  AOI211_X1 U19918 ( .C1(n16758), .C2(n16733), .A(n16732), .B(n16731), .ZN(
        n16734) );
  OAI21_X1 U19919 ( .B1(n16953), .B2(n16735), .A(n16734), .ZN(P3_U2652) );
  AOI211_X1 U19920 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16749), .A(n16736), .B(
        n16952), .ZN(n16737) );
  AOI21_X1 U19921 ( .B1(n16900), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16737), .ZN(n16744) );
  OAI21_X1 U19922 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17677), .A(
        n16738), .ZN(n17692) );
  INV_X1 U19923 ( .A(n16759), .ZN(n16746) );
  AOI21_X1 U19924 ( .B1(n17677), .B2(n16746), .A(n16918), .ZN(n16739) );
  XNOR2_X1 U19925 ( .A(n17692), .B(n16739), .ZN(n16741) );
  AOI21_X1 U19926 ( .B1(n16741), .B2(n16946), .A(n16740), .ZN(n16743) );
  AOI22_X1 U19927 ( .A1(n16965), .A2(P3_EBX_REG_18__SCAN_IN), .B1(
        P3_REIP_REG_18__SCAN_IN), .B2(n16754), .ZN(n16742) );
  NAND4_X1 U19928 ( .A1(n16744), .A2(n16743), .A3(n16742), .A4(n18253), .ZN(
        P3_U2653) );
  NAND4_X1 U19929 ( .A1(n16920), .A2(n16782), .A3(P3_REIP_REG_14__SCAN_IN), 
        .A4(P3_REIP_REG_13__SCAN_IN), .ZN(n16780) );
  OAI21_X1 U19930 ( .B1(n16765), .B2(n16780), .A(n20986), .ZN(n16753) );
  AOI21_X1 U19931 ( .B1(n17678), .B2(n16745), .A(n17677), .ZN(n17707) );
  INV_X1 U19932 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17733) );
  NOR2_X1 U19933 ( .A1(n17918), .A2(n17742), .ZN(n16793) );
  NAND2_X1 U19934 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16793), .ZN(
        n17714) );
  NOR2_X1 U19935 ( .A1(n17733), .A2(n17714), .ZN(n16770) );
  OAI21_X1 U19936 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16770), .A(
        n16745), .ZN(n17715) );
  AOI21_X1 U19937 ( .B1(n16746), .B2(n17715), .A(n16918), .ZN(n16748) );
  AOI21_X1 U19938 ( .B1(n17707), .B2(n16748), .A(n18767), .ZN(n16747) );
  OAI21_X1 U19939 ( .B1(n17707), .B2(n16748), .A(n16747), .ZN(n16751) );
  OAI211_X1 U19940 ( .C1(n16757), .C2(n16756), .A(n16964), .B(n16749), .ZN(
        n16750) );
  OAI211_X1 U19941 ( .C1(n16947), .C2(n17678), .A(n16751), .B(n16750), .ZN(
        n16752) );
  AOI21_X1 U19942 ( .B1(n16754), .B2(n16753), .A(n16752), .ZN(n16755) );
  OAI211_X1 U19943 ( .C1(n16953), .C2(n16756), .A(n16755), .B(n18253), .ZN(
        P3_U2654) );
  AOI21_X1 U19944 ( .B1(n16920), .B2(n16781), .A(n16961), .ZN(n16779) );
  INV_X1 U19945 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18819) );
  AOI211_X1 U19946 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16772), .A(n16757), .B(
        n16952), .ZN(n16764) );
  INV_X1 U19947 ( .A(n16758), .ZN(n16906) );
  NAND2_X1 U19948 ( .A1(n16949), .A2(n16759), .ZN(n16760) );
  NAND2_X1 U19949 ( .A1(n17715), .A2(n16760), .ZN(n16761) );
  AOI221_X1 U19950 ( .B1(n17715), .B2(n16761), .C1(n16760), .C2(n16761), .A(
        n9587), .ZN(n16762) );
  OAI22_X1 U19951 ( .A1(n16906), .A2(n16762), .B1(n16953), .B2(n17121), .ZN(
        n16763) );
  AOI211_X1 U19952 ( .C1(n16900), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16764), .B(n16763), .ZN(n16768) );
  INV_X1 U19953 ( .A(n16780), .ZN(n16766) );
  OAI211_X1 U19954 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16766), .B(n16765), .ZN(n16767) );
  OAI211_X1 U19955 ( .C1(n16779), .C2(n18819), .A(n16768), .B(n16767), .ZN(
        P3_U2655) );
  INV_X1 U19956 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18817) );
  OAI22_X1 U19957 ( .A1(n17733), .A2(n16947), .B1(n16953), .B2(n16773), .ZN(
        n16777) );
  NOR2_X1 U19958 ( .A1(n16769), .A2(n16918), .ZN(n16771) );
  AOI21_X1 U19959 ( .B1(n17733), .B2(n17714), .A(n16770), .ZN(n17736) );
  XNOR2_X1 U19960 ( .A(n16771), .B(n17736), .ZN(n16775) );
  OAI211_X1 U19961 ( .C1(n16783), .C2(n16773), .A(n16964), .B(n16772), .ZN(
        n16774) );
  OAI21_X1 U19962 ( .B1(n18767), .B2(n16775), .A(n16774), .ZN(n16776) );
  NOR3_X1 U19963 ( .A1(n9587), .A2(n16777), .A3(n16776), .ZN(n16778) );
  OAI221_X1 U19964 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16780), .C1(n18817), 
        .C2(n16779), .A(n16778), .ZN(P3_U2656) );
  NOR2_X1 U19965 ( .A1(n16961), .A2(n16781), .ZN(n16792) );
  NAND2_X1 U19966 ( .A1(n16932), .A2(n16959), .ZN(n16963) );
  AND2_X1 U19967 ( .A1(n16920), .A2(n16782), .ZN(n16799) );
  AOI22_X1 U19968 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16963), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16799), .ZN(n16791) );
  AOI211_X1 U19969 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16800), .A(n16783), .B(
        n16952), .ZN(n16789) );
  OAI21_X1 U19970 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16793), .A(
        n17714), .ZN(n17753) );
  OAI21_X1 U19971 ( .B1(n17742), .B2(n16908), .A(n16949), .ZN(n16785) );
  AOI21_X1 U19972 ( .B1(n17753), .B2(n16785), .A(n18767), .ZN(n16784) );
  OAI21_X1 U19973 ( .B1(n17753), .B2(n16785), .A(n16784), .ZN(n16786) );
  OAI211_X1 U19974 ( .C1(n16953), .C2(n16787), .A(n18253), .B(n16786), .ZN(
        n16788) );
  AOI211_X1 U19975 ( .C1(n16900), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16789), .B(n16788), .ZN(n16790) );
  OAI21_X1 U19976 ( .B1(n16792), .B2(n16791), .A(n16790), .ZN(P3_U2657) );
  INV_X1 U19977 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16796) );
  INV_X1 U19978 ( .A(n16857), .ZN(n17823) );
  NAND2_X1 U19979 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17823), .ZN(
        n16879) );
  NOR2_X1 U19980 ( .A1(n17784), .A2(n16879), .ZN(n16828) );
  NAND2_X1 U19981 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16828), .ZN(
        n17754) );
  INV_X1 U19982 ( .A(n17754), .ZN(n16806) );
  NAND2_X1 U19983 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16806), .ZN(
        n16805) );
  AOI21_X1 U19984 ( .B1(n16796), .B2(n16805), .A(n16793), .ZN(n17757) );
  OAI21_X1 U19985 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16805), .A(
        n16949), .ZN(n16795) );
  OAI21_X1 U19986 ( .B1(n17757), .B2(n16795), .A(n18253), .ZN(n16794) );
  AOI21_X1 U19987 ( .B1(n17757), .B2(n16795), .A(n16794), .ZN(n16804) );
  INV_X1 U19988 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18813) );
  AOI21_X1 U19989 ( .B1(n16920), .B2(n16811), .A(n16961), .ZN(n16826) );
  OAI21_X1 U19990 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16959), .A(n16826), 
        .ZN(n16798) );
  OAI22_X1 U19991 ( .A1(n16796), .A2(n16947), .B1(n16953), .B2(n16801), .ZN(
        n16797) );
  AOI221_X1 U19992 ( .B1(n16799), .B2(n18813), .C1(n16798), .C2(
        P3_REIP_REG_13__SCAN_IN), .A(n16797), .ZN(n16803) );
  OAI211_X1 U19993 ( .C1(n16809), .C2(n16801), .A(n16964), .B(n16800), .ZN(
        n16802) );
  OAI211_X1 U19994 ( .C1(n16906), .C2(n16804), .A(n16803), .B(n16802), .ZN(
        P3_U2658) );
  INV_X1 U19995 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17770) );
  OAI21_X1 U19996 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16806), .A(
        n16805), .ZN(n17779) );
  NAND2_X1 U19997 ( .A1(n17823), .A2(n16937), .ZN(n16866) );
  OAI21_X1 U19998 ( .B1(n17784), .B2(n16866), .A(n16949), .ZN(n16818) );
  OAI21_X1 U19999 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16918), .A(
        n16818), .ZN(n16807) );
  XNOR2_X1 U20000 ( .A(n17779), .B(n16807), .ZN(n16808) );
  AOI21_X1 U20001 ( .B1(n16808), .B2(n16946), .A(n9587), .ZN(n16815) );
  AOI211_X1 U20002 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16821), .A(n16809), .B(
        n16952), .ZN(n16813) );
  NAND2_X1 U20003 ( .A1(n16920), .A2(n18812), .ZN(n16810) );
  OAI22_X1 U20004 ( .A1(n16826), .A2(n18812), .B1(n16811), .B2(n16810), .ZN(
        n16812) );
  AOI211_X1 U20005 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16965), .A(n16813), .B(
        n16812), .ZN(n16814) );
  OAI211_X1 U20006 ( .C1(n17770), .C2(n16947), .A(n16815), .B(n16814), .ZN(
        P3_U2659) );
  NAND2_X1 U20007 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16835) );
  INV_X1 U20008 ( .A(n16835), .ZN(n16817) );
  INV_X1 U20009 ( .A(n16816), .ZN(n16851) );
  NOR2_X1 U20010 ( .A1(n16959), .A2(n16851), .ZN(n16847) );
  AOI21_X1 U20011 ( .B1(n16817), .B2(n16847), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16825) );
  OAI21_X1 U20012 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16828), .A(
        n17754), .ZN(n17787) );
  XNOR2_X1 U20013 ( .A(n17787), .B(n16818), .ZN(n16819) );
  OAI22_X1 U20014 ( .A1(n16953), .A2(n16822), .B1(n18767), .B2(n16819), .ZN(
        n16820) );
  AOI211_X1 U20015 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16900), .A(
        n9587), .B(n16820), .ZN(n16824) );
  OAI211_X1 U20016 ( .C1(n16827), .C2(n16822), .A(n16964), .B(n16821), .ZN(
        n16823) );
  OAI211_X1 U20017 ( .C1(n16826), .C2(n16825), .A(n16824), .B(n16823), .ZN(
        P3_U2660) );
  AOI21_X1 U20018 ( .B1(n16920), .B2(n16851), .A(n16961), .ZN(n16854) );
  INV_X1 U20019 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18807) );
  AOI211_X1 U20020 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16842), .A(n16827), .B(
        n16952), .ZN(n16834) );
  INV_X1 U20021 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17796) );
  NOR2_X1 U20022 ( .A1(n17797), .A2(n16879), .ZN(n16838) );
  INV_X1 U20023 ( .A(n16838), .ZN(n16858) );
  NOR2_X1 U20024 ( .A1(n17796), .A2(n16858), .ZN(n16830) );
  INV_X1 U20025 ( .A(n16828), .ZN(n16829) );
  OAI21_X1 U20026 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16830), .A(
        n16829), .ZN(n17798) );
  INV_X1 U20027 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17842) );
  NOR2_X1 U20028 ( .A1(n17842), .A2(n16866), .ZN(n16859) );
  NAND2_X1 U20029 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16859), .ZN(
        n16840) );
  OAI21_X1 U20030 ( .B1(n17796), .B2(n16840), .A(n16949), .ZN(n16839) );
  AOI21_X1 U20031 ( .B1(n17798), .B2(n16839), .A(n18767), .ZN(n16831) );
  OAI21_X1 U20032 ( .B1(n17798), .B2(n16839), .A(n16831), .ZN(n16832) );
  OAI211_X1 U20033 ( .C1(n16953), .C2(n17205), .A(n18253), .B(n16832), .ZN(
        n16833) );
  AOI211_X1 U20034 ( .C1(n16900), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16834), .B(n16833), .ZN(n16837) );
  OAI211_X1 U20035 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16847), .B(n16835), .ZN(n16836) );
  OAI211_X1 U20036 ( .C1(n16854), .C2(n18807), .A(n16837), .B(n16836), .ZN(
        P3_U2661) );
  INV_X1 U20037 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18805) );
  AOI22_X1 U20038 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16900), .B1(
        n16965), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16849) );
  OAI22_X1 U20039 ( .A1(n17796), .A2(n16838), .B1(n16858), .B2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16841) );
  AOI211_X1 U20040 ( .C1(n16841), .C2(n16840), .A(n18767), .B(n16839), .ZN(
        n16846) );
  INV_X1 U20041 ( .A(n16841), .ZN(n17813) );
  NAND2_X1 U20042 ( .A1(n16946), .A2(n16918), .ZN(n16939) );
  OAI211_X1 U20043 ( .C1(n16850), .C2(n16843), .A(n16964), .B(n16842), .ZN(
        n16844) );
  OAI211_X1 U20044 ( .C1(n17813), .C2(n16939), .A(n18253), .B(n16844), .ZN(
        n16845) );
  AOI211_X1 U20045 ( .C1(n16847), .C2(n18805), .A(n16846), .B(n16845), .ZN(
        n16848) );
  OAI211_X1 U20046 ( .C1(n16854), .C2(n18805), .A(n16849), .B(n16848), .ZN(
        P3_U2662) );
  AOI211_X1 U20047 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16872), .A(n16850), .B(
        n16952), .ZN(n16856) );
  NAND2_X1 U20048 ( .A1(n16920), .A2(n16851), .ZN(n16852) );
  OAI22_X1 U20049 ( .A1(n16854), .A2(n18804), .B1(n16853), .B2(n16852), .ZN(
        n16855) );
  AOI211_X1 U20050 ( .C1(n16900), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16856), .B(n16855), .ZN(n16863) );
  NOR3_X1 U20051 ( .A1(n17918), .A2(n16857), .A3(n17842), .ZN(n16865) );
  OAI21_X1 U20052 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16865), .A(
        n16858), .ZN(n17826) );
  NOR2_X1 U20053 ( .A1(n16859), .A2(n16918), .ZN(n16860) );
  XNOR2_X1 U20054 ( .A(n17826), .B(n16860), .ZN(n16861) );
  AOI21_X1 U20055 ( .B1(n16861), .B2(n16946), .A(n9587), .ZN(n16862) );
  OAI211_X1 U20056 ( .C1(n17262), .C2(n16953), .A(n16863), .B(n16862), .ZN(
        P3_U2663) );
  AOI21_X1 U20057 ( .B1(n16920), .B2(n16864), .A(n16961), .ZN(n16889) );
  OR3_X1 U20058 ( .A1(n16959), .A2(n16864), .A3(P3_REIP_REG_6__SCAN_IN), .ZN(
        n16885) );
  INV_X1 U20059 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18801) );
  AOI21_X1 U20060 ( .B1(n16889), .B2(n16885), .A(n18801), .ZN(n16871) );
  AOI21_X1 U20061 ( .B1(n17842), .B2(n16879), .A(n16865), .ZN(n17846) );
  NAND2_X1 U20062 ( .A1(n16949), .A2(n16866), .ZN(n16878) );
  XOR2_X1 U20063 ( .A(n17846), .B(n16878), .Z(n16869) );
  NAND3_X1 U20064 ( .A1(n16920), .A2(n16867), .A3(n18801), .ZN(n16868) );
  OAI211_X1 U20065 ( .C1(n16869), .C2(n18767), .A(n18253), .B(n16868), .ZN(
        n16870) );
  AOI211_X1 U20066 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16965), .A(n16871), .B(
        n16870), .ZN(n16875) );
  OAI211_X1 U20067 ( .C1(n16876), .C2(n16873), .A(n16964), .B(n16872), .ZN(
        n16874) );
  OAI211_X1 U20068 ( .C1(n16947), .C2(n17842), .A(n16875), .B(n16874), .ZN(
        P3_U2664) );
  INV_X1 U20069 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16887) );
  AOI211_X1 U20070 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16892), .A(n16876), .B(
        n16952), .ZN(n16884) );
  AND2_X1 U20071 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17855), .ZN(
        n16894) );
  INV_X1 U20072 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16960) );
  OAI221_X1 U20073 ( .B1(n16918), .B2(n16894), .C1(n16918), .C2(n16960), .A(
        n16946), .ZN(n16877) );
  INV_X1 U20074 ( .A(n16877), .ZN(n16881) );
  NOR2_X1 U20075 ( .A1(n18767), .A2(n16878), .ZN(n16880) );
  OAI21_X1 U20076 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16894), .A(
        n16879), .ZN(n17858) );
  MUX2_X1 U20077 ( .A(n16881), .B(n16880), .S(n17858), .Z(n16883) );
  OAI22_X1 U20078 ( .A1(n16953), .A2(n17267), .B1(n18799), .B2(n16889), .ZN(
        n16882) );
  NOR4_X1 U20079 ( .A1(n9587), .A2(n16884), .A3(n16883), .A4(n16882), .ZN(
        n16886) );
  OAI211_X1 U20080 ( .C1(n16947), .C2(n16887), .A(n16886), .B(n16885), .ZN(
        P3_U2665) );
  AOI21_X1 U20081 ( .B1(n16920), .B2(n16888), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16890) );
  OAI22_X1 U20082 ( .A1(n16890), .A2(n16889), .B1(n17865), .B2(n16947), .ZN(
        n16891) );
  AOI21_X1 U20083 ( .B1(n16965), .B2(P3_EBX_REG_5__SCAN_IN), .A(n16891), .ZN(
        n16899) );
  OAI211_X1 U20084 ( .C1(n16910), .C2(n16893), .A(n16964), .B(n16892), .ZN(
        n16898) );
  OR2_X1 U20085 ( .A1(n17918), .A2(n17866), .ZN(n16902) );
  AOI21_X1 U20086 ( .B1(n17865), .B2(n16902), .A(n16894), .ZN(n16896) );
  OAI21_X1 U20087 ( .B1(n17866), .B2(n16908), .A(n16949), .ZN(n16895) );
  INV_X1 U20088 ( .A(n16895), .ZN(n16904) );
  INV_X1 U20089 ( .A(n16896), .ZN(n17871) );
  OAI221_X1 U20090 ( .B1(n16896), .B2(n16904), .C1(n17871), .C2(n16895), .A(
        n16946), .ZN(n16897) );
  NAND4_X1 U20091 ( .A1(n16899), .A2(n18253), .A3(n16898), .A4(n16897), .ZN(
        P3_U2666) );
  AOI21_X1 U20092 ( .B1(n16920), .B2(n16909), .A(n16961), .ZN(n16921) );
  AOI22_X1 U20093 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16900), .B1(
        n16965), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16916) );
  INV_X1 U20094 ( .A(n18914), .ZN(n18930) );
  NOR2_X1 U20095 ( .A1(n18269), .A2(n18930), .ZN(n16945) );
  INV_X1 U20096 ( .A(n16945), .ZN(n18932) );
  AOI21_X1 U20097 ( .B1(n9649), .B2(n16901), .A(n18932), .ZN(n16914) );
  NOR2_X1 U20098 ( .A1(n17918), .A2(n16905), .ZN(n16917) );
  OAI21_X1 U20099 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16917), .A(
        n16902), .ZN(n17884) );
  INV_X1 U20100 ( .A(n17884), .ZN(n16903) );
  AOI221_X1 U20101 ( .B1(n16904), .B2(n17884), .C1(n16918), .C2(n16903), .A(
        n9587), .ZN(n16907) );
  OR2_X1 U20102 ( .A1(n16905), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17876) );
  AOI221_X1 U20103 ( .B1(n16908), .B2(n16907), .C1(n17876), .C2(n16907), .A(
        n16906), .ZN(n16913) );
  NOR3_X1 U20104 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16959), .A3(n16909), .ZN(
        n16912) );
  AOI211_X1 U20105 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16925), .A(n16910), .B(
        n16952), .ZN(n16911) );
  NOR4_X1 U20106 ( .A1(n16914), .A2(n16913), .A3(n16912), .A4(n16911), .ZN(
        n16915) );
  OAI211_X1 U20107 ( .C1(n18795), .C2(n16921), .A(n16916), .B(n16915), .ZN(
        P3_U2667) );
  NAND2_X1 U20108 ( .A1(n18726), .A2(n18715), .ZN(n18713) );
  AOI21_X1 U20109 ( .B1(n18868), .B2(n18713), .A(n17258), .ZN(n18866) );
  INV_X1 U20110 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17892) );
  NAND2_X1 U20111 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16935) );
  AOI21_X1 U20112 ( .B1(n17892), .B2(n16935), .A(n16917), .ZN(n17896) );
  AOI21_X1 U20113 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16937), .A(
        n16918), .ZN(n16936) );
  OAI21_X1 U20114 ( .B1(n17896), .B2(n16936), .A(n16946), .ZN(n16919) );
  AOI21_X1 U20115 ( .B1(n17896), .B2(n16936), .A(n16919), .ZN(n16924) );
  INV_X1 U20116 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18791) );
  NOR2_X1 U20117 ( .A1(n18895), .A2(n18791), .ZN(n16929) );
  AOI21_X1 U20118 ( .B1(n16920), .B2(n16929), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n16922) );
  OAI22_X1 U20119 ( .A1(n16922), .A2(n16921), .B1(n17892), .B2(n16947), .ZN(
        n16923) );
  AOI211_X1 U20120 ( .C1(n16945), .C2(n18866), .A(n16924), .B(n16923), .ZN(
        n16927) );
  OAI211_X1 U20121 ( .C1(n16934), .C2(n16928), .A(n16964), .B(n16925), .ZN(
        n16926) );
  OAI211_X1 U20122 ( .C1(n16928), .C2(n16953), .A(n16927), .B(n16926), .ZN(
        P3_U2668) );
  INV_X1 U20123 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17909) );
  AOI211_X1 U20124 ( .C1(n18895), .C2(n18791), .A(n16929), .B(n16959), .ZN(
        n16930) );
  AOI21_X1 U20125 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n16965), .A(n16930), .ZN(
        n16943) );
  AOI22_X1 U20126 ( .A1(n18715), .A2(n18726), .B1(n18878), .B2(n18731), .ZN(
        n18874) );
  NOR2_X1 U20127 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16950) );
  OAI21_X1 U20128 ( .B1(n16950), .B2(n16931), .A(n16964), .ZN(n16933) );
  OAI22_X1 U20129 ( .A1(n16934), .A2(n16933), .B1(n18791), .B2(n16932), .ZN(
        n16941) );
  OAI21_X1 U20130 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16935), .ZN(n17904) );
  OAI211_X1 U20131 ( .C1(n16937), .C2(n17904), .A(n16946), .B(n16936), .ZN(
        n16938) );
  OAI21_X1 U20132 ( .B1(n16939), .B2(n17904), .A(n16938), .ZN(n16940) );
  AOI211_X1 U20133 ( .C1(n18874), .C2(n16945), .A(n16941), .B(n16940), .ZN(
        n16942) );
  OAI211_X1 U20134 ( .C1(n17909), .C2(n16947), .A(n16943), .B(n16942), .ZN(
        P3_U2669) );
  INV_X1 U20135 ( .A(n18731), .ZN(n18717) );
  NOR2_X1 U20136 ( .A1(n18717), .A2(n16944), .ZN(n18882) );
  AOI22_X1 U20137 ( .A1(n16961), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18882), 
        .B2(n16945), .ZN(n16958) );
  NAND2_X1 U20138 ( .A1(n16949), .A2(n16946), .ZN(n16948) );
  OAI211_X1 U20139 ( .C1(n16960), .C2(n16948), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n16947), .ZN(n16956) );
  AOI21_X1 U20140 ( .B1(n16949), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18767), .ZN(n16955) );
  INV_X1 U20141 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17292) );
  INV_X1 U20142 ( .A(n16950), .ZN(n16951) );
  NAND2_X1 U20143 ( .A1(n16951), .A2(n17285), .ZN(n17293) );
  OAI22_X1 U20144 ( .A1(n16953), .A2(n17292), .B1(n16952), .B2(n17293), .ZN(
        n16954) );
  AOI221_X1 U20145 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16956), .C1(
        n16955), .C2(n16956), .A(n16954), .ZN(n16957) );
  OAI211_X1 U20146 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n16959), .A(n16958), .B(
        n16957), .ZN(P3_U2670) );
  NOR3_X1 U20147 ( .A1(n18889), .A2(n16961), .A3(n16960), .ZN(n16962) );
  AOI21_X1 U20148 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n16963), .A(n16962), .ZN(
        n16967) );
  OAI21_X1 U20149 ( .B1(n16965), .B2(n16964), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16966) );
  OAI211_X1 U20150 ( .C1(n18726), .C2(n18932), .A(n16967), .B(n16966), .ZN(
        P3_U2671) );
  NOR4_X1 U20151 ( .A1(n16969), .A2(n16968), .A3(n20891), .A4(n17061), .ZN(
        n16972) );
  INV_X1 U20152 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U20153 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .ZN(n16970) );
  NOR4_X1 U20154 ( .A1(n17008), .A2(n17047), .A3(n17090), .A4(n16970), .ZN(
        n16971) );
  NAND4_X1 U20155 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n16972), .A4(n16971), .ZN(n16975) );
  NAND2_X1 U20156 ( .A1(n9582), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16974) );
  NAND2_X1 U20157 ( .A1(n17003), .A2(n17425), .ZN(n16973) );
  OAI22_X1 U20158 ( .A1(n17003), .A2(n16974), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16973), .ZN(P3_U2672) );
  NAND2_X1 U20159 ( .A1(n16976), .A2(n16975), .ZN(n16977) );
  NAND2_X1 U20160 ( .A1(n16977), .A2(n9582), .ZN(n17002) );
  AOI22_X1 U20161 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16987) );
  INV_X1 U20162 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20163 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20164 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16978) );
  OAI211_X1 U20165 ( .C1(n9649), .C2(n17141), .A(n16979), .B(n16978), .ZN(
        n16985) );
  AOI22_X1 U20166 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20167 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U20168 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16981) );
  NAND2_X1 U20169 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n16980) );
  NAND4_X1 U20170 ( .A1(n16983), .A2(n16982), .A3(n16981), .A4(n16980), .ZN(
        n16984) );
  AOI211_X1 U20171 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n16985), .B(n16984), .ZN(n16986) );
  OAI211_X1 U20172 ( .C1(n17199), .C2(n16988), .A(n16987), .B(n16986), .ZN(
        n17001) );
  AOI22_X1 U20173 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20174 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20175 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16997) );
  OAI22_X1 U20176 ( .A1(n10131), .A2(n17158), .B1(n17142), .B2(n16989), .ZN(
        n16995) );
  AOI22_X1 U20177 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20178 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20179 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16991) );
  NAND2_X1 U20180 ( .A1(n10178), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n16990) );
  NAND4_X1 U20181 ( .A1(n16993), .A2(n16992), .A3(n16991), .A4(n16990), .ZN(
        n16994) );
  AOI211_X1 U20182 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n16995), .B(n16994), .ZN(n16996) );
  NAND4_X1 U20183 ( .A1(n16999), .A2(n16998), .A3(n16997), .A4(n16996), .ZN(
        n17007) );
  NAND3_X1 U20184 ( .A1(n17007), .A2(n17004), .A3(n17005), .ZN(n17000) );
  XOR2_X1 U20185 ( .A(n17001), .B(n17000), .Z(n17312) );
  OAI22_X1 U20186 ( .A1(n17003), .A2(n17002), .B1(n17312), .B2(n9582), .ZN(
        P3_U2673) );
  NAND2_X1 U20187 ( .A1(n17005), .A2(n17004), .ZN(n17006) );
  XOR2_X1 U20188 ( .A(n17007), .B(n17006), .Z(n17316) );
  AOI22_X1 U20189 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17010), .B1(n17009), 
        .B2(n17008), .ZN(n17011) );
  OAI21_X1 U20190 ( .B1(n9582), .B2(n17316), .A(n17011), .ZN(P3_U2674) );
  OAI21_X1 U20191 ( .B1(n17014), .B2(n17013), .A(n17012), .ZN(n17326) );
  NAND3_X1 U20192 ( .A1(n17016), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n9582), .ZN(
        n17015) );
  OAI221_X1 U20193 ( .B1(n17016), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n9582), 
        .C2(n17326), .A(n17015), .ZN(P3_U2676) );
  AOI21_X1 U20194 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n9582), .A(n17024), .ZN(
        n17018) );
  XNOR2_X1 U20195 ( .A(n17017), .B(n17020), .ZN(n17331) );
  OAI22_X1 U20196 ( .A1(n17019), .A2(n17018), .B1(n9582), .B2(n17331), .ZN(
        P3_U2677) );
  AOI22_X1 U20197 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n9582), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n17032), .ZN(n17023) );
  OAI21_X1 U20198 ( .B1(n17022), .B2(n17021), .A(n17020), .ZN(n17336) );
  OAI22_X1 U20199 ( .A1(n17024), .A2(n17023), .B1(n9582), .B2(n17336), .ZN(
        P3_U2678) );
  XNOR2_X1 U20200 ( .A(n17025), .B(n17028), .ZN(n17341) );
  NAND3_X1 U20201 ( .A1(n17027), .A2(P3_EBX_REG_24__SCAN_IN), .A3(n9582), .ZN(
        n17026) );
  OAI221_X1 U20202 ( .B1(n17027), .B2(P3_EBX_REG_24__SCAN_IN), .C1(n9582), 
        .C2(n17341), .A(n17026), .ZN(P3_U2679) );
  AOI21_X1 U20203 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n9582), .A(n17046), .ZN(
        n17031) );
  OAI21_X1 U20204 ( .B1(n17030), .B2(n17029), .A(n17028), .ZN(n17346) );
  OAI22_X1 U20205 ( .A1(n17032), .A2(n17031), .B1(n9582), .B2(n17346), .ZN(
        P3_U2680) );
  AOI21_X1 U20206 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n9582), .A(n17033), .ZN(
        n17045) );
  AOI22_X1 U20207 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20208 ( .A1(n10178), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20209 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17034) );
  OAI211_X1 U20210 ( .C1(n9616), .C2(n17157), .A(n17035), .B(n17034), .ZN(
        n17041) );
  AOI22_X1 U20211 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20212 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20213 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17037) );
  NAND2_X1 U20214 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n17036) );
  NAND4_X1 U20215 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17040) );
  AOI211_X1 U20216 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17041), .B(n17040), .ZN(n17042) );
  OAI211_X1 U20217 ( .C1(n17224), .C2(n17269), .A(n17043), .B(n17042), .ZN(
        n17347) );
  INV_X1 U20218 ( .A(n17347), .ZN(n17044) );
  OAI22_X1 U20219 ( .A1(n17046), .A2(n17045), .B1(n17044), .B2(n9582), .ZN(
        P3_U2681) );
  OAI21_X1 U20220 ( .B1(n17047), .B2(n17090), .A(n9582), .ZN(n17075) );
  AOI22_X1 U20221 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20222 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20223 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17048) );
  OAI211_X1 U20224 ( .C1(n9616), .C2(n17050), .A(n17049), .B(n17048), .ZN(
        n17056) );
  AOI22_X1 U20225 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20226 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20227 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U20228 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n17051) );
  NAND4_X1 U20229 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n17051), .ZN(
        n17055) );
  AOI211_X1 U20230 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n17056), .B(n17055), .ZN(n17057) );
  OAI211_X1 U20231 ( .C1(n10102), .C2(n17059), .A(n17058), .B(n17057), .ZN(
        n17353) );
  NAND2_X1 U20232 ( .A1(n17295), .A2(n17353), .ZN(n17060) );
  OAI221_X1 U20233 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17062), .C1(n17061), 
        .C2(n17075), .A(n17060), .ZN(P3_U2682) );
  AOI22_X1 U20234 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17073) );
  INV_X1 U20235 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20236 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20237 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17063) );
  OAI211_X1 U20238 ( .C1(n9649), .C2(n17065), .A(n17064), .B(n17063), .ZN(
        n17071) );
  AOI22_X1 U20239 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20240 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20241 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17067) );
  NAND2_X1 U20242 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n17066) );
  NAND4_X1 U20243 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n17070) );
  AOI211_X1 U20244 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17071), .B(n17070), .ZN(n17072) );
  OAI211_X1 U20245 ( .C1(n17224), .C2(n17279), .A(n17073), .B(n17072), .ZN(
        n17358) );
  INV_X1 U20246 ( .A(n17358), .ZN(n17077) );
  NOR2_X1 U20247 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17074), .ZN(n17076) );
  OAI22_X1 U20248 ( .A1(n17077), .A2(n9582), .B1(n17076), .B2(n17075), .ZN(
        P3_U2683) );
  AOI22_X1 U20249 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17078) );
  OAI21_X1 U20250 ( .B1(n10102), .B2(n17079), .A(n17078), .ZN(n17089) );
  AOI22_X1 U20251 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20252 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17258), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17080) );
  OAI21_X1 U20253 ( .B1(n17224), .B2(n17282), .A(n17080), .ZN(n17084) );
  AOI22_X1 U20254 ( .A1(n10178), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20255 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17081) );
  OAI211_X1 U20256 ( .C1(n9616), .C2(n17189), .A(n17082), .B(n17081), .ZN(
        n17083) );
  AOI211_X1 U20257 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17084), .B(n17083), .ZN(n17085) );
  OAI211_X1 U20258 ( .C1(n9651), .C2(n17087), .A(n17086), .B(n17085), .ZN(
        n17088) );
  AOI211_X1 U20259 ( .C1(n17250), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17089), .B(n17088), .ZN(n17366) );
  OAI21_X1 U20260 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n9637), .A(n17090), .ZN(
        n17091) );
  AOI22_X1 U20261 ( .A1(n17295), .A2(n17366), .B1(n17091), .B2(n9582), .ZN(
        P3_U2684) );
  AOI21_X1 U20262 ( .B1(n20919), .B2(n17119), .A(n17295), .ZN(n17092) );
  INV_X1 U20263 ( .A(n17092), .ZN(n17105) );
  AOI22_X1 U20264 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20265 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20266 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17093) );
  OAI211_X1 U20267 ( .C1(n9616), .C2(n17095), .A(n17094), .B(n17093), .ZN(
        n17101) );
  AOI22_X1 U20268 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20269 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20270 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17097) );
  NAND2_X1 U20271 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n17096) );
  NAND4_X1 U20272 ( .A1(n17099), .A2(n17098), .A3(n17097), .A4(n17096), .ZN(
        n17100) );
  AOI211_X1 U20273 ( .C1(n10247), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17101), .B(n17100), .ZN(n17102) );
  OAI211_X1 U20274 ( .C1(n17224), .C2(n17289), .A(n17103), .B(n17102), .ZN(
        n17367) );
  INV_X1 U20275 ( .A(n17367), .ZN(n17104) );
  OAI22_X1 U20276 ( .A1(n9637), .A2(n17105), .B1(n17104), .B2(n9582), .ZN(
        P3_U2685) );
  OAI22_X1 U20277 ( .A1(n17224), .A2(n17290), .B1(n18597), .B2(n9722), .ZN(
        n17118) );
  AOI22_X1 U20278 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17250), .ZN(n17116) );
  AOI22_X1 U20279 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17171), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17211), .ZN(n17115) );
  OAI22_X1 U20280 ( .A1(n17107), .A2(n9616), .B1(n17199), .B2(n17106), .ZN(
        n17113) );
  AOI22_X1 U20281 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17251), .ZN(n17111) );
  AOI22_X1 U20282 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n9586), .ZN(n17110) );
  AOI22_X1 U20283 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17258), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17109) );
  NAND3_X1 U20284 ( .A1(n17111), .A2(n17110), .A3(n17109), .ZN(n17112) );
  AOI211_X1 U20285 ( .C1(n9610), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17113), .B(n17112), .ZN(n17114) );
  NAND3_X1 U20286 ( .A1(n17116), .A2(n17115), .A3(n17114), .ZN(n17117) );
  AOI211_X1 U20287 ( .C1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .C2(n10178), .A(
        n17118), .B(n17117), .ZN(n17377) );
  OAI21_X1 U20288 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17135), .A(n17119), .ZN(
        n17120) );
  AOI22_X1 U20289 ( .A1(n17295), .A2(n17377), .B1(n17120), .B2(n9582), .ZN(
        P3_U2686) );
  AOI21_X1 U20290 ( .B1(n17121), .B2(n17151), .A(n17295), .ZN(n17122) );
  INV_X1 U20291 ( .A(n17122), .ZN(n17134) );
  AOI22_X1 U20292 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17132) );
  INV_X1 U20293 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20933) );
  AOI22_X1 U20294 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20295 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17123) );
  OAI211_X1 U20296 ( .C1(n9649), .C2(n20933), .A(n17124), .B(n17123), .ZN(
        n17130) );
  AOI22_X1 U20297 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20298 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20299 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17126) );
  NAND2_X1 U20300 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n17125) );
  NAND4_X1 U20301 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17129) );
  AOI211_X1 U20302 ( .C1(n9622), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17130), .B(n17129), .ZN(n17131) );
  OAI211_X1 U20303 ( .C1(n17224), .C2(n20925), .A(n17132), .B(n17131), .ZN(
        n17378) );
  INV_X1 U20304 ( .A(n17378), .ZN(n17133) );
  OAI22_X1 U20305 ( .A1(n17135), .A2(n17134), .B1(n17133), .B2(n9582), .ZN(
        P3_U2687) );
  AOI22_X1 U20306 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17136) );
  OAI21_X1 U20307 ( .B1(n9612), .B2(n17264), .A(n17136), .ZN(n17150) );
  INV_X1 U20308 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20309 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20310 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17258), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17138) );
  OAI21_X1 U20311 ( .B1(n17199), .B2(n20949), .A(n17138), .ZN(n17144) );
  AOI22_X1 U20312 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17250), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20313 ( .A1(n10178), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17139) );
  OAI211_X1 U20314 ( .C1(n17142), .C2(n17141), .A(n17140), .B(n17139), .ZN(
        n17143) );
  AOI211_X1 U20315 ( .C1(n9622), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17144), .B(n17143), .ZN(n17145) );
  OAI211_X1 U20316 ( .C1(n17148), .C2(n17147), .A(n17146), .B(n17145), .ZN(
        n17149) );
  AOI211_X1 U20317 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n17150), .B(n17149), .ZN(n17388) );
  OAI21_X1 U20318 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17170), .A(n17151), .ZN(
        n17152) );
  AOI22_X1 U20319 ( .A1(n17295), .A2(n17388), .B1(n17152), .B2(n9582), .ZN(
        P3_U2688) );
  AOI21_X1 U20320 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n9582), .A(n17153), .ZN(
        n17169) );
  AOI22_X1 U20321 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U20322 ( .B1(n17156), .B2(n17155), .A(n17154), .ZN(n17168) );
  INV_X1 U20323 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20324 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10247), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17165) );
  OAI22_X1 U20325 ( .A1(n17224), .A2(n17158), .B1(n9722), .B2(n17157), .ZN(
        n17163) );
  AOI22_X1 U20326 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20327 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20328 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17159) );
  NAND3_X1 U20329 ( .A1(n17161), .A2(n17160), .A3(n17159), .ZN(n17162) );
  AOI211_X1 U20330 ( .C1(n17238), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17163), .B(n17162), .ZN(n17164) );
  OAI211_X1 U20331 ( .C1(n10102), .C2(n17166), .A(n17165), .B(n17164), .ZN(
        n17167) );
  AOI211_X1 U20332 ( .C1(n9576), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17168), .B(n17167), .ZN(n17393) );
  OAI22_X1 U20333 ( .A1(n17170), .A2(n17169), .B1(n17393), .B2(n9582), .ZN(
        P3_U2689) );
  AOI22_X1 U20334 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20335 ( .B1(n10102), .B2(n17173), .A(n17172), .ZN(n17184) );
  AOI22_X1 U20336 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20337 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17258), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17174) );
  INV_X1 U20338 ( .A(n17174), .ZN(n17179) );
  AOI22_X1 U20339 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20340 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20341 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17175) );
  NAND3_X1 U20342 ( .A1(n17177), .A2(n17176), .A3(n17175), .ZN(n17178) );
  AOI211_X1 U20343 ( .C1(n10142), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n17179), .B(n17178), .ZN(n17180) );
  OAI211_X1 U20344 ( .C1(n17224), .C2(n17182), .A(n17181), .B(n17180), .ZN(
        n17183) );
  AOI211_X1 U20345 ( .C1(n9586), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17184), .B(n17183), .ZN(n17399) );
  AOI21_X1 U20346 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n9582), .A(n17185), .ZN(
        n17186) );
  OAI22_X1 U20347 ( .A1(n17399), .A2(n9582), .B1(n17187), .B2(n17186), .ZN(
        P3_U2691) );
  AOI22_X1 U20348 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17188) );
  OAI21_X1 U20349 ( .B1(n9722), .B2(n17189), .A(n17188), .ZN(n17201) );
  INV_X1 U20350 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20351 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20352 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17190) );
  INV_X1 U20353 ( .A(n17190), .ZN(n17195) );
  AOI22_X1 U20354 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20355 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20356 ( .A1(n17258), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17191) );
  NAND3_X1 U20357 ( .A1(n17193), .A2(n17192), .A3(n17191), .ZN(n17194) );
  AOI211_X1 U20358 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n17195), .B(n17194), .ZN(n17196) );
  OAI211_X1 U20359 ( .C1(n17199), .C2(n17198), .A(n17197), .B(n17196), .ZN(
        n17200) );
  AOI211_X1 U20360 ( .C1(n17250), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17201), .B(n17200), .ZN(n17403) );
  OAI21_X1 U20361 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17204), .A(n17202), .ZN(
        n17203) );
  AOI22_X1 U20362 ( .A1(n17295), .A2(n17403), .B1(n17203), .B2(n9582), .ZN(
        P3_U2692) );
  AOI21_X1 U20363 ( .B1(n17205), .B2(n17239), .A(n17295), .ZN(n17221) );
  INV_X1 U20364 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18601) );
  AOI22_X1 U20365 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17220) );
  INV_X1 U20366 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20367 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20368 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17208) );
  OAI211_X1 U20369 ( .C1(n9616), .C2(n17210), .A(n17209), .B(n17208), .ZN(
        n17218) );
  AOI22_X1 U20370 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20371 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20372 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10247), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U20373 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n17213) );
  NAND4_X1 U20374 ( .A1(n17216), .A2(n17215), .A3(n17214), .A4(n17213), .ZN(
        n17217) );
  AOI211_X1 U20375 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17218), .B(n17217), .ZN(n17219) );
  OAI211_X1 U20376 ( .C1(n10131), .C2(n18601), .A(n17220), .B(n17219), .ZN(
        n17410) );
  AOI22_X1 U20377 ( .A1(n9817), .A2(n17221), .B1(n17410), .B2(n17295), .ZN(
        n17222) );
  INV_X1 U20378 ( .A(n17222), .ZN(P3_U2693) );
  AOI22_X1 U20379 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17251), .B1(
        n10178), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17223) );
  OAI21_X1 U20380 ( .B1(n10131), .B2(n18597), .A(n17223), .ZN(n17237) );
  INV_X1 U20381 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20382 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10142), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17233) );
  OAI22_X1 U20383 ( .A1(n17225), .A2(n9652), .B1(n17224), .B2(n20941), .ZN(
        n17231) );
  AOI22_X1 U20384 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9586), .ZN(n17229) );
  AOI22_X1 U20385 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17243), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20386 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9622), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17258), .ZN(n17227) );
  NAND3_X1 U20387 ( .A1(n17229), .A2(n17228), .A3(n17227), .ZN(n17230) );
  AOI211_X1 U20388 ( .C1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .C2(n10247), .A(
        n17231), .B(n17230), .ZN(n17232) );
  OAI211_X1 U20389 ( .C1(n10102), .C2(n17234), .A(n17233), .B(n17232), .ZN(
        n17236) );
  AOI211_X1 U20390 ( .C1(n17238), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n17237), .B(n17236), .ZN(n17416) );
  OAI21_X1 U20391 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17240), .A(n17239), .ZN(
        n17241) );
  AOI22_X1 U20392 ( .A1(n17295), .A2(n17416), .B1(n17241), .B2(n9582), .ZN(
        P3_U2694) );
  NAND3_X1 U20393 ( .A1(n17425), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n17271), .ZN(
        n17263) );
  NAND2_X1 U20394 ( .A1(n9582), .A2(n17242), .ZN(n17265) );
  AOI22_X1 U20395 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17260) );
  INV_X1 U20396 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20397 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20398 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17246) );
  OAI211_X1 U20399 ( .C1(n9616), .C2(n17248), .A(n17247), .B(n17246), .ZN(
        n17257) );
  AOI22_X1 U20400 ( .A1(n17250), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20401 ( .A1(n10178), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20402 ( .A1(n10142), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17253) );
  NAND2_X1 U20403 ( .A1(n10247), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n17252) );
  NAND4_X1 U20404 ( .A1(n17255), .A2(n17254), .A3(n17253), .A4(n17252), .ZN(
        n17256) );
  AOI211_X1 U20405 ( .C1(n17258), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17257), .B(n17256), .ZN(n17259) );
  OAI211_X1 U20406 ( .C1(n9652), .C2(n20973), .A(n17260), .B(n17259), .ZN(
        n17420) );
  NAND2_X1 U20407 ( .A1(n17295), .A2(n17420), .ZN(n17261) );
  OAI221_X1 U20408 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17263), .C1(n17262), 
        .C2(n17265), .A(n17261), .ZN(P3_U2695) );
  NOR2_X1 U20409 ( .A1(n17271), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17266) );
  OAI22_X1 U20410 ( .A1(n17266), .A2(n17265), .B1(n17264), .B2(n9582), .ZN(
        P3_U2696) );
  AOI21_X1 U20411 ( .B1(n17267), .B2(n17272), .A(n17295), .ZN(n17268) );
  INV_X1 U20412 ( .A(n17268), .ZN(n17270) );
  OAI22_X1 U20413 ( .A1(n17271), .A2(n17270), .B1(n17269), .B2(n9582), .ZN(
        P3_U2697) );
  OAI21_X1 U20414 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17273), .A(n17272), .ZN(
        n17274) );
  AOI22_X1 U20415 ( .A1(n17295), .A2(n17275), .B1(n17274), .B2(n9582), .ZN(
        P3_U2698) );
  INV_X1 U20416 ( .A(n17276), .ZN(n17277) );
  NAND2_X1 U20417 ( .A1(n17425), .A2(n17291), .ZN(n17297) );
  NOR2_X1 U20418 ( .A1(n17277), .A2(n17297), .ZN(n17287) );
  AND2_X1 U20419 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17287), .ZN(n17284) );
  AOI21_X1 U20420 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n9582), .A(n17284), .ZN(
        n17281) );
  NOR2_X1 U20421 ( .A1(n17278), .A2(n17297), .ZN(n17280) );
  OAI22_X1 U20422 ( .A1(n17281), .A2(n17280), .B1(n17279), .B2(n9582), .ZN(
        P3_U2699) );
  AOI21_X1 U20423 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n9582), .A(n17287), .ZN(
        n17283) );
  OAI22_X1 U20424 ( .A1(n17284), .A2(n17283), .B1(n17282), .B2(n9582), .ZN(
        P3_U2700) );
  AOI21_X1 U20425 ( .B1(n17425), .B2(n17285), .A(n17294), .ZN(n17286) );
  NOR2_X1 U20426 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17286), .ZN(n17288) );
  AOI211_X1 U20427 ( .C1(n17295), .C2(n17289), .A(n17288), .B(n17287), .ZN(
        P3_U2701) );
  OAI222_X1 U20428 ( .A1(n17297), .A2(n17293), .B1(n17292), .B2(n17291), .C1(
        n17290), .C2(n9582), .ZN(P3_U2702) );
  AOI22_X1 U20429 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17295), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17294), .ZN(n17296) );
  OAI21_X1 U20430 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17297), .A(n17296), .ZN(
        P3_U2703) );
  INV_X1 U20431 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17521) );
  INV_X1 U20432 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20910) );
  INV_X1 U20433 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20950) );
  NAND2_X1 U20434 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17454), .ZN(n17452) );
  NAND2_X1 U20435 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17426) );
  NAND4_X1 U20436 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17298) );
  NOR3_X2 U20437 ( .A1(n17452), .A2(n17426), .A3(n17298), .ZN(n17422) );
  NAND2_X1 U20438 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17422), .ZN(n17421) );
  INV_X1 U20439 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17546) );
  INV_X1 U20440 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17544) );
  NOR2_X1 U20441 ( .A1(n17546), .A2(n17544), .ZN(n17299) );
  NAND4_X1 U20442 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(n17299), .ZN(n17389) );
  NOR2_X2 U20443 ( .A1(n17421), .A2(n17389), .ZN(n17390) );
  NAND2_X1 U20444 ( .A1(n17390), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n17385) );
  NOR2_X2 U20445 ( .A1(n20950), .A2(n17385), .ZN(n17384) );
  INV_X1 U20446 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20983) );
  INV_X1 U20447 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17507) );
  NOR2_X1 U20448 ( .A1(n20983), .A2(n17507), .ZN(n17300) );
  NAND4_X1 U20449 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17300), .ZN(n17348) );
  INV_X1 U20450 ( .A(n17348), .ZN(n17301) );
  INV_X1 U20451 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17510) );
  NAND2_X1 U20452 ( .A1(n17301), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17302) );
  NAND2_X1 U20453 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17343), .ZN(n17342) );
  NAND2_X1 U20454 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17319), .ZN(n17313) );
  NAND2_X1 U20455 ( .A1(n17309), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17308) );
  NOR2_X2 U20456 ( .A1(n17303), .A2(n17453), .ZN(n17379) );
  OAI22_X1 U20457 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17304), .B1(n17414), 
        .B2(n17309), .ZN(n17305) );
  AOI22_X1 U20458 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17379), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17305), .ZN(n17306) );
  OAI21_X1 U20459 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17308), .A(n17306), .ZN(
        P3_U2704) );
  NAND2_X1 U20460 ( .A1(n17307), .A2(n17414), .ZN(n17383) );
  AOI22_X1 U20461 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17379), .ZN(n17311) );
  OAI211_X1 U20462 ( .C1(n17309), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17453), .B(
        n17308), .ZN(n17310) );
  OAI211_X1 U20463 ( .C1(n17312), .C2(n17447), .A(n17311), .B(n17310), .ZN(
        P3_U2705) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17379), .ZN(n17315) );
  OAI211_X1 U20465 ( .C1(n17319), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17453), .B(
        n17313), .ZN(n17314) );
  OAI211_X1 U20466 ( .C1(n17447), .C2(n17316), .A(n17315), .B(n17314), .ZN(
        P3_U2706) );
  AOI22_X1 U20467 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17372), .B1(n17317), .B2(
        n17450), .ZN(n17318) );
  INV_X1 U20468 ( .A(n17318), .ZN(n17321) );
  AOI211_X1 U20469 ( .C1(n17521), .C2(n17323), .A(n17319), .B(n17414), .ZN(
        n17320) );
  AOI211_X1 U20470 ( .C1(n17379), .C2(BUF2_REG_28__SCAN_IN), .A(n17321), .B(
        n17320), .ZN(n17322) );
  INV_X1 U20471 ( .A(n17322), .ZN(P3_U2707) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17379), .ZN(n17325) );
  OAI211_X1 U20473 ( .C1(n17327), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17453), .B(
        n17323), .ZN(n17324) );
  OAI211_X1 U20474 ( .C1(n17326), .C2(n17447), .A(n17325), .B(n17324), .ZN(
        P3_U2708) );
  AOI22_X1 U20475 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17379), .ZN(n17330) );
  AOI211_X1 U20476 ( .C1(n20910), .C2(n17332), .A(n17327), .B(n17414), .ZN(
        n17328) );
  INV_X1 U20477 ( .A(n17328), .ZN(n17329) );
  OAI211_X1 U20478 ( .C1(n17331), .C2(n17447), .A(n17330), .B(n17329), .ZN(
        P3_U2709) );
  AOI22_X1 U20479 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17379), .ZN(n17335) );
  OAI211_X1 U20480 ( .C1(n17333), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17453), .B(
        n17332), .ZN(n17334) );
  OAI211_X1 U20481 ( .C1(n17336), .C2(n17447), .A(n17335), .B(n17334), .ZN(
        P3_U2710) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17379), .ZN(n17340) );
  OAI211_X1 U20483 ( .C1(n17338), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17453), .B(
        n17337), .ZN(n17339) );
  OAI211_X1 U20484 ( .C1(n17341), .C2(n17447), .A(n17340), .B(n17339), .ZN(
        P3_U2711) );
  AOI22_X1 U20485 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17379), .ZN(n17345) );
  OAI211_X1 U20486 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17343), .A(n17453), .B(
        n17342), .ZN(n17344) );
  OAI211_X1 U20487 ( .C1(n17346), .C2(n17447), .A(n17345), .B(n17344), .ZN(
        P3_U2712) );
  AOI22_X1 U20488 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17379), .B1(n17450), .B2(
        n17347), .ZN(n17352) );
  OR3_X1 U20489 ( .A1(n18299), .A2(n17380), .A3(n17348), .ZN(n17350) );
  INV_X1 U20490 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17505) );
  NAND2_X1 U20491 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17374), .ZN(n17373) );
  NAND2_X1 U20492 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17362), .ZN(n17359) );
  AND2_X1 U20493 ( .A1(n17453), .A2(n17359), .ZN(n17355) );
  NOR2_X1 U20494 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17359), .ZN(n17354) );
  NOR2_X1 U20495 ( .A1(n17355), .A2(n17354), .ZN(n17349) );
  MUX2_X1 U20496 ( .A(n17350), .B(n17349), .S(P3_EAX_REG_22__SCAN_IN), .Z(
        n17351) );
  OAI211_X1 U20497 ( .C1(n18296), .C2(n17383), .A(n17352), .B(n17351), .ZN(
        P3_U2713) );
  AOI22_X1 U20498 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17379), .B1(n17450), .B2(
        n17353), .ZN(n17357) );
  AOI21_X1 U20499 ( .B1(n17355), .B2(P3_EAX_REG_21__SCAN_IN), .A(n17354), .ZN(
        n17356) );
  OAI211_X1 U20500 ( .C1(n18292), .C2(n17383), .A(n17357), .B(n17356), .ZN(
        P3_U2714) );
  INV_X1 U20501 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18288) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17379), .B1(n17450), .B2(
        n17358), .ZN(n17361) );
  OAI211_X1 U20503 ( .C1(n17362), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17453), .B(
        n17359), .ZN(n17360) );
  OAI211_X1 U20504 ( .C1(n17383), .C2(n18288), .A(n17361), .B(n17360), .ZN(
        P3_U2715) );
  AOI22_X1 U20505 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17379), .ZN(n17365) );
  AOI211_X1 U20506 ( .C1(n17505), .C2(n17368), .A(n17362), .B(n17414), .ZN(
        n17363) );
  INV_X1 U20507 ( .A(n17363), .ZN(n17364) );
  OAI211_X1 U20508 ( .C1(n17366), .C2(n17447), .A(n17365), .B(n17364), .ZN(
        P3_U2716) );
  INV_X1 U20509 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U20510 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17379), .B1(n17450), .B2(
        n17367), .ZN(n17371) );
  OAI211_X1 U20511 ( .C1(n17369), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17453), .B(
        n17368), .ZN(n17370) );
  OAI211_X1 U20512 ( .C1(n17383), .C2(n18281), .A(n17371), .B(n17370), .ZN(
        P3_U2717) );
  AOI22_X1 U20513 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17372), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17379), .ZN(n17376) );
  OAI211_X1 U20514 ( .C1(n17374), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17453), .B(
        n17373), .ZN(n17375) );
  OAI211_X1 U20515 ( .C1(n17377), .C2(n17447), .A(n17376), .B(n17375), .ZN(
        P3_U2718) );
  INV_X1 U20516 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U20517 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17379), .B1(n17450), .B2(
        n17378), .ZN(n17382) );
  OAI211_X1 U20518 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17384), .A(n17453), .B(
        n17380), .ZN(n17381) );
  OAI211_X1 U20519 ( .C1(n17383), .C2(n18270), .A(n17382), .B(n17381), .ZN(
        P3_U2719) );
  AOI211_X1 U20520 ( .C1(n20950), .C2(n17385), .A(n17414), .B(n17384), .ZN(
        n17386) );
  AOI21_X1 U20521 ( .B1(n17451), .B2(BUF2_REG_15__SCAN_IN), .A(n17386), .ZN(
        n17387) );
  OAI21_X1 U20522 ( .B1(n17388), .B2(n17447), .A(n17387), .ZN(P3_U2720) );
  AND2_X1 U20523 ( .A1(n17425), .A2(n17422), .ZN(n17429) );
  NAND2_X1 U20524 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17429), .ZN(n17413) );
  NOR2_X1 U20525 ( .A1(n17389), .A2(n17413), .ZN(n17395) );
  INV_X1 U20526 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U20527 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17451), .B1(n17395), .B2(
        n17557), .ZN(n17392) );
  OR3_X1 U20528 ( .A1(n17557), .A2(n17414), .A3(n17390), .ZN(n17391) );
  OAI211_X1 U20529 ( .C1(n17393), .C2(n17447), .A(n17392), .B(n17391), .ZN(
        P3_U2721) );
  INV_X1 U20530 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17397) );
  INV_X1 U20531 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17551) );
  NOR2_X1 U20532 ( .A1(n17544), .A2(n17413), .ZN(n17418) );
  INV_X1 U20533 ( .A(n17418), .ZN(n17408) );
  NAND2_X1 U20534 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17407), .ZN(n17398) );
  NOR2_X1 U20535 ( .A1(n17551), .A2(n17398), .ZN(n17401) );
  AOI21_X1 U20536 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17453), .A(n17401), .ZN(
        n17396) );
  OAI222_X1 U20537 ( .A1(n17448), .A2(n17397), .B1(n17396), .B2(n17395), .C1(
        n17447), .C2(n17394), .ZN(P3_U2722) );
  INV_X1 U20538 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17402) );
  INV_X1 U20539 ( .A(n17398), .ZN(n17405) );
  AOI21_X1 U20540 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17453), .A(n17405), .ZN(
        n17400) );
  OAI222_X1 U20541 ( .A1(n17448), .A2(n17402), .B1(n17401), .B2(n17400), .C1(
        n17447), .C2(n17399), .ZN(P3_U2723) );
  INV_X1 U20542 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17406) );
  AOI21_X1 U20543 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17453), .A(n17407), .ZN(
        n17404) );
  OAI222_X1 U20544 ( .A1(n17448), .A2(n17406), .B1(n17405), .B2(n17404), .C1(
        n17447), .C2(n17403), .ZN(P3_U2724) );
  INV_X1 U20545 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17412) );
  AOI211_X1 U20546 ( .C1(n17546), .C2(n17408), .A(n17414), .B(n17407), .ZN(
        n17409) );
  AOI21_X1 U20547 ( .B1(n17450), .B2(n17410), .A(n17409), .ZN(n17411) );
  OAI21_X1 U20548 ( .B1(n17412), .B2(n17448), .A(n17411), .ZN(P3_U2725) );
  INV_X1 U20549 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17419) );
  OAI21_X1 U20550 ( .B1(n17544), .B2(n17414), .A(n17413), .ZN(n17415) );
  INV_X1 U20551 ( .A(n17415), .ZN(n17417) );
  OAI222_X1 U20552 ( .A1(n17448), .A2(n17419), .B1(n17418), .B2(n17417), .C1(
        n17447), .C2(n17416), .ZN(P3_U2726) );
  AOI22_X1 U20553 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17451), .B1(n17450), .B2(
        n17420), .ZN(n17424) );
  OAI211_X1 U20554 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17422), .A(n17453), .B(
        n17421), .ZN(n17423) );
  NAND2_X1 U20555 ( .A1(n17424), .A2(n17423), .ZN(P3_U2727) );
  INV_X1 U20556 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18301) );
  INV_X1 U20557 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17533) );
  INV_X1 U20558 ( .A(n17452), .ZN(n17443) );
  NAND3_X1 U20559 ( .A1(n17425), .A2(n17443), .A3(P3_EAX_REG_2__SCAN_IN), .ZN(
        n17442) );
  NOR2_X1 U20560 ( .A1(n17533), .A2(n17442), .ZN(n17437) );
  NAND2_X1 U20561 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17437), .ZN(n17433) );
  NOR2_X1 U20562 ( .A1(n17426), .A2(n17433), .ZN(n17431) );
  AOI21_X1 U20563 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17453), .A(n17431), .ZN(
        n17428) );
  OAI222_X1 U20564 ( .A1(n17448), .A2(n18301), .B1(n17429), .B2(n17428), .C1(
        n17447), .C2(n17427), .ZN(P3_U2728) );
  INV_X1 U20565 ( .A(n17433), .ZN(n17440) );
  AOI22_X1 U20566 ( .A1(n17440), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17453), .ZN(n17432) );
  OAI222_X1 U20567 ( .A1(n17448), .A2(n18296), .B1(n17432), .B2(n17431), .C1(
        n17447), .C2(n17430), .ZN(P3_U2729) );
  AOI21_X1 U20568 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17453), .A(n17440), .ZN(
        n17436) );
  INV_X1 U20569 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17536) );
  NOR2_X1 U20570 ( .A1(n17536), .A2(n17433), .ZN(n17435) );
  OAI222_X1 U20571 ( .A1(n17448), .A2(n18292), .B1(n17436), .B2(n17435), .C1(
        n17447), .C2(n17434), .ZN(P3_U2730) );
  AOI21_X1 U20572 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17453), .A(n17437), .ZN(
        n17439) );
  OAI222_X1 U20573 ( .A1(n18288), .A2(n17448), .B1(n17440), .B2(n17439), .C1(
        n17447), .C2(n17438), .ZN(P3_U2731) );
  NAND2_X1 U20574 ( .A1(n17453), .A2(n17442), .ZN(n17445) );
  AOI22_X1 U20575 ( .A1(n17451), .A2(BUF2_REG_3__SCAN_IN), .B1(n17450), .B2(
        n10128), .ZN(n17441) );
  OAI221_X1 U20576 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17442), .C1(n17533), 
        .C2(n17445), .A(n17441), .ZN(P3_U2732) );
  NOR2_X1 U20577 ( .A1(n17443), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n17444) );
  OAI222_X1 U20578 ( .A1(n17448), .A2(n18281), .B1(n17447), .B2(n17446), .C1(
        n17445), .C2(n17444), .ZN(P3_U2733) );
  AOI22_X1 U20579 ( .A1(n17451), .A2(BUF2_REG_1__SCAN_IN), .B1(n17450), .B2(
        n17449), .ZN(n17456) );
  OAI211_X1 U20580 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17454), .A(n17453), .B(
        n17452), .ZN(n17455) );
  NAND2_X1 U20581 ( .A1(n17456), .A2(n17455), .ZN(P3_U2734) );
  NOR2_X4 U20582 ( .A1(n17492), .A2(n17476), .ZN(n17485) );
  AND2_X1 U20583 ( .A1(n17485), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20584 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20585 ( .A1(n17492), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20586 ( .B1(n17525), .B2(n17474), .A(n17459), .ZN(P3_U2737) );
  INV_X1 U20587 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17523) );
  AOI22_X1 U20588 ( .A1(n17492), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20589 ( .B1(n17523), .B2(n17474), .A(n17460), .ZN(P3_U2738) );
  AOI22_X1 U20590 ( .A1(n17492), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U20591 ( .B1(n17521), .B2(n17474), .A(n17461), .ZN(P3_U2739) );
  INV_X1 U20592 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20593 ( .A1(n17492), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U20594 ( .B1(n17519), .B2(n17474), .A(n17462), .ZN(P3_U2740) );
  AOI22_X1 U20595 ( .A1(n17492), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20596 ( .B1(n20910), .B2(n17474), .A(n17463), .ZN(P3_U2741) );
  INV_X1 U20597 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17516) );
  AOI22_X1 U20598 ( .A1(n17492), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20599 ( .B1(n17516), .B2(n17474), .A(n17464), .ZN(P3_U2742) );
  INV_X1 U20600 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17514) );
  INV_X2 U20601 ( .A(n18911), .ZN(n17492) );
  AOI22_X1 U20602 ( .A1(n17492), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20603 ( .B1(n17514), .B2(n17474), .A(n17465), .ZN(P3_U2743) );
  INV_X1 U20604 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20605 ( .A1(n17492), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20606 ( .B1(n17512), .B2(n17474), .A(n17466), .ZN(P3_U2744) );
  AOI22_X1 U20607 ( .A1(n17492), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20608 ( .B1(n17510), .B2(n17474), .A(n17467), .ZN(P3_U2745) );
  AOI22_X1 U20609 ( .A1(n17492), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U20610 ( .B1(n20983), .B2(n17474), .A(n17468), .ZN(P3_U2746) );
  AOI22_X1 U20611 ( .A1(n17492), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20612 ( .B1(n17507), .B2(n17474), .A(n17469), .ZN(P3_U2747) );
  AOI22_X1 U20613 ( .A1(n17492), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17470) );
  OAI21_X1 U20614 ( .B1(n17505), .B2(n17474), .A(n17470), .ZN(P3_U2748) );
  INV_X1 U20615 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20616 ( .A1(n17492), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20617 ( .B1(n17503), .B2(n17474), .A(n17471), .ZN(P3_U2749) );
  INV_X1 U20618 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17501) );
  AOI22_X1 U20619 ( .A1(n17492), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17472) );
  OAI21_X1 U20620 ( .B1(n17501), .B2(n17474), .A(n17472), .ZN(P3_U2750) );
  INV_X1 U20621 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U20622 ( .A1(n17492), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U20623 ( .B1(n17499), .B2(n17474), .A(n17473), .ZN(P3_U2751) );
  INV_X1 U20624 ( .A(P3_LWORD_REG_15__SCAN_IN), .ZN(n20944) );
  AOI22_X1 U20625 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17476), .B1(n17485), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20626 ( .B1(n18911), .B2(n20944), .A(n17475), .ZN(P3_U2752) );
  AOI22_X1 U20627 ( .A1(n17492), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20628 ( .B1(n17557), .B2(n17494), .A(n17477), .ZN(P3_U2753) );
  INV_X1 U20629 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20630 ( .A1(n17492), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U20631 ( .B1(n17554), .B2(n17494), .A(n17478), .ZN(P3_U2754) );
  AOI22_X1 U20632 ( .A1(n17492), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17479) );
  OAI21_X1 U20633 ( .B1(n17551), .B2(n17494), .A(n17479), .ZN(P3_U2755) );
  INV_X1 U20634 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U20635 ( .A1(n17492), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17480) );
  OAI21_X1 U20636 ( .B1(n17548), .B2(n17494), .A(n17480), .ZN(P3_U2756) );
  AOI22_X1 U20637 ( .A1(n17492), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20638 ( .B1(n17546), .B2(n17494), .A(n17481), .ZN(P3_U2757) );
  AOI22_X1 U20639 ( .A1(n17492), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17482) );
  OAI21_X1 U20640 ( .B1(n17544), .B2(n17494), .A(n17482), .ZN(P3_U2758) );
  INV_X1 U20641 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U20642 ( .A1(n17492), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20643 ( .B1(n17542), .B2(n17494), .A(n17483), .ZN(P3_U2759) );
  INV_X1 U20644 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17540) );
  AOI22_X1 U20645 ( .A1(n17492), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17484) );
  OAI21_X1 U20646 ( .B1(n17540), .B2(n17494), .A(n17484), .ZN(P3_U2760) );
  INV_X1 U20647 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U20648 ( .A1(n17492), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17486) );
  OAI21_X1 U20649 ( .B1(n17538), .B2(n17494), .A(n17486), .ZN(P3_U2761) );
  AOI22_X1 U20650 ( .A1(n17492), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17487) );
  OAI21_X1 U20651 ( .B1(n17536), .B2(n17494), .A(n17487), .ZN(P3_U2762) );
  INV_X1 U20652 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20875) );
  AOI22_X1 U20653 ( .A1(n17492), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17488) );
  OAI21_X1 U20654 ( .B1(n20875), .B2(n17494), .A(n17488), .ZN(P3_U2763) );
  AOI22_X1 U20655 ( .A1(n17492), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17489) );
  OAI21_X1 U20656 ( .B1(n17533), .B2(n17494), .A(n17489), .ZN(P3_U2764) );
  INV_X1 U20657 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20658 ( .A1(n17492), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17490) );
  OAI21_X1 U20659 ( .B1(n17531), .B2(n17494), .A(n17490), .ZN(P3_U2765) );
  INV_X1 U20660 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17529) );
  AOI22_X1 U20661 ( .A1(n17492), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U20662 ( .B1(n17529), .B2(n17494), .A(n17491), .ZN(P3_U2766) );
  AOI22_X1 U20663 ( .A1(n17492), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17485), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U20664 ( .B1(n17527), .B2(n17494), .A(n17493), .ZN(P3_U2767) );
  NOR2_X1 U20665 ( .A1(n18277), .A2(n17495), .ZN(n18751) );
  NAND2_X2 U20666 ( .A1(n17496), .A2(n18751), .ZN(n17556) );
  AOI22_X1 U20667 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17560), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17559), .ZN(n17498) );
  OAI21_X1 U20668 ( .B1(n17499), .B2(n17556), .A(n17498), .ZN(P3_U2768) );
  AOI22_X1 U20669 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17560), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17559), .ZN(n17500) );
  OAI21_X1 U20670 ( .B1(n17501), .B2(n17556), .A(n17500), .ZN(P3_U2769) );
  AOI22_X1 U20671 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17560), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17559), .ZN(n17502) );
  OAI21_X1 U20672 ( .B1(n17503), .B2(n17556), .A(n17502), .ZN(P3_U2770) );
  AOI22_X1 U20673 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17559), .ZN(n17504) );
  OAI21_X1 U20674 ( .B1(n17505), .B2(n17556), .A(n17504), .ZN(P3_U2771) );
  AOI22_X1 U20675 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17559), .ZN(n17506) );
  OAI21_X1 U20676 ( .B1(n17507), .B2(n17556), .A(n17506), .ZN(P3_U2772) );
  AOI22_X1 U20677 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17559), .ZN(n17508) );
  OAI21_X1 U20678 ( .B1(n20983), .B2(n17556), .A(n17508), .ZN(P3_U2773) );
  AOI22_X1 U20679 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17559), .ZN(n17509) );
  OAI21_X1 U20680 ( .B1(n17510), .B2(n17556), .A(n17509), .ZN(P3_U2774) );
  AOI22_X1 U20681 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17559), .ZN(n17511) );
  OAI21_X1 U20682 ( .B1(n17512), .B2(n17556), .A(n17511), .ZN(P3_U2775) );
  AOI22_X1 U20683 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17559), .ZN(n17513) );
  OAI21_X1 U20684 ( .B1(n17514), .B2(n17556), .A(n17513), .ZN(P3_U2776) );
  AOI22_X1 U20685 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17559), .ZN(n17515) );
  OAI21_X1 U20686 ( .B1(n17516), .B2(n17556), .A(n17515), .ZN(P3_U2777) );
  AOI22_X1 U20687 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17559), .ZN(n17517) );
  OAI21_X1 U20688 ( .B1(n20910), .B2(n17556), .A(n17517), .ZN(P3_U2778) );
  AOI22_X1 U20689 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17559), .ZN(n17518) );
  OAI21_X1 U20690 ( .B1(n17519), .B2(n17556), .A(n17518), .ZN(P3_U2779) );
  AOI22_X1 U20691 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17560), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17559), .ZN(n17520) );
  OAI21_X1 U20692 ( .B1(n17521), .B2(n17556), .A(n17520), .ZN(P3_U2780) );
  AOI22_X1 U20693 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17560), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17559), .ZN(n17522) );
  OAI21_X1 U20694 ( .B1(n17523), .B2(n17556), .A(n17522), .ZN(P3_U2781) );
  AOI22_X1 U20695 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17560), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17559), .ZN(n17524) );
  OAI21_X1 U20696 ( .B1(n17525), .B2(n17556), .A(n17524), .ZN(P3_U2782) );
  AOI22_X1 U20697 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17559), .ZN(n17526) );
  OAI21_X1 U20698 ( .B1(n17527), .B2(n17556), .A(n17526), .ZN(P3_U2783) );
  AOI22_X1 U20699 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17559), .ZN(n17528) );
  OAI21_X1 U20700 ( .B1(n17529), .B2(n17556), .A(n17528), .ZN(P3_U2784) );
  AOI22_X1 U20701 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17552), .ZN(n17530) );
  OAI21_X1 U20702 ( .B1(n17531), .B2(n17556), .A(n17530), .ZN(P3_U2785) );
  AOI22_X1 U20703 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17552), .ZN(n17532) );
  OAI21_X1 U20704 ( .B1(n17533), .B2(n17556), .A(n17532), .ZN(P3_U2786) );
  AOI22_X1 U20705 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17552), .ZN(n17534) );
  OAI21_X1 U20706 ( .B1(n20875), .B2(n17556), .A(n17534), .ZN(P3_U2787) );
  AOI22_X1 U20707 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17552), .ZN(n17535) );
  OAI21_X1 U20708 ( .B1(n17536), .B2(n17556), .A(n17535), .ZN(P3_U2788) );
  AOI22_X1 U20709 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17552), .ZN(n17537) );
  OAI21_X1 U20710 ( .B1(n17538), .B2(n17556), .A(n17537), .ZN(P3_U2789) );
  AOI22_X1 U20711 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17552), .ZN(n17539) );
  OAI21_X1 U20712 ( .B1(n17540), .B2(n17556), .A(n17539), .ZN(P3_U2790) );
  AOI22_X1 U20713 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17552), .ZN(n17541) );
  OAI21_X1 U20714 ( .B1(n17542), .B2(n17556), .A(n17541), .ZN(P3_U2791) );
  AOI22_X1 U20715 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17552), .ZN(n17543) );
  OAI21_X1 U20716 ( .B1(n17544), .B2(n17556), .A(n17543), .ZN(P3_U2792) );
  AOI22_X1 U20717 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17559), .ZN(n17545) );
  OAI21_X1 U20718 ( .B1(n17546), .B2(n17556), .A(n17545), .ZN(P3_U2793) );
  AOI22_X1 U20719 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17552), .ZN(n17547) );
  OAI21_X1 U20720 ( .B1(n17548), .B2(n17556), .A(n17547), .ZN(P3_U2794) );
  AOI22_X1 U20721 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17559), .ZN(n17550) );
  OAI21_X1 U20722 ( .B1(n17551), .B2(n17556), .A(n17550), .ZN(P3_U2795) );
  AOI22_X1 U20723 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17552), .ZN(n17553) );
  OAI21_X1 U20724 ( .B1(n17554), .B2(n17556), .A(n17553), .ZN(P3_U2796) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17560), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17559), .ZN(n17555) );
  OAI21_X1 U20726 ( .B1(n17557), .B2(n17556), .A(n17555), .ZN(P3_U2797) );
  AOI222_X1 U20727 ( .A1(n17560), .A2(BUF2_REG_15__SCAN_IN), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17559), .C1(P3_EAX_REG_15__SCAN_IN), 
        .C2(n17558), .ZN(n17561) );
  INV_X1 U20728 ( .A(n17561), .ZN(P3_U2798) );
  NAND2_X1 U20729 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17562), .ZN(
        n17577) );
  NOR2_X1 U20730 ( .A1(n17911), .A2(n17791), .ZN(n17670) );
  NOR3_X1 U20731 ( .A1(n17670), .A2(n17563), .A3(n17562), .ZN(n17570) );
  OAI211_X1 U20732 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17565), .B(n17564), .ZN(n17567) );
  OAI211_X1 U20733 ( .C1(n17780), .C2(n17568), .A(n17567), .B(n17566), .ZN(
        n17569) );
  AOI211_X1 U20734 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17571), .A(
        n17570), .B(n17569), .ZN(n17576) );
  OAI211_X1 U20735 ( .C1(n17574), .C2(n17573), .A(n17834), .B(n17572), .ZN(
        n17575) );
  OAI211_X1 U20736 ( .C1(n17578), .C2(n17577), .A(n17576), .B(n17575), .ZN(
        P3_U2802) );
  AOI21_X1 U20737 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17580), .A(
        n17579), .ZN(n17948) );
  NAND3_X1 U20738 ( .A1(n18648), .A2(n17582), .A3(n17581), .ZN(n17584) );
  AOI21_X1 U20739 ( .B1(n17585), .B2(n17584), .A(n17583), .ZN(n17588) );
  AOI21_X1 U20740 ( .B1(n17780), .B2(n17702), .A(n17586), .ZN(n17587) );
  AOI211_X1 U20741 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n9587), .A(n17588), .B(
        n17587), .ZN(n17592) );
  NOR3_X1 U20742 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n20894), .A3(
        n17950), .ZN(n17942) );
  NAND2_X1 U20743 ( .A1(n17589), .A2(n17708), .ZN(n17618) );
  INV_X1 U20744 ( .A(n17618), .ZN(n17631) );
  AOI22_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17590), .B1(
        n17942), .B2(n17631), .ZN(n17591) );
  OAI211_X1 U20746 ( .C1(n17948), .C2(n17807), .A(n17592), .B(n17591), .ZN(
        P3_U2804) );
  INV_X1 U20747 ( .A(n18065), .ZN(n17644) );
  NOR2_X1 U20748 ( .A1(n17644), .A2(n17600), .ZN(n17963) );
  NAND2_X1 U20749 ( .A1(n17963), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17593) );
  XOR2_X1 U20750 ( .A(n17593), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17961) );
  OAI21_X1 U20751 ( .B1(n17623), .B2(n18771), .A(n17922), .ZN(n17594) );
  AOI21_X1 U20752 ( .B1(n18648), .B2(n17595), .A(n17594), .ZN(n17628) );
  OAI21_X1 U20753 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17702), .A(
        n17628), .ZN(n17612) );
  NOR2_X1 U20754 ( .A1(n18253), .A2(n18836), .ZN(n17956) );
  OAI21_X1 U20755 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17596), .ZN(n17597) );
  OAI22_X1 U20756 ( .A1(n17780), .A2(n17598), .B1(n17609), .B2(n17597), .ZN(
        n17599) );
  AOI211_X1 U20757 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17612), .A(
        n17956), .B(n17599), .ZN(n17606) );
  INV_X1 U20758 ( .A(n18064), .ZN(n17645) );
  NOR2_X1 U20759 ( .A1(n17645), .A2(n17600), .ZN(n17962) );
  NAND2_X1 U20760 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17962), .ZN(
        n17601) );
  XOR2_X1 U20761 ( .A(n20894), .B(n17601), .Z(n17958) );
  OAI21_X1 U20762 ( .B1(n17729), .B2(n17603), .A(n17602), .ZN(n17604) );
  XOR2_X1 U20763 ( .A(n17604), .B(n20894), .Z(n17957) );
  AOI22_X1 U20764 ( .A1(n9574), .A2(n17958), .B1(n17834), .B2(n17957), .ZN(
        n17605) );
  OAI211_X1 U20765 ( .C1(n17837), .C2(n17961), .A(n17606), .B(n17605), .ZN(
        P3_U2805) );
  NAND2_X1 U20766 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17974), .ZN(
        n17617) );
  NOR2_X1 U20767 ( .A1(n18253), .A2(n18834), .ZN(n17611) );
  INV_X1 U20768 ( .A(n17607), .ZN(n17608) );
  OAI22_X1 U20769 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17609), .B1(
        n17608), .B2(n17780), .ZN(n17610) );
  AOI211_X1 U20770 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17612), .A(
        n17611), .B(n17610), .ZN(n17616) );
  OAI22_X1 U20771 ( .A1(n17963), .A2(n17837), .B1(n17962), .B2(n17926), .ZN(
        n17630) );
  OAI21_X1 U20772 ( .B1(n17614), .B2(n17974), .A(n17613), .ZN(n17973) );
  AOI22_X1 U20773 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17630), .B1(
        n17834), .B2(n17973), .ZN(n17615) );
  OAI211_X1 U20774 ( .C1(n17618), .C2(n17617), .A(n17616), .B(n17615), .ZN(
        P3_U2806) );
  OAI22_X1 U20775 ( .A1(n17833), .A2(n17649), .B1(n17647), .B2(n17619), .ZN(
        n17620) );
  NOR2_X1 U20776 ( .A1(n17620), .A2(n17671), .ZN(n17621) );
  XOR2_X1 U20777 ( .A(n17621), .B(n17967), .Z(n17981) );
  AOI21_X1 U20778 ( .B1(n17622), .B2(n18648), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17627) );
  NOR2_X1 U20779 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17702), .ZN(
        n17624) );
  AOI22_X1 U20780 ( .A1(n17758), .A2(n17625), .B1(n17624), .B2(n17623), .ZN(
        n17626) );
  NAND2_X1 U20781 ( .A1(n9587), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17980) );
  OAI211_X1 U20782 ( .C1(n17628), .C2(n17627), .A(n17626), .B(n17980), .ZN(
        n17629) );
  AOI221_X1 U20783 ( .B1(n17631), .B2(n17967), .C1(n17630), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17629), .ZN(n17632) );
  OAI21_X1 U20784 ( .B1(n17807), .B2(n17981), .A(n17632), .ZN(P3_U2807) );
  INV_X1 U20785 ( .A(n17676), .ZN(n17881) );
  OAI21_X1 U20786 ( .B1(n17635), .B2(n17881), .A(n17922), .ZN(n17633) );
  AOI21_X1 U20787 ( .B1(n17755), .B2(n17634), .A(n17633), .ZN(n17666) );
  OAI21_X1 U20788 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17702), .A(
        n17666), .ZN(n17656) );
  NAND2_X1 U20789 ( .A1(n17635), .A2(n17763), .ZN(n17654) );
  AOI221_X1 U20790 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17637), .C2(n17636), .A(
        n17654), .ZN(n17641) );
  INV_X1 U20791 ( .A(n17638), .ZN(n17639) );
  NAND2_X1 U20792 ( .A1(n9587), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17996) );
  OAI21_X1 U20793 ( .B1(n17639), .B2(n17780), .A(n17996), .ZN(n17640) );
  AOI211_X1 U20794 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17656), .A(
        n17641), .B(n17640), .ZN(n17652) );
  INV_X1 U20795 ( .A(n17642), .ZN(n18037) );
  NAND2_X1 U20796 ( .A1(n18037), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17989) );
  NOR2_X1 U20797 ( .A1(n17643), .A2(n17989), .ZN(n17986) );
  AOI22_X1 U20798 ( .A1(n9574), .A2(n17645), .B1(n17791), .B2(n17644), .ZN(
        n17722) );
  OAI21_X1 U20799 ( .B1(n17670), .B2(n17986), .A(n17722), .ZN(n17661) );
  INV_X1 U20800 ( .A(n17671), .ZN(n17646) );
  OAI221_X1 U20801 ( .B1(n17647), .B2(n17994), .C1(n17647), .C2(n17657), .A(
        n17646), .ZN(n17648) );
  XOR2_X1 U20802 ( .A(n17649), .B(n17648), .Z(n17995) );
  AOI22_X1 U20803 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17661), .B1(
        n17834), .B2(n17995), .ZN(n17651) );
  NAND3_X1 U20804 ( .A1(n17708), .A2(n17986), .A3(n17649), .ZN(n17650) );
  NAND3_X1 U20805 ( .A1(n17652), .A2(n17651), .A3(n17650), .ZN(P3_U2808) );
  INV_X1 U20806 ( .A(n18005), .ZN(n17990) );
  NAND2_X1 U20807 ( .A1(n17990), .A2(n20969), .ZN(n18011) );
  NOR2_X1 U20808 ( .A1(n18253), .A2(n18829), .ZN(n18008) );
  OAI22_X1 U20809 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17654), .B1(
        n17653), .B2(n17780), .ZN(n17655) );
  AOI211_X1 U20810 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17656), .A(
        n18008), .B(n17655), .ZN(n17663) );
  NAND3_X1 U20811 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17833), .A3(
        n17657), .ZN(n17685) );
  INV_X1 U20812 ( .A(n17658), .ZN(n17697) );
  OAI22_X1 U20813 ( .A1(n18005), .A2(n17685), .B1(n17659), .B2(n17697), .ZN(
        n17660) );
  XNOR2_X1 U20814 ( .A(n20969), .B(n17660), .ZN(n18009) );
  AOI22_X1 U20815 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17661), .B1(
        n17834), .B2(n18009), .ZN(n17662) );
  OAI211_X1 U20816 ( .C1(n18011), .C2(n17690), .A(n17663), .B(n17662), .ZN(
        P3_U2809) );
  NAND2_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17984), .ZN(
        n18023) );
  INV_X1 U20818 ( .A(n17702), .ZN(n17668) );
  NOR2_X1 U20819 ( .A1(n18587), .A2(n17679), .ZN(n17703) );
  AOI21_X1 U20820 ( .B1(n17664), .B2(n17703), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17665) );
  NAND2_X1 U20821 ( .A1(n9587), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18020) );
  OAI21_X1 U20822 ( .B1(n17666), .B2(n17665), .A(n18020), .ZN(n17667) );
  AOI221_X1 U20823 ( .B1(n17758), .B2(n17669), .C1(n17668), .C2(n17669), .A(
        n17667), .ZN(n17674) );
  INV_X1 U20824 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20929) );
  NOR2_X1 U20825 ( .A1(n20929), .A2(n17989), .ZN(n18014) );
  OAI21_X1 U20826 ( .B1(n17670), .B2(n18014), .A(n17722), .ZN(n17687) );
  AOI221_X1 U20827 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17685), 
        .C1(n20929), .C2(n17696), .A(n17671), .ZN(n17672) );
  XOR2_X1 U20828 ( .A(n17672), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18018) );
  AOI22_X1 U20829 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17687), .B1(
        n17834), .B2(n18018), .ZN(n17673) );
  OAI211_X1 U20830 ( .C1(n17690), .C2(n18023), .A(n17674), .B(n17673), .ZN(
        P3_U2810) );
  OR2_X1 U20831 ( .A1(n17679), .A2(n17678), .ZN(n17675) );
  AOI21_X1 U20832 ( .B1(n17676), .B2(n17675), .A(n17893), .ZN(n17705) );
  OAI21_X1 U20833 ( .B1(n17677), .B2(n18771), .A(n17705), .ZN(n17694) );
  INV_X1 U20834 ( .A(n17763), .ZN(n17680) );
  NOR3_X1 U20835 ( .A1(n17680), .A2(n17679), .A3(n17678), .ZN(n17695) );
  OAI211_X1 U20836 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17695), .B(n17681), .ZN(n17682) );
  NAND2_X1 U20837 ( .A1(n9587), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18026) );
  OAI211_X1 U20838 ( .C1(n17780), .C2(n17683), .A(n17682), .B(n18026), .ZN(
        n17684) );
  AOI21_X1 U20839 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17694), .A(
        n17684), .ZN(n17689) );
  OAI21_X1 U20840 ( .B1(n17696), .B2(n17697), .A(n17685), .ZN(n17686) );
  XOR2_X1 U20841 ( .A(n17686), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18025) );
  AOI22_X1 U20842 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17687), .B1(
        n17834), .B2(n18025), .ZN(n17688) );
  OAI211_X1 U20843 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17690), .A(
        n17689), .B(n17688), .ZN(P3_U2811) );
  NAND2_X1 U20844 ( .A1(n17691), .A2(n18001), .ZN(n18044) );
  INV_X1 U20845 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20902) );
  NAND2_X1 U20846 ( .A1(n9587), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18042) );
  OAI21_X1 U20847 ( .B1(n17780), .B2(n17692), .A(n18042), .ZN(n17693) );
  AOI221_X1 U20848 ( .B1(n17695), .B2(n20902), .C1(n17694), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17693), .ZN(n17700) );
  OAI21_X1 U20849 ( .B1(n18001), .B2(n17729), .A(n17696), .ZN(n17698) );
  XOR2_X1 U20850 ( .A(n17698), .B(n17697), .Z(n18040) );
  OAI211_X1 U20851 ( .C1(n17820), .C2(n18044), .A(n17700), .B(n17699), .ZN(
        P3_U2812) );
  AOI21_X1 U20852 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17701), .A(
        n9701), .ZN(n18051) );
  NOR2_X1 U20853 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17703), .ZN(
        n17704) );
  NAND2_X1 U20854 ( .A1(n9587), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18049) );
  OAI21_X1 U20855 ( .B1(n17705), .B2(n17704), .A(n18049), .ZN(n17706) );
  AOI21_X1 U20856 ( .B1(n17707), .B2(n17914), .A(n17706), .ZN(n17711) );
  NOR2_X1 U20857 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18059), .ZN(
        n18047) );
  AOI22_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17709), .B1(
        n17708), .B2(n18047), .ZN(n17710) );
  OAI211_X1 U20859 ( .C1(n18051), .C2(n17807), .A(n17711), .B(n17710), .ZN(
        P3_U2813) );
  NAND2_X1 U20860 ( .A1(n17833), .A2(n18126), .ZN(n17782) );
  INV_X1 U20861 ( .A(n17782), .ZN(n17808) );
  AOI22_X1 U20862 ( .A1(n17808), .A2(n17988), .B1(n17712), .B2(n17729), .ZN(
        n17713) );
  XOR2_X1 U20863 ( .A(n18059), .B(n17713), .Z(n18061) );
  OAI21_X1 U20864 ( .B1(n17731), .B2(n17881), .A(n17922), .ZN(n17744) );
  AOI21_X1 U20865 ( .B1(n17755), .B2(n17714), .A(n17744), .ZN(n17732) );
  INV_X1 U20866 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17716) );
  OAI22_X1 U20867 ( .A1(n17732), .A2(n17716), .B1(n17780), .B2(n17715), .ZN(
        n17720) );
  NOR2_X1 U20868 ( .A1(n17733), .A2(n17716), .ZN(n17718) );
  OAI211_X1 U20869 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17731), .B(n17763), .ZN(n17717) );
  OAI22_X1 U20870 ( .A1(n17718), .A2(n17717), .B1(n18253), .B2(n18819), .ZN(
        n17719) );
  AOI211_X1 U20871 ( .C1(n17834), .C2(n18061), .A(n17720), .B(n17719), .ZN(
        n17721) );
  OAI221_X1 U20872 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17723), 
        .C1(n18059), .C2(n17722), .A(n17721), .ZN(P3_U2814) );
  NOR2_X1 U20873 ( .A1(n17833), .A2(n17724), .ZN(n17809) );
  NAND2_X1 U20874 ( .A1(n17725), .A2(n17809), .ZN(n17781) );
  NOR2_X1 U20875 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17781), .ZN(
        n17772) );
  INV_X1 U20876 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18096) );
  NOR4_X1 U20877 ( .A1(n18114), .A2(n18106), .A3(n18096), .A4(n17726), .ZN(
        n17727) );
  AOI21_X1 U20878 ( .B1(n17772), .B2(n18106), .A(n17727), .ZN(n17728) );
  AOI221_X1 U20879 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18113), 
        .C1(n17729), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17728), .ZN(
        n17730) );
  XOR2_X1 U20880 ( .A(n18078), .B(n17730), .Z(n18071) );
  NAND2_X1 U20881 ( .A1(n17731), .A2(n17763), .ZN(n17734) );
  NAND2_X1 U20882 ( .A1(n9587), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18076) );
  OAI221_X1 U20883 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17734), .C1(
        n17733), .C2(n17732), .A(n18076), .ZN(n17735) );
  AOI21_X1 U20884 ( .B1(n17758), .B2(n17736), .A(n17735), .ZN(n17740) );
  NOR2_X1 U20885 ( .A1(n18065), .A2(n17837), .ZN(n17738) );
  NAND2_X1 U20886 ( .A1(n18078), .A2(n17749), .ZN(n18069) );
  NOR2_X1 U20887 ( .A1(n18064), .A2(n17926), .ZN(n17737) );
  NAND2_X1 U20888 ( .A1(n17747), .A2(n18078), .ZN(n18074) );
  AOI22_X1 U20889 ( .A1(n17738), .A2(n18069), .B1(n17737), .B2(n18074), .ZN(
        n17739) );
  OAI211_X1 U20890 ( .C1(n17807), .C2(n18071), .A(n17740), .B(n17739), .ZN(
        P3_U2815) );
  OAI21_X1 U20891 ( .B1(n17742), .B2(n18587), .A(n17741), .ZN(n17743) );
  AOI22_X1 U20892 ( .A1(n9587), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17744), 
        .B2(n17743), .ZN(n17752) );
  NOR3_X1 U20893 ( .A1(n18114), .A2(n18113), .A3(n17782), .ZN(n17759) );
  AND2_X1 U20894 ( .A1(n18113), .A2(n17772), .ZN(n17745) );
  AOI22_X1 U20895 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17759), .B1(
        n17745), .B2(n18106), .ZN(n17746) );
  XOR2_X1 U20896 ( .A(n18096), .B(n17746), .Z(n18093) );
  OAI21_X1 U20897 ( .B1(n17748), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17747), .ZN(n18091) );
  OAI221_X1 U20898 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18079), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18126), .A(n17749), .ZN(
        n18090) );
  OAI22_X1 U20899 ( .A1(n17926), .A2(n18091), .B1(n17837), .B2(n18090), .ZN(
        n17750) );
  AOI21_X1 U20900 ( .B1(n17834), .B2(n18093), .A(n17750), .ZN(n17751) );
  OAI211_X1 U20901 ( .C1(n17905), .C2(n17753), .A(n17752), .B(n17751), .ZN(
        P3_U2816) );
  AOI21_X1 U20902 ( .B1(n17755), .B2(n17754), .A(n17893), .ZN(n17756) );
  OAI21_X1 U20903 ( .B1(n17786), .B2(n17881), .A(n17756), .ZN(n17769) );
  AOI22_X1 U20904 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17769), .B1(
        n17758), .B2(n17757), .ZN(n17767) );
  AOI21_X1 U20905 ( .B1(n17772), .B2(n18113), .A(n17759), .ZN(n17760) );
  XOR2_X1 U20906 ( .A(n18106), .B(n17760), .Z(n18109) );
  NAND2_X1 U20907 ( .A1(n18083), .A2(n18106), .ZN(n18112) );
  NOR2_X1 U20908 ( .A1(n18123), .A2(n18082), .ZN(n18105) );
  INV_X1 U20909 ( .A(n18105), .ZN(n17761) );
  NAND2_X1 U20910 ( .A1(n18083), .A2(n18126), .ZN(n18100) );
  AOI22_X1 U20911 ( .A1(n9574), .A2(n17761), .B1(n17791), .B2(n18100), .ZN(
        n17774) );
  OAI22_X1 U20912 ( .A1(n17820), .A2(n18112), .B1(n17774), .B2(n18106), .ZN(
        n17762) );
  AOI21_X1 U20913 ( .B1(n17834), .B2(n18109), .A(n17762), .ZN(n17766) );
  NAND2_X1 U20914 ( .A1(n9587), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18110) );
  AND2_X1 U20915 ( .A1(n17763), .A2(n17786), .ZN(n17771) );
  NAND2_X1 U20916 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17764) );
  OAI211_X1 U20917 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17771), .B(n17764), .ZN(n17765) );
  NAND4_X1 U20918 ( .A1(n17767), .A2(n17766), .A3(n18110), .A4(n17765), .ZN(
        P3_U2817) );
  NOR2_X1 U20919 ( .A1(n18253), .A2(n18812), .ZN(n17768) );
  AOI221_X1 U20920 ( .B1(n17771), .B2(n17770), .C1(n17769), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17768), .ZN(n17778) );
  NOR2_X1 U20921 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17820), .ZN(
        n17776) );
  INV_X1 U20922 ( .A(n18114), .ZN(n18099) );
  AOI21_X1 U20923 ( .B1(n18099), .B2(n17808), .A(n17772), .ZN(n17773) );
  XNOR2_X1 U20924 ( .A(n18113), .B(n17773), .ZN(n18120) );
  OAI22_X1 U20925 ( .A1(n18120), .A2(n17807), .B1(n17774), .B2(n18113), .ZN(
        n17775) );
  AOI21_X1 U20926 ( .B1(n17776), .B2(n18099), .A(n17775), .ZN(n17777) );
  OAI211_X1 U20927 ( .C1(n17780), .C2(n17779), .A(n17778), .B(n17777), .ZN(
        P3_U2818) );
  INV_X1 U20928 ( .A(n17790), .ZN(n18129) );
  OR2_X1 U20929 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18134) );
  OAI21_X1 U20930 ( .B1(n17782), .B2(n18129), .A(n17781), .ZN(n17783) );
  XOR2_X1 U20931 ( .A(n17783), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18121) );
  INV_X1 U20932 ( .A(n17919), .ZN(n17812) );
  NAND3_X1 U20933 ( .A1(n18648), .A2(n17855), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17811) );
  NOR2_X1 U20934 ( .A1(n17784), .A2(n17811), .ZN(n17800) );
  AOI21_X1 U20935 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17812), .A(
        n17800), .ZN(n17785) );
  AOI21_X1 U20936 ( .B1(n17786), .B2(n18648), .A(n17785), .ZN(n17789) );
  INV_X1 U20937 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18809) );
  OAI22_X1 U20938 ( .A1(n17905), .A2(n17787), .B1(n18253), .B2(n18809), .ZN(
        n17788) );
  AOI211_X1 U20939 ( .C1(n17834), .C2(n18121), .A(n17789), .B(n17788), .ZN(
        n17794) );
  NOR2_X1 U20940 ( .A1(n17790), .A2(n17820), .ZN(n17803) );
  AOI22_X1 U20941 ( .A1(n17792), .A2(n17791), .B1(n17911), .B2(n18123), .ZN(
        n17819) );
  INV_X1 U20942 ( .A(n17819), .ZN(n17804) );
  OAI21_X1 U20943 ( .B1(n17803), .B2(n17804), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17793) );
  OAI211_X1 U20944 ( .C1(n17820), .C2(n18134), .A(n17794), .B(n17793), .ZN(
        P3_U2819) );
  AOI22_X1 U20945 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17808), .B1(
        n17809), .B2(n18155), .ZN(n17795) );
  XNOR2_X1 U20946 ( .A(n18138), .B(n17795), .ZN(n18145) );
  NOR3_X1 U20947 ( .A1(n17797), .A2(n17796), .A3(n17811), .ZN(n17815) );
  AOI21_X1 U20948 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17812), .A(
        n17815), .ZN(n17799) );
  OAI22_X1 U20949 ( .A1(n17800), .A2(n17799), .B1(n17905), .B2(n17798), .ZN(
        n17801) );
  AOI21_X1 U20950 ( .B1(n9587), .B2(P3_REIP_REG_10__SCAN_IN), .A(n17801), .ZN(
        n17806) );
  AOI22_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17804), .B1(
        n17803), .B2(n17802), .ZN(n17805) );
  OAI211_X1 U20952 ( .C1(n18145), .C2(n17807), .A(n17806), .B(n17805), .ZN(
        P3_U2820) );
  NOR2_X1 U20953 ( .A1(n17809), .A2(n17808), .ZN(n17810) );
  XOR2_X1 U20954 ( .A(n17810), .B(n18155), .Z(n18152) );
  NOR2_X1 U20955 ( .A1(n18253), .A2(n18805), .ZN(n17817) );
  INV_X1 U20956 ( .A(n17811), .ZN(n17843) );
  AOI22_X1 U20957 ( .A1(n17821), .A2(n17843), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17812), .ZN(n17814) );
  OAI22_X1 U20958 ( .A1(n17815), .A2(n17814), .B1(n17905), .B2(n17813), .ZN(
        n17816) );
  AOI211_X1 U20959 ( .C1(n17834), .C2(n18152), .A(n17817), .B(n17816), .ZN(
        n17818) );
  OAI221_X1 U20960 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17820), .C1(
        n18155), .C2(n17819), .A(n17818), .ZN(P3_U2821) );
  INV_X1 U20961 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17824) );
  NAND2_X1 U20962 ( .A1(n17823), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17822) );
  AOI211_X1 U20963 ( .C1(n17824), .C2(n17822), .A(n17821), .B(n18587), .ZN(
        n17828) );
  OAI21_X1 U20964 ( .B1(n17881), .B2(n17823), .A(n17922), .ZN(n17841) );
  INV_X1 U20965 ( .A(n17841), .ZN(n17825) );
  OAI22_X1 U20966 ( .A1(n17905), .A2(n17826), .B1(n17825), .B2(n17824), .ZN(
        n17827) );
  AOI211_X1 U20967 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n9587), .A(n17828), .B(
        n17827), .ZN(n17836) );
  AOI21_X1 U20968 ( .B1(n17830), .B2(n18165), .A(n17829), .ZN(n18169) );
  OAI21_X1 U20969 ( .B1(n17833), .B2(n17832), .A(n17831), .ZN(n18167) );
  AOI22_X1 U20970 ( .A1(n17911), .A2(n18169), .B1(n17834), .B2(n18167), .ZN(
        n17835) );
  OAI211_X1 U20971 ( .C1(n17837), .C2(n18173), .A(n17836), .B(n17835), .ZN(
        P3_U2822) );
  NAND2_X1 U20972 ( .A1(n17839), .A2(n17838), .ZN(n17840) );
  XOR2_X1 U20973 ( .A(n17840), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18183) );
  NOR2_X1 U20974 ( .A1(n18253), .A2(n18801), .ZN(n18174) );
  AOI221_X1 U20975 ( .B1(n17843), .B2(n17842), .C1(n17841), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18174), .ZN(n17848) );
  AOI21_X1 U20976 ( .B1(n18177), .B2(n17845), .A(n17844), .ZN(n18179) );
  AOI22_X1 U20977 ( .A1(n17915), .A2(n18179), .B1(n17846), .B2(n17914), .ZN(
        n17847) );
  OAI211_X1 U20978 ( .C1(n17926), .C2(n18183), .A(n17848), .B(n17847), .ZN(
        P3_U2823) );
  AOI21_X1 U20979 ( .B1(n17850), .B2(n17849), .A(n9717), .ZN(n18187) );
  NAND2_X1 U20980 ( .A1(n18648), .A2(n17855), .ZN(n17851) );
  OAI22_X1 U20981 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17851), .B1(
        n18253), .B2(n18799), .ZN(n17852) );
  AOI21_X1 U20982 ( .B1(n17915), .B2(n18187), .A(n17852), .ZN(n17857) );
  AOI21_X1 U20983 ( .B1(n17854), .B2(n18178), .A(n17853), .ZN(n18188) );
  AOI21_X1 U20984 ( .B1(n17855), .B2(n18648), .A(n17919), .ZN(n17868) );
  AOI22_X1 U20985 ( .A1(n9574), .A2(n18188), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17868), .ZN(n17856) );
  OAI211_X1 U20986 ( .C1(n17905), .C2(n17858), .A(n17857), .B(n17856), .ZN(
        P3_U2824) );
  AOI21_X1 U20987 ( .B1(n17861), .B2(n17860), .A(n17859), .ZN(n18194) );
  AOI22_X1 U20988 ( .A1(n17915), .A2(n18194), .B1(n9587), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17870) );
  AOI21_X1 U20989 ( .B1(n17864), .B2(n17863), .A(n17862), .ZN(n18193) );
  OAI21_X1 U20990 ( .B1(n17893), .B2(n17866), .A(n17865), .ZN(n17867) );
  AOI22_X1 U20991 ( .A1(n17911), .A2(n18193), .B1(n17868), .B2(n17867), .ZN(
        n17869) );
  OAI211_X1 U20992 ( .C1(n17905), .C2(n17871), .A(n17870), .B(n17869), .ZN(
        P3_U2825) );
  OAI21_X1 U20993 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n17875) );
  XOR2_X1 U20994 ( .A(n17875), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18209) );
  OAI22_X1 U20995 ( .A1(n17926), .A2(n18209), .B1(n18587), .B2(n17876), .ZN(
        n17877) );
  AOI21_X1 U20996 ( .B1(n9587), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17877), .ZN(
        n17883) );
  AOI21_X1 U20997 ( .B1(n17880), .B2(n17879), .A(n17878), .ZN(n18199) );
  OAI21_X1 U20998 ( .B1(n9905), .B2(n17881), .A(n17922), .ZN(n17895) );
  AOI22_X1 U20999 ( .A1(n17915), .A2(n18199), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17895), .ZN(n17882) );
  OAI211_X1 U21000 ( .C1(n17905), .C2(n17884), .A(n17883), .B(n17882), .ZN(
        P3_U2826) );
  OAI21_X1 U21001 ( .B1(n17887), .B2(n17886), .A(n17885), .ZN(n17888) );
  XOR2_X1 U21002 ( .A(n17888), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18219) );
  AOI21_X1 U21003 ( .B1(n17891), .B2(n17890), .A(n17889), .ZN(n18216) );
  AOI22_X1 U21004 ( .A1(n9574), .A2(n18216), .B1(n9587), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17898) );
  OAI21_X1 U21005 ( .B1(n17893), .B2(n17909), .A(n17892), .ZN(n17894) );
  AOI22_X1 U21006 ( .A1(n17896), .A2(n17914), .B1(n17895), .B2(n17894), .ZN(
        n17897) );
  OAI211_X1 U21007 ( .C1(n17925), .C2(n18219), .A(n17898), .B(n17897), .ZN(
        P3_U2827) );
  AOI21_X1 U21008 ( .B1(n17901), .B2(n17900), .A(n17899), .ZN(n18231) );
  NAND2_X1 U21009 ( .A1(n9587), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18233) );
  INV_X1 U21010 ( .A(n18233), .ZN(n17907) );
  XNOR2_X1 U21011 ( .A(n17903), .B(n17902), .ZN(n18230) );
  OAI22_X1 U21012 ( .A1(n17905), .A2(n17904), .B1(n17925), .B2(n18230), .ZN(
        n17906) );
  AOI211_X1 U21013 ( .C1(n17911), .C2(n18231), .A(n17907), .B(n17906), .ZN(
        n17908) );
  OAI221_X1 U21014 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18587), .C1(
        n17909), .C2(n17922), .A(n17908), .ZN(P3_U2828) );
  NOR2_X1 U21015 ( .A1(n17921), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17910) );
  XNOR2_X1 U21016 ( .A(n17910), .B(n17913), .ZN(n18243) );
  AOI22_X1 U21017 ( .A1(n17911), .A2(n18243), .B1(n9587), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17917) );
  AOI21_X1 U21018 ( .B1(n17913), .B2(n17920), .A(n17912), .ZN(n18236) );
  AOI22_X1 U21019 ( .A1(n17915), .A2(n18236), .B1(n17918), .B2(n17914), .ZN(
        n17916) );
  OAI211_X1 U21020 ( .C1(n17919), .C2(n17918), .A(n17917), .B(n17916), .ZN(
        P3_U2829) );
  OAI21_X1 U21021 ( .B1(n17921), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17920), .ZN(n18249) );
  INV_X1 U21022 ( .A(n18249), .ZN(n18251) );
  NAND3_X1 U21023 ( .A1(n18871), .A2(n18771), .A3(n17922), .ZN(n17923) );
  AOI22_X1 U21024 ( .A1(n9587), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17923), .ZN(n17924) );
  OAI221_X1 U21025 ( .B1(n18251), .B2(n17926), .C1(n18249), .C2(n17925), .A(
        n17924), .ZN(P3_U2830) );
  OAI21_X1 U21026 ( .B1(n18254), .B2(n17928), .A(n17927), .ZN(n17937) );
  NOR2_X1 U21027 ( .A1(n18224), .A2(n17929), .ZN(n17964) );
  AOI21_X1 U21028 ( .B1(n17952), .B2(n17964), .A(n18222), .ZN(n17949) );
  OAI22_X1 U21029 ( .A1(n18716), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18723), .B2(n17930), .ZN(n17934) );
  OAI22_X1 U21030 ( .A1(n17932), .A2(n18104), .B1(n17931), .B2(n18125), .ZN(
        n17933) );
  NOR4_X1 U21031 ( .A1(n17935), .A2(n17949), .A3(n17934), .A4(n17933), .ZN(
        n17941) );
  OAI211_X1 U21032 ( .C1(n18716), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17941), .ZN(n17936) );
  AOI22_X1 U21033 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18211), .B1(
        n17937), .B2(n17936), .ZN(n17939) );
  OAI211_X1 U21034 ( .C1(n17940), .C2(n18144), .A(n17939), .B(n17938), .ZN(
        P3_U2835) );
  INV_X1 U21035 ( .A(n17941), .ZN(n17943) );
  AOI22_X1 U21036 ( .A1(n17943), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n17978), .B2(n17942), .ZN(n17944) );
  INV_X1 U21037 ( .A(n17944), .ZN(n17945) );
  AOI22_X1 U21038 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18211), .B1(
        n18238), .B2(n17945), .ZN(n17947) );
  NAND2_X1 U21039 ( .A1(n9587), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17946) );
  OAI211_X1 U21040 ( .C1(n17948), .C2(n18144), .A(n17947), .B(n17946), .ZN(
        P3_U2836) );
  AOI221_X1 U21041 ( .B1(n17950), .B2(n18707), .C1(n17968), .C2(n18707), .A(
        n17949), .ZN(n17954) );
  NAND2_X1 U21042 ( .A1(n17952), .A2(n17951), .ZN(n17953) );
  AOI221_X1 U21043 ( .B1(n17954), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17953), .C2(n20894), .A(n18254), .ZN(n17955) );
  AOI211_X1 U21044 ( .C1(n18211), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17956), .B(n17955), .ZN(n17960) );
  AOI22_X1 U21045 ( .A1(n18250), .A2(n17958), .B1(n9572), .B2(n17957), .ZN(
        n17959) );
  OAI211_X1 U21046 ( .C1(n18172), .C2(n17961), .A(n17960), .B(n17959), .ZN(
        P3_U2837) );
  INV_X1 U21047 ( .A(n17962), .ZN(n17966) );
  OAI22_X1 U21048 ( .A1(n18222), .A2(n17964), .B1(n17963), .B2(n18125), .ZN(
        n17965) );
  AOI211_X1 U21049 ( .C1(n18705), .C2(n17966), .A(n18211), .B(n17965), .ZN(
        n17970) );
  AOI21_X1 U21050 ( .B1(n18707), .B2(n17968), .A(n17967), .ZN(n17969) );
  AOI21_X1 U21051 ( .B1(n17970), .B2(n17969), .A(n9587), .ZN(n17977) );
  INV_X1 U21052 ( .A(n18162), .ZN(n17971) );
  AOI21_X1 U21053 ( .B1(n17971), .B2(n17970), .A(n17974), .ZN(n17972) );
  AOI22_X1 U21054 ( .A1(n9572), .A2(n17973), .B1(n17977), .B2(n17972), .ZN(
        n17976) );
  NAND4_X1 U21055 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18238), .A3(
        n17978), .A4(n17974), .ZN(n17975) );
  OAI211_X1 U21056 ( .C1(n18834), .C2(n18253), .A(n17976), .B(n17975), .ZN(
        P3_U2838) );
  OAI221_X1 U21057 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17978), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18239), .A(n17977), .ZN(
        n17979) );
  OAI211_X1 U21058 ( .C1(n17981), .C2(n18144), .A(n17980), .B(n17979), .ZN(
        P3_U2839) );
  OAI22_X1 U21059 ( .A1(n18064), .A2(n18104), .B1(n18065), .B2(n18125), .ZN(
        n18002) );
  NAND2_X1 U21060 ( .A1(n18104), .A2(n18125), .ZN(n18128) );
  INV_X1 U21061 ( .A(n18128), .ZN(n18036) );
  OAI21_X1 U21062 ( .B1(n18001), .B2(n18039), .A(n18707), .ZN(n17982) );
  OAI221_X1 U21063 ( .B1(n18716), .B2(n17983), .C1(n18716), .C2(n18014), .A(
        n17982), .ZN(n18016) );
  AOI21_X1 U21064 ( .B1(n18725), .B2(n17984), .A(n18016), .ZN(n17985) );
  OAI21_X1 U21065 ( .B1(n17986), .B2(n18036), .A(n17985), .ZN(n18004) );
  OAI22_X1 U21066 ( .A1(n18057), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18723), .B2(n17987), .ZN(n17992) );
  NAND2_X1 U21067 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18135), .ZN(
        n18080) );
  INV_X1 U21068 ( .A(n18080), .ZN(n18149) );
  NAND2_X1 U21069 ( .A1(n17988), .A2(n18149), .ZN(n18053) );
  OAI21_X1 U21070 ( .B1(n17989), .B2(n18053), .A(n18081), .ZN(n18003) );
  OAI211_X1 U21071 ( .C1(n17990), .C2(n18736), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18003), .ZN(n17991) );
  NOR4_X1 U21072 ( .A1(n18002), .A2(n18004), .A3(n17992), .A4(n17991), .ZN(
        n17999) );
  INV_X1 U21073 ( .A(n18000), .ZN(n17993) );
  OAI221_X1 U21074 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17994), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17993), .A(n18238), .ZN(
        n17998) );
  AOI22_X1 U21075 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18211), .B1(
        n9572), .B2(n17995), .ZN(n17997) );
  OAI211_X1 U21076 ( .C1(n17999), .C2(n17998), .A(n17997), .B(n17996), .ZN(
        P3_U2840) );
  NOR3_X1 U21077 ( .A1(n18001), .A2(n18254), .A3(n18000), .ZN(n18024) );
  INV_X1 U21078 ( .A(n18024), .ZN(n18022) );
  NAND2_X1 U21079 ( .A1(n18723), .A2(n18736), .ZN(n18237) );
  NOR2_X1 U21080 ( .A1(n18254), .A2(n18002), .ZN(n18033) );
  NAND2_X1 U21081 ( .A1(n18033), .A2(n18003), .ZN(n18012) );
  AOI211_X1 U21082 ( .C1(n18005), .C2(n18237), .A(n18004), .B(n18012), .ZN(
        n18006) );
  NOR3_X1 U21083 ( .A1(n9587), .A2(n18006), .A3(n20969), .ZN(n18007) );
  AOI211_X1 U21084 ( .C1(n9572), .C2(n18009), .A(n18008), .B(n18007), .ZN(
        n18010) );
  OAI21_X1 U21085 ( .B1(n18011), .B2(n18022), .A(n18010), .ZN(P3_U2841) );
  NAND3_X1 U21086 ( .A1(n20929), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18237), 
        .ZN(n18017) );
  INV_X1 U21087 ( .A(n18012), .ZN(n18013) );
  OAI21_X1 U21088 ( .B1(n18014), .B2(n18036), .A(n18013), .ZN(n18015) );
  OAI21_X1 U21089 ( .B1(n18016), .B2(n18015), .A(n18253), .ZN(n18028) );
  NAND2_X1 U21090 ( .A1(n18017), .A2(n18028), .ZN(n18019) );
  AOI22_X1 U21091 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18019), .B1(
        n9572), .B2(n18018), .ZN(n18021) );
  OAI211_X1 U21092 ( .C1(n18023), .C2(n18022), .A(n18021), .B(n18020), .ZN(
        P3_U2842) );
  AOI22_X1 U21093 ( .A1(n9572), .A2(n18025), .B1(n18024), .B2(n20929), .ZN(
        n18027) );
  OAI211_X1 U21094 ( .C1(n20929), .C2(n18028), .A(n18027), .B(n18026), .ZN(
        P3_U2843) );
  OAI22_X1 U21095 ( .A1(n18227), .A2(n18736), .B1(n18202), .B2(n18220), .ZN(
        n18192) );
  INV_X1 U21096 ( .A(n18192), .ZN(n18214) );
  NOR2_X1 U21097 ( .A1(n18029), .A2(n18214), .ZN(n18184) );
  NAND2_X1 U21098 ( .A1(n18030), .A2(n18184), .ZN(n18087) );
  INV_X1 U21099 ( .A(n18087), .ZN(n18032) );
  INV_X1 U21100 ( .A(n18033), .ZN(n18058) );
  NOR3_X1 U21101 ( .A1(n18224), .A2(n18059), .A3(n18034), .ZN(n18035) );
  OAI22_X1 U21102 ( .A1(n18037), .A2(n18036), .B1(n18222), .B2(n18035), .ZN(
        n18038) );
  AOI211_X1 U21103 ( .C1(n18707), .C2(n18039), .A(n18058), .B(n18038), .ZN(
        n18045) );
  AOI221_X1 U21104 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18045), 
        .C1(n18222), .C2(n18045), .A(n9587), .ZN(n18041) );
  AOI22_X1 U21105 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18041), .B1(
        n9572), .B2(n18040), .ZN(n18043) );
  OAI211_X1 U21106 ( .C1(n18156), .C2(n18044), .A(n18043), .B(n18042), .ZN(
        P3_U2844) );
  NOR2_X1 U21107 ( .A1(n9587), .A2(n18045), .ZN(n18048) );
  NOR2_X1 U21108 ( .A1(n18046), .A2(n18156), .ZN(n18060) );
  AOI22_X1 U21109 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18048), .B1(
        n18060), .B2(n18047), .ZN(n18050) );
  OAI211_X1 U21110 ( .C1(n18051), .C2(n18144), .A(n18050), .B(n18049), .ZN(
        P3_U2845) );
  NOR2_X1 U21111 ( .A1(n18052), .A2(n18736), .ZN(n18122) );
  AOI21_X1 U21112 ( .B1(n18157), .B2(n18161), .A(n18716), .ZN(n18151) );
  AOI211_X1 U21113 ( .C1(n18725), .C2(n18165), .A(n18122), .B(n18151), .ZN(
        n18055) );
  OAI21_X1 U21114 ( .B1(n18078), .B2(n18081), .A(n18053), .ZN(n18054) );
  OAI211_X1 U21115 ( .C1(n18057), .C2(n18056), .A(n18055), .B(n18054), .ZN(
        n18068) );
  OAI221_X1 U21116 ( .B1(n18058), .B2(n18162), .C1(n18058), .C2(n18068), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U21117 ( .A1(n9572), .A2(n18061), .B1(n18060), .B2(n18059), .ZN(
        n18062) );
  OAI221_X1 U21118 ( .B1(n9587), .B2(n18063), .C1(n18253), .C2(n18819), .A(
        n18062), .ZN(P3_U2846) );
  NOR2_X1 U21119 ( .A1(n18064), .A2(n18210), .ZN(n18075) );
  NOR2_X1 U21120 ( .A1(n18065), .A2(n18125), .ZN(n18070) );
  OAI21_X1 U21121 ( .B1(n18066), .B2(n18087), .A(n18078), .ZN(n18067) );
  AOI22_X1 U21122 ( .A1(n18070), .A2(n18069), .B1(n18068), .B2(n18067), .ZN(
        n18072) );
  OAI22_X1 U21123 ( .A1(n18072), .A2(n18254), .B1(n18144), .B2(n18071), .ZN(
        n18073) );
  AOI21_X1 U21124 ( .B1(n18075), .B2(n18074), .A(n18073), .ZN(n18077) );
  OAI211_X1 U21125 ( .C1(n18239), .C2(n18078), .A(n18077), .B(n18076), .ZN(
        P3_U2847) );
  AOI21_X1 U21126 ( .B1(n18079), .B2(n18135), .A(n18716), .ZN(n18085) );
  AOI221_X1 U21127 ( .B1(n18082), .B2(n18081), .C1(n18080), .C2(n18081), .A(
        n18122), .ZN(n18103) );
  OAI211_X1 U21128 ( .C1(n18083), .C2(n18736), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18103), .ZN(n18084) );
  AOI211_X1 U21129 ( .C1(n18106), .C2(n18237), .A(n18085), .B(n18084), .ZN(
        n18086) );
  AOI221_X1 U21130 ( .B1(n18088), .B2(n18096), .C1(n18087), .C2(n18096), .A(
        n18086), .ZN(n18089) );
  AOI22_X1 U21131 ( .A1(n9587), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18238), 
        .B2(n18089), .ZN(n18095) );
  OAI22_X1 U21132 ( .A1(n18210), .A2(n18091), .B1(n18172), .B2(n18090), .ZN(
        n18092) );
  AOI21_X1 U21133 ( .B1(n9572), .B2(n18093), .A(n18092), .ZN(n18094) );
  OAI211_X1 U21134 ( .C1(n18096), .C2(n18239), .A(n18095), .B(n18094), .ZN(
        P3_U2848) );
  OAI21_X1 U21135 ( .B1(n18716), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18117) );
  OAI21_X1 U21136 ( .B1(n18129), .B2(n18097), .A(n18725), .ZN(n18098) );
  OAI21_X1 U21137 ( .B1(n18099), .B2(n18736), .A(n18098), .ZN(n18131) );
  AOI21_X1 U21138 ( .B1(n18101), .B2(n18100), .A(n18131), .ZN(n18102) );
  OAI211_X1 U21139 ( .C1(n18105), .C2(n18104), .A(n18103), .B(n18102), .ZN(
        n18116) );
  AOI211_X1 U21140 ( .C1(n18136), .C2(n18117), .A(n18254), .B(n18116), .ZN(
        n18107) );
  NOR3_X1 U21141 ( .A1(n9587), .A2(n18107), .A3(n18106), .ZN(n18108) );
  AOI21_X1 U21142 ( .B1(n9572), .B2(n18109), .A(n18108), .ZN(n18111) );
  OAI211_X1 U21143 ( .C1(n18156), .C2(n18112), .A(n18111), .B(n18110), .ZN(
        P3_U2849) );
  AOI22_X1 U21144 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18211), .B1(
        n9587), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n18119) );
  OAI22_X1 U21145 ( .A1(n18114), .A2(n18156), .B1(n18113), .B2(n18254), .ZN(
        n18115) );
  OAI21_X1 U21146 ( .B1(n18117), .B2(n18116), .A(n18115), .ZN(n18118) );
  OAI211_X1 U21147 ( .C1(n18120), .C2(n18144), .A(n18119), .B(n18118), .ZN(
        P3_U2850) );
  AOI22_X1 U21148 ( .A1(n9587), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n9572), .B2(
        n18121), .ZN(n18133) );
  AOI21_X1 U21149 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18149), .A(
        n18723), .ZN(n18127) );
  AOI211_X1 U21150 ( .C1(n18123), .C2(n18705), .A(n18122), .B(n18254), .ZN(
        n18124) );
  OAI21_X1 U21151 ( .B1(n18126), .B2(n18125), .A(n18124), .ZN(n18146) );
  AOI211_X1 U21152 ( .C1(n18129), .C2(n18128), .A(n18127), .B(n18146), .ZN(
        n18140) );
  OAI21_X1 U21153 ( .B1(n18723), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18140), .ZN(n18130) );
  OAI211_X1 U21154 ( .C1(n18131), .C2(n18130), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18253), .ZN(n18132) );
  OAI211_X1 U21155 ( .C1(n18134), .C2(n18156), .A(n18133), .B(n18132), .ZN(
        P3_U2851) );
  NOR2_X1 U21156 ( .A1(n18716), .A2(n18135), .ZN(n18137) );
  OAI21_X1 U21157 ( .B1(n18137), .B2(n18155), .A(n18136), .ZN(n18139) );
  AOI21_X1 U21158 ( .B1(n18140), .B2(n18139), .A(n18138), .ZN(n18142) );
  NOR3_X1 U21159 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18155), .A3(
        n18156), .ZN(n18141) );
  AOI221_X1 U21160 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9587), .C1(n18142), 
        .C2(n18253), .A(n18141), .ZN(n18143) );
  OAI21_X1 U21161 ( .B1(n18145), .B2(n18144), .A(n18143), .ZN(P3_U2852) );
  NAND2_X1 U21162 ( .A1(n18725), .A2(n18165), .ZN(n18148) );
  INV_X1 U21163 ( .A(n18146), .ZN(n18147) );
  OAI211_X1 U21164 ( .C1(n18149), .C2(n18723), .A(n18148), .B(n18147), .ZN(
        n18150) );
  OAI21_X1 U21165 ( .B1(n18151), .B2(n18150), .A(n18253), .ZN(n18154) );
  AOI22_X1 U21166 ( .A1(n9587), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n9572), .B2(
        n18152), .ZN(n18153) );
  OAI221_X1 U21167 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18156), .C1(
        n18155), .C2(n18154), .A(n18153), .ZN(P3_U2853) );
  INV_X1 U21168 ( .A(n18157), .ZN(n18158) );
  INV_X1 U21169 ( .A(n18184), .ZN(n18176) );
  NOR3_X1 U21170 ( .A1(n18254), .A2(n18158), .A3(n18176), .ZN(n18166) );
  AOI21_X1 U21171 ( .B1(n18707), .B2(n18159), .A(n18224), .ZN(n18160) );
  OAI21_X1 U21172 ( .B1(n18222), .B2(n18161), .A(n18160), .ZN(n18185) );
  AOI211_X1 U21173 ( .C1(n18162), .C2(n18178), .A(n18177), .B(n18185), .ZN(
        n18175) );
  OAI21_X1 U21174 ( .B1(n18175), .B2(n18240), .A(n18239), .ZN(n18164) );
  NOR2_X1 U21175 ( .A1(n18253), .A2(n18804), .ZN(n18163) );
  AOI221_X1 U21176 ( .B1(n18166), .B2(n18165), .C1(n18164), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18163), .ZN(n18171) );
  AOI22_X1 U21177 ( .A1(n18250), .A2(n18169), .B1(n9572), .B2(n18167), .ZN(
        n18170) );
  OAI211_X1 U21178 ( .C1(n18173), .C2(n18172), .A(n18171), .B(n18170), .ZN(
        P3_U2854) );
  AOI21_X1 U21179 ( .B1(n18211), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18174), .ZN(n18182) );
  AOI221_X1 U21180 ( .B1(n18178), .B2(n18177), .C1(n18176), .C2(n18177), .A(
        n18175), .ZN(n18180) );
  AOI22_X1 U21181 ( .A1(n18238), .A2(n18180), .B1(n18252), .B2(n18179), .ZN(
        n18181) );
  OAI211_X1 U21182 ( .C1(n18210), .C2(n18183), .A(n18182), .B(n18181), .ZN(
        P3_U2855) );
  NAND2_X1 U21183 ( .A1(n18238), .A2(n18184), .ZN(n18191) );
  OAI21_X1 U21184 ( .B1(n18254), .B2(n18185), .A(n18253), .ZN(n18186) );
  INV_X1 U21185 ( .A(n18186), .ZN(n18195) );
  AOI22_X1 U21186 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18195), .B1(
        n9587), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18190) );
  AOI22_X1 U21187 ( .A1(n18250), .A2(n18188), .B1(n18252), .B2(n18187), .ZN(
        n18189) );
  OAI211_X1 U21188 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18191), .A(
        n18190), .B(n18189), .ZN(P3_U2856) );
  NAND4_X1 U21189 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n18238), .A4(n18192), .ZN(
        n18198) );
  AOI22_X1 U21190 ( .A1(n9587), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18250), .B2(
        n18193), .ZN(n18197) );
  AOI22_X1 U21191 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18195), .B1(
        n18252), .B2(n18194), .ZN(n18196) );
  OAI211_X1 U21192 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18198), .A(
        n18197), .B(n18196), .ZN(P3_U2857) );
  AOI22_X1 U21193 ( .A1(n9587), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18252), .B2(
        n18199), .ZN(n18208) );
  INV_X1 U21194 ( .A(n18227), .ZN(n18200) );
  OAI21_X1 U21195 ( .B1(n18736), .B2(n18200), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18201) );
  AOI211_X1 U21196 ( .C1(n18203), .C2(n18202), .A(n18224), .B(n18201), .ZN(
        n18212) );
  OAI21_X1 U21197 ( .B1(n18212), .B2(n18240), .A(n18239), .ZN(n18206) );
  NOR3_X1 U21198 ( .A1(n18214), .A2(n18254), .A3(n18213), .ZN(n18205) );
  AOI22_X1 U21199 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18206), .B1(
        n18205), .B2(n18204), .ZN(n18207) );
  OAI211_X1 U21200 ( .C1(n18210), .C2(n18209), .A(n18208), .B(n18207), .ZN(
        P3_U2858) );
  AOI22_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18211), .B1(
        n9587), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18218) );
  AOI211_X1 U21202 ( .C1(n18214), .C2(n18213), .A(n18212), .B(n18254), .ZN(
        n18215) );
  AOI21_X1 U21203 ( .B1(n18216), .B2(n18250), .A(n18215), .ZN(n18217) );
  OAI211_X1 U21204 ( .C1(n18246), .C2(n18219), .A(n18218), .B(n18217), .ZN(
        P3_U2859) );
  OR2_X1 U21205 ( .A1(n18872), .A2(n18220), .ZN(n18226) );
  NAND2_X1 U21206 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18221) );
  OAI22_X1 U21207 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18222), .B1(
        n18736), .B2(n18221), .ZN(n18223) );
  NOR2_X1 U21208 ( .A1(n18224), .A2(n18223), .ZN(n18225) );
  MUX2_X1 U21209 ( .A(n18226), .B(n18225), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18229) );
  NAND2_X1 U21210 ( .A1(n18707), .A2(n18227), .ZN(n18228) );
  OAI211_X1 U21211 ( .C1(n18230), .C2(n18700), .A(n18229), .B(n18228), .ZN(
        n18232) );
  AOI22_X1 U21212 ( .A1(n18238), .A2(n18232), .B1(n18250), .B2(n18231), .ZN(
        n18234) );
  OAI211_X1 U21213 ( .C1(n18239), .C2(n18235), .A(n18234), .B(n18233), .ZN(
        P3_U2860) );
  INV_X1 U21214 ( .A(n18236), .ZN(n18247) );
  NAND3_X1 U21215 ( .A1(n18238), .A2(n18890), .A3(n18237), .ZN(n18256) );
  AOI21_X1 U21216 ( .B1(n18239), .B2(n18256), .A(n18872), .ZN(n18242) );
  AOI211_X1 U21217 ( .C1(n18716), .C2(n18890), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18240), .ZN(n18241) );
  AOI211_X1 U21218 ( .C1(n18250), .C2(n18243), .A(n18242), .B(n18241), .ZN(
        n18245) );
  NAND2_X1 U21219 ( .A1(n9587), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18244) );
  OAI211_X1 U21220 ( .C1(n18247), .C2(n18246), .A(n18245), .B(n18244), .ZN(
        P3_U2861) );
  INV_X1 U21221 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18901) );
  NOR2_X1 U21222 ( .A1(n18253), .A2(n18901), .ZN(n18248) );
  AOI221_X1 U21223 ( .B1(n18252), .B2(n18251), .C1(n18250), .C2(n18249), .A(
        n18248), .ZN(n18257) );
  OAI211_X1 U21224 ( .C1(n18725), .C2(n18254), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18253), .ZN(n18255) );
  NAND3_X1 U21225 ( .A1(n18257), .A2(n18256), .A3(n18255), .ZN(P3_U2862) );
  INV_X1 U21226 ( .A(n18265), .ZN(n18261) );
  OAI211_X1 U21227 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18258), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18760)
         );
  OAI21_X1 U21228 ( .B1(n18261), .B2(n18259), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18260) );
  OAI221_X1 U21229 ( .B1(n18261), .B2(n18760), .C1(n18261), .C2(n18307), .A(
        n18260), .ZN(P3_U2863) );
  INV_X1 U21230 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18742) );
  NAND2_X1 U21231 ( .A1(n18271), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18536) );
  INV_X1 U21232 ( .A(n18536), .ZN(n18559) );
  NAND2_X1 U21233 ( .A1(n18742), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18443) );
  INV_X1 U21234 ( .A(n18443), .ZN(n18445) );
  NOR2_X1 U21235 ( .A1(n18559), .A2(n18445), .ZN(n18263) );
  OAI22_X1 U21236 ( .A1(n18264), .A2(n18742), .B1(n18263), .B2(n18262), .ZN(
        P3_U2866) );
  NOR2_X1 U21237 ( .A1(n18266), .A2(n18265), .ZN(P3_U2867) );
  NOR2_X1 U21238 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U21239 ( .A1(n18271), .A2(n18742), .ZN(n18396) );
  INV_X1 U21240 ( .A(n18396), .ZN(n18350) );
  NAND2_X1 U21241 ( .A1(n18728), .A2(n18350), .ZN(n18328) );
  NOR2_X1 U21242 ( .A1(n18268), .A2(n18267), .ZN(n18300) );
  NAND2_X1 U21243 ( .A1(n18300), .A2(n18269), .ZN(n18652) );
  NOR2_X2 U21244 ( .A1(n18372), .A2(n18270), .ZN(n18643) );
  INV_X1 U21245 ( .A(n18589), .ZN(n18761) );
  NAND2_X1 U21246 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18537) );
  INV_X1 U21247 ( .A(n18537), .ZN(n18727) );
  NOR2_X1 U21248 ( .A1(n18271), .A2(n18742), .ZN(n18272) );
  NAND2_X1 U21249 ( .A1(n18727), .A2(n18272), .ZN(n18699) );
  NAND2_X1 U21250 ( .A1(n18699), .A2(n18328), .ZN(n18329) );
  AND2_X1 U21251 ( .A1(n18761), .A2(n18329), .ZN(n18302) );
  AND2_X1 U21252 ( .A1(n18648), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18649) );
  NOR2_X1 U21253 ( .A1(n18397), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18512) );
  NAND2_X1 U21254 ( .A1(n18272), .A2(n18512), .ZN(n18642) );
  INV_X1 U21255 ( .A(n18642), .ZN(n18324) );
  AOI22_X1 U21256 ( .A1(n18643), .A2(n18302), .B1(n18649), .B2(n18324), .ZN(
        n18276) );
  NOR2_X1 U21257 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18273), .ZN(
        n18488) );
  NOR2_X1 U21258 ( .A1(n18512), .A2(n18488), .ZN(n18562) );
  INV_X1 U21259 ( .A(n18272), .ZN(n18274) );
  NOR2_X1 U21260 ( .A1(n18562), .A2(n18274), .ZN(n18622) );
  OAI21_X1 U21261 ( .B1(n18273), .B2(n18862), .A(n18564), .ZN(n18420) );
  INV_X1 U21262 ( .A(n18420), .ZN(n18619) );
  AOI22_X1 U21263 ( .A1(n18648), .A2(n18622), .B1(n18619), .B2(n18329), .ZN(
        n18304) );
  NOR2_X1 U21264 ( .A1(n18274), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18647) );
  NAND2_X1 U21265 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18647), .ZN(
        n18618) );
  INV_X1 U21266 ( .A(n18618), .ZN(n18692) );
  AND2_X1 U21267 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18648), .ZN(n18644) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18304), .B1(
        n18692), .B2(n18644), .ZN(n18275) );
  OAI211_X1 U21269 ( .C1(n18328), .C2(n18652), .A(n18276), .B(n18275), .ZN(
        P3_U2868) );
  NAND2_X1 U21270 ( .A1(n18300), .A2(n18277), .ZN(n18658) );
  AND2_X1 U21271 ( .A1(n18564), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18653) );
  AND2_X1 U21272 ( .A1(n18648), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18654) );
  AOI22_X1 U21273 ( .A1(n18302), .A2(n18653), .B1(n18324), .B2(n18654), .ZN(
        n18279) );
  AND2_X1 U21274 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18648), .ZN(n18655) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18304), .B1(
        n18692), .B2(n18655), .ZN(n18278) );
  OAI211_X1 U21276 ( .C1(n18328), .C2(n18658), .A(n18279), .B(n18278), .ZN(
        P3_U2869) );
  NAND2_X1 U21277 ( .A1(n18300), .A2(n18280), .ZN(n18664) );
  NOR2_X2 U21278 ( .A1(n14947), .A2(n18587), .ZN(n18661) );
  NOR2_X2 U21279 ( .A1(n18372), .A2(n18281), .ZN(n18659) );
  AOI22_X1 U21280 ( .A1(n18692), .A2(n18661), .B1(n18302), .B2(n18659), .ZN(
        n18283) );
  AND2_X1 U21281 ( .A1(n18648), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18660) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18660), .ZN(n18282) );
  OAI211_X1 U21283 ( .C1(n18328), .C2(n18664), .A(n18283), .B(n18282), .ZN(
        P3_U2870) );
  NAND2_X1 U21284 ( .A1(n18300), .A2(n18284), .ZN(n18670) );
  AND2_X1 U21285 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18648), .ZN(n18666) );
  AND2_X1 U21286 ( .A1(n18564), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18665) );
  AOI22_X1 U21287 ( .A1(n18692), .A2(n18666), .B1(n18302), .B2(n18665), .ZN(
        n18286) );
  AND2_X1 U21288 ( .A1(n18648), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18667) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18667), .ZN(n18285) );
  OAI211_X1 U21290 ( .C1(n18328), .C2(n18670), .A(n18286), .B(n18285), .ZN(
        P3_U2871) );
  NAND2_X1 U21291 ( .A1(n18300), .A2(n18287), .ZN(n18676) );
  AND2_X1 U21292 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18648), .ZN(n18671) );
  NOR2_X2 U21293 ( .A1(n18372), .A2(n18288), .ZN(n18672) );
  AOI22_X1 U21294 ( .A1(n18692), .A2(n18671), .B1(n18302), .B2(n18672), .ZN(
        n18290) );
  AND2_X1 U21295 ( .A1(n18648), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18673) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18673), .ZN(n18289) );
  OAI211_X1 U21297 ( .C1(n18328), .C2(n18676), .A(n18290), .B(n18289), .ZN(
        P3_U2872) );
  NAND2_X1 U21298 ( .A1(n18300), .A2(n18291), .ZN(n18682) );
  NOR2_X2 U21299 ( .A1(n18292), .A2(n18372), .ZN(n18677) );
  AND2_X1 U21300 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18648), .ZN(n18678) );
  AOI22_X1 U21301 ( .A1(n18302), .A2(n18677), .B1(n18324), .B2(n18678), .ZN(
        n18294) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18304), .B1(
        n18692), .B2(n18679), .ZN(n18293) );
  OAI211_X1 U21303 ( .C1(n18328), .C2(n18682), .A(n18294), .B(n18293), .ZN(
        P3_U2873) );
  NAND2_X1 U21304 ( .A1(n18300), .A2(n18295), .ZN(n18688) );
  NOR2_X2 U21305 ( .A1(n18296), .A2(n18372), .ZN(n18683) );
  AND2_X1 U21306 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18648), .ZN(n18684) );
  AOI22_X1 U21307 ( .A1(n18302), .A2(n18683), .B1(n18324), .B2(n18684), .ZN(
        n18298) );
  AND2_X1 U21308 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18648), .ZN(n18685) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18304), .B1(
        n18692), .B2(n18685), .ZN(n18297) );
  OAI211_X1 U21310 ( .C1(n18328), .C2(n18688), .A(n18298), .B(n18297), .ZN(
        P3_U2874) );
  NAND2_X1 U21311 ( .A1(n18300), .A2(n18299), .ZN(n18698) );
  NOR2_X2 U21312 ( .A1(n18301), .A2(n18372), .ZN(n18690) );
  AND2_X1 U21313 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18648), .ZN(n18691) );
  AOI22_X1 U21314 ( .A1(n18302), .A2(n18690), .B1(n18324), .B2(n18691), .ZN(
        n18306) );
  NOR2_X2 U21315 ( .A1(n18587), .A2(n18303), .ZN(n18694) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18304), .B1(
        n18692), .B2(n18694), .ZN(n18305) );
  OAI211_X1 U21317 ( .C1(n18328), .C2(n18698), .A(n18306), .B(n18305), .ZN(
        P3_U2875) );
  NAND2_X1 U21318 ( .A1(n18350), .A2(n18488), .ZN(n18351) );
  NAND2_X1 U21319 ( .A1(n18397), .A2(n18761), .ZN(n18489) );
  NOR2_X1 U21320 ( .A1(n18396), .A2(n18489), .ZN(n18323) );
  AOI22_X1 U21321 ( .A1(n18644), .A2(n18324), .B1(n18643), .B2(n18323), .ZN(
        n18310) );
  NOR2_X1 U21322 ( .A1(n18742), .A2(n18490), .ZN(n18645) );
  INV_X1 U21323 ( .A(n18307), .ZN(n18308) );
  NOR2_X1 U21324 ( .A1(n18372), .A2(n18308), .ZN(n18646) );
  INV_X1 U21325 ( .A(n18646), .ZN(n18585) );
  NOR2_X1 U21326 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18585), .ZN(
        n18398) );
  AOI22_X1 U21327 ( .A1(n18648), .A2(n18645), .B1(n18350), .B2(n18398), .ZN(
        n18325) );
  INV_X1 U21328 ( .A(n18699), .ZN(n18346) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18649), .ZN(n18309) );
  OAI211_X1 U21330 ( .C1(n18652), .C2(n18351), .A(n18310), .B(n18309), .ZN(
        P3_U2876) );
  AOI22_X1 U21331 ( .A1(n18346), .A2(n18654), .B1(n18653), .B2(n18323), .ZN(
        n18312) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18655), .ZN(n18311) );
  OAI211_X1 U21333 ( .C1(n18658), .C2(n18351), .A(n18312), .B(n18311), .ZN(
        P3_U2877) );
  AOI22_X1 U21334 ( .A1(n18324), .A2(n18661), .B1(n18659), .B2(n18323), .ZN(
        n18314) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18660), .ZN(n18313) );
  OAI211_X1 U21336 ( .C1(n18664), .C2(n18351), .A(n18314), .B(n18313), .ZN(
        P3_U2878) );
  AOI22_X1 U21337 ( .A1(n18346), .A2(n18667), .B1(n18665), .B2(n18323), .ZN(
        n18316) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18666), .ZN(n18315) );
  OAI211_X1 U21339 ( .C1(n18670), .C2(n18351), .A(n18316), .B(n18315), .ZN(
        P3_U2879) );
  AOI22_X1 U21340 ( .A1(n18324), .A2(n18671), .B1(n18672), .B2(n18323), .ZN(
        n18318) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18673), .ZN(n18317) );
  OAI211_X1 U21342 ( .C1(n18676), .C2(n18351), .A(n18318), .B(n18317), .ZN(
        P3_U2880) );
  AOI22_X1 U21343 ( .A1(n18324), .A2(n18679), .B1(n18677), .B2(n18323), .ZN(
        n18320) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18678), .ZN(n18319) );
  OAI211_X1 U21345 ( .C1(n18682), .C2(n18351), .A(n18320), .B(n18319), .ZN(
        P3_U2881) );
  AOI22_X1 U21346 ( .A1(n18324), .A2(n18685), .B1(n18683), .B2(n18323), .ZN(
        n18322) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18684), .ZN(n18321) );
  OAI211_X1 U21348 ( .C1(n18688), .C2(n18351), .A(n18322), .B(n18321), .ZN(
        P3_U2882) );
  AOI22_X1 U21349 ( .A1(n18324), .A2(n18694), .B1(n18690), .B2(n18323), .ZN(
        n18327) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18691), .ZN(n18326) );
  OAI211_X1 U21351 ( .C1(n18698), .C2(n18351), .A(n18327), .B(n18326), .ZN(
        P3_U2883) );
  NAND2_X1 U21352 ( .A1(n18350), .A2(n18512), .ZN(n18375) );
  INV_X1 U21353 ( .A(n18328), .ZN(n18367) );
  NAND2_X1 U21354 ( .A1(n18351), .A2(n18375), .ZN(n18330) );
  INV_X1 U21355 ( .A(n18330), .ZN(n18373) );
  NOR2_X1 U21356 ( .A1(n18589), .A2(n18373), .ZN(n18345) );
  AOI22_X1 U21357 ( .A1(n18367), .A2(n18649), .B1(n18643), .B2(n18345), .ZN(
        n18332) );
  OAI221_X1 U21358 ( .B1(n18330), .B2(n18621), .C1(n18330), .C2(n18329), .A(
        n18619), .ZN(n18347) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18347), .B1(
        n18644), .B2(n18346), .ZN(n18331) );
  OAI211_X1 U21360 ( .C1(n18652), .C2(n18375), .A(n18332), .B(n18331), .ZN(
        P3_U2884) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18347), .B1(
        n18653), .B2(n18345), .ZN(n18334) );
  AOI22_X1 U21362 ( .A1(n18346), .A2(n18655), .B1(n18367), .B2(n18654), .ZN(
        n18333) );
  OAI211_X1 U21363 ( .C1(n18658), .C2(n18375), .A(n18334), .B(n18333), .ZN(
        P3_U2885) );
  AOI22_X1 U21364 ( .A1(n18367), .A2(n18660), .B1(n18659), .B2(n18345), .ZN(
        n18336) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18661), .ZN(n18335) );
  OAI211_X1 U21366 ( .C1(n18664), .C2(n18375), .A(n18336), .B(n18335), .ZN(
        P3_U2886) );
  AOI22_X1 U21367 ( .A1(n18367), .A2(n18667), .B1(n18665), .B2(n18345), .ZN(
        n18338) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18666), .ZN(n18337) );
  OAI211_X1 U21369 ( .C1(n18670), .C2(n18375), .A(n18338), .B(n18337), .ZN(
        P3_U2887) );
  AOI22_X1 U21370 ( .A1(n18346), .A2(n18671), .B1(n18672), .B2(n18345), .ZN(
        n18340) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18347), .B1(
        n18367), .B2(n18673), .ZN(n18339) );
  OAI211_X1 U21372 ( .C1(n18676), .C2(n18375), .A(n18340), .B(n18339), .ZN(
        P3_U2888) );
  AOI22_X1 U21373 ( .A1(n18346), .A2(n18679), .B1(n18677), .B2(n18345), .ZN(
        n18342) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18347), .B1(
        n18367), .B2(n18678), .ZN(n18341) );
  OAI211_X1 U21375 ( .C1(n18682), .C2(n18375), .A(n18342), .B(n18341), .ZN(
        P3_U2889) );
  AOI22_X1 U21376 ( .A1(n18367), .A2(n18684), .B1(n18683), .B2(n18345), .ZN(
        n18344) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18685), .ZN(n18343) );
  OAI211_X1 U21378 ( .C1(n18688), .C2(n18375), .A(n18344), .B(n18343), .ZN(
        P3_U2890) );
  AOI22_X1 U21379 ( .A1(n18367), .A2(n18691), .B1(n18690), .B2(n18345), .ZN(
        n18349) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18694), .ZN(n18348) );
  OAI211_X1 U21381 ( .C1(n18698), .C2(n18375), .A(n18349), .B(n18348), .ZN(
        P3_U2891) );
  NOR2_X2 U21382 ( .A1(n18537), .A2(n18396), .ZN(n18438) );
  INV_X1 U21383 ( .A(n18438), .ZN(n18371) );
  AOI22_X1 U21384 ( .A1(n18644), .A2(n18367), .B1(n18643), .B2(n18366), .ZN(
        n18353) );
  AOI21_X1 U21385 ( .B1(n18397), .B2(n18513), .A(n18585), .ZN(n18444) );
  NAND2_X1 U21386 ( .A1(n18350), .A2(n18444), .ZN(n18368) );
  INV_X1 U21387 ( .A(n18351), .ZN(n18391) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18368), .B1(
        n18649), .B2(n18391), .ZN(n18352) );
  OAI211_X1 U21389 ( .C1(n18652), .C2(n18371), .A(n18353), .B(n18352), .ZN(
        P3_U2892) );
  AOI22_X1 U21390 ( .A1(n18367), .A2(n18655), .B1(n18653), .B2(n18366), .ZN(
        n18355) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18368), .B1(
        n18654), .B2(n18391), .ZN(n18354) );
  OAI211_X1 U21392 ( .C1(n18658), .C2(n18371), .A(n18355), .B(n18354), .ZN(
        P3_U2893) );
  AOI22_X1 U21393 ( .A1(n18660), .A2(n18391), .B1(n18659), .B2(n18366), .ZN(
        n18357) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18368), .B1(
        n18367), .B2(n18661), .ZN(n18356) );
  OAI211_X1 U21395 ( .C1(n18664), .C2(n18371), .A(n18357), .B(n18356), .ZN(
        P3_U2894) );
  AOI22_X1 U21396 ( .A1(n18667), .A2(n18391), .B1(n18665), .B2(n18366), .ZN(
        n18359) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18368), .B1(
        n18367), .B2(n18666), .ZN(n18358) );
  OAI211_X1 U21398 ( .C1(n18670), .C2(n18371), .A(n18359), .B(n18358), .ZN(
        P3_U2895) );
  AOI22_X1 U21399 ( .A1(n18673), .A2(n18391), .B1(n18672), .B2(n18366), .ZN(
        n18361) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18368), .B1(
        n18367), .B2(n18671), .ZN(n18360) );
  OAI211_X1 U21401 ( .C1(n18676), .C2(n18371), .A(n18361), .B(n18360), .ZN(
        P3_U2896) );
  AOI22_X1 U21402 ( .A1(n18678), .A2(n18391), .B1(n18677), .B2(n18366), .ZN(
        n18363) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18368), .B1(
        n18367), .B2(n18679), .ZN(n18362) );
  OAI211_X1 U21404 ( .C1(n18682), .C2(n18371), .A(n18363), .B(n18362), .ZN(
        P3_U2897) );
  AOI22_X1 U21405 ( .A1(n18684), .A2(n18391), .B1(n18683), .B2(n18366), .ZN(
        n18365) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18368), .B1(
        n18367), .B2(n18685), .ZN(n18364) );
  OAI211_X1 U21407 ( .C1(n18688), .C2(n18371), .A(n18365), .B(n18364), .ZN(
        P3_U2898) );
  AOI22_X1 U21408 ( .A1(n18367), .A2(n18694), .B1(n18690), .B2(n18366), .ZN(
        n18370) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18368), .B1(
        n18691), .B2(n18391), .ZN(n18369) );
  OAI211_X1 U21410 ( .C1(n18698), .C2(n18371), .A(n18370), .B(n18369), .ZN(
        P3_U2899) );
  NAND2_X1 U21411 ( .A1(n18728), .A2(n18445), .ZN(n18395) );
  NOR2_X1 U21412 ( .A1(n18438), .A2(n18461), .ZN(n18421) );
  NOR2_X1 U21413 ( .A1(n18589), .A2(n18421), .ZN(n18390) );
  AOI22_X1 U21414 ( .A1(n18644), .A2(n18391), .B1(n18643), .B2(n18390), .ZN(
        n18377) );
  OAI22_X1 U21415 ( .A1(n18373), .A2(n18587), .B1(n18421), .B2(n18372), .ZN(
        n18374) );
  OAI21_X1 U21416 ( .B1(n18461), .B2(n18862), .A(n18374), .ZN(n18392) );
  INV_X1 U21417 ( .A(n18375), .ZN(n18415) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18392), .B1(
        n18649), .B2(n18415), .ZN(n18376) );
  OAI211_X1 U21419 ( .C1(n18652), .C2(n18395), .A(n18377), .B(n18376), .ZN(
        P3_U2900) );
  AOI22_X1 U21420 ( .A1(n18653), .A2(n18390), .B1(n18654), .B2(n18415), .ZN(
        n18379) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18392), .B1(
        n18655), .B2(n18391), .ZN(n18378) );
  OAI211_X1 U21422 ( .C1(n18658), .C2(n18395), .A(n18379), .B(n18378), .ZN(
        P3_U2901) );
  AOI22_X1 U21423 ( .A1(n18660), .A2(n18415), .B1(n18659), .B2(n18390), .ZN(
        n18381) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18392), .B1(
        n18661), .B2(n18391), .ZN(n18380) );
  OAI211_X1 U21425 ( .C1(n18664), .C2(n18395), .A(n18381), .B(n18380), .ZN(
        P3_U2902) );
  AOI22_X1 U21426 ( .A1(n18666), .A2(n18391), .B1(n18665), .B2(n18390), .ZN(
        n18383) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18392), .B1(
        n18667), .B2(n18415), .ZN(n18382) );
  OAI211_X1 U21428 ( .C1(n18670), .C2(n18395), .A(n18383), .B(n18382), .ZN(
        P3_U2903) );
  AOI22_X1 U21429 ( .A1(n18672), .A2(n18390), .B1(n18671), .B2(n18391), .ZN(
        n18385) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18392), .B1(
        n18673), .B2(n18415), .ZN(n18384) );
  OAI211_X1 U21431 ( .C1(n18676), .C2(n18395), .A(n18385), .B(n18384), .ZN(
        P3_U2904) );
  AOI22_X1 U21432 ( .A1(n18679), .A2(n18391), .B1(n18677), .B2(n18390), .ZN(
        n18387) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18392), .B1(
        n18678), .B2(n18415), .ZN(n18386) );
  OAI211_X1 U21434 ( .C1(n18682), .C2(n18395), .A(n18387), .B(n18386), .ZN(
        P3_U2905) );
  AOI22_X1 U21435 ( .A1(n18684), .A2(n18415), .B1(n18683), .B2(n18390), .ZN(
        n18389) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18392), .B1(
        n18685), .B2(n18391), .ZN(n18388) );
  OAI211_X1 U21437 ( .C1(n18688), .C2(n18395), .A(n18389), .B(n18388), .ZN(
        P3_U2906) );
  AOI22_X1 U21438 ( .A1(n18694), .A2(n18391), .B1(n18690), .B2(n18390), .ZN(
        n18394) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18392), .B1(
        n18691), .B2(n18415), .ZN(n18393) );
  OAI211_X1 U21440 ( .C1(n18698), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        P3_U2907) );
  NAND2_X1 U21441 ( .A1(n18445), .A2(n18488), .ZN(n18419) );
  NOR2_X1 U21442 ( .A1(n18443), .A2(n18489), .ZN(n18414) );
  AOI22_X1 U21443 ( .A1(n18644), .A2(n18415), .B1(n18643), .B2(n18414), .ZN(
        n18401) );
  NOR2_X1 U21444 ( .A1(n18397), .A2(n18396), .ZN(n18399) );
  AOI22_X1 U21445 ( .A1(n18648), .A2(n18399), .B1(n18445), .B2(n18398), .ZN(
        n18416) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18416), .B1(
        n18649), .B2(n18438), .ZN(n18400) );
  OAI211_X1 U21447 ( .C1(n18652), .C2(n18419), .A(n18401), .B(n18400), .ZN(
        P3_U2908) );
  AOI22_X1 U21448 ( .A1(n18655), .A2(n18415), .B1(n18653), .B2(n18414), .ZN(
        n18403) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18416), .B1(
        n18654), .B2(n18438), .ZN(n18402) );
  OAI211_X1 U21450 ( .C1(n18658), .C2(n18419), .A(n18403), .B(n18402), .ZN(
        P3_U2909) );
  AOI22_X1 U21451 ( .A1(n18660), .A2(n18438), .B1(n18659), .B2(n18414), .ZN(
        n18405) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18416), .B1(
        n18661), .B2(n18415), .ZN(n18404) );
  OAI211_X1 U21453 ( .C1(n18664), .C2(n18419), .A(n18405), .B(n18404), .ZN(
        P3_U2910) );
  AOI22_X1 U21454 ( .A1(n18667), .A2(n18438), .B1(n18665), .B2(n18414), .ZN(
        n18407) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18416), .B1(
        n18666), .B2(n18415), .ZN(n18406) );
  OAI211_X1 U21456 ( .C1(n18670), .C2(n18419), .A(n18407), .B(n18406), .ZN(
        P3_U2911) );
  AOI22_X1 U21457 ( .A1(n18672), .A2(n18414), .B1(n18671), .B2(n18415), .ZN(
        n18409) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18416), .B1(
        n18673), .B2(n18438), .ZN(n18408) );
  OAI211_X1 U21459 ( .C1(n18676), .C2(n18419), .A(n18409), .B(n18408), .ZN(
        P3_U2912) );
  AOI22_X1 U21460 ( .A1(n18679), .A2(n18415), .B1(n18677), .B2(n18414), .ZN(
        n18411) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18416), .B1(
        n18678), .B2(n18438), .ZN(n18410) );
  OAI211_X1 U21462 ( .C1(n18682), .C2(n18419), .A(n18411), .B(n18410), .ZN(
        P3_U2913) );
  AOI22_X1 U21463 ( .A1(n18685), .A2(n18415), .B1(n18683), .B2(n18414), .ZN(
        n18413) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18416), .B1(
        n18684), .B2(n18438), .ZN(n18412) );
  OAI211_X1 U21465 ( .C1(n18688), .C2(n18419), .A(n18413), .B(n18412), .ZN(
        P3_U2914) );
  AOI22_X1 U21466 ( .A1(n18691), .A2(n18438), .B1(n18690), .B2(n18414), .ZN(
        n18418) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18416), .B1(
        n18694), .B2(n18415), .ZN(n18417) );
  OAI211_X1 U21468 ( .C1(n18698), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        P3_U2915) );
  NAND2_X1 U21469 ( .A1(n18445), .A2(n18512), .ZN(n18442) );
  INV_X1 U21470 ( .A(n18419), .ZN(n18483) );
  NOR2_X1 U21471 ( .A1(n18483), .A2(n18508), .ZN(n18466) );
  NOR2_X1 U21472 ( .A1(n18589), .A2(n18466), .ZN(n18437) );
  AOI22_X1 U21473 ( .A1(n18644), .A2(n18438), .B1(n18643), .B2(n18437), .ZN(
        n18424) );
  AOI221_X1 U21474 ( .B1(n18466), .B2(n18513), .C1(n18466), .C2(n18421), .A(
        n18420), .ZN(n18422) );
  INV_X1 U21475 ( .A(n18422), .ZN(n18439) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18439), .B1(
        n18649), .B2(n18461), .ZN(n18423) );
  OAI211_X1 U21477 ( .C1(n18652), .C2(n18442), .A(n18424), .B(n18423), .ZN(
        P3_U2916) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18439), .B1(
        n18653), .B2(n18437), .ZN(n18426) );
  AOI22_X1 U21479 ( .A1(n18655), .A2(n18438), .B1(n18654), .B2(n18461), .ZN(
        n18425) );
  OAI211_X1 U21480 ( .C1(n18658), .C2(n18442), .A(n18426), .B(n18425), .ZN(
        P3_U2917) );
  AOI22_X1 U21481 ( .A1(n18660), .A2(n18461), .B1(n18659), .B2(n18437), .ZN(
        n18428) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18439), .B1(
        n18661), .B2(n18438), .ZN(n18427) );
  OAI211_X1 U21483 ( .C1(n18664), .C2(n18442), .A(n18428), .B(n18427), .ZN(
        P3_U2918) );
  AOI22_X1 U21484 ( .A1(n18667), .A2(n18461), .B1(n18665), .B2(n18437), .ZN(
        n18430) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18439), .B1(
        n18666), .B2(n18438), .ZN(n18429) );
  OAI211_X1 U21486 ( .C1(n18670), .C2(n18442), .A(n18430), .B(n18429), .ZN(
        P3_U2919) );
  AOI22_X1 U21487 ( .A1(n18672), .A2(n18437), .B1(n18671), .B2(n18438), .ZN(
        n18432) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18439), .B1(
        n18673), .B2(n18461), .ZN(n18431) );
  OAI211_X1 U21489 ( .C1(n18676), .C2(n18442), .A(n18432), .B(n18431), .ZN(
        P3_U2920) );
  AOI22_X1 U21490 ( .A1(n18679), .A2(n18438), .B1(n18677), .B2(n18437), .ZN(
        n18434) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18439), .B1(
        n18678), .B2(n18461), .ZN(n18433) );
  OAI211_X1 U21492 ( .C1(n18682), .C2(n18442), .A(n18434), .B(n18433), .ZN(
        P3_U2921) );
  AOI22_X1 U21493 ( .A1(n18685), .A2(n18438), .B1(n18683), .B2(n18437), .ZN(
        n18436) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18439), .B1(
        n18684), .B2(n18461), .ZN(n18435) );
  OAI211_X1 U21495 ( .C1(n18688), .C2(n18442), .A(n18436), .B(n18435), .ZN(
        P3_U2922) );
  AOI22_X1 U21496 ( .A1(n18691), .A2(n18461), .B1(n18690), .B2(n18437), .ZN(
        n18441) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18439), .B1(
        n18694), .B2(n18438), .ZN(n18440) );
  OAI211_X1 U21498 ( .C1(n18698), .C2(n18442), .A(n18441), .B(n18440), .ZN(
        P3_U2923) );
  NOR2_X2 U21499 ( .A1(n18537), .A2(n18443), .ZN(n18531) );
  INV_X1 U21500 ( .A(n18531), .ZN(n18465) );
  AOI22_X1 U21501 ( .A1(n18644), .A2(n18461), .B1(n18643), .B2(n18460), .ZN(
        n18447) );
  NAND2_X1 U21502 ( .A1(n18445), .A2(n18444), .ZN(n18462) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18462), .B1(
        n18649), .B2(n18483), .ZN(n18446) );
  OAI211_X1 U21504 ( .C1(n18652), .C2(n18465), .A(n18447), .B(n18446), .ZN(
        P3_U2924) );
  AOI22_X1 U21505 ( .A1(n18655), .A2(n18461), .B1(n18653), .B2(n18460), .ZN(
        n18449) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18462), .B1(
        n18654), .B2(n18483), .ZN(n18448) );
  OAI211_X1 U21507 ( .C1(n18658), .C2(n18465), .A(n18449), .B(n18448), .ZN(
        P3_U2925) );
  AOI22_X1 U21508 ( .A1(n18660), .A2(n18483), .B1(n18659), .B2(n18460), .ZN(
        n18451) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18462), .B1(
        n18661), .B2(n18461), .ZN(n18450) );
  OAI211_X1 U21510 ( .C1(n18664), .C2(n18465), .A(n18451), .B(n18450), .ZN(
        P3_U2926) );
  AOI22_X1 U21511 ( .A1(n18666), .A2(n18461), .B1(n18665), .B2(n18460), .ZN(
        n18453) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18462), .B1(
        n18667), .B2(n18483), .ZN(n18452) );
  OAI211_X1 U21513 ( .C1(n18670), .C2(n18465), .A(n18453), .B(n18452), .ZN(
        P3_U2927) );
  AOI22_X1 U21514 ( .A1(n18672), .A2(n18460), .B1(n18671), .B2(n18461), .ZN(
        n18455) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18462), .B1(
        n18673), .B2(n18483), .ZN(n18454) );
  OAI211_X1 U21516 ( .C1(n18676), .C2(n18465), .A(n18455), .B(n18454), .ZN(
        P3_U2928) );
  AOI22_X1 U21517 ( .A1(n18679), .A2(n18461), .B1(n18677), .B2(n18460), .ZN(
        n18457) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18462), .B1(
        n18678), .B2(n18483), .ZN(n18456) );
  OAI211_X1 U21519 ( .C1(n18682), .C2(n18465), .A(n18457), .B(n18456), .ZN(
        P3_U2929) );
  AOI22_X1 U21520 ( .A1(n18685), .A2(n18461), .B1(n18683), .B2(n18460), .ZN(
        n18459) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18462), .B1(
        n18684), .B2(n18483), .ZN(n18458) );
  OAI211_X1 U21522 ( .C1(n18688), .C2(n18465), .A(n18459), .B(n18458), .ZN(
        P3_U2930) );
  AOI22_X1 U21523 ( .A1(n18691), .A2(n18483), .B1(n18690), .B2(n18460), .ZN(
        n18464) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18462), .B1(
        n18694), .B2(n18461), .ZN(n18463) );
  OAI211_X1 U21525 ( .C1(n18698), .C2(n18465), .A(n18464), .B(n18463), .ZN(
        P3_U2931) );
  NAND2_X1 U21526 ( .A1(n18728), .A2(n18559), .ZN(n18487) );
  AOI21_X1 U21527 ( .B1(n18465), .B2(n18487), .A(n18589), .ZN(n18482) );
  AOI22_X1 U21528 ( .A1(n18643), .A2(n18482), .B1(n18649), .B2(n18508), .ZN(
        n18469) );
  AOI221_X1 U21529 ( .B1(n18466), .B2(n18465), .C1(n18513), .C2(n18465), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18467) );
  OAI21_X1 U21530 ( .B1(n18554), .B2(n18467), .A(n18564), .ZN(n18484) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18484), .B1(
        n18644), .B2(n18483), .ZN(n18468) );
  OAI211_X1 U21532 ( .C1(n18652), .C2(n18487), .A(n18469), .B(n18468), .ZN(
        P3_U2932) );
  AOI22_X1 U21533 ( .A1(n18653), .A2(n18482), .B1(n18654), .B2(n18508), .ZN(
        n18471) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18484), .B1(
        n18655), .B2(n18483), .ZN(n18470) );
  OAI211_X1 U21535 ( .C1(n18658), .C2(n18487), .A(n18471), .B(n18470), .ZN(
        P3_U2933) );
  AOI22_X1 U21536 ( .A1(n18659), .A2(n18482), .B1(n18661), .B2(n18483), .ZN(
        n18473) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18484), .B1(
        n18660), .B2(n18508), .ZN(n18472) );
  OAI211_X1 U21538 ( .C1(n18664), .C2(n18487), .A(n18473), .B(n18472), .ZN(
        P3_U2934) );
  AOI22_X1 U21539 ( .A1(n18666), .A2(n18483), .B1(n18665), .B2(n18482), .ZN(
        n18475) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18484), .B1(
        n18667), .B2(n18508), .ZN(n18474) );
  OAI211_X1 U21541 ( .C1(n18670), .C2(n18487), .A(n18475), .B(n18474), .ZN(
        P3_U2935) );
  AOI22_X1 U21542 ( .A1(n18672), .A2(n18482), .B1(n18671), .B2(n18483), .ZN(
        n18477) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18484), .B1(
        n18673), .B2(n18508), .ZN(n18476) );
  OAI211_X1 U21544 ( .C1(n18676), .C2(n18487), .A(n18477), .B(n18476), .ZN(
        P3_U2936) );
  AOI22_X1 U21545 ( .A1(n18678), .A2(n18508), .B1(n18677), .B2(n18482), .ZN(
        n18479) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18484), .B1(
        n18679), .B2(n18483), .ZN(n18478) );
  OAI211_X1 U21547 ( .C1(n18682), .C2(n18487), .A(n18479), .B(n18478), .ZN(
        P3_U2937) );
  AOI22_X1 U21548 ( .A1(n18684), .A2(n18508), .B1(n18683), .B2(n18482), .ZN(
        n18481) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18484), .B1(
        n18685), .B2(n18483), .ZN(n18480) );
  OAI211_X1 U21550 ( .C1(n18688), .C2(n18487), .A(n18481), .B(n18480), .ZN(
        P3_U2938) );
  AOI22_X1 U21551 ( .A1(n18691), .A2(n18508), .B1(n18690), .B2(n18482), .ZN(
        n18486) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18484), .B1(
        n18694), .B2(n18483), .ZN(n18485) );
  OAI211_X1 U21553 ( .C1(n18698), .C2(n18487), .A(n18486), .B(n18485), .ZN(
        P3_U2939) );
  NAND2_X1 U21554 ( .A1(n18559), .A2(n18488), .ZN(n18538) );
  NOR2_X1 U21555 ( .A1(n18536), .A2(n18489), .ZN(n18507) );
  AOI22_X1 U21556 ( .A1(n18643), .A2(n18507), .B1(n18649), .B2(n18531), .ZN(
        n18494) );
  NOR2_X1 U21557 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18490), .ZN(
        n18492) );
  NOR2_X1 U21558 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18536), .ZN(
        n18491) );
  AOI22_X1 U21559 ( .A1(n18648), .A2(n18492), .B1(n18646), .B2(n18491), .ZN(
        n18509) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18509), .B1(
        n18644), .B2(n18508), .ZN(n18493) );
  OAI211_X1 U21561 ( .C1(n18652), .C2(n18538), .A(n18494), .B(n18493), .ZN(
        P3_U2940) );
  AOI22_X1 U21562 ( .A1(n18653), .A2(n18507), .B1(n18654), .B2(n18531), .ZN(
        n18496) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18509), .B1(
        n18655), .B2(n18508), .ZN(n18495) );
  OAI211_X1 U21564 ( .C1(n18658), .C2(n18538), .A(n18496), .B(n18495), .ZN(
        P3_U2941) );
  AOI22_X1 U21565 ( .A1(n18660), .A2(n18531), .B1(n18659), .B2(n18507), .ZN(
        n18498) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18509), .B1(
        n18661), .B2(n18508), .ZN(n18497) );
  OAI211_X1 U21567 ( .C1(n18664), .C2(n18538), .A(n18498), .B(n18497), .ZN(
        P3_U2942) );
  AOI22_X1 U21568 ( .A1(n18667), .A2(n18531), .B1(n18665), .B2(n18507), .ZN(
        n18500) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18509), .B1(
        n18666), .B2(n18508), .ZN(n18499) );
  OAI211_X1 U21570 ( .C1(n18670), .C2(n18538), .A(n18500), .B(n18499), .ZN(
        P3_U2943) );
  AOI22_X1 U21571 ( .A1(n18673), .A2(n18531), .B1(n18672), .B2(n18507), .ZN(
        n18502) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18509), .B1(
        n18671), .B2(n18508), .ZN(n18501) );
  OAI211_X1 U21573 ( .C1(n18676), .C2(n18538), .A(n18502), .B(n18501), .ZN(
        P3_U2944) );
  AOI22_X1 U21574 ( .A1(n18678), .A2(n18531), .B1(n18677), .B2(n18507), .ZN(
        n18504) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18509), .B1(
        n18679), .B2(n18508), .ZN(n18503) );
  OAI211_X1 U21576 ( .C1(n18682), .C2(n18538), .A(n18504), .B(n18503), .ZN(
        P3_U2945) );
  AOI22_X1 U21577 ( .A1(n18684), .A2(n18531), .B1(n18683), .B2(n18507), .ZN(
        n18506) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18509), .B1(
        n18685), .B2(n18508), .ZN(n18505) );
  OAI211_X1 U21579 ( .C1(n18688), .C2(n18538), .A(n18506), .B(n18505), .ZN(
        P3_U2946) );
  AOI22_X1 U21580 ( .A1(n18691), .A2(n18531), .B1(n18690), .B2(n18507), .ZN(
        n18511) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18509), .B1(
        n18694), .B2(n18508), .ZN(n18510) );
  OAI211_X1 U21582 ( .C1(n18698), .C2(n18538), .A(n18511), .B(n18510), .ZN(
        P3_U2947) );
  NAND2_X1 U21583 ( .A1(n18559), .A2(n18512), .ZN(n18535) );
  AOI22_X1 U21584 ( .A1(n18643), .A2(n18530), .B1(n18649), .B2(n18554), .ZN(
        n18517) );
  INV_X1 U21585 ( .A(n18535), .ZN(n18614) );
  NOR2_X1 U21586 ( .A1(n18531), .A2(n18554), .ZN(n18514) );
  AOI221_X1 U21587 ( .B1(n18514), .B2(n18538), .C1(n18513), .C2(n18538), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18515) );
  OAI21_X1 U21588 ( .B1(n18614), .B2(n18515), .A(n18564), .ZN(n18532) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18532), .B1(
        n18644), .B2(n18531), .ZN(n18516) );
  OAI211_X1 U21590 ( .C1(n18652), .C2(n18535), .A(n18517), .B(n18516), .ZN(
        P3_U2948) );
  AOI22_X1 U21591 ( .A1(n18653), .A2(n18530), .B1(n18654), .B2(n18554), .ZN(
        n18519) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18532), .B1(
        n18655), .B2(n18531), .ZN(n18518) );
  OAI211_X1 U21593 ( .C1(n18658), .C2(n18535), .A(n18519), .B(n18518), .ZN(
        P3_U2949) );
  AOI22_X1 U21594 ( .A1(n18660), .A2(n18554), .B1(n18659), .B2(n18530), .ZN(
        n18521) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18532), .B1(
        n18661), .B2(n18531), .ZN(n18520) );
  OAI211_X1 U21596 ( .C1(n18664), .C2(n18535), .A(n18521), .B(n18520), .ZN(
        P3_U2950) );
  AOI22_X1 U21597 ( .A1(n18666), .A2(n18531), .B1(n18665), .B2(n18530), .ZN(
        n18523) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18532), .B1(
        n18667), .B2(n18554), .ZN(n18522) );
  OAI211_X1 U21599 ( .C1(n18670), .C2(n18535), .A(n18523), .B(n18522), .ZN(
        P3_U2951) );
  AOI22_X1 U21600 ( .A1(n18673), .A2(n18554), .B1(n18672), .B2(n18530), .ZN(
        n18525) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18532), .B1(
        n18671), .B2(n18531), .ZN(n18524) );
  OAI211_X1 U21602 ( .C1(n18676), .C2(n18535), .A(n18525), .B(n18524), .ZN(
        P3_U2952) );
  AOI22_X1 U21603 ( .A1(n18679), .A2(n18531), .B1(n18677), .B2(n18530), .ZN(
        n18527) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18532), .B1(
        n18678), .B2(n18554), .ZN(n18526) );
  OAI211_X1 U21605 ( .C1(n18682), .C2(n18535), .A(n18527), .B(n18526), .ZN(
        P3_U2953) );
  AOI22_X1 U21606 ( .A1(n18685), .A2(n18531), .B1(n18683), .B2(n18530), .ZN(
        n18529) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18532), .B1(
        n18684), .B2(n18554), .ZN(n18528) );
  OAI211_X1 U21608 ( .C1(n18688), .C2(n18535), .A(n18529), .B(n18528), .ZN(
        P3_U2954) );
  AOI22_X1 U21609 ( .A1(n18694), .A2(n18531), .B1(n18690), .B2(n18530), .ZN(
        n18534) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18532), .B1(
        n18691), .B2(n18554), .ZN(n18533) );
  OAI211_X1 U21611 ( .C1(n18698), .C2(n18535), .A(n18534), .B(n18533), .ZN(
        P3_U2955) );
  NOR2_X2 U21612 ( .A1(n18537), .A2(n18536), .ZN(n18638) );
  INV_X1 U21613 ( .A(n18638), .ZN(n18558) );
  NAND2_X1 U21614 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18559), .ZN(
        n18586) );
  NOR2_X1 U21615 ( .A1(n18589), .A2(n18586), .ZN(n18553) );
  INV_X1 U21616 ( .A(n18538), .ZN(n18581) );
  AOI22_X1 U21617 ( .A1(n18643), .A2(n18553), .B1(n18649), .B2(n18581), .ZN(
        n18540) );
  OAI211_X1 U21618 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18648), .A(
        n18646), .B(n18559), .ZN(n18555) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18555), .B1(
        n18644), .B2(n18554), .ZN(n18539) );
  OAI211_X1 U21620 ( .C1(n18652), .C2(n18558), .A(n18540), .B(n18539), .ZN(
        P3_U2956) );
  AOI22_X1 U21621 ( .A1(n18655), .A2(n18554), .B1(n18653), .B2(n18553), .ZN(
        n18542) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18555), .B1(
        n18654), .B2(n18581), .ZN(n18541) );
  OAI211_X1 U21623 ( .C1(n18658), .C2(n18558), .A(n18542), .B(n18541), .ZN(
        P3_U2957) );
  AOI22_X1 U21624 ( .A1(n18659), .A2(n18553), .B1(n18661), .B2(n18554), .ZN(
        n18544) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18555), .B1(
        n18660), .B2(n18581), .ZN(n18543) );
  OAI211_X1 U21626 ( .C1(n18664), .C2(n18558), .A(n18544), .B(n18543), .ZN(
        P3_U2958) );
  AOI22_X1 U21627 ( .A1(n18666), .A2(n18554), .B1(n18665), .B2(n18553), .ZN(
        n18546) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18555), .B1(
        n18667), .B2(n18581), .ZN(n18545) );
  OAI211_X1 U21629 ( .C1(n18670), .C2(n18558), .A(n18546), .B(n18545), .ZN(
        P3_U2959) );
  AOI22_X1 U21630 ( .A1(n18673), .A2(n18581), .B1(n18672), .B2(n18553), .ZN(
        n18548) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18555), .B1(
        n18671), .B2(n18554), .ZN(n18547) );
  OAI211_X1 U21632 ( .C1(n18676), .C2(n18558), .A(n18548), .B(n18547), .ZN(
        P3_U2960) );
  AOI22_X1 U21633 ( .A1(n18678), .A2(n18581), .B1(n18677), .B2(n18553), .ZN(
        n18550) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18555), .B1(
        n18679), .B2(n18554), .ZN(n18549) );
  OAI211_X1 U21635 ( .C1(n18682), .C2(n18558), .A(n18550), .B(n18549), .ZN(
        P3_U2961) );
  AOI22_X1 U21636 ( .A1(n18684), .A2(n18581), .B1(n18683), .B2(n18553), .ZN(
        n18552) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18555), .B1(
        n18685), .B2(n18554), .ZN(n18551) );
  OAI211_X1 U21638 ( .C1(n18688), .C2(n18558), .A(n18552), .B(n18551), .ZN(
        P3_U2962) );
  AOI22_X1 U21639 ( .A1(n18691), .A2(n18581), .B1(n18690), .B2(n18553), .ZN(
        n18557) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18555), .B1(
        n18694), .B2(n18554), .ZN(n18556) );
  OAI211_X1 U21641 ( .C1(n18698), .C2(n18558), .A(n18557), .B(n18556), .ZN(
        P3_U2963) );
  INV_X1 U21642 ( .A(n18647), .ZN(n18588) );
  NOR2_X2 U21643 ( .A1(n18588), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18693) );
  NAND2_X1 U21644 ( .A1(n18558), .A2(n18584), .ZN(n18620) );
  INV_X1 U21645 ( .A(n18620), .ZN(n18560) );
  NOR2_X1 U21646 ( .A1(n18589), .A2(n18560), .ZN(n18579) );
  AOI22_X1 U21647 ( .A1(n18643), .A2(n18579), .B1(n18649), .B2(n18614), .ZN(
        n18566) );
  NAND2_X1 U21648 ( .A1(n18621), .A2(n18559), .ZN(n18561) );
  OAI21_X1 U21649 ( .B1(n18562), .B2(n18561), .A(n18560), .ZN(n18563) );
  OAI211_X1 U21650 ( .C1(n18693), .C2(n18862), .A(n18564), .B(n18563), .ZN(
        n18580) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18580), .B1(
        n18644), .B2(n18581), .ZN(n18565) );
  OAI211_X1 U21652 ( .C1(n18652), .C2(n18584), .A(n18566), .B(n18565), .ZN(
        P3_U2964) );
  AOI22_X1 U21653 ( .A1(n18655), .A2(n18581), .B1(n18653), .B2(n18579), .ZN(
        n18568) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18580), .B1(
        n18654), .B2(n18614), .ZN(n18567) );
  OAI211_X1 U21655 ( .C1(n18658), .C2(n18584), .A(n18568), .B(n18567), .ZN(
        P3_U2965) );
  AOI22_X1 U21656 ( .A1(n18659), .A2(n18579), .B1(n18661), .B2(n18581), .ZN(
        n18570) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18580), .B1(
        n18660), .B2(n18614), .ZN(n18569) );
  OAI211_X1 U21658 ( .C1(n18664), .C2(n18584), .A(n18570), .B(n18569), .ZN(
        P3_U2966) );
  AOI22_X1 U21659 ( .A1(n18666), .A2(n18581), .B1(n18665), .B2(n18579), .ZN(
        n18572) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18580), .B1(
        n18667), .B2(n18614), .ZN(n18571) );
  OAI211_X1 U21661 ( .C1(n18670), .C2(n18584), .A(n18572), .B(n18571), .ZN(
        P3_U2967) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18580), .B1(
        n18672), .B2(n18579), .ZN(n18574) );
  AOI22_X1 U21663 ( .A1(n18673), .A2(n18614), .B1(n18671), .B2(n18581), .ZN(
        n18573) );
  OAI211_X1 U21664 ( .C1(n18676), .C2(n18584), .A(n18574), .B(n18573), .ZN(
        P3_U2968) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18580), .B1(
        n18677), .B2(n18579), .ZN(n18576) );
  AOI22_X1 U21666 ( .A1(n18679), .A2(n18581), .B1(n18678), .B2(n18614), .ZN(
        n18575) );
  OAI211_X1 U21667 ( .C1(n18682), .C2(n18584), .A(n18576), .B(n18575), .ZN(
        P3_U2969) );
  AOI22_X1 U21668 ( .A1(n18685), .A2(n18581), .B1(n18683), .B2(n18579), .ZN(
        n18578) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18580), .B1(
        n18684), .B2(n18614), .ZN(n18577) );
  OAI211_X1 U21670 ( .C1(n18688), .C2(n18584), .A(n18578), .B(n18577), .ZN(
        P3_U2970) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18580), .B1(
        n18690), .B2(n18579), .ZN(n18583) );
  AOI22_X1 U21672 ( .A1(n18694), .A2(n18581), .B1(n18691), .B2(n18614), .ZN(
        n18582) );
  OAI211_X1 U21673 ( .C1(n18698), .C2(n18584), .A(n18583), .B(n18582), .ZN(
        P3_U2971) );
  OAI22_X1 U21674 ( .A1(n18587), .A2(n18586), .B1(n18588), .B2(n18585), .ZN(
        n18606) );
  NOR2_X1 U21675 ( .A1(n18589), .A2(n18588), .ZN(n18613) );
  AOI22_X1 U21676 ( .A1(n18643), .A2(n18613), .B1(n18649), .B2(n18638), .ZN(
        n18592) );
  INV_X1 U21677 ( .A(n18652), .ZN(n18590) );
  AOI22_X1 U21678 ( .A1(n18692), .A2(n18590), .B1(n18644), .B2(n18614), .ZN(
        n18591) );
  OAI211_X1 U21679 ( .C1(n18593), .C2(n18606), .A(n18592), .B(n18591), .ZN(
        P3_U2972) );
  AOI22_X1 U21680 ( .A1(n18655), .A2(n18614), .B1(n18653), .B2(n18613), .ZN(
        n18596) );
  INV_X1 U21681 ( .A(n18658), .ZN(n18594) );
  AOI22_X1 U21682 ( .A1(n18692), .A2(n18594), .B1(n18654), .B2(n18638), .ZN(
        n18595) );
  OAI211_X1 U21683 ( .C1(n18597), .C2(n18606), .A(n18596), .B(n18595), .ZN(
        P3_U2973) );
  AOI22_X1 U21684 ( .A1(n18659), .A2(n18613), .B1(n18661), .B2(n18614), .ZN(
        n18600) );
  INV_X1 U21685 ( .A(n18664), .ZN(n18598) );
  AOI22_X1 U21686 ( .A1(n18692), .A2(n18598), .B1(n18660), .B2(n18638), .ZN(
        n18599) );
  OAI211_X1 U21687 ( .C1(n18601), .C2(n18606), .A(n18600), .B(n18599), .ZN(
        P3_U2974) );
  AOI22_X1 U21688 ( .A1(n18666), .A2(n18614), .B1(n18665), .B2(n18613), .ZN(
        n18604) );
  INV_X1 U21689 ( .A(n18670), .ZN(n18602) );
  AOI22_X1 U21690 ( .A1(n18692), .A2(n18602), .B1(n18667), .B2(n18638), .ZN(
        n18603) );
  OAI211_X1 U21691 ( .C1(n18605), .C2(n18606), .A(n18604), .B(n18603), .ZN(
        P3_U2975) );
  AOI22_X1 U21692 ( .A1(n18673), .A2(n18638), .B1(n18672), .B2(n18613), .ZN(
        n18608) );
  INV_X1 U21693 ( .A(n18606), .ZN(n18615) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18615), .B1(
        n18671), .B2(n18614), .ZN(n18607) );
  OAI211_X1 U21695 ( .C1(n18618), .C2(n18676), .A(n18608), .B(n18607), .ZN(
        P3_U2976) );
  AOI22_X1 U21696 ( .A1(n18679), .A2(n18614), .B1(n18677), .B2(n18613), .ZN(
        n18610) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18615), .B1(
        n18678), .B2(n18638), .ZN(n18609) );
  OAI211_X1 U21698 ( .C1(n18618), .C2(n18682), .A(n18610), .B(n18609), .ZN(
        P3_U2977) );
  AOI22_X1 U21699 ( .A1(n18684), .A2(n18638), .B1(n18683), .B2(n18613), .ZN(
        n18612) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18615), .B1(
        n18685), .B2(n18614), .ZN(n18611) );
  OAI211_X1 U21701 ( .C1(n18618), .C2(n18688), .A(n18612), .B(n18611), .ZN(
        P3_U2978) );
  AOI22_X1 U21702 ( .A1(n18691), .A2(n18638), .B1(n18690), .B2(n18613), .ZN(
        n18617) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18615), .B1(
        n18694), .B2(n18614), .ZN(n18616) );
  OAI211_X1 U21704 ( .C1(n18618), .C2(n18698), .A(n18617), .B(n18616), .ZN(
        P3_U2979) );
  AND2_X1 U21705 ( .A1(n18761), .A2(n18622), .ZN(n18637) );
  AOI22_X1 U21706 ( .A1(n18643), .A2(n18637), .B1(n18649), .B2(n18693), .ZN(
        n18624) );
  OAI221_X1 U21707 ( .B1(n18622), .B2(n18621), .C1(n18622), .C2(n18620), .A(
        n18619), .ZN(n18639) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18639), .B1(
        n18644), .B2(n18638), .ZN(n18623) );
  OAI211_X1 U21709 ( .C1(n18652), .C2(n18642), .A(n18624), .B(n18623), .ZN(
        P3_U2980) );
  AOI22_X1 U21710 ( .A1(n18653), .A2(n18637), .B1(n18654), .B2(n18693), .ZN(
        n18626) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18639), .B1(
        n18655), .B2(n18638), .ZN(n18625) );
  OAI211_X1 U21712 ( .C1(n18642), .C2(n18658), .A(n18626), .B(n18625), .ZN(
        P3_U2981) );
  AOI22_X1 U21713 ( .A1(n18660), .A2(n18693), .B1(n18659), .B2(n18637), .ZN(
        n18628) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18639), .B1(
        n18661), .B2(n18638), .ZN(n18627) );
  OAI211_X1 U21715 ( .C1(n18642), .C2(n18664), .A(n18628), .B(n18627), .ZN(
        P3_U2982) );
  AOI22_X1 U21716 ( .A1(n18666), .A2(n18638), .B1(n18665), .B2(n18637), .ZN(
        n18630) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18639), .B1(
        n18667), .B2(n18693), .ZN(n18629) );
  OAI211_X1 U21718 ( .C1(n18642), .C2(n18670), .A(n18630), .B(n18629), .ZN(
        P3_U2983) );
  AOI22_X1 U21719 ( .A1(n18673), .A2(n18693), .B1(n18672), .B2(n18637), .ZN(
        n18632) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18639), .B1(
        n18671), .B2(n18638), .ZN(n18631) );
  OAI211_X1 U21721 ( .C1(n18642), .C2(n18676), .A(n18632), .B(n18631), .ZN(
        P3_U2984) );
  AOI22_X1 U21722 ( .A1(n18678), .A2(n18693), .B1(n18677), .B2(n18637), .ZN(
        n18634) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18639), .B1(
        n18679), .B2(n18638), .ZN(n18633) );
  OAI211_X1 U21724 ( .C1(n18642), .C2(n18682), .A(n18634), .B(n18633), .ZN(
        P3_U2985) );
  AOI22_X1 U21725 ( .A1(n18684), .A2(n18693), .B1(n18683), .B2(n18637), .ZN(
        n18636) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18639), .B1(
        n18685), .B2(n18638), .ZN(n18635) );
  OAI211_X1 U21727 ( .C1(n18642), .C2(n18688), .A(n18636), .B(n18635), .ZN(
        P3_U2986) );
  AOI22_X1 U21728 ( .A1(n18694), .A2(n18638), .B1(n18690), .B2(n18637), .ZN(
        n18641) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18639), .B1(
        n18691), .B2(n18693), .ZN(n18640) );
  OAI211_X1 U21730 ( .C1(n18642), .C2(n18698), .A(n18641), .B(n18640), .ZN(
        P3_U2987) );
  AND2_X1 U21731 ( .A1(n18761), .A2(n18645), .ZN(n18689) );
  AOI22_X1 U21732 ( .A1(n18644), .A2(n18693), .B1(n18643), .B2(n18689), .ZN(
        n18651) );
  AOI22_X1 U21733 ( .A1(n18648), .A2(n18647), .B1(n18646), .B2(n18645), .ZN(
        n18695) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18695), .B1(
        n18692), .B2(n18649), .ZN(n18650) );
  OAI211_X1 U21735 ( .C1(n18699), .C2(n18652), .A(n18651), .B(n18650), .ZN(
        P3_U2988) );
  AOI22_X1 U21736 ( .A1(n18692), .A2(n18654), .B1(n18653), .B2(n18689), .ZN(
        n18657) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18695), .B1(
        n18655), .B2(n18693), .ZN(n18656) );
  OAI211_X1 U21738 ( .C1(n18699), .C2(n18658), .A(n18657), .B(n18656), .ZN(
        P3_U2989) );
  AOI22_X1 U21739 ( .A1(n18692), .A2(n18660), .B1(n18659), .B2(n18689), .ZN(
        n18663) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18695), .B1(
        n18661), .B2(n18693), .ZN(n18662) );
  OAI211_X1 U21741 ( .C1(n18699), .C2(n18664), .A(n18663), .B(n18662), .ZN(
        P3_U2990) );
  AOI22_X1 U21742 ( .A1(n18666), .A2(n18693), .B1(n18665), .B2(n18689), .ZN(
        n18669) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18695), .B1(
        n18692), .B2(n18667), .ZN(n18668) );
  OAI211_X1 U21744 ( .C1(n18699), .C2(n18670), .A(n18669), .B(n18668), .ZN(
        P3_U2991) );
  AOI22_X1 U21745 ( .A1(n18672), .A2(n18689), .B1(n18671), .B2(n18693), .ZN(
        n18675) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18695), .B1(
        n18692), .B2(n18673), .ZN(n18674) );
  OAI211_X1 U21747 ( .C1(n18699), .C2(n18676), .A(n18675), .B(n18674), .ZN(
        P3_U2992) );
  AOI22_X1 U21748 ( .A1(n18692), .A2(n18678), .B1(n18677), .B2(n18689), .ZN(
        n18681) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18695), .B1(
        n18679), .B2(n18693), .ZN(n18680) );
  OAI211_X1 U21750 ( .C1(n18699), .C2(n18682), .A(n18681), .B(n18680), .ZN(
        P3_U2993) );
  AOI22_X1 U21751 ( .A1(n18692), .A2(n18684), .B1(n18683), .B2(n18689), .ZN(
        n18687) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18695), .B1(
        n18685), .B2(n18693), .ZN(n18686) );
  OAI211_X1 U21753 ( .C1(n18699), .C2(n18688), .A(n18687), .B(n18686), .ZN(
        P3_U2994) );
  AOI22_X1 U21754 ( .A1(n18692), .A2(n18691), .B1(n18690), .B2(n18689), .ZN(
        n18697) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18695), .B1(
        n18694), .B2(n18693), .ZN(n18696) );
  OAI211_X1 U21756 ( .C1(n18699), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        P3_U2995) );
  OAI22_X1 U21757 ( .A1(n18703), .A2(n18702), .B1(n18701), .B2(n18700), .ZN(
        n18704) );
  AOI221_X1 U21758 ( .B1(n18707), .B2(n18706), .C1(n18705), .C2(n18706), .A(
        n18704), .ZN(n18907) );
  AOI211_X1 U21759 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18738), .A(
        n18709), .B(n18708), .ZN(n18749) );
  OAI21_X1 U21760 ( .B1(n18712), .B2(n18711), .A(n18710), .ZN(n18730) );
  AOI22_X1 U21761 ( .A1(n18878), .A2(n18731), .B1(n18730), .B2(n18713), .ZN(
        n18714) );
  OAI21_X1 U21762 ( .B1(n18715), .B2(n18716), .A(n18714), .ZN(n18867) );
  NOR2_X1 U21763 ( .A1(n18738), .A2(n18867), .ZN(n18721) );
  OAI21_X1 U21764 ( .B1(n18893), .B2(n18723), .A(n18716), .ZN(n18733) );
  INV_X1 U21765 ( .A(n18733), .ZN(n18719) );
  NOR2_X1 U21766 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18717), .ZN(
        n18718) );
  OAI22_X1 U21767 ( .A1(n18719), .A2(n18732), .B1(n18718), .B2(n18736), .ZN(
        n18864) );
  NAND2_X1 U21768 ( .A1(n18868), .A2(n18864), .ZN(n18720) );
  OAI22_X1 U21769 ( .A1(n18721), .A2(n18868), .B1(n18738), .B2(n18720), .ZN(
        n18745) );
  NAND2_X1 U21770 ( .A1(n18723), .A2(n18722), .ZN(n18724) );
  AOI22_X1 U21771 ( .A1(n18882), .A2(n18724), .B1(n18885), .B2(n18733), .ZN(
        n18879) );
  AOI22_X1 U21772 ( .A1(n18726), .A2(n18725), .B1(n18724), .B2(n18893), .ZN(
        n18886) );
  AOI222_X1 U21773 ( .A1(n18879), .A2(n18886), .B1(n18879), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18886), .C2(n18727), .ZN(
        n18729) );
  INV_X1 U21774 ( .A(n18738), .ZN(n18737) );
  AOI21_X1 U21775 ( .B1(n18729), .B2(n18737), .A(n18728), .ZN(n18740) );
  NAND3_X1 U21776 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18731), .A3(
        n18730), .ZN(n18735) );
  OAI211_X1 U21777 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18733), .B(n18732), .ZN(
        n18734) );
  OAI211_X1 U21778 ( .C1(n18874), .C2(n18736), .A(n18735), .B(n18734), .ZN(
        n18876) );
  AOI22_X1 U21779 ( .A1(n18738), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18876), .B2(n18737), .ZN(n18741) );
  OR2_X1 U21780 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18741), .ZN(
        n18739) );
  AOI221_X1 U21781 ( .B1(n18740), .B2(n18739), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18741), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18744) );
  OAI21_X1 U21782 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18741), .ZN(n18743) );
  AOI222_X1 U21783 ( .A1(n18745), .A2(n18744), .B1(n18745), .B2(n18743), .C1(
        n18744), .C2(n18742), .ZN(n18748) );
  OAI21_X1 U21784 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18746), .ZN(n18747) );
  NAND4_X1 U21785 ( .A1(n18907), .A2(n18749), .A3(n18748), .A4(n18747), .ZN(
        n18758) );
  AOI211_X1 U21786 ( .C1(n18752), .C2(n18751), .A(n18750), .B(n18758), .ZN(
        n18860) );
  AOI21_X1 U21787 ( .B1(n18912), .B2(n18753), .A(n18860), .ZN(n18762) );
  NOR2_X1 U21788 ( .A1(n18754), .A2(n18761), .ZN(n18757) );
  NAND2_X1 U21789 ( .A1(n18912), .A2(n17492), .ZN(n18766) );
  INV_X1 U21790 ( .A(n18766), .ZN(n18755) );
  AOI211_X1 U21791 ( .C1(n18887), .C2(n18920), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18755), .ZN(n18756) );
  AOI211_X1 U21792 ( .C1(n18910), .C2(n18758), .A(n18757), .B(n18756), .ZN(
        n18759) );
  OAI221_X1 U21793 ( .B1(n18859), .B2(n18762), .C1(n18859), .C2(n18760), .A(
        n18759), .ZN(P3_U2996) );
  NOR4_X1 U21794 ( .A1(n18859), .A2(n18871), .A3(n18918), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18769) );
  INV_X1 U21795 ( .A(n18769), .ZN(n18765) );
  NAND3_X1 U21796 ( .A1(n18763), .A2(n18762), .A3(n18761), .ZN(n18764) );
  NAND4_X1 U21797 ( .A1(n18767), .A2(n18766), .A3(n18765), .A4(n18764), .ZN(
        P3_U2997) );
  OAI21_X1 U21798 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18768), .ZN(n18770) );
  AOI21_X1 U21799 ( .B1(n18771), .B2(n18770), .A(n18769), .ZN(P3_U2998) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18772), .ZN(
        P3_U2999) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18772), .ZN(
        P3_U3000) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18772), .ZN(
        P3_U3001) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18772), .ZN(
        P3_U3002) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18772), .ZN(
        P3_U3003) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18772), .ZN(
        P3_U3004) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18772), .ZN(
        P3_U3005) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18772), .ZN(
        P3_U3006) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18772), .ZN(
        P3_U3007) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18772), .ZN(
        P3_U3008) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18772), .ZN(
        P3_U3009) );
  AND2_X1 U21811 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18772), .ZN(
        P3_U3010) );
  AND2_X1 U21812 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18772), .ZN(
        P3_U3011) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18772), .ZN(
        P3_U3012) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18772), .ZN(
        P3_U3013) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18772), .ZN(
        P3_U3014) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18772), .ZN(
        P3_U3015) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18772), .ZN(
        P3_U3016) );
  AND2_X1 U21818 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18772), .ZN(
        P3_U3017) );
  AND2_X1 U21819 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18772), .ZN(
        P3_U3018) );
  AND2_X1 U21820 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18772), .ZN(
        P3_U3019) );
  AND2_X1 U21821 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18772), .ZN(
        P3_U3020) );
  AND2_X1 U21822 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18772), .ZN(P3_U3021) );
  AND2_X1 U21823 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18772), .ZN(P3_U3022) );
  AND2_X1 U21824 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18772), .ZN(P3_U3023) );
  AND2_X1 U21825 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18772), .ZN(P3_U3024) );
  AND2_X1 U21826 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18772), .ZN(P3_U3025) );
  AND2_X1 U21827 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18772), .ZN(P3_U3026) );
  AND2_X1 U21828 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18772), .ZN(P3_U3027) );
  AND2_X1 U21829 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18772), .ZN(P3_U3028) );
  INV_X1 U21830 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18777) );
  NOR2_X1 U21831 ( .A1(n18789), .A2(n20782), .ZN(n18785) );
  INV_X1 U21832 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18773) );
  NOR2_X1 U21833 ( .A1(n18785), .A2(n18773), .ZN(n18779) );
  OAI21_X1 U21834 ( .B1(n18777), .B2(n20782), .A(n18779), .ZN(n18774) );
  AOI22_X1 U21835 ( .A1(n18787), .A2(n18789), .B1(n18926), .B2(n18774), .ZN(
        n18775) );
  NAND3_X1 U21836 ( .A1(NA), .A2(n18787), .A3(n18777), .ZN(n18782) );
  OAI211_X1 U21837 ( .C1(n18918), .C2(n18776), .A(n18775), .B(n18782), .ZN(
        P3_U3029) );
  NOR2_X1 U21838 ( .A1(n18777), .A2(n20782), .ZN(n18778) );
  AOI22_X1 U21839 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18779), .B1(n18778), 
        .B2(n18789), .ZN(n18780) );
  NAND2_X1 U21840 ( .A1(n18912), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18783) );
  NAND3_X1 U21841 ( .A1(n18780), .A2(n18915), .A3(n18783), .ZN(P3_U3030) );
  INV_X1 U21842 ( .A(n18783), .ZN(n18781) );
  AOI21_X1 U21843 ( .B1(n18787), .B2(n18782), .A(n18781), .ZN(n18788) );
  OAI22_X1 U21844 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18783), .ZN(n18784) );
  OAI22_X1 U21845 ( .A1(n18785), .A2(n18784), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18786) );
  OAI22_X1 U21846 ( .A1(n18788), .A2(n18789), .B1(n18787), .B2(n18786), .ZN(
        P3_U3031) );
  OAI222_X1 U21847 ( .A1(n18895), .A2(n18850), .B1(n18790), .B2(n18925), .C1(
        n18791), .C2(n18846), .ZN(P3_U3032) );
  INV_X1 U21848 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18793) );
  OAI222_X1 U21849 ( .A1(n18846), .A2(n18793), .B1(n18792), .B2(n18925), .C1(
        n18791), .C2(n18850), .ZN(P3_U3033) );
  OAI222_X1 U21850 ( .A1(n18846), .A2(n18795), .B1(n18794), .B2(n18925), .C1(
        n18793), .C2(n18850), .ZN(P3_U3034) );
  INV_X1 U21851 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18797) );
  OAI222_X1 U21852 ( .A1(n18846), .A2(n18797), .B1(n18796), .B2(n18925), .C1(
        n18795), .C2(n18850), .ZN(P3_U3035) );
  OAI222_X1 U21853 ( .A1(n18846), .A2(n18799), .B1(n18798), .B2(n18925), .C1(
        n18797), .C2(n18850), .ZN(P3_U3036) );
  OAI222_X1 U21854 ( .A1(n18846), .A2(n18801), .B1(n18800), .B2(n18925), .C1(
        n18799), .C2(n18850), .ZN(P3_U3037) );
  OAI222_X1 U21855 ( .A1(n18846), .A2(n18804), .B1(n18802), .B2(n18925), .C1(
        n18801), .C2(n18850), .ZN(P3_U3038) );
  OAI222_X1 U21856 ( .A1(n18804), .A2(n18850), .B1(n18803), .B2(n18925), .C1(
        n18805), .C2(n18846), .ZN(P3_U3039) );
  OAI222_X1 U21857 ( .A1(n18846), .A2(n18807), .B1(n18806), .B2(n18925), .C1(
        n18805), .C2(n18850), .ZN(P3_U3040) );
  OAI222_X1 U21858 ( .A1(n18846), .A2(n18809), .B1(n18808), .B2(n18925), .C1(
        n18807), .C2(n18850), .ZN(P3_U3041) );
  OAI222_X1 U21859 ( .A1(n18846), .A2(n18812), .B1(n18810), .B2(n18925), .C1(
        n18809), .C2(n18850), .ZN(P3_U3042) );
  OAI222_X1 U21860 ( .A1(n18812), .A2(n18850), .B1(n18811), .B2(n18925), .C1(
        n18813), .C2(n18846), .ZN(P3_U3043) );
  INV_X1 U21861 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18816) );
  OAI222_X1 U21862 ( .A1(n18846), .A2(n18816), .B1(n18814), .B2(n18925), .C1(
        n18813), .C2(n18850), .ZN(P3_U3044) );
  OAI222_X1 U21863 ( .A1(n18816), .A2(n18850), .B1(n18815), .B2(n18925), .C1(
        n18817), .C2(n18846), .ZN(P3_U3045) );
  OAI222_X1 U21864 ( .A1(n18846), .A2(n18819), .B1(n18818), .B2(n18925), .C1(
        n18817), .C2(n18850), .ZN(P3_U3046) );
  OAI222_X1 U21865 ( .A1(n18846), .A2(n20986), .B1(n18820), .B2(n18925), .C1(
        n18819), .C2(n18850), .ZN(P3_U3047) );
  OAI222_X1 U21866 ( .A1(n18846), .A2(n18822), .B1(n18821), .B2(n18925), .C1(
        n20986), .C2(n18850), .ZN(P3_U3048) );
  OAI222_X1 U21867 ( .A1(n18846), .A2(n18825), .B1(n18823), .B2(n18925), .C1(
        n18822), .C2(n18850), .ZN(P3_U3049) );
  INV_X1 U21868 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18826) );
  OAI222_X1 U21869 ( .A1(n18825), .A2(n18850), .B1(n18824), .B2(n18925), .C1(
        n18826), .C2(n18846), .ZN(P3_U3050) );
  OAI222_X1 U21870 ( .A1(n18846), .A2(n18829), .B1(n18827), .B2(n18925), .C1(
        n18826), .C2(n18850), .ZN(P3_U3051) );
  OAI222_X1 U21871 ( .A1(n18829), .A2(n18850), .B1(n18828), .B2(n18925), .C1(
        n18830), .C2(n18846), .ZN(P3_U3052) );
  OAI222_X1 U21872 ( .A1(n18846), .A2(n18833), .B1(n18831), .B2(n18925), .C1(
        n18830), .C2(n18850), .ZN(P3_U3053) );
  OAI222_X1 U21873 ( .A1(n18833), .A2(n18850), .B1(n18832), .B2(n18925), .C1(
        n18834), .C2(n18846), .ZN(P3_U3054) );
  OAI222_X1 U21874 ( .A1(n18846), .A2(n18836), .B1(n18835), .B2(n18925), .C1(
        n18834), .C2(n18850), .ZN(P3_U3055) );
  INV_X1 U21875 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18838) );
  OAI222_X1 U21876 ( .A1(n18846), .A2(n18838), .B1(n18837), .B2(n18925), .C1(
        n18836), .C2(n18850), .ZN(P3_U3056) );
  OAI222_X1 U21877 ( .A1(n18846), .A2(n18840), .B1(n18839), .B2(n18925), .C1(
        n18838), .C2(n18850), .ZN(P3_U3057) );
  INV_X1 U21878 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18843) );
  OAI222_X1 U21879 ( .A1(n18846), .A2(n18843), .B1(n18841), .B2(n18925), .C1(
        n18840), .C2(n18850), .ZN(P3_U3058) );
  OAI222_X1 U21880 ( .A1(n18843), .A2(n18850), .B1(n18842), .B2(n18925), .C1(
        n18844), .C2(n18846), .ZN(P3_U3059) );
  OAI222_X1 U21881 ( .A1(n18846), .A2(n18849), .B1(n18845), .B2(n18925), .C1(
        n18844), .C2(n18850), .ZN(P3_U3060) );
  OAI222_X1 U21882 ( .A1(n18850), .A2(n18849), .B1(n18848), .B2(n18925), .C1(
        n18847), .C2(n18846), .ZN(P3_U3061) );
  OAI22_X1 U21883 ( .A1(n18926), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18925), .ZN(n18851) );
  INV_X1 U21884 ( .A(n18851), .ZN(P3_U3274) );
  OAI22_X1 U21885 ( .A1(n18926), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18925), .ZN(n18852) );
  INV_X1 U21886 ( .A(n18852), .ZN(P3_U3275) );
  OAI22_X1 U21887 ( .A1(n18926), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18925), .ZN(n18853) );
  INV_X1 U21888 ( .A(n18853), .ZN(P3_U3276) );
  OAI22_X1 U21889 ( .A1(n18926), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18925), .ZN(n18854) );
  INV_X1 U21890 ( .A(n18854), .ZN(P3_U3277) );
  OAI21_X1 U21891 ( .B1(n18858), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18856), 
        .ZN(n18855) );
  INV_X1 U21892 ( .A(n18855), .ZN(P3_U3280) );
  OAI21_X1 U21893 ( .B1(n18858), .B2(n18857), .A(n18856), .ZN(P3_U3281) );
  NOR2_X1 U21894 ( .A1(n18860), .A2(n18859), .ZN(n18863) );
  OAI21_X1 U21895 ( .B1(n18863), .B2(n18862), .A(n18861), .ZN(P3_U3282) );
  INV_X1 U21896 ( .A(n18891), .ZN(n18894) );
  NOR2_X1 U21897 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18928), .ZN(
        n18865) );
  AOI22_X1 U21898 ( .A1(n18887), .A2(n18866), .B1(n18865), .B2(n18864), .ZN(
        n18870) );
  AOI21_X1 U21899 ( .B1(n18889), .B2(n18867), .A(n18894), .ZN(n18869) );
  OAI22_X1 U21900 ( .A1(n18894), .A2(n18870), .B1(n18869), .B2(n18868), .ZN(
        P3_U3285) );
  NOR2_X1 U21901 ( .A1(n18871), .A2(n18890), .ZN(n18880) );
  OAI22_X1 U21902 ( .A1(n18873), .A2(n18872), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18881) );
  INV_X1 U21903 ( .A(n18881), .ZN(n18875) );
  AOI222_X1 U21904 ( .A1(n18876), .A2(n18889), .B1(n18880), .B2(n18875), .C1(
        n18887), .C2(n18874), .ZN(n18877) );
  AOI22_X1 U21905 ( .A1(n18894), .A2(n18878), .B1(n18877), .B2(n18891), .ZN(
        P3_U3288) );
  INV_X1 U21906 ( .A(n18879), .ZN(n18883) );
  AOI222_X1 U21907 ( .A1(n18883), .A2(n18889), .B1(n18887), .B2(n18882), .C1(
        n18881), .C2(n18880), .ZN(n18884) );
  AOI22_X1 U21908 ( .A1(n18894), .A2(n18885), .B1(n18884), .B2(n18891), .ZN(
        P3_U3289) );
  INV_X1 U21909 ( .A(n18886), .ZN(n18888) );
  AOI222_X1 U21910 ( .A1(n18890), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18889), 
        .B2(n18888), .C1(n18893), .C2(n18887), .ZN(n18892) );
  AOI22_X1 U21911 ( .A1(n18894), .A2(n18893), .B1(n18892), .B2(n18891), .ZN(
        P3_U3290) );
  AOI21_X1 U21912 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18896) );
  AOI22_X1 U21913 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18896), .B2(n18895), .ZN(n18898) );
  INV_X1 U21914 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18897) );
  AOI22_X1 U21915 ( .A1(n18899), .A2(n18898), .B1(n18897), .B2(n18902), .ZN(
        P3_U3292) );
  INV_X1 U21916 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18903) );
  NOR2_X1 U21917 ( .A1(n18902), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18900) );
  AOI22_X1 U21918 ( .A1(n18903), .A2(n18902), .B1(n18901), .B2(n18900), .ZN(
        P3_U3293) );
  INV_X1 U21919 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18904) );
  AOI22_X1 U21920 ( .A1(n18925), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18904), 
        .B2(n18926), .ZN(P3_U3294) );
  INV_X1 U21921 ( .A(n18905), .ZN(n18908) );
  NAND2_X1 U21922 ( .A1(n18908), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18906) );
  OAI21_X1 U21923 ( .B1(n18908), .B2(n18907), .A(n18906), .ZN(P3_U3295) );
  OAI22_X1 U21924 ( .A1(n18912), .A2(n18911), .B1(n18910), .B2(n18909), .ZN(
        n18913) );
  NOR2_X1 U21925 ( .A1(n18914), .A2(n18913), .ZN(n18924) );
  AOI21_X1 U21926 ( .B1(n18917), .B2(n18916), .A(n18915), .ZN(n18919) );
  OAI211_X1 U21927 ( .C1(n18929), .C2(n18919), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18918), .ZN(n18921) );
  AOI21_X1 U21928 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18921), .A(n18920), 
        .ZN(n18923) );
  NAND2_X1 U21929 ( .A1(n18924), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18922) );
  OAI21_X1 U21930 ( .B1(n18924), .B2(n18923), .A(n18922), .ZN(P3_U3296) );
  OAI22_X1 U21931 ( .A1(n18926), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18925), .ZN(n18927) );
  INV_X1 U21932 ( .A(n18927), .ZN(P3_U3297) );
  OAI21_X1 U21933 ( .B1(n18928), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18930), 
        .ZN(n18933) );
  OAI22_X1 U21934 ( .A1(n18933), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18930), 
        .B2(n18929), .ZN(n18931) );
  INV_X1 U21935 ( .A(n18931), .ZN(P3_U3298) );
  OAI21_X1 U21936 ( .B1(n18933), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18932), 
        .ZN(n18934) );
  INV_X1 U21937 ( .A(n18934), .ZN(P3_U3299) );
  INV_X1 U21938 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19802) );
  NAND2_X1 U21939 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19802), .ZN(n19795) );
  OR2_X1 U21940 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19792) );
  OAI21_X1 U21941 ( .B1(n19791), .B2(n19795), .A(n19792), .ZN(n19864) );
  AOI21_X1 U21942 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19864), .ZN(n18935) );
  INV_X1 U21943 ( .A(n18935), .ZN(P2_U2815) );
  INV_X1 U21944 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18937) );
  OAI22_X1 U21945 ( .A1(n21033), .A2(n18937), .B1(n19866), .B2(n18936), .ZN(
        P2_U2816) );
  INV_X1 U21946 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n18939) );
  AOI21_X1 U21947 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n18937), .A(n18940), 
        .ZN(n18938) );
  OAI22_X1 U21948 ( .A1(n19909), .A2(n18939), .B1(P2_STATE_REG_0__SCAN_IN), 
        .B2(n18938), .ZN(P2_U2817) );
  OAI21_X1 U21949 ( .B1(n18940), .B2(BS16), .A(n19864), .ZN(n19862) );
  OAI21_X1 U21950 ( .B1(n19864), .B2(n19467), .A(n19862), .ZN(P2_U2818) );
  NOR4_X1 U21951 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18944) );
  NOR4_X1 U21952 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18943) );
  NOR4_X1 U21953 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18942) );
  NOR4_X1 U21954 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18941) );
  NAND4_X1 U21955 ( .A1(n18944), .A2(n18943), .A3(n18942), .A4(n18941), .ZN(
        n18950) );
  NOR4_X1 U21956 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18948) );
  AOI211_X1 U21957 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18947) );
  NOR4_X1 U21958 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18946) );
  NOR4_X1 U21959 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18945) );
  NAND4_X1 U21960 ( .A1(n18948), .A2(n18947), .A3(n18946), .A4(n18945), .ZN(
        n18949) );
  NOR2_X1 U21961 ( .A1(n18950), .A2(n18949), .ZN(n18960) );
  INV_X1 U21962 ( .A(n18960), .ZN(n18958) );
  NOR2_X1 U21963 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18958), .ZN(n18953) );
  INV_X1 U21964 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18951) );
  AOI22_X1 U21965 ( .A1(n18953), .A2(n10738), .B1(n18958), .B2(n18951), .ZN(
        P2_U2820) );
  OR3_X1 U21966 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18957) );
  INV_X1 U21967 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18952) );
  AOI22_X1 U21968 ( .A1(n18953), .A2(n18957), .B1(n18952), .B2(n18958), .ZN(
        P2_U2821) );
  INV_X1 U21969 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19863) );
  NAND2_X1 U21970 ( .A1(n18953), .A2(n19863), .ZN(n18956) );
  OAI21_X1 U21971 ( .B1(n13003), .B2(n10738), .A(n18960), .ZN(n18954) );
  OAI21_X1 U21972 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18960), .A(n18954), 
        .ZN(n18955) );
  OAI221_X1 U21973 ( .B1(n18956), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18956), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18955), .ZN(P2_U2822) );
  INV_X1 U21974 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18959) );
  OAI221_X1 U21975 ( .B1(n18960), .B2(n18959), .C1(n18958), .C2(n18957), .A(
        n18956), .ZN(P2_U2823) );
  NOR2_X1 U21976 ( .A1(n18961), .A2(n18962), .ZN(n18963) );
  OAI22_X1 U21977 ( .A1(n18964), .A2(n18963), .B1(n19013), .B2(n18962), .ZN(
        n18969) );
  INV_X1 U21978 ( .A(n18965), .ZN(n18967) );
  AOI22_X1 U21979 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19109), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19116), .ZN(n18966) );
  OAI21_X1 U21980 ( .B1(n18967), .B2(n19112), .A(n18966), .ZN(n18968) );
  AOI211_X1 U21981 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n19110), .A(n18969), .B(
        n18968), .ZN(n18974) );
  NOR2_X1 U21982 ( .A1(n18970), .A2(n19127), .ZN(n18971) );
  AOI21_X1 U21983 ( .B1(n18972), .B2(n19122), .A(n18971), .ZN(n18973) );
  NAND2_X1 U21984 ( .A1(n18974), .A2(n18973), .ZN(P2_U2835) );
  NAND2_X1 U21985 ( .A1(n19118), .A2(n18975), .ZN(n18976) );
  XOR2_X1 U21986 ( .A(n18977), .B(n18976), .Z(n18987) );
  OAI21_X1 U21987 ( .B1(n19833), .B2(n19096), .A(n11494), .ZN(n18981) );
  OAI22_X1 U21988 ( .A1(n18979), .A2(n19112), .B1(n19084), .B2(n18978), .ZN(
        n18980) );
  AOI211_X1 U21989 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19110), .A(n18981), .B(
        n18980), .ZN(n18986) );
  OAI22_X1 U21990 ( .A1(n18983), .A2(n19090), .B1(n18982), .B2(n19127), .ZN(
        n18984) );
  INV_X1 U21991 ( .A(n18984), .ZN(n18985) );
  OAI211_X1 U21992 ( .C1(n19782), .C2(n18987), .A(n18986), .B(n18985), .ZN(
        P2_U2836) );
  NOR2_X1 U21993 ( .A1(n19102), .A2(n18988), .ZN(n19002) );
  XOR2_X1 U21994 ( .A(n19002), .B(n18989), .Z(n18999) );
  INV_X1 U21995 ( .A(n18990), .ZN(n18992) );
  AOI22_X1 U21996 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19109), .ZN(n18991) );
  OAI21_X1 U21997 ( .B1(n18992), .B2(n19112), .A(n18991), .ZN(n18993) );
  AOI211_X1 U21998 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19116), .A(n19115), 
        .B(n18993), .ZN(n18998) );
  OAI22_X1 U21999 ( .A1(n18995), .A2(n19090), .B1(n18994), .B2(n19127), .ZN(
        n18996) );
  INV_X1 U22000 ( .A(n18996), .ZN(n18997) );
  OAI211_X1 U22001 ( .C1(n19782), .C2(n18999), .A(n18998), .B(n18997), .ZN(
        P2_U2837) );
  INV_X1 U22002 ( .A(n19000), .ZN(n19006) );
  INV_X1 U22003 ( .A(n19001), .ZN(n19003) );
  OAI211_X1 U22004 ( .C1(n19003), .C2(n19014), .A(n19123), .B(n19002), .ZN(
        n19005) );
  AOI22_X1 U22005 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19109), .ZN(n19004) );
  OAI211_X1 U22006 ( .C1(n19006), .C2(n19112), .A(n19005), .B(n19004), .ZN(
        n19007) );
  AOI211_X1 U22007 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19116), .A(n19115), 
        .B(n19007), .ZN(n19012) );
  OAI22_X1 U22008 ( .A1(n19009), .A2(n19090), .B1(n19008), .B2(n19127), .ZN(
        n19010) );
  INV_X1 U22009 ( .A(n19010), .ZN(n19011) );
  OAI211_X1 U22010 ( .C1(n19014), .C2(n19013), .A(n19012), .B(n19011), .ZN(
        P2_U2838) );
  OAI21_X1 U22011 ( .B1(n19827), .B2(n19096), .A(n11494), .ZN(n19018) );
  OAI22_X1 U22012 ( .A1(n19016), .A2(n19112), .B1(n19015), .B2(n19097), .ZN(
        n19017) );
  AOI211_X1 U22013 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19109), .A(
        n19018), .B(n19017), .ZN(n19025) );
  NAND2_X1 U22014 ( .A1(n19118), .A2(n19019), .ZN(n19021) );
  XNOR2_X1 U22015 ( .A(n19021), .B(n19020), .ZN(n19023) );
  AOI22_X1 U22016 ( .A1(n19023), .A2(n19123), .B1(n19022), .B2(n19122), .ZN(
        n19024) );
  OAI211_X1 U22017 ( .C1(n19175), .C2(n19127), .A(n19025), .B(n19024), .ZN(
        P2_U2840) );
  NOR2_X1 U22018 ( .A1(n19102), .A2(n19026), .ZN(n19028) );
  XOR2_X1 U22019 ( .A(n19028), .B(n19027), .Z(n19037) );
  INV_X1 U22020 ( .A(n19029), .ZN(n19031) );
  AOI22_X1 U22021 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19109), .ZN(n19030) );
  OAI21_X1 U22022 ( .B1(n19031), .B2(n19112), .A(n19030), .ZN(n19032) );
  AOI211_X1 U22023 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19116), .A(n19115), 
        .B(n19032), .ZN(n19036) );
  INV_X1 U22024 ( .A(n19033), .ZN(n19178) );
  OAI22_X1 U22025 ( .A1(n19136), .A2(n19090), .B1(n19178), .B2(n19127), .ZN(
        n19034) );
  INV_X1 U22026 ( .A(n19034), .ZN(n19035) );
  OAI211_X1 U22027 ( .C1(n19782), .C2(n19037), .A(n19036), .B(n19035), .ZN(
        P2_U2841) );
  INV_X1 U22028 ( .A(n19038), .ZN(n19040) );
  AOI22_X1 U22029 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19109), .ZN(n19039) );
  OAI21_X1 U22030 ( .B1(n19040), .B2(n19112), .A(n19039), .ZN(n19041) );
  AOI211_X1 U22031 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19116), .A(n19115), 
        .B(n19041), .ZN(n19048) );
  NAND2_X1 U22032 ( .A1(n19118), .A2(n19042), .ZN(n19044) );
  XNOR2_X1 U22033 ( .A(n19044), .B(n19043), .ZN(n19046) );
  AOI22_X1 U22034 ( .A1(n19046), .A2(n19123), .B1(n19045), .B2(n19122), .ZN(
        n19047) );
  OAI211_X1 U22035 ( .C1(n19180), .C2(n19127), .A(n19048), .B(n19047), .ZN(
        P2_U2842) );
  NAND2_X1 U22036 ( .A1(n19118), .A2(n19049), .ZN(n19051) );
  XOR2_X1 U22037 ( .A(n19051), .B(n19050), .Z(n19059) );
  INV_X1 U22038 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19821) );
  INV_X1 U22039 ( .A(n19052), .ZN(n19053) );
  AOI22_X1 U22040 ( .A1(n19053), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19109), .ZN(n19054) );
  OAI211_X1 U22041 ( .C1(n19821), .C2(n19096), .A(n19054), .B(n19088), .ZN(
        n19057) );
  OAI22_X1 U22042 ( .A1(n19055), .A2(n19090), .B1(n19185), .B2(n19127), .ZN(
        n19056) );
  AOI211_X1 U22043 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19110), .A(n19057), .B(
        n19056), .ZN(n19058) );
  OAI21_X1 U22044 ( .B1(n19059), .B2(n19782), .A(n19058), .ZN(P2_U2844) );
  AOI22_X1 U22045 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19109), .ZN(n19060) );
  OAI21_X1 U22046 ( .B1(n19061), .B2(n19112), .A(n19060), .ZN(n19062) );
  AOI211_X1 U22047 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19116), .A(n19115), 
        .B(n19062), .ZN(n19069) );
  NOR2_X1 U22048 ( .A1(n19102), .A2(n19063), .ZN(n19065) );
  XNOR2_X1 U22049 ( .A(n19065), .B(n19064), .ZN(n19067) );
  AOI22_X1 U22050 ( .A1(n19067), .A2(n19123), .B1(n19066), .B2(n19122), .ZN(
        n19068) );
  OAI211_X1 U22051 ( .C1(n19188), .C2(n19127), .A(n19069), .B(n19068), .ZN(
        P2_U2845) );
  NAND2_X1 U22052 ( .A1(n19118), .A2(n19070), .ZN(n19072) );
  XOR2_X1 U22053 ( .A(n19072), .B(n19071), .Z(n19079) );
  AOI22_X1 U22054 ( .A1(n19073), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19109), .ZN(n19074) );
  OAI211_X1 U22055 ( .C1(n20975), .C2(n19096), .A(n19074), .B(n19088), .ZN(
        n19077) );
  OAI22_X1 U22056 ( .A1(n19075), .A2(n19090), .B1(n19191), .B2(n19127), .ZN(
        n19076) );
  AOI211_X1 U22057 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19110), .A(n19077), .B(
        n19076), .ZN(n19078) );
  OAI21_X1 U22058 ( .B1(n19079), .B2(n19782), .A(n19078), .ZN(P2_U2846) );
  NAND2_X1 U22059 ( .A1(n19118), .A2(n19080), .ZN(n19082) );
  XOR2_X1 U22060 ( .A(n19082), .B(n19081), .Z(n19095) );
  NOR2_X1 U22061 ( .A1(n19084), .A2(n19083), .ZN(n19085) );
  AOI21_X1 U22062 ( .B1(n19087), .B2(n19086), .A(n19085), .ZN(n19089) );
  OAI211_X1 U22063 ( .C1(n19814), .C2(n19096), .A(n19089), .B(n19088), .ZN(
        n19093) );
  OAI22_X1 U22064 ( .A1(n19091), .A2(n19090), .B1(n19195), .B2(n19127), .ZN(
        n19092) );
  AOI211_X1 U22065 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19110), .A(n19093), .B(
        n19092), .ZN(n19094) );
  OAI21_X1 U22066 ( .B1(n19095), .B2(n19782), .A(n19094), .ZN(P2_U2848) );
  INV_X1 U22067 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19812) );
  OAI21_X1 U22068 ( .B1(n19812), .B2(n19096), .A(n11494), .ZN(n19100) );
  OAI22_X1 U22069 ( .A1(n19098), .A2(n19112), .B1(n19097), .B2(n11182), .ZN(
        n19099) );
  AOI211_X1 U22070 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19109), .A(
        n19100), .B(n19099), .ZN(n19108) );
  NOR2_X1 U22071 ( .A1(n19102), .A2(n19101), .ZN(n19104) );
  XNOR2_X1 U22072 ( .A(n19104), .B(n19103), .ZN(n19106) );
  AOI22_X1 U22073 ( .A1(n19106), .A2(n19123), .B1(n19122), .B2(n19105), .ZN(
        n19107) );
  OAI211_X1 U22074 ( .C1(n19127), .C2(n19197), .A(n19108), .B(n19107), .ZN(
        P2_U2849) );
  AOI22_X1 U22075 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19109), .ZN(n19111) );
  OAI21_X1 U22076 ( .B1(n19113), .B2(n19112), .A(n19111), .ZN(n19114) );
  AOI211_X1 U22077 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19116), .A(n19115), .B(
        n19114), .ZN(n19126) );
  NAND2_X1 U22078 ( .A1(n19118), .A2(n19117), .ZN(n19119) );
  XNOR2_X1 U22079 ( .A(n19120), .B(n19119), .ZN(n19124) );
  AOI22_X1 U22080 ( .A1(n19124), .A2(n19123), .B1(n19122), .B2(n19121), .ZN(
        n19125) );
  OAI211_X1 U22081 ( .C1(n19127), .C2(n19204), .A(n19126), .B(n19125), .ZN(
        P2_U2850) );
  OAI21_X1 U22082 ( .B1(n14901), .B2(n19128), .A(n14895), .ZN(n19129) );
  INV_X1 U22083 ( .A(n19129), .ZN(n19169) );
  AOI22_X1 U22084 ( .A1(n19169), .A2(n19156), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19153), .ZN(n19130) );
  OAI21_X1 U22085 ( .B1(n19153), .B2(n19131), .A(n19130), .ZN(P2_U2871) );
  XOR2_X1 U22086 ( .A(n19133), .B(n19132), .Z(n19134) );
  AOI22_X1 U22087 ( .A1(n19134), .A2(n19156), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19153), .ZN(n19135) );
  OAI21_X1 U22088 ( .B1(n19136), .B2(n19153), .A(n19135), .ZN(P2_U2873) );
  XOR2_X1 U22089 ( .A(n19138), .B(n19137), .Z(n19139) );
  AOI22_X1 U22090 ( .A1(n19139), .A2(n19156), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19153), .ZN(n19140) );
  OAI21_X1 U22091 ( .B1(n19141), .B2(n19153), .A(n19140), .ZN(P2_U2875) );
  XOR2_X1 U22092 ( .A(n13830), .B(n19142), .Z(n19143) );
  AOI22_X1 U22093 ( .A1(n19143), .A2(n19156), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19153), .ZN(n19144) );
  OAI21_X1 U22094 ( .B1(n19145), .B2(n19153), .A(n19144), .ZN(P2_U2877) );
  INV_X1 U22095 ( .A(n19146), .ZN(n19149) );
  AOI211_X1 U22096 ( .C1(n19150), .C2(n19149), .A(n19148), .B(n19147), .ZN(
        n19151) );
  AOI21_X1 U22097 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19153), .A(n19151), .ZN(
        n19152) );
  OAI21_X1 U22098 ( .B1(n19154), .B2(n19153), .A(n19152), .ZN(P2_U2879) );
  INV_X1 U22099 ( .A(n19200), .ZN(n19157) );
  AOI22_X1 U22100 ( .A1(n19157), .A2(n19156), .B1(n19159), .B2(n19155), .ZN(
        n19158) );
  OAI21_X1 U22101 ( .B1(n19159), .B2(n11172), .A(n19158), .ZN(P2_U2883) );
  AOI22_X1 U22102 ( .A1(n19160), .A2(n19214), .B1(n19165), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19162) );
  AOI22_X1 U22103 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19213), .B1(n19166), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19161) );
  NAND2_X1 U22104 ( .A1(n19162), .A2(n19161), .ZN(P2_U2888) );
  AOI22_X1 U22105 ( .A1(n19164), .A2(n19163), .B1(n19213), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19172) );
  AOI22_X1 U22106 ( .A1(n19166), .A2(BUF1_REG_16__SCAN_IN), .B1(n19165), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19171) );
  AOI22_X1 U22107 ( .A1(n19169), .A2(n19168), .B1(n19214), .B2(n19167), .ZN(
        n19170) );
  NAND3_X1 U22108 ( .A1(n19172), .A2(n19171), .A3(n19170), .ZN(P2_U2903) );
  OAI222_X1 U22109 ( .A1(n19175), .A2(n19205), .B1(n13139), .B2(n19196), .C1(
        n19174), .C2(n19222), .ZN(P2_U2904) );
  AOI22_X1 U22110 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19213), .B1(n19176), 
        .B2(n19198), .ZN(n19177) );
  OAI21_X1 U22111 ( .B1(n19205), .B2(n19178), .A(n19177), .ZN(P2_U2905) );
  INV_X1 U22112 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19229) );
  OAI222_X1 U22113 ( .A1(n19180), .A2(n19205), .B1(n19229), .B2(n19196), .C1(
        n19222), .C2(n19179), .ZN(P2_U2906) );
  INV_X1 U22114 ( .A(n19181), .ZN(n19183) );
  INV_X1 U22115 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19231) );
  OAI222_X1 U22116 ( .A1(n19183), .A2(n19205), .B1(n19231), .B2(n19196), .C1(
        n19222), .C2(n19182), .ZN(P2_U2907) );
  INV_X1 U22117 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19233) );
  OAI222_X1 U22118 ( .A1(n19185), .A2(n19205), .B1(n19233), .B2(n19196), .C1(
        n19222), .C2(n19184), .ZN(P2_U2908) );
  AOI22_X1 U22119 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19213), .B1(n19186), 
        .B2(n19198), .ZN(n19187) );
  OAI21_X1 U22120 ( .B1(n19205), .B2(n19188), .A(n19187), .ZN(P2_U2909) );
  AOI22_X1 U22121 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19213), .B1(n19189), .B2(
        n19198), .ZN(n19190) );
  OAI21_X1 U22122 ( .B1(n19205), .B2(n19191), .A(n19190), .ZN(P2_U2910) );
  AOI22_X1 U22123 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19213), .B1(n19192), .B2(
        n19198), .ZN(n19193) );
  OAI21_X1 U22124 ( .B1(n19205), .B2(n19194), .A(n19193), .ZN(P2_U2911) );
  INV_X1 U22125 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20905) );
  OAI222_X1 U22126 ( .A1(n19195), .A2(n19205), .B1(n20905), .B2(n19196), .C1(
        n19222), .C2(n19311), .ZN(P2_U2912) );
  INV_X1 U22127 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19242) );
  OAI222_X1 U22128 ( .A1(n19197), .A2(n19205), .B1(n19242), .B2(n19196), .C1(
        n19222), .C2(n19303), .ZN(P2_U2913) );
  AOI22_X1 U22129 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19213), .B1(n19199), .B2(
        n19198), .ZN(n19203) );
  OR3_X1 U22130 ( .A1(n19201), .A2(n19200), .A3(n19218), .ZN(n19202) );
  OAI211_X1 U22131 ( .C1(n19205), .C2(n19204), .A(n19203), .B(n19202), .ZN(
        P2_U2914) );
  INV_X1 U22132 ( .A(n19206), .ZN(n19870) );
  AOI22_X1 U22133 ( .A1(n19870), .A2(n19214), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19213), .ZN(n19212) );
  AOI21_X1 U22134 ( .B1(n19209), .B2(n19208), .A(n19207), .ZN(n19210) );
  OR2_X1 U22135 ( .A1(n19210), .A2(n19218), .ZN(n19211) );
  OAI211_X1 U22136 ( .C1(n19293), .C2(n19222), .A(n19212), .B(n19211), .ZN(
        P2_U2916) );
  AOI22_X1 U22137 ( .A1(n19214), .A2(n19889), .B1(n19213), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19221) );
  AOI21_X1 U22138 ( .B1(n19217), .B2(n19216), .A(n19215), .ZN(n19219) );
  OR2_X1 U22139 ( .A1(n19219), .A2(n19218), .ZN(n19220) );
  OAI211_X1 U22140 ( .C1(n19223), .C2(n19222), .A(n19221), .B(n19220), .ZN(
        P2_U2918) );
  AND2_X1 U22141 ( .A1(n19243), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22142 ( .A1(n21034), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19225) );
  OAI21_X1 U22143 ( .B1(n13139), .B2(n19254), .A(n19225), .ZN(P2_U2936) );
  AOI22_X1 U22144 ( .A1(n21034), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19226) );
  OAI21_X1 U22145 ( .B1(n19227), .B2(n19254), .A(n19226), .ZN(P2_U2937) );
  AOI22_X1 U22146 ( .A1(n21034), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19228) );
  OAI21_X1 U22147 ( .B1(n19229), .B2(n19254), .A(n19228), .ZN(P2_U2938) );
  AOI22_X1 U22148 ( .A1(n21034), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19230) );
  OAI21_X1 U22149 ( .B1(n19231), .B2(n19254), .A(n19230), .ZN(P2_U2939) );
  AOI22_X1 U22150 ( .A1(n21034), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19232) );
  OAI21_X1 U22151 ( .B1(n19233), .B2(n19254), .A(n19232), .ZN(P2_U2940) );
  AOI22_X1 U22152 ( .A1(n21034), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19234) );
  OAI21_X1 U22153 ( .B1(n19235), .B2(n19254), .A(n19234), .ZN(P2_U2941) );
  AOI22_X1 U22154 ( .A1(n21034), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19236) );
  OAI21_X1 U22155 ( .B1(n19237), .B2(n19254), .A(n19236), .ZN(P2_U2942) );
  AOI22_X1 U22156 ( .A1(n21034), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19238) );
  OAI21_X1 U22157 ( .B1(n19239), .B2(n19254), .A(n19238), .ZN(P2_U2943) );
  AOI22_X1 U22158 ( .A1(n21034), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19240) );
  OAI21_X1 U22159 ( .B1(n20905), .B2(n19254), .A(n19240), .ZN(P2_U2944) );
  AOI22_X1 U22160 ( .A1(n21034), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19241) );
  OAI21_X1 U22161 ( .B1(n19242), .B2(n19254), .A(n19241), .ZN(P2_U2945) );
  INV_X1 U22162 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20955) );
  AOI22_X1 U22163 ( .A1(n21034), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19244) );
  OAI21_X1 U22164 ( .B1(n20955), .B2(n19254), .A(n19244), .ZN(P2_U2946) );
  INV_X1 U22165 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19246) );
  AOI22_X1 U22166 ( .A1(n21034), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19245) );
  OAI21_X1 U22167 ( .B1(n19246), .B2(n19254), .A(n19245), .ZN(P2_U2947) );
  INV_X1 U22168 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19248) );
  AOI22_X1 U22169 ( .A1(n21034), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19247) );
  OAI21_X1 U22170 ( .B1(n19248), .B2(n19254), .A(n19247), .ZN(P2_U2948) );
  AOI22_X1 U22171 ( .A1(n21034), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19249) );
  OAI21_X1 U22172 ( .B1(n19250), .B2(n19254), .A(n19249), .ZN(P2_U2949) );
  INV_X1 U22173 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19252) );
  AOI22_X1 U22174 ( .A1(n21034), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22175 ( .B1(n19252), .B2(n19254), .A(n19251), .ZN(P2_U2950) );
  AOI22_X1 U22176 ( .A1(n21034), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19243), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19253) );
  OAI21_X1 U22177 ( .B1(n13135), .B2(n19254), .A(n19253), .ZN(P2_U2951) );
  INV_X1 U22178 ( .A(n19256), .ZN(n19268) );
  OAI22_X1 U22179 ( .A1(n19260), .A2(n19259), .B1(n19258), .B2(n19257), .ZN(
        n19267) );
  NAND2_X1 U22180 ( .A1(n19879), .A2(n19261), .ZN(n19263) );
  OAI211_X1 U22181 ( .C1(n19265), .C2(n19264), .A(n19263), .B(n19262), .ZN(
        n19266) );
  AOI211_X1 U22182 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n19268), .A(
        n19267), .B(n19266), .ZN(n19274) );
  INV_X1 U22183 ( .A(n19269), .ZN(n19272) );
  OAI21_X1 U22184 ( .B1(n19272), .B2(n19271), .A(n19270), .ZN(n19273) );
  OAI211_X1 U22185 ( .C1(n19276), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3044) );
  NAND2_X1 U22186 ( .A1(n19279), .A2(n19495), .ZN(n19758) );
  NAND2_X1 U22187 ( .A1(n19874), .A2(n19881), .ZN(n19374) );
  INV_X1 U22188 ( .A(n19374), .ZN(n19376) );
  NAND2_X1 U22189 ( .A1(n19376), .A2(n19891), .ZN(n19320) );
  NOR2_X1 U22190 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19320), .ZN(
        n19310) );
  AOI22_X1 U22191 ( .A1(n19652), .A2(n19771), .B1(n19718), .B2(n19310), .ZN(
        n19288) );
  AOI21_X1 U22192 ( .B1(n19758), .B2(n19323), .A(n19467), .ZN(n19280) );
  NOR2_X1 U22193 ( .A1(n19280), .A2(n19722), .ZN(n19283) );
  AOI21_X1 U22194 ( .B1(n19284), .B2(n19678), .A(n19869), .ZN(n19281) );
  AOI21_X1 U22195 ( .B1(n19283), .B2(n19723), .A(n19281), .ZN(n19282) );
  OAI21_X1 U22196 ( .B1(n19282), .B2(n19310), .A(n19726), .ZN(n19313) );
  INV_X1 U22197 ( .A(n19723), .ZN(n19767) );
  OAI21_X1 U22198 ( .B1(n19767), .B2(n19310), .A(n19283), .ZN(n19286) );
  OAI21_X1 U22199 ( .B1(n19284), .B2(n19310), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19285) );
  NAND2_X1 U22200 ( .A1(n19286), .A2(n19285), .ZN(n19312) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19313), .B1(
        n13454), .B2(n19312), .ZN(n19287) );
  OAI211_X1 U22202 ( .C1(n19507), .C2(n19323), .A(n19288), .B(n19287), .ZN(
        P2_U3048) );
  AOI22_X1 U22203 ( .A1(n19732), .A2(n19771), .B1(n13381), .B2(n19310), .ZN(
        n19290) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19313), .B1(
        n13380), .B2(n19312), .ZN(n19289) );
  OAI211_X1 U22205 ( .C1(n19735), .C2(n19323), .A(n19290), .B(n19289), .ZN(
        P2_U3049) );
  AOI22_X1 U22206 ( .A1(n19737), .A2(n19771), .B1(n19736), .B2(n19310), .ZN(
        n19292) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19313), .B1(
        n13449), .B2(n19312), .ZN(n19291) );
  OAI211_X1 U22208 ( .C1(n19740), .C2(n19323), .A(n19292), .B(n19291), .ZN(
        P2_U3050) );
  AOI22_X1 U22209 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19306), .ZN(n19564) );
  AOI22_X1 U22210 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19306), .ZN(n19745) );
  INV_X1 U22211 ( .A(n19745), .ZN(n19609) );
  NOR2_X2 U22212 ( .A1(n10714), .A2(n19308), .ZN(n19741) );
  AOI22_X1 U22213 ( .A1(n19609), .A2(n19771), .B1(n19741), .B2(n19310), .ZN(
        n19296) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19313), .B1(
        n19294), .B2(n19312), .ZN(n19295) );
  OAI211_X1 U22215 ( .C1(n19564), .C2(n19323), .A(n19296), .B(n19295), .ZN(
        P2_U3051) );
  AOI22_X1 U22216 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19306), .ZN(n19700) );
  AOI22_X1 U22217 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19306), .ZN(n19751) );
  NOR2_X2 U22218 ( .A1(n10704), .A2(n19308), .ZN(n19746) );
  AOI22_X1 U22219 ( .A1(n19697), .A2(n19771), .B1(n19746), .B2(n19310), .ZN(
        n19299) );
  NOR2_X2 U22220 ( .A1(n19297), .A2(n19680), .ZN(n19747) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19313), .B1(
        n19747), .B2(n19312), .ZN(n19298) );
  OAI211_X1 U22222 ( .C1(n19700), .C2(n19323), .A(n19299), .B(n19298), .ZN(
        P2_U3052) );
  AOI22_X1 U22223 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19306), .ZN(n19759) );
  AOI22_X1 U22224 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19306), .ZN(n19643) );
  NOR2_X2 U22225 ( .A1(n11593), .A2(n19308), .ZN(n19752) );
  AOI22_X1 U22226 ( .A1(n19754), .A2(n19771), .B1(n19752), .B2(n19310), .ZN(
        n19302) );
  NOR2_X2 U22227 ( .A1(n19300), .A2(n19680), .ZN(n19753) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19313), .B1(
        n19753), .B2(n19312), .ZN(n19301) );
  OAI211_X1 U22229 ( .C1(n19759), .C2(n19323), .A(n19302), .B(n19301), .ZN(
        P2_U3053) );
  AOI22_X1 U22230 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19306), .ZN(n19620) );
  AOI22_X1 U22231 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19306), .ZN(n19765) );
  INV_X1 U22232 ( .A(n19765), .ZN(n19616) );
  NOR2_X2 U22233 ( .A1(n10609), .A2(n19308), .ZN(n19760) );
  AOI22_X1 U22234 ( .A1(n19616), .A2(n19771), .B1(n19760), .B2(n19310), .ZN(
        n19305) );
  NOR2_X2 U22235 ( .A1(n19303), .A2(n19680), .ZN(n19761) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19313), .B1(
        n19761), .B2(n19312), .ZN(n19304) );
  OAI211_X1 U22237 ( .C1(n19620), .C2(n19323), .A(n19305), .B(n19304), .ZN(
        P2_U3054) );
  AOI22_X1 U22238 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19306), .ZN(n19713) );
  AOI22_X1 U22239 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19307), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19306), .ZN(n19776) );
  NOR2_X2 U22240 ( .A1(n19309), .A2(n19308), .ZN(n19766) );
  AOI22_X1 U22241 ( .A1(n19708), .A2(n19771), .B1(n19766), .B2(n19310), .ZN(
        n19315) );
  NOR2_X2 U22242 ( .A1(n19311), .A2(n19680), .ZN(n19768) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19313), .B1(
        n19768), .B2(n19312), .ZN(n19314) );
  OAI211_X1 U22244 ( .C1(n19713), .C2(n19323), .A(n19315), .B(n19314), .ZN(
        P2_U3055) );
  NOR2_X1 U22245 ( .A1(n19316), .A2(n19374), .ZN(n19338) );
  NOR3_X1 U22246 ( .A1(n19317), .A2(n19338), .A3(n19676), .ZN(n19319) );
  AOI211_X2 U22247 ( .C1(n19320), .C2(n19676), .A(n19497), .B(n19319), .ZN(
        n19339) );
  AOI22_X1 U22248 ( .A1(n19339), .A2(n13454), .B1(n19718), .B2(n19338), .ZN(
        n19325) );
  NAND2_X1 U22249 ( .A1(n19499), .A2(n19318), .ZN(n19321) );
  AOI21_X1 U22250 ( .B1(n19321), .B2(n19320), .A(n19319), .ZN(n19322) );
  OAI211_X1 U22251 ( .C1(n19338), .C2(n19678), .A(n19322), .B(n19726), .ZN(
        n19341) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19652), .ZN(n19324) );
  OAI211_X1 U22253 ( .C1(n19507), .C2(n19373), .A(n19325), .B(n19324), .ZN(
        P2_U3056) );
  AOI22_X1 U22254 ( .A1(n19339), .A2(n13380), .B1(n13381), .B2(n19338), .ZN(
        n19327) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19732), .ZN(n19326) );
  OAI211_X1 U22256 ( .C1(n19735), .C2(n19373), .A(n19327), .B(n19326), .ZN(
        P2_U3057) );
  AOI22_X1 U22257 ( .A1(n19339), .A2(n13449), .B1(n19736), .B2(n19338), .ZN(
        n19329) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19737), .ZN(n19328) );
  OAI211_X1 U22259 ( .C1(n19740), .C2(n19373), .A(n19329), .B(n19328), .ZN(
        P2_U3058) );
  AOI22_X1 U22260 ( .A1(n19339), .A2(n19294), .B1(n19741), .B2(n19338), .ZN(
        n19331) );
  AOI22_X1 U22261 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19609), .ZN(n19330) );
  OAI211_X1 U22262 ( .C1(n19564), .C2(n19373), .A(n19331), .B(n19330), .ZN(
        P2_U3059) );
  AOI22_X1 U22263 ( .A1(n19339), .A2(n19747), .B1(n19746), .B2(n19338), .ZN(
        n19333) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19697), .ZN(n19332) );
  OAI211_X1 U22265 ( .C1(n19700), .C2(n19373), .A(n19333), .B(n19332), .ZN(
        P2_U3060) );
  AOI22_X1 U22266 ( .A1(n19339), .A2(n19753), .B1(n19752), .B2(n19338), .ZN(
        n19335) );
  AOI22_X1 U22267 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19754), .ZN(n19334) );
  OAI211_X1 U22268 ( .C1(n19759), .C2(n19373), .A(n19335), .B(n19334), .ZN(
        P2_U3061) );
  AOI22_X1 U22269 ( .A1(n19339), .A2(n19761), .B1(n19760), .B2(n19338), .ZN(
        n19337) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19616), .ZN(n19336) );
  OAI211_X1 U22271 ( .C1(n19620), .C2(n19373), .A(n19337), .B(n19336), .ZN(
        P2_U3062) );
  AOI22_X1 U22272 ( .A1(n19339), .A2(n19768), .B1(n19766), .B2(n19338), .ZN(
        n19343) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19341), .B1(
        n19340), .B2(n19708), .ZN(n19342) );
  OAI211_X1 U22274 ( .C1(n19713), .C2(n19373), .A(n19343), .B(n19342), .ZN(
        P2_U3063) );
  INV_X1 U22275 ( .A(n19347), .ZN(n19344) );
  NOR2_X1 U22276 ( .A1(n19891), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19578) );
  AND2_X1 U22277 ( .A1(n19578), .A2(n19376), .ZN(n19368) );
  OAI21_X1 U22278 ( .B1(n19344), .B2(n19368), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19345) );
  OR2_X1 U22279 ( .A1(n19581), .A2(n19374), .ZN(n19349) );
  NAND2_X1 U22280 ( .A1(n19345), .A2(n19349), .ZN(n19369) );
  AOI22_X1 U22281 ( .A1(n19369), .A2(n13454), .B1(n19718), .B2(n19368), .ZN(
        n19355) );
  INV_X1 U22282 ( .A(n19368), .ZN(n19346) );
  OAI21_X1 U22283 ( .B1(n19347), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19346), 
        .ZN(n19352) );
  INV_X1 U22284 ( .A(n19373), .ZN(n19348) );
  OAI21_X1 U22285 ( .B1(n19396), .B2(n19348), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19350) );
  NAND2_X1 U22286 ( .A1(n19350), .A2(n19349), .ZN(n19351) );
  MUX2_X1 U22287 ( .A(n19352), .B(n19351), .S(n19869), .Z(n19353) );
  NAND2_X1 U22288 ( .A1(n19353), .A2(n19726), .ZN(n19370) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19728), .ZN(n19354) );
  OAI211_X1 U22290 ( .C1(n19731), .C2(n19373), .A(n19355), .B(n19354), .ZN(
        P2_U3064) );
  AOI22_X1 U22291 ( .A1(n19369), .A2(n13380), .B1(n13381), .B2(n19368), .ZN(
        n19357) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19689), .ZN(n19356) );
  OAI211_X1 U22293 ( .C1(n19692), .C2(n19373), .A(n19357), .B(n19356), .ZN(
        P2_U3065) );
  AOI22_X1 U22294 ( .A1(n19369), .A2(n13449), .B1(n19736), .B2(n19368), .ZN(
        n19359) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19631), .ZN(n19358) );
  OAI211_X1 U22296 ( .C1(n19634), .C2(n19373), .A(n19359), .B(n19358), .ZN(
        P2_U3066) );
  AOI22_X1 U22297 ( .A1(n19369), .A2(n19294), .B1(n19741), .B2(n19368), .ZN(
        n19361) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19742), .ZN(n19360) );
  OAI211_X1 U22299 ( .C1(n19745), .C2(n19373), .A(n19361), .B(n19360), .ZN(
        P2_U3067) );
  AOI22_X1 U22300 ( .A1(n19369), .A2(n19747), .B1(n19746), .B2(n19368), .ZN(
        n19363) );
  INV_X1 U22301 ( .A(n19700), .ZN(n19748) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19748), .ZN(n19362) );
  OAI211_X1 U22303 ( .C1(n19751), .C2(n19373), .A(n19363), .B(n19362), .ZN(
        P2_U3068) );
  AOI22_X1 U22304 ( .A1(n19369), .A2(n19753), .B1(n19752), .B2(n19368), .ZN(
        n19365) );
  INV_X1 U22305 ( .A(n19759), .ZN(n19640) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19640), .ZN(n19364) );
  OAI211_X1 U22307 ( .C1(n19643), .C2(n19373), .A(n19365), .B(n19364), .ZN(
        P2_U3069) );
  AOI22_X1 U22308 ( .A1(n19369), .A2(n19761), .B1(n19760), .B2(n19368), .ZN(
        n19367) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19762), .ZN(n19366) );
  OAI211_X1 U22310 ( .C1(n19765), .C2(n19373), .A(n19367), .B(n19366), .ZN(
        P2_U3070) );
  AOI22_X1 U22311 ( .A1(n19369), .A2(n19768), .B1(n19766), .B2(n19368), .ZN(
        n19372) );
  INV_X1 U22312 ( .A(n19713), .ZN(n19770) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19370), .B1(
        n19396), .B2(n19770), .ZN(n19371) );
  OAI211_X1 U22314 ( .C1(n19776), .C2(n19373), .A(n19372), .B(n19371), .ZN(
        P2_U3071) );
  NOR2_X1 U22315 ( .A1(n19375), .A2(n19374), .ZN(n19400) );
  AOI22_X1 U22316 ( .A1(n19652), .A2(n19396), .B1(n19718), .B2(n19400), .ZN(
        n19385) );
  AOI21_X1 U22317 ( .B1(n10884), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19378) );
  AOI21_X1 U22318 ( .B1(n19499), .B2(n19865), .A(n19722), .ZN(n19379) );
  NAND2_X1 U22319 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19376), .ZN(
        n19382) );
  NAND2_X1 U22320 ( .A1(n19379), .A2(n19382), .ZN(n19377) );
  OAI211_X1 U22321 ( .C1(n19400), .C2(n19378), .A(n19377), .B(n19726), .ZN(
        n19402) );
  INV_X1 U22322 ( .A(n19379), .ZN(n19383) );
  OAI21_X1 U22323 ( .B1(n19380), .B2(n19400), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19381) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19402), .B1(
        n13454), .B2(n19401), .ZN(n19384) );
  OAI211_X1 U22325 ( .C1(n19507), .C2(n19399), .A(n19385), .B(n19384), .ZN(
        P2_U3072) );
  AOI22_X1 U22326 ( .A1(n19732), .A2(n19396), .B1(n13381), .B2(n19400), .ZN(
        n19387) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19402), .B1(
        n13380), .B2(n19401), .ZN(n19386) );
  OAI211_X1 U22328 ( .C1(n19735), .C2(n19399), .A(n19387), .B(n19386), .ZN(
        P2_U3073) );
  AOI22_X1 U22329 ( .A1(n19737), .A2(n19396), .B1(n19736), .B2(n19400), .ZN(
        n19389) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19402), .B1(
        n13449), .B2(n19401), .ZN(n19388) );
  OAI211_X1 U22331 ( .C1(n19740), .C2(n19399), .A(n19389), .B(n19388), .ZN(
        P2_U3074) );
  AOI22_X1 U22332 ( .A1(n19609), .A2(n19396), .B1(n19400), .B2(n19741), .ZN(
        n19391) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19402), .B1(
        n19294), .B2(n19401), .ZN(n19390) );
  OAI211_X1 U22334 ( .C1(n19564), .C2(n19399), .A(n19391), .B(n19390), .ZN(
        P2_U3075) );
  AOI22_X1 U22335 ( .A1(n19697), .A2(n19396), .B1(n19400), .B2(n19746), .ZN(
        n19393) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19402), .B1(
        n19747), .B2(n19401), .ZN(n19392) );
  OAI211_X1 U22337 ( .C1(n19700), .C2(n19399), .A(n19393), .B(n19392), .ZN(
        P2_U3076) );
  INV_X1 U22338 ( .A(n19396), .ZN(n19405) );
  AOI22_X1 U22339 ( .A1(n19640), .A2(n19429), .B1(n19400), .B2(n19752), .ZN(
        n19395) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19402), .B1(
        n19753), .B2(n19401), .ZN(n19394) );
  OAI211_X1 U22341 ( .C1(n19643), .C2(n19405), .A(n19395), .B(n19394), .ZN(
        P2_U3077) );
  AOI22_X1 U22342 ( .A1(n19616), .A2(n19396), .B1(n19400), .B2(n19760), .ZN(
        n19398) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19402), .B1(
        n19761), .B2(n19401), .ZN(n19397) );
  OAI211_X1 U22344 ( .C1(n19620), .C2(n19399), .A(n19398), .B(n19397), .ZN(
        P2_U3078) );
  AOI22_X1 U22345 ( .A1(n19770), .A2(n19429), .B1(n19400), .B2(n19766), .ZN(
        n19404) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19402), .B1(
        n19768), .B2(n19401), .ZN(n19403) );
  OAI211_X1 U22347 ( .C1(n19776), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P2_U3079) );
  NAND2_X1 U22348 ( .A1(n19406), .A2(n19874), .ZN(n19411) );
  NAND3_X1 U22349 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19874), .A3(
        n19891), .ZN(n19440) );
  NOR2_X1 U22350 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19440), .ZN(
        n19427) );
  OAI21_X1 U22351 ( .B1(n19408), .B2(n19427), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19407) );
  OAI21_X1 U22352 ( .B1(n19411), .B2(n19722), .A(n19407), .ZN(n19428) );
  AOI22_X1 U22353 ( .A1(n19428), .A2(n13454), .B1(n19718), .B2(n19427), .ZN(
        n19414) );
  OAI21_X1 U22354 ( .B1(n19429), .B2(n19457), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19410) );
  AOI211_X1 U22355 ( .C1(n19408), .C2(n19678), .A(n19427), .B(n19869), .ZN(
        n19409) );
  AOI211_X1 U22356 ( .C1(n19411), .C2(n19410), .A(n19680), .B(n19409), .ZN(
        n19412) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19652), .ZN(n19413) );
  OAI211_X1 U22358 ( .C1(n19507), .C2(n19456), .A(n19414), .B(n19413), .ZN(
        P2_U3080) );
  AOI22_X1 U22359 ( .A1(n19428), .A2(n13380), .B1(n13381), .B2(n19427), .ZN(
        n19416) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19732), .ZN(n19415) );
  OAI211_X1 U22361 ( .C1(n19735), .C2(n19456), .A(n19416), .B(n19415), .ZN(
        P2_U3081) );
  AOI22_X1 U22362 ( .A1(n19428), .A2(n13449), .B1(n19736), .B2(n19427), .ZN(
        n19418) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19737), .ZN(n19417) );
  OAI211_X1 U22364 ( .C1(n19740), .C2(n19456), .A(n19418), .B(n19417), .ZN(
        P2_U3082) );
  AOI22_X1 U22365 ( .A1(n19428), .A2(n19294), .B1(n19741), .B2(n19427), .ZN(
        n19420) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19609), .ZN(n19419) );
  OAI211_X1 U22367 ( .C1(n19564), .C2(n19456), .A(n19420), .B(n19419), .ZN(
        P2_U3083) );
  AOI22_X1 U22368 ( .A1(n19428), .A2(n19747), .B1(n19746), .B2(n19427), .ZN(
        n19422) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19697), .ZN(n19421) );
  OAI211_X1 U22370 ( .C1(n19700), .C2(n19456), .A(n19422), .B(n19421), .ZN(
        P2_U3084) );
  AOI22_X1 U22371 ( .A1(n19428), .A2(n19753), .B1(n19752), .B2(n19427), .ZN(
        n19424) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19754), .ZN(n19423) );
  OAI211_X1 U22373 ( .C1(n19759), .C2(n19456), .A(n19424), .B(n19423), .ZN(
        P2_U3085) );
  AOI22_X1 U22374 ( .A1(n19428), .A2(n19761), .B1(n19760), .B2(n19427), .ZN(
        n19426) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19616), .ZN(n19425) );
  OAI211_X1 U22376 ( .C1(n19620), .C2(n19456), .A(n19426), .B(n19425), .ZN(
        P2_U3086) );
  AOI22_X1 U22377 ( .A1(n19428), .A2(n19768), .B1(n19766), .B2(n19427), .ZN(
        n19432) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19708), .ZN(n19431) );
  OAI211_X1 U22379 ( .C1(n19713), .C2(n19456), .A(n19432), .B(n19431), .ZN(
        P2_U3087) );
  NOR2_X1 U22380 ( .A1(n19900), .A2(n19440), .ZN(n19469) );
  AOI22_X1 U22381 ( .A1(n19652), .A2(n19457), .B1(n19718), .B2(n19469), .ZN(
        n19443) );
  AOI21_X1 U22382 ( .B1(n19499), .B2(n19433), .A(n19722), .ZN(n19437) );
  INV_X1 U22383 ( .A(n19469), .ZN(n19434) );
  NOR2_X1 U22384 ( .A1(n19438), .A2(n19676), .ZN(n19435) );
  AOI21_X1 U22385 ( .B1(n19437), .B2(n19440), .A(n19435), .ZN(n19436) );
  OAI211_X1 U22386 ( .C1(n19469), .C2(n19678), .A(n19436), .B(n19726), .ZN(
        n19459) );
  INV_X1 U22387 ( .A(n19437), .ZN(n19441) );
  INV_X1 U22388 ( .A(n19438), .ZN(n19439) );
  OAI22_X1 U22389 ( .A1(n19441), .A2(n19440), .B1(n19439), .B2(n19676), .ZN(
        n19458) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19459), .B1(
        n13454), .B2(n19458), .ZN(n19442) );
  OAI211_X1 U22391 ( .C1(n19507), .C2(n19486), .A(n19443), .B(n19442), .ZN(
        P2_U3088) );
  AOI22_X1 U22392 ( .A1(n19689), .A2(n19489), .B1(n13381), .B2(n19469), .ZN(
        n19445) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19459), .B1(
        n13380), .B2(n19458), .ZN(n19444) );
  OAI211_X1 U22394 ( .C1(n19692), .C2(n19456), .A(n19445), .B(n19444), .ZN(
        P2_U3089) );
  AOI22_X1 U22395 ( .A1(n19737), .A2(n19457), .B1(n19736), .B2(n19469), .ZN(
        n19447) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19459), .B1(
        n13449), .B2(n19458), .ZN(n19446) );
  OAI211_X1 U22397 ( .C1(n19740), .C2(n19486), .A(n19447), .B(n19446), .ZN(
        P2_U3090) );
  AOI22_X1 U22398 ( .A1(n19742), .A2(n19489), .B1(n19469), .B2(n19741), .ZN(
        n19449) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19459), .B1(
        n19294), .B2(n19458), .ZN(n19448) );
  OAI211_X1 U22400 ( .C1(n19745), .C2(n19456), .A(n19449), .B(n19448), .ZN(
        P2_U3091) );
  AOI22_X1 U22401 ( .A1(n19748), .A2(n19489), .B1(n19469), .B2(n19746), .ZN(
        n19451) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19459), .B1(
        n19747), .B2(n19458), .ZN(n19450) );
  OAI211_X1 U22403 ( .C1(n19751), .C2(n19456), .A(n19451), .B(n19450), .ZN(
        P2_U3092) );
  AOI22_X1 U22404 ( .A1(n19754), .A2(n19457), .B1(n19469), .B2(n19752), .ZN(
        n19453) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19459), .B1(
        n19753), .B2(n19458), .ZN(n19452) );
  OAI211_X1 U22406 ( .C1(n19759), .C2(n19486), .A(n19453), .B(n19452), .ZN(
        P2_U3093) );
  AOI22_X1 U22407 ( .A1(n19762), .A2(n19489), .B1(n19469), .B2(n19760), .ZN(
        n19455) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19459), .B1(
        n19761), .B2(n19458), .ZN(n19454) );
  OAI211_X1 U22409 ( .C1(n19765), .C2(n19456), .A(n19455), .B(n19454), .ZN(
        P2_U3094) );
  AOI22_X1 U22410 ( .A1(n19708), .A2(n19457), .B1(n19469), .B2(n19766), .ZN(
        n19461) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19459), .B1(
        n19768), .B2(n19458), .ZN(n19460) );
  OAI211_X1 U22412 ( .C1(n19713), .C2(n19486), .A(n19461), .B(n19460), .ZN(
        P2_U3095) );
  NAND2_X1 U22413 ( .A1(n19462), .A2(n19495), .ZN(n19493) );
  NAND2_X1 U22414 ( .A1(n19874), .A2(n19714), .ZN(n19498) );
  NOR2_X1 U22415 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19498), .ZN(
        n19487) );
  NOR2_X1 U22416 ( .A1(n19469), .A2(n19487), .ZN(n19463) );
  OR2_X1 U22417 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19463), .ZN(n19466) );
  INV_X1 U22418 ( .A(n19464), .ZN(n19465) );
  NOR3_X1 U22419 ( .A1(n19465), .A2(n19487), .A3(n19676), .ZN(n19470) );
  AOI21_X1 U22420 ( .B1(n19676), .B2(n19466), .A(n19470), .ZN(n19488) );
  AOI22_X1 U22421 ( .A1(n19488), .A2(n13454), .B1(n19718), .B2(n19487), .ZN(
        n19473) );
  AOI21_X1 U22422 ( .B1(n19486), .B2(n19493), .A(n19467), .ZN(n19468) );
  AOI221_X1 U22423 ( .B1(n19678), .B2(n19469), .C1(n19678), .C2(n19468), .A(
        n19487), .ZN(n19471) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19652), .ZN(n19472) );
  OAI211_X1 U22425 ( .C1(n19507), .C2(n19493), .A(n19473), .B(n19472), .ZN(
        P2_U3096) );
  AOI22_X1 U22426 ( .A1(n19488), .A2(n13380), .B1(n13381), .B2(n19487), .ZN(
        n19475) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19490), .B1(
        n19521), .B2(n19689), .ZN(n19474) );
  OAI211_X1 U22428 ( .C1(n19692), .C2(n19486), .A(n19475), .B(n19474), .ZN(
        P2_U3097) );
  AOI22_X1 U22429 ( .A1(n19488), .A2(n13449), .B1(n19736), .B2(n19487), .ZN(
        n19477) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19737), .ZN(n19476) );
  OAI211_X1 U22431 ( .C1(n19740), .C2(n19493), .A(n19477), .B(n19476), .ZN(
        P2_U3098) );
  AOI22_X1 U22432 ( .A1(n19488), .A2(n19294), .B1(n19741), .B2(n19487), .ZN(
        n19479) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19609), .ZN(n19478) );
  OAI211_X1 U22434 ( .C1(n19564), .C2(n19493), .A(n19479), .B(n19478), .ZN(
        P2_U3099) );
  AOI22_X1 U22435 ( .A1(n19488), .A2(n19747), .B1(n19746), .B2(n19487), .ZN(
        n19481) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19697), .ZN(n19480) );
  OAI211_X1 U22437 ( .C1(n19700), .C2(n19493), .A(n19481), .B(n19480), .ZN(
        P2_U3100) );
  AOI22_X1 U22438 ( .A1(n19488), .A2(n19753), .B1(n19752), .B2(n19487), .ZN(
        n19483) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19490), .B1(
        n19521), .B2(n19640), .ZN(n19482) );
  OAI211_X1 U22440 ( .C1(n19643), .C2(n19486), .A(n19483), .B(n19482), .ZN(
        P2_U3101) );
  AOI22_X1 U22441 ( .A1(n19488), .A2(n19761), .B1(n19760), .B2(n19487), .ZN(
        n19485) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19490), .B1(
        n19521), .B2(n19762), .ZN(n19484) );
  OAI211_X1 U22443 ( .C1(n19765), .C2(n19486), .A(n19485), .B(n19484), .ZN(
        P2_U3102) );
  AOI22_X1 U22444 ( .A1(n19488), .A2(n19768), .B1(n19766), .B2(n19487), .ZN(
        n19492) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19708), .ZN(n19491) );
  OAI211_X1 U22446 ( .C1(n19713), .C2(n19493), .A(n19492), .B(n19491), .ZN(
        P2_U3103) );
  INV_X1 U22447 ( .A(n10881), .ZN(n19496) );
  NOR2_X1 U22448 ( .A1(n19900), .A2(n19498), .ZN(n19528) );
  NOR3_X1 U22449 ( .A1(n19496), .A2(n19528), .A3(n19676), .ZN(n19501) );
  AOI211_X2 U22450 ( .C1(n19498), .C2(n19676), .A(n19497), .B(n19501), .ZN(
        n19520) );
  AOI22_X1 U22451 ( .A1(n19520), .A2(n13454), .B1(n19718), .B2(n19528), .ZN(
        n19506) );
  INV_X1 U22452 ( .A(n19498), .ZN(n19504) );
  INV_X1 U22453 ( .A(n19499), .ZN(n19500) );
  NOR2_X1 U22454 ( .A1(n19500), .A2(n19720), .ZN(n19868) );
  INV_X1 U22455 ( .A(n19528), .ZN(n19502) );
  AOI211_X1 U22456 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19502), .A(n19680), 
        .B(n19501), .ZN(n19503) );
  OAI21_X1 U22457 ( .B1(n19504), .B2(n19868), .A(n19503), .ZN(n19522) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19652), .ZN(n19505) );
  OAI211_X1 U22459 ( .C1(n19507), .C2(n19555), .A(n19506), .B(n19505), .ZN(
        P2_U3104) );
  AOI22_X1 U22460 ( .A1(n19520), .A2(n13380), .B1(n13381), .B2(n19528), .ZN(
        n19509) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19732), .ZN(n19508) );
  OAI211_X1 U22462 ( .C1(n19735), .C2(n19555), .A(n19509), .B(n19508), .ZN(
        P2_U3105) );
  AOI22_X1 U22463 ( .A1(n19520), .A2(n13449), .B1(n19736), .B2(n19528), .ZN(
        n19511) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19737), .ZN(n19510) );
  OAI211_X1 U22465 ( .C1(n19740), .C2(n19555), .A(n19511), .B(n19510), .ZN(
        P2_U3106) );
  AOI22_X1 U22466 ( .A1(n19520), .A2(n19294), .B1(n19741), .B2(n19528), .ZN(
        n19513) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19609), .ZN(n19512) );
  OAI211_X1 U22468 ( .C1(n19564), .C2(n19555), .A(n19513), .B(n19512), .ZN(
        P2_U3107) );
  AOI22_X1 U22469 ( .A1(n19520), .A2(n19747), .B1(n19746), .B2(n19528), .ZN(
        n19515) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19697), .ZN(n19514) );
  OAI211_X1 U22471 ( .C1(n19700), .C2(n19555), .A(n19515), .B(n19514), .ZN(
        P2_U3108) );
  AOI22_X1 U22472 ( .A1(n19520), .A2(n19753), .B1(n19752), .B2(n19528), .ZN(
        n19517) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19754), .ZN(n19516) );
  OAI211_X1 U22474 ( .C1(n19759), .C2(n19555), .A(n19517), .B(n19516), .ZN(
        P2_U3109) );
  AOI22_X1 U22475 ( .A1(n19520), .A2(n19761), .B1(n19760), .B2(n19528), .ZN(
        n19519) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19616), .ZN(n19518) );
  OAI211_X1 U22477 ( .C1(n19620), .C2(n19555), .A(n19519), .B(n19518), .ZN(
        P2_U3110) );
  AOI22_X1 U22478 ( .A1(n19520), .A2(n19768), .B1(n19766), .B2(n19528), .ZN(
        n19524) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19522), .B1(
        n19521), .B2(n19708), .ZN(n19523) );
  OAI211_X1 U22480 ( .C1(n19713), .C2(n19555), .A(n19524), .B(n19523), .ZN(
        P2_U3111) );
  NOR2_X1 U22481 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19525), .ZN(
        n19550) );
  AOI22_X1 U22482 ( .A1(n19728), .A2(n19572), .B1(n19718), .B2(n19550), .ZN(
        n19537) );
  INV_X1 U22483 ( .A(n19555), .ZN(n19526) );
  OAI21_X1 U22484 ( .B1(n19572), .B2(n19526), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19527) );
  NAND2_X1 U22485 ( .A1(n19527), .A2(n19869), .ZN(n19535) );
  NOR2_X1 U22486 ( .A1(n19550), .A2(n19528), .ZN(n19533) );
  INV_X1 U22487 ( .A(n19533), .ZN(n19531) );
  INV_X1 U22488 ( .A(n19550), .ZN(n19529) );
  OAI211_X1 U22489 ( .C1(n10895), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19529), 
        .B(n19722), .ZN(n19530) );
  OAI211_X1 U22490 ( .C1(n19535), .C2(n19531), .A(n19726), .B(n19530), .ZN(
        n19552) );
  INV_X1 U22491 ( .A(n10895), .ZN(n19532) );
  OAI21_X1 U22492 ( .B1(n19532), .B2(n19550), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19534) );
  AOI22_X1 U22493 ( .A1(n19535), .A2(n19534), .B1(n19533), .B2(n19676), .ZN(
        n19551) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19552), .B1(
        n13454), .B2(n19551), .ZN(n19536) );
  OAI211_X1 U22495 ( .C1(n19731), .C2(n19555), .A(n19537), .B(n19536), .ZN(
        P2_U3112) );
  AOI22_X1 U22496 ( .A1(n19689), .A2(n19572), .B1(n13381), .B2(n19550), .ZN(
        n19539) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19552), .B1(
        n13380), .B2(n19551), .ZN(n19538) );
  OAI211_X1 U22498 ( .C1(n19692), .C2(n19555), .A(n19539), .B(n19538), .ZN(
        P2_U3113) );
  AOI22_X1 U22499 ( .A1(n19631), .A2(n19572), .B1(n19736), .B2(n19550), .ZN(
        n19541) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19552), .B1(
        n13449), .B2(n19551), .ZN(n19540) );
  OAI211_X1 U22501 ( .C1(n19634), .C2(n19555), .A(n19541), .B(n19540), .ZN(
        P2_U3114) );
  AOI22_X1 U22502 ( .A1(n19742), .A2(n19572), .B1(n19741), .B2(n19550), .ZN(
        n19543) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19552), .B1(
        n19294), .B2(n19551), .ZN(n19542) );
  OAI211_X1 U22504 ( .C1(n19745), .C2(n19555), .A(n19543), .B(n19542), .ZN(
        P2_U3115) );
  AOI22_X1 U22505 ( .A1(n19748), .A2(n19572), .B1(n19746), .B2(n19550), .ZN(
        n19545) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19552), .B1(
        n19747), .B2(n19551), .ZN(n19544) );
  OAI211_X1 U22507 ( .C1(n19751), .C2(n19555), .A(n19545), .B(n19544), .ZN(
        P2_U3116) );
  AOI22_X1 U22508 ( .A1(n19640), .A2(n19572), .B1(n19752), .B2(n19550), .ZN(
        n19547) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19552), .B1(
        n19753), .B2(n19551), .ZN(n19546) );
  OAI211_X1 U22510 ( .C1(n19643), .C2(n19555), .A(n19547), .B(n19546), .ZN(
        P2_U3117) );
  AOI22_X1 U22511 ( .A1(n19762), .A2(n19572), .B1(n19760), .B2(n19550), .ZN(
        n19549) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19552), .B1(
        n19761), .B2(n19551), .ZN(n19548) );
  OAI211_X1 U22513 ( .C1(n19765), .C2(n19555), .A(n19549), .B(n19548), .ZN(
        P2_U3118) );
  AOI22_X1 U22514 ( .A1(n19770), .A2(n19572), .B1(n19766), .B2(n19550), .ZN(
        n19554) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19552), .B1(
        n19768), .B2(n19551), .ZN(n19553) );
  OAI211_X1 U22516 ( .C1(n19776), .C2(n19555), .A(n19554), .B(n19553), .ZN(
        P2_U3119) );
  AOI22_X1 U22517 ( .A1(n19728), .A2(n19584), .B1(n19718), .B2(n19583), .ZN(
        n19557) );
  AOI22_X1 U22518 ( .A1(n13454), .A2(n19573), .B1(n19572), .B2(n19652), .ZN(
        n19556) );
  OAI211_X1 U22519 ( .C1(n19559), .C2(n19558), .A(n19557), .B(n19556), .ZN(
        P2_U3120) );
  AOI22_X1 U22520 ( .A1(n19631), .A2(n19584), .B1(n19736), .B2(n19583), .ZN(
        n19561) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19574), .B1(
        n13449), .B2(n19573), .ZN(n19560) );
  OAI211_X1 U22522 ( .C1(n19634), .C2(n19567), .A(n19561), .B(n19560), .ZN(
        P2_U3122) );
  AOI22_X1 U22523 ( .A1(n19609), .A2(n19572), .B1(n19583), .B2(n19741), .ZN(
        n19563) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19574), .B1(
        n19294), .B2(n19573), .ZN(n19562) );
  OAI211_X1 U22525 ( .C1(n19564), .C2(n19606), .A(n19563), .B(n19562), .ZN(
        P2_U3123) );
  AOI22_X1 U22526 ( .A1(n19748), .A2(n19584), .B1(n19583), .B2(n19746), .ZN(
        n19566) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19574), .B1(
        n19747), .B2(n19573), .ZN(n19565) );
  OAI211_X1 U22528 ( .C1(n19751), .C2(n19567), .A(n19566), .B(n19565), .ZN(
        P2_U3124) );
  AOI22_X1 U22529 ( .A1(n19754), .A2(n19572), .B1(n19583), .B2(n19752), .ZN(
        n19569) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19574), .B1(
        n19753), .B2(n19573), .ZN(n19568) );
  OAI211_X1 U22531 ( .C1(n19759), .C2(n19606), .A(n19569), .B(n19568), .ZN(
        P2_U3125) );
  AOI22_X1 U22532 ( .A1(n19616), .A2(n19572), .B1(n19583), .B2(n19760), .ZN(
        n19571) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19574), .B1(
        n19761), .B2(n19573), .ZN(n19570) );
  OAI211_X1 U22534 ( .C1(n19620), .C2(n19606), .A(n19571), .B(n19570), .ZN(
        P2_U3126) );
  AOI22_X1 U22535 ( .A1(n19708), .A2(n19572), .B1(n19583), .B2(n19766), .ZN(
        n19576) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19574), .B1(
        n19768), .B2(n19573), .ZN(n19575) );
  OAI211_X1 U22537 ( .C1(n19713), .C2(n19606), .A(n19576), .B(n19575), .ZN(
        P2_U3127) );
  INV_X1 U22538 ( .A(n10892), .ZN(n19579) );
  AND2_X1 U22539 ( .A1(n19578), .A2(n19577), .ZN(n19601) );
  OAI21_X1 U22540 ( .B1(n19579), .B2(n19601), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19580) );
  OAI21_X1 U22541 ( .B1(n19582), .B2(n19581), .A(n19580), .ZN(n19602) );
  AOI22_X1 U22542 ( .A1(n19602), .A2(n13454), .B1(n19718), .B2(n19601), .ZN(
        n19588) );
  AOI221_X1 U22543 ( .B1(n19584), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19623), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19583), .ZN(n19585) );
  AOI211_X1 U22544 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n10892), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19585), .ZN(n19586) );
  OAI21_X1 U22545 ( .B1(n19586), .B2(n19601), .A(n19726), .ZN(n19603) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19728), .ZN(n19587) );
  OAI211_X1 U22547 ( .C1(n19731), .C2(n19606), .A(n19588), .B(n19587), .ZN(
        P2_U3128) );
  AOI22_X1 U22548 ( .A1(n19602), .A2(n13380), .B1(n13381), .B2(n19601), .ZN(
        n19590) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19689), .ZN(n19589) );
  OAI211_X1 U22550 ( .C1(n19692), .C2(n19606), .A(n19590), .B(n19589), .ZN(
        P2_U3129) );
  AOI22_X1 U22551 ( .A1(n19602), .A2(n13449), .B1(n19736), .B2(n19601), .ZN(
        n19592) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19631), .ZN(n19591) );
  OAI211_X1 U22553 ( .C1(n19634), .C2(n19606), .A(n19592), .B(n19591), .ZN(
        P2_U3130) );
  AOI22_X1 U22554 ( .A1(n19602), .A2(n19294), .B1(n19741), .B2(n19601), .ZN(
        n19594) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19742), .ZN(n19593) );
  OAI211_X1 U22556 ( .C1(n19745), .C2(n19606), .A(n19594), .B(n19593), .ZN(
        P2_U3131) );
  AOI22_X1 U22557 ( .A1(n19602), .A2(n19747), .B1(n19746), .B2(n19601), .ZN(
        n19596) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19748), .ZN(n19595) );
  OAI211_X1 U22559 ( .C1(n19751), .C2(n19606), .A(n19596), .B(n19595), .ZN(
        P2_U3132) );
  AOI22_X1 U22560 ( .A1(n19602), .A2(n19753), .B1(n19752), .B2(n19601), .ZN(
        n19598) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19640), .ZN(n19597) );
  OAI211_X1 U22562 ( .C1(n19643), .C2(n19606), .A(n19598), .B(n19597), .ZN(
        P2_U3133) );
  AOI22_X1 U22563 ( .A1(n19602), .A2(n19761), .B1(n19760), .B2(n19601), .ZN(
        n19600) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19762), .ZN(n19599) );
  OAI211_X1 U22565 ( .C1(n19765), .C2(n19606), .A(n19600), .B(n19599), .ZN(
        P2_U3134) );
  AOI22_X1 U22566 ( .A1(n19602), .A2(n19768), .B1(n19766), .B2(n19601), .ZN(
        n19605) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19603), .B1(
        n19623), .B2(n19770), .ZN(n19604) );
  OAI211_X1 U22568 ( .C1(n19776), .C2(n19606), .A(n19605), .B(n19604), .ZN(
        P2_U3135) );
  AOI22_X1 U22569 ( .A1(n19622), .A2(n13380), .B1(n19621), .B2(n13381), .ZN(
        n19608) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19732), .ZN(n19607) );
  OAI211_X1 U22571 ( .C1(n19735), .C2(n19651), .A(n19608), .B(n19607), .ZN(
        P2_U3137) );
  AOI22_X1 U22572 ( .A1(n19622), .A2(n19294), .B1(n19621), .B2(n19741), .ZN(
        n19611) );
  AOI22_X1 U22573 ( .A1(n19623), .A2(n19609), .B1(n19637), .B2(n19742), .ZN(
        n19610) );
  OAI211_X1 U22574 ( .C1(n19627), .C2(n20876), .A(n19611), .B(n19610), .ZN(
        P2_U3139) );
  AOI22_X1 U22575 ( .A1(n19622), .A2(n19747), .B1(n19621), .B2(n19746), .ZN(
        n19613) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19697), .ZN(n19612) );
  OAI211_X1 U22577 ( .C1(n19700), .C2(n19651), .A(n19613), .B(n19612), .ZN(
        P2_U3140) );
  AOI22_X1 U22578 ( .A1(n19622), .A2(n19753), .B1(n19621), .B2(n19752), .ZN(
        n19615) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19754), .ZN(n19614) );
  OAI211_X1 U22580 ( .C1(n19759), .C2(n19651), .A(n19615), .B(n19614), .ZN(
        P2_U3141) );
  AOI22_X1 U22581 ( .A1(n19622), .A2(n19761), .B1(n19621), .B2(n19760), .ZN(
        n19619) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19616), .ZN(n19618) );
  OAI211_X1 U22583 ( .C1(n19620), .C2(n19651), .A(n19619), .B(n19618), .ZN(
        P2_U3142) );
  INV_X1 U22584 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19626) );
  AOI22_X1 U22585 ( .A1(n19622), .A2(n19768), .B1(n19621), .B2(n19766), .ZN(
        n19625) );
  AOI22_X1 U22586 ( .A1(n19623), .A2(n19708), .B1(n19637), .B2(n19770), .ZN(
        n19624) );
  OAI211_X1 U22587 ( .C1(n19627), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P2_U3143) );
  AOI22_X1 U22588 ( .A1(n19647), .A2(n13380), .B1(n19646), .B2(n13381), .ZN(
        n19630) );
  INV_X1 U22589 ( .A(n19628), .ZN(n19648) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19648), .B1(
        n19670), .B2(n19689), .ZN(n19629) );
  OAI211_X1 U22591 ( .C1(n19692), .C2(n19651), .A(n19630), .B(n19629), .ZN(
        P2_U3145) );
  AOI22_X1 U22592 ( .A1(n19647), .A2(n13449), .B1(n19646), .B2(n19736), .ZN(
        n19633) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19648), .B1(
        n19670), .B2(n19631), .ZN(n19632) );
  OAI211_X1 U22594 ( .C1(n19634), .C2(n19651), .A(n19633), .B(n19632), .ZN(
        P2_U3146) );
  AOI22_X1 U22595 ( .A1(n19647), .A2(n19294), .B1(n19646), .B2(n19741), .ZN(
        n19636) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19648), .B1(
        n19670), .B2(n19742), .ZN(n19635) );
  OAI211_X1 U22597 ( .C1(n19745), .C2(n19651), .A(n19636), .B(n19635), .ZN(
        P2_U3147) );
  AOI22_X1 U22598 ( .A1(n19647), .A2(n19747), .B1(n19646), .B2(n19746), .ZN(
        n19639) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19648), .B1(
        n19637), .B2(n19697), .ZN(n19638) );
  OAI211_X1 U22600 ( .C1(n19700), .C2(n19668), .A(n19639), .B(n19638), .ZN(
        P2_U3148) );
  AOI22_X1 U22601 ( .A1(n19647), .A2(n19753), .B1(n19646), .B2(n19752), .ZN(
        n19642) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19648), .B1(
        n19670), .B2(n19640), .ZN(n19641) );
  OAI211_X1 U22603 ( .C1(n19643), .C2(n19651), .A(n19642), .B(n19641), .ZN(
        P2_U3149) );
  AOI22_X1 U22604 ( .A1(n19647), .A2(n19761), .B1(n19646), .B2(n19760), .ZN(
        n19645) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19648), .B1(
        n19670), .B2(n19762), .ZN(n19644) );
  OAI211_X1 U22606 ( .C1(n19765), .C2(n19651), .A(n19645), .B(n19644), .ZN(
        P2_U3150) );
  AOI22_X1 U22607 ( .A1(n19647), .A2(n19768), .B1(n19646), .B2(n19766), .ZN(
        n19650) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19648), .B1(
        n19670), .B2(n19770), .ZN(n19649) );
  OAI211_X1 U22609 ( .C1(n19776), .C2(n19651), .A(n19650), .B(n19649), .ZN(
        P2_U3151) );
  AOI22_X1 U22610 ( .A1(n19669), .A2(n13454), .B1(n19718), .B2(n19682), .ZN(
        n19654) );
  AOI22_X1 U22611 ( .A1(n19670), .A2(n19652), .B1(n19707), .B2(n19728), .ZN(
        n19653) );
  OAI211_X1 U22612 ( .C1(n19663), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3152) );
  AOI22_X1 U22613 ( .A1(n19669), .A2(n13449), .B1(n19736), .B2(n19682), .ZN(
        n19657) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19737), .ZN(n19656) );
  OAI211_X1 U22615 ( .C1(n19740), .C2(n19705), .A(n19657), .B(n19656), .ZN(
        P2_U3154) );
  AOI22_X1 U22616 ( .A1(n19669), .A2(n19294), .B1(n19682), .B2(n19741), .ZN(
        n19659) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19671), .B1(
        n19707), .B2(n19742), .ZN(n19658) );
  OAI211_X1 U22618 ( .C1(n19745), .C2(n19668), .A(n19659), .B(n19658), .ZN(
        P2_U3155) );
  AOI22_X1 U22619 ( .A1(n19669), .A2(n19747), .B1(n19682), .B2(n19746), .ZN(
        n19661) );
  AOI22_X1 U22620 ( .A1(n19670), .A2(n19697), .B1(n19707), .B2(n19748), .ZN(
        n19660) );
  OAI211_X1 U22621 ( .C1(n19663), .C2(n19662), .A(n19661), .B(n19660), .ZN(
        P2_U3156) );
  AOI22_X1 U22622 ( .A1(n19669), .A2(n19753), .B1(n19682), .B2(n19752), .ZN(
        n19665) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19754), .ZN(n19664) );
  OAI211_X1 U22624 ( .C1(n19759), .C2(n19705), .A(n19665), .B(n19664), .ZN(
        P2_U3157) );
  AOI22_X1 U22625 ( .A1(n19669), .A2(n19761), .B1(n19682), .B2(n19760), .ZN(
        n19667) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19671), .B1(
        n19707), .B2(n19762), .ZN(n19666) );
  OAI211_X1 U22627 ( .C1(n19765), .C2(n19668), .A(n19667), .B(n19666), .ZN(
        P2_U3158) );
  AOI22_X1 U22628 ( .A1(n19669), .A2(n19768), .B1(n19682), .B2(n19766), .ZN(
        n19673) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19708), .ZN(n19672) );
  OAI211_X1 U22630 ( .C1(n19713), .C2(n19705), .A(n19673), .B(n19672), .ZN(
        P2_U3159) );
  INV_X1 U22631 ( .A(n19714), .ZN(n19719) );
  NOR3_X2 U22632 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19874), .A3(
        n19719), .ZN(n19706) );
  AOI22_X1 U22633 ( .A1(n19728), .A2(n19755), .B1(n19718), .B2(n19706), .ZN(
        n19688) );
  INV_X1 U22634 ( .A(n19675), .ZN(n19683) );
  NOR3_X1 U22635 ( .A1(n19683), .A2(n19706), .A3(n19676), .ZN(n19681) );
  OAI21_X1 U22636 ( .B1(n19755), .B2(n19707), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19677) );
  NAND2_X1 U22637 ( .A1(n19677), .A2(n19869), .ZN(n19686) );
  AOI221_X1 U22638 ( .B1(n19678), .B2(n19686), .C1(n19678), .C2(n19682), .A(
        n19706), .ZN(n19679) );
  NOR2_X1 U22639 ( .A1(n19706), .A2(n19682), .ZN(n19685) );
  OAI21_X1 U22640 ( .B1(n19683), .B2(n19706), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19684) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19710), .B1(
        n13454), .B2(n19709), .ZN(n19687) );
  OAI211_X1 U22642 ( .C1(n19731), .C2(n19705), .A(n19688), .B(n19687), .ZN(
        P2_U3160) );
  AOI22_X1 U22643 ( .A1(n19689), .A2(n19755), .B1(n13381), .B2(n19706), .ZN(
        n19691) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19710), .B1(
        n13380), .B2(n19709), .ZN(n19690) );
  OAI211_X1 U22645 ( .C1(n19692), .C2(n19705), .A(n19691), .B(n19690), .ZN(
        P2_U3161) );
  AOI22_X1 U22646 ( .A1(n19737), .A2(n19707), .B1(n19736), .B2(n19706), .ZN(
        n19694) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19710), .B1(
        n13449), .B2(n19709), .ZN(n19693) );
  OAI211_X1 U22648 ( .C1(n19740), .C2(n19775), .A(n19694), .B(n19693), .ZN(
        P2_U3162) );
  AOI22_X1 U22649 ( .A1(n19742), .A2(n19755), .B1(n19741), .B2(n19706), .ZN(
        n19696) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19710), .B1(
        n19294), .B2(n19709), .ZN(n19695) );
  OAI211_X1 U22651 ( .C1(n19745), .C2(n19705), .A(n19696), .B(n19695), .ZN(
        P2_U3163) );
  AOI22_X1 U22652 ( .A1(n19697), .A2(n19707), .B1(n19746), .B2(n19706), .ZN(
        n19699) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19710), .B1(
        n19747), .B2(n19709), .ZN(n19698) );
  OAI211_X1 U22654 ( .C1(n19700), .C2(n19775), .A(n19699), .B(n19698), .ZN(
        P2_U3164) );
  AOI22_X1 U22655 ( .A1(n19754), .A2(n19707), .B1(n19752), .B2(n19706), .ZN(
        n19702) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19710), .B1(
        n19753), .B2(n19709), .ZN(n19701) );
  OAI211_X1 U22657 ( .C1(n19759), .C2(n19775), .A(n19702), .B(n19701), .ZN(
        P2_U3165) );
  AOI22_X1 U22658 ( .A1(n19762), .A2(n19755), .B1(n19760), .B2(n19706), .ZN(
        n19704) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19710), .B1(
        n19761), .B2(n19709), .ZN(n19703) );
  OAI211_X1 U22660 ( .C1(n19765), .C2(n19705), .A(n19704), .B(n19703), .ZN(
        P2_U3166) );
  AOI22_X1 U22661 ( .A1(n19708), .A2(n19707), .B1(n19766), .B2(n19706), .ZN(
        n19712) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19710), .B1(
        n19768), .B2(n19709), .ZN(n19711) );
  OAI211_X1 U22663 ( .C1(n19713), .C2(n19775), .A(n19712), .B(n19711), .ZN(
        P2_U3167) );
  NAND2_X1 U22664 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19714), .ZN(
        n19717) );
  INV_X1 U22665 ( .A(n19724), .ZN(n19715) );
  OAI21_X1 U22666 ( .B1(n19715), .B2(n19767), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19716) );
  OAI21_X1 U22667 ( .B1(n19717), .B2(n19722), .A(n19716), .ZN(n19769) );
  AOI22_X1 U22668 ( .A1(n19769), .A2(n13454), .B1(n19767), .B2(n19718), .ZN(
        n19730) );
  OAI22_X1 U22669 ( .A1(n19721), .A2(n19720), .B1(n19719), .B2(n19874), .ZN(
        n19727) );
  OAI211_X1 U22670 ( .C1(n19724), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19723), 
        .B(n19722), .ZN(n19725) );
  NAND3_X1 U22671 ( .A1(n19727), .A2(n19726), .A3(n19725), .ZN(n19772) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19728), .ZN(n19729) );
  OAI211_X1 U22673 ( .C1(n19731), .C2(n19775), .A(n19730), .B(n19729), .ZN(
        P2_U3168) );
  AOI22_X1 U22674 ( .A1(n19769), .A2(n13380), .B1(n19767), .B2(n13381), .ZN(
        n19734) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19772), .B1(
        n19755), .B2(n19732), .ZN(n19733) );
  OAI211_X1 U22676 ( .C1(n19735), .C2(n19758), .A(n19734), .B(n19733), .ZN(
        P2_U3169) );
  AOI22_X1 U22677 ( .A1(n19769), .A2(n13449), .B1(n19767), .B2(n19736), .ZN(
        n19739) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19772), .B1(
        n19755), .B2(n19737), .ZN(n19738) );
  OAI211_X1 U22679 ( .C1(n19740), .C2(n19758), .A(n19739), .B(n19738), .ZN(
        P2_U3170) );
  AOI22_X1 U22680 ( .A1(n19769), .A2(n19294), .B1(n19767), .B2(n19741), .ZN(
        n19744) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19742), .ZN(n19743) );
  OAI211_X1 U22682 ( .C1(n19745), .C2(n19775), .A(n19744), .B(n19743), .ZN(
        P2_U3171) );
  AOI22_X1 U22683 ( .A1(n19769), .A2(n19747), .B1(n19767), .B2(n19746), .ZN(
        n19750) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19748), .ZN(n19749) );
  OAI211_X1 U22685 ( .C1(n19751), .C2(n19775), .A(n19750), .B(n19749), .ZN(
        P2_U3172) );
  AOI22_X1 U22686 ( .A1(n19769), .A2(n19753), .B1(n19767), .B2(n19752), .ZN(
        n19757) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19772), .B1(
        n19755), .B2(n19754), .ZN(n19756) );
  OAI211_X1 U22688 ( .C1(n19759), .C2(n19758), .A(n19757), .B(n19756), .ZN(
        P2_U3173) );
  AOI22_X1 U22689 ( .A1(n19769), .A2(n19761), .B1(n19767), .B2(n19760), .ZN(
        n19764) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19762), .ZN(n19763) );
  OAI211_X1 U22691 ( .C1(n19765), .C2(n19775), .A(n19764), .B(n19763), .ZN(
        P2_U3174) );
  AOI22_X1 U22692 ( .A1(n19769), .A2(n19768), .B1(n19767), .B2(n19766), .ZN(
        n19774) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19772), .B1(
        n19771), .B2(n19770), .ZN(n19773) );
  OAI211_X1 U22694 ( .C1(n19776), .C2(n19775), .A(n19774), .B(n19773), .ZN(
        P2_U3175) );
  AOI21_X1 U22695 ( .B1(n19779), .B2(n19778), .A(n19777), .ZN(n19783) );
  OAI211_X1 U22696 ( .C1(n19784), .C2(n19780), .A(n19786), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19781) );
  OAI211_X1 U22697 ( .C1(n19784), .C2(n19783), .A(n19782), .B(n19781), .ZN(
        P2_U3177) );
  AND2_X1 U22698 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19785), .ZN(
        P2_U3179) );
  AND2_X1 U22699 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19785), .ZN(
        P2_U3180) );
  AND2_X1 U22700 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19785), .ZN(
        P2_U3181) );
  AND2_X1 U22701 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19785), .ZN(
        P2_U3182) );
  AND2_X1 U22702 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19785), .ZN(
        P2_U3183) );
  AND2_X1 U22703 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19785), .ZN(
        P2_U3184) );
  AND2_X1 U22704 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19785), .ZN(
        P2_U3185) );
  AND2_X1 U22705 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19785), .ZN(
        P2_U3186) );
  AND2_X1 U22706 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19785), .ZN(
        P2_U3187) );
  AND2_X1 U22707 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19785), .ZN(
        P2_U3188) );
  AND2_X1 U22708 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19785), .ZN(
        P2_U3189) );
  AND2_X1 U22709 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19785), .ZN(
        P2_U3190) );
  AND2_X1 U22710 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19785), .ZN(
        P2_U3191) );
  AND2_X1 U22711 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19785), .ZN(
        P2_U3192) );
  AND2_X1 U22712 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19785), .ZN(
        P2_U3193) );
  AND2_X1 U22713 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19785), .ZN(
        P2_U3194) );
  AND2_X1 U22714 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19785), .ZN(
        P2_U3195) );
  AND2_X1 U22715 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19785), .ZN(
        P2_U3196) );
  AND2_X1 U22716 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19785), .ZN(
        P2_U3197) );
  AND2_X1 U22717 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19785), .ZN(
        P2_U3198) );
  AND2_X1 U22718 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19785), .ZN(
        P2_U3199) );
  AND2_X1 U22719 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19785), .ZN(
        P2_U3200) );
  AND2_X1 U22720 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19785), .ZN(P2_U3201) );
  AND2_X1 U22721 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19785), .ZN(P2_U3202) );
  AND2_X1 U22722 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19785), .ZN(P2_U3203) );
  AND2_X1 U22723 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19785), .ZN(P2_U3204) );
  AND2_X1 U22724 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19785), .ZN(P2_U3205) );
  AND2_X1 U22725 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19785), .ZN(P2_U3206) );
  AND2_X1 U22726 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19785), .ZN(P2_U3207) );
  AND2_X1 U22727 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19785), .ZN(P2_U3208) );
  INV_X1 U22728 ( .A(NA), .ZN(n20787) );
  OAI21_X1 U22729 ( .B1(n20787), .B2(n19792), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19801) );
  INV_X1 U22730 ( .A(n19801), .ZN(n19789) );
  NAND2_X1 U22731 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19786), .ZN(n19799) );
  INV_X1 U22732 ( .A(n19799), .ZN(n19790) );
  INV_X1 U22733 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21048) );
  NOR3_X1 U22734 ( .A1(n19790), .A2(n21048), .A3(n19791), .ZN(n19788) );
  OAI21_X1 U22735 ( .B1(HOLD), .B2(n21048), .A(n19796), .ZN(n19787) );
  OAI22_X1 U22736 ( .A1(n19789), .A2(n19788), .B1(n19909), .B2(n19787), .ZN(
        P2_U3209) );
  NOR2_X1 U22737 ( .A1(n21041), .A2(n19790), .ZN(n19794) );
  NOR2_X1 U22738 ( .A1(HOLD), .A2(n19791), .ZN(n19800) );
  OAI211_X1 U22739 ( .C1(n19800), .C2(n19802), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19792), .ZN(n19793) );
  OAI211_X1 U22740 ( .C1(n19795), .C2(n20782), .A(n19794), .B(n19793), .ZN(
        P2_U3210) );
  OAI22_X1 U22741 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19796), .B1(NA), 
        .B2(n19799), .ZN(n19797) );
  OAI211_X1 U22742 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19797), .ZN(n19798) );
  OAI221_X1 U22743 ( .B1(n19801), .B2(n19800), .C1(n19801), .C2(n19799), .A(
        n19798), .ZN(P2_U3211) );
  OAI222_X1 U22744 ( .A1(n19857), .A2(n19804), .B1(n19803), .B2(n19909), .C1(
        n13003), .C2(n19855), .ZN(P2_U3212) );
  OAI222_X1 U22745 ( .A1(n19857), .A2(n19806), .B1(n19805), .B2(n19909), .C1(
        n19804), .C2(n19855), .ZN(P2_U3213) );
  OAI222_X1 U22746 ( .A1(n19857), .A2(n19808), .B1(n19807), .B2(n19909), .C1(
        n19806), .C2(n19855), .ZN(P2_U3214) );
  INV_X1 U22747 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19810) );
  OAI222_X1 U22748 ( .A1(n19857), .A2(n19810), .B1(n19809), .B2(n19909), .C1(
        n19808), .C2(n19855), .ZN(P2_U3215) );
  OAI222_X1 U22749 ( .A1(n19857), .A2(n19812), .B1(n19811), .B2(n19909), .C1(
        n19810), .C2(n19855), .ZN(P2_U3216) );
  OAI222_X1 U22750 ( .A1(n19857), .A2(n19814), .B1(n19813), .B2(n19909), .C1(
        n19812), .C2(n19855), .ZN(P2_U3217) );
  INV_X1 U22751 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19816) );
  OAI222_X1 U22752 ( .A1(n19857), .A2(n19816), .B1(n19815), .B2(n19909), .C1(
        n19814), .C2(n19855), .ZN(P2_U3218) );
  OAI222_X1 U22753 ( .A1(n19857), .A2(n20975), .B1(n19817), .B2(n19909), .C1(
        n19816), .C2(n19855), .ZN(P2_U3219) );
  OAI222_X1 U22754 ( .A1(n19857), .A2(n19819), .B1(n19818), .B2(n19909), .C1(
        n20975), .C2(n19855), .ZN(P2_U3220) );
  OAI222_X1 U22755 ( .A1(n19857), .A2(n19821), .B1(n19820), .B2(n19909), .C1(
        n19819), .C2(n19855), .ZN(P2_U3221) );
  OAI222_X1 U22756 ( .A1(n19857), .A2(n19823), .B1(n19822), .B2(n19909), .C1(
        n19821), .C2(n19855), .ZN(P2_U3222) );
  OAI222_X1 U22757 ( .A1(n19857), .A2(n15193), .B1(n19824), .B2(n19909), .C1(
        n19823), .C2(n19855), .ZN(P2_U3223) );
  OAI222_X1 U22758 ( .A1(n19857), .A2(n15182), .B1(n19825), .B2(n19909), .C1(
        n15193), .C2(n19855), .ZN(P2_U3224) );
  OAI222_X1 U22759 ( .A1(n19857), .A2(n19827), .B1(n19826), .B2(n19909), .C1(
        n15182), .C2(n19855), .ZN(P2_U3225) );
  OAI222_X1 U22760 ( .A1(n19857), .A2(n15153), .B1(n19828), .B2(n19909), .C1(
        n19827), .C2(n19855), .ZN(P2_U3226) );
  OAI222_X1 U22761 ( .A1(n19857), .A2(n19830), .B1(n19829), .B2(n19909), .C1(
        n15153), .C2(n19855), .ZN(P2_U3227) );
  OAI222_X1 U22762 ( .A1(n19857), .A2(n15135), .B1(n19831), .B2(n19909), .C1(
        n19830), .C2(n19855), .ZN(P2_U3228) );
  OAI222_X1 U22763 ( .A1(n19857), .A2(n19833), .B1(n19832), .B2(n19909), .C1(
        n15135), .C2(n19855), .ZN(P2_U3229) );
  OAI222_X1 U22764 ( .A1(n19857), .A2(n19835), .B1(n19834), .B2(n19909), .C1(
        n19833), .C2(n19855), .ZN(P2_U3230) );
  OAI222_X1 U22765 ( .A1(n19857), .A2(n19837), .B1(n19836), .B2(n19909), .C1(
        n19835), .C2(n19855), .ZN(P2_U3231) );
  INV_X1 U22766 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19839) );
  OAI222_X1 U22767 ( .A1(n19857), .A2(n19839), .B1(n19838), .B2(n19909), .C1(
        n19837), .C2(n19855), .ZN(P2_U3232) );
  OAI222_X1 U22768 ( .A1(n19857), .A2(n19841), .B1(n19840), .B2(n19909), .C1(
        n19839), .C2(n19855), .ZN(P2_U3233) );
  OAI222_X1 U22769 ( .A1(n19857), .A2(n19843), .B1(n19842), .B2(n19909), .C1(
        n19841), .C2(n19855), .ZN(P2_U3234) );
  OAI222_X1 U22770 ( .A1(n19857), .A2(n19845), .B1(n19844), .B2(n19909), .C1(
        n19843), .C2(n19855), .ZN(P2_U3235) );
  OAI222_X1 U22771 ( .A1(n19857), .A2(n19847), .B1(n19846), .B2(n19909), .C1(
        n19845), .C2(n19855), .ZN(P2_U3236) );
  OAI222_X1 U22772 ( .A1(n19857), .A2(n19850), .B1(n19848), .B2(n19909), .C1(
        n19847), .C2(n19855), .ZN(P2_U3237) );
  OAI222_X1 U22773 ( .A1(n19855), .A2(n19850), .B1(n19849), .B2(n19909), .C1(
        n19851), .C2(n19857), .ZN(P2_U3238) );
  OAI222_X1 U22774 ( .A1(n19857), .A2(n19853), .B1(n19852), .B2(n19909), .C1(
        n19851), .C2(n19855), .ZN(P2_U3239) );
  OAI222_X1 U22775 ( .A1(n19857), .A2(n11609), .B1(n19854), .B2(n19909), .C1(
        n19853), .C2(n19855), .ZN(P2_U3240) );
  OAI222_X1 U22776 ( .A1(n19857), .A2(n20991), .B1(n19856), .B2(n19909), .C1(
        n11609), .C2(n19855), .ZN(P2_U3241) );
  OAI22_X1 U22777 ( .A1(n19910), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19909), .ZN(n19858) );
  INV_X1 U22778 ( .A(n19858), .ZN(P2_U3585) );
  MUX2_X1 U22779 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19910), .Z(P2_U3586) );
  OAI22_X1 U22780 ( .A1(n19910), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19909), .ZN(n19859) );
  INV_X1 U22781 ( .A(n19859), .ZN(P2_U3587) );
  OAI22_X1 U22782 ( .A1(n19910), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19909), .ZN(n19860) );
  INV_X1 U22783 ( .A(n19860), .ZN(P2_U3588) );
  OAI21_X1 U22784 ( .B1(n19864), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19862), 
        .ZN(n19861) );
  INV_X1 U22785 ( .A(n19861), .ZN(P2_U3591) );
  OAI21_X1 U22786 ( .B1(n19864), .B2(n19863), .A(n19862), .ZN(P2_U3592) );
  AND2_X1 U22787 ( .A1(n19869), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19882) );
  NAND2_X1 U22788 ( .A1(n19865), .A2(n19882), .ZN(n19875) );
  NAND3_X1 U22789 ( .A1(n19887), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19866), 
        .ZN(n19867) );
  NAND2_X1 U22790 ( .A1(n19867), .A2(n19892), .ZN(n19876) );
  NAND2_X1 U22791 ( .A1(n19875), .A2(n19876), .ZN(n19872) );
  AOI222_X1 U22792 ( .A1(n19872), .A2(n19871), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19870), .C1(n19869), .C2(n19868), .ZN(n19873) );
  INV_X1 U22793 ( .A(n19901), .ZN(n19898) );
  AOI22_X1 U22794 ( .A1(n19901), .A2(n19874), .B1(n19873), .B2(n19898), .ZN(
        P2_U3602) );
  OAI21_X1 U22795 ( .B1(n19877), .B2(n19876), .A(n19875), .ZN(n19878) );
  AOI21_X1 U22796 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19879), .A(n19878), 
        .ZN(n19880) );
  AOI22_X1 U22797 ( .A1(n19901), .A2(n19881), .B1(n19880), .B2(n19898), .ZN(
        P2_U3603) );
  INV_X1 U22798 ( .A(n19882), .ZN(n19886) );
  INV_X1 U22799 ( .A(n19883), .ZN(n19884) );
  NAND3_X1 U22800 ( .A1(n19887), .A2(n19892), .A3(n19884), .ZN(n19885) );
  OAI21_X1 U22801 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(n19888) );
  AOI21_X1 U22802 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19889), .A(n19888), 
        .ZN(n19890) );
  AOI22_X1 U22803 ( .A1(n19901), .A2(n19891), .B1(n19890), .B2(n19898), .ZN(
        P2_U3604) );
  INV_X1 U22804 ( .A(n19892), .ZN(n19893) );
  OAI22_X1 U22805 ( .A1(n19894), .A2(n19893), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19678), .ZN(n19895) );
  AOI21_X1 U22806 ( .B1(n19897), .B2(n19896), .A(n19895), .ZN(n19899) );
  AOI22_X1 U22807 ( .A1(n19901), .A2(n19900), .B1(n19899), .B2(n19898), .ZN(
        P2_U3605) );
  INV_X1 U22808 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19902) );
  AOI22_X1 U22809 ( .A1(n19909), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19902), 
        .B2(n19910), .ZN(P2_U3608) );
  AOI21_X1 U22810 ( .B1(n19905), .B2(n19904), .A(n19903), .ZN(n19907) );
  NAND2_X1 U22811 ( .A1(n19908), .A2(P2_MORE_REG_SCAN_IN), .ZN(n19906) );
  OAI21_X1 U22812 ( .B1(n19908), .B2(n19907), .A(n19906), .ZN(P2_U3609) );
  OAI22_X1 U22813 ( .A1(n19910), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19909), .ZN(n19911) );
  INV_X1 U22814 ( .A(n19911), .ZN(P2_U3611) );
  AOI21_X1 U22815 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20794), .A(n20970), 
        .ZN(n19918) );
  INV_X1 U22816 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19912) );
  NAND2_X2 U22817 ( .A1(n20970), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20869) );
  AOI21_X1 U22818 ( .B1(n19918), .B2(n19912), .A(n20868), .ZN(P1_U2802) );
  OAI21_X1 U22819 ( .B1(n19914), .B2(n19913), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19915) );
  OAI21_X1 U22820 ( .B1(n19916), .B2(n20777), .A(n19915), .ZN(P1_U2803) );
  NOR2_X1 U22821 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19919) );
  OAI21_X1 U22822 ( .B1(n19919), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20869), .ZN(
        n19917) );
  OAI21_X1 U22823 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20869), .A(n19917), 
        .ZN(P1_U2804) );
  NOR2_X1 U22824 ( .A1(n20868), .A2(n19918), .ZN(n20845) );
  OAI21_X1 U22825 ( .B1(BS16), .B2(n19919), .A(n20845), .ZN(n20843) );
  OAI21_X1 U22826 ( .B1(n20845), .B2(n20857), .A(n20843), .ZN(P1_U2805) );
  OAI21_X1 U22827 ( .B1(n19922), .B2(n19921), .A(n19920), .ZN(P1_U2806) );
  NOR4_X1 U22828 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19932) );
  NOR4_X1 U22829 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19931) );
  INV_X1 U22830 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20850) );
  INV_X1 U22831 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20844) );
  NOR4_X1 U22832 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19923) );
  OAI21_X1 U22833 ( .B1(n20850), .B2(n20844), .A(n19923), .ZN(n19929) );
  NOR4_X1 U22834 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19927) );
  NOR4_X1 U22835 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19926) );
  NOR4_X1 U22836 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19925) );
  NOR4_X1 U22837 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19924) );
  NAND4_X1 U22838 ( .A1(n19927), .A2(n19926), .A3(n19925), .A4(n19924), .ZN(
        n19928) );
  NOR4_X1 U22839 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(n19929), .A4(n19928), .ZN(n19930) );
  NAND3_X1 U22840 ( .A1(n19932), .A2(n19931), .A3(n19930), .ZN(n19933) );
  NOR2_X1 U22841 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n19933), .ZN(n19935) );
  INV_X1 U22842 ( .A(n19933), .ZN(n20853) );
  NOR2_X1 U22843 ( .A1(n20853), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19934)
         );
  NOR2_X1 U22844 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n19933), .ZN(n20846) );
  NAND3_X1 U22845 ( .A1(n20846), .A2(n20850), .A3(n20844), .ZN(n19936) );
  OAI21_X1 U22846 ( .B1(n19935), .B2(n19934), .A(n19936), .ZN(P1_U2807) );
  INV_X1 U22847 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19937) );
  NAND2_X1 U22848 ( .A1(n19935), .A2(n20844), .ZN(n20851) );
  OAI211_X1 U22849 ( .C1(n20853), .C2(n19937), .A(n19936), .B(n20851), .ZN(
        P1_U2808) );
  AOI21_X1 U22850 ( .B1(n19962), .B2(n19938), .A(n19961), .ZN(n19953) );
  AOI22_X1 U22851 ( .A1(n19963), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19987), .B2(
        n19939), .ZN(n19940) );
  OAI211_X1 U22852 ( .C1(n19949), .C2(n19941), .A(n19940), .B(n20101), .ZN(
        n19942) );
  AOI21_X1 U22853 ( .B1(n19977), .B2(n20006), .A(n19942), .ZN(n19946) );
  INV_X1 U22854 ( .A(n19943), .ZN(n20007) );
  AOI22_X1 U22855 ( .A1(n20007), .A2(n12623), .B1(n19944), .B2(n13771), .ZN(
        n19945) );
  OAI211_X1 U22856 ( .C1(n19953), .C2(n13771), .A(n19946), .B(n19945), .ZN(
        P1_U2831) );
  NAND2_X1 U22857 ( .A1(n19963), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n19947) );
  OAI211_X1 U22858 ( .C1(n19949), .C2(n19948), .A(n19947), .B(n20101), .ZN(
        n19950) );
  AOI21_X1 U22859 ( .B1(n19951), .B2(n19977), .A(n19950), .ZN(n19960) );
  NOR3_X1 U22860 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19952), .A3(n19981), .ZN(
        n19957) );
  OAI22_X1 U22861 ( .A1(n19955), .A2(n19954), .B1(n13724), .B2(n19953), .ZN(
        n19956) );
  AOI211_X1 U22862 ( .C1(n19987), .C2(n19958), .A(n19957), .B(n19956), .ZN(
        n19959) );
  NAND2_X1 U22863 ( .A1(n19960), .A2(n19959), .ZN(P1_U2832) );
  NAND2_X1 U22864 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19966) );
  AOI21_X1 U22865 ( .B1(n19962), .B2(n19966), .A(n19961), .ZN(n19986) );
  INV_X1 U22866 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19972) );
  AOI22_X1 U22867 ( .A1(n19963), .A2(P1_EBX_REG_7__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19989), .ZN(n19964) );
  INV_X1 U22868 ( .A(n19964), .ZN(n19965) );
  AOI211_X1 U22869 ( .C1(n19977), .C2(n9704), .A(n12840), .B(n19965), .ZN(
        n19971) );
  NOR3_X1 U22870 ( .A1(n19981), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n19966), .ZN(
        n19969) );
  NOR2_X1 U22871 ( .A1(n19974), .A2(n19967), .ZN(n19968) );
  AOI211_X1 U22872 ( .C1(n20011), .C2(n12623), .A(n19969), .B(n19968), .ZN(
        n19970) );
  OAI211_X1 U22873 ( .C1(n19986), .C2(n19972), .A(n19971), .B(n19970), .ZN(
        P1_U2833) );
  INV_X1 U22874 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20801) );
  NAND2_X1 U22875 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20801), .ZN(n19982) );
  AOI21_X1 U22876 ( .B1(n19989), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n12840), .ZN(n19973) );
  OAI21_X1 U22877 ( .B1(n19975), .B2(n19974), .A(n19973), .ZN(n19976) );
  AOI21_X1 U22878 ( .B1(n19963), .B2(P1_EBX_REG_6__SCAN_IN), .A(n19976), .ZN(
        n19980) );
  NAND2_X1 U22879 ( .A1(n19978), .A2(n19977), .ZN(n19979) );
  OAI211_X1 U22880 ( .C1(n19982), .C2(n19981), .A(n19980), .B(n19979), .ZN(
        n19983) );
  AOI21_X1 U22881 ( .B1(n19984), .B2(n12623), .A(n19983), .ZN(n19985) );
  OAI21_X1 U22882 ( .B1(n19986), .B2(n20801), .A(n19985), .ZN(P1_U2834) );
  AOI22_X1 U22883 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19989), .B1(
        n19988), .B2(n19987), .ZN(n20003) );
  INV_X1 U22884 ( .A(n19990), .ZN(n20000) );
  INV_X1 U22885 ( .A(n19991), .ZN(n19998) );
  INV_X1 U22886 ( .A(n19992), .ZN(n19996) );
  OAI21_X1 U22887 ( .B1(n19994), .B2(n20946), .A(n19993), .ZN(n19995) );
  AOI22_X1 U22888 ( .A1(n19996), .A2(n19995), .B1(n19963), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n19997) );
  OAI21_X1 U22889 ( .B1(n20564), .B2(n19998), .A(n19997), .ZN(n19999) );
  AOI21_X1 U22890 ( .B1(n20001), .B2(n20000), .A(n19999), .ZN(n20002) );
  OAI211_X1 U22891 ( .C1(n20005), .C2(n20004), .A(n20003), .B(n20002), .ZN(
        P1_U2838) );
  AOI22_X1 U22892 ( .A1(n20007), .A2(n20010), .B1(n12863), .B2(n20006), .ZN(
        n20008) );
  OAI21_X1 U22893 ( .B1(n20014), .B2(n20009), .A(n20008), .ZN(P1_U2863) );
  AOI22_X1 U22894 ( .A1(n20011), .A2(n20010), .B1(n12863), .B2(n9704), .ZN(
        n20012) );
  OAI21_X1 U22895 ( .B1(n20014), .B2(n20013), .A(n20012), .ZN(P1_U2865) );
  AOI22_X1 U22896 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20016) );
  OAI21_X1 U22897 ( .B1(n13333), .B2(n20046), .A(n20016), .ZN(P1_U2921) );
  INV_X1 U22898 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20018) );
  AOI22_X1 U22899 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20017) );
  OAI21_X1 U22900 ( .B1(n20018), .B2(n20046), .A(n20017), .ZN(P1_U2922) );
  INV_X1 U22901 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20020) );
  AOI22_X1 U22902 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20019) );
  OAI21_X1 U22903 ( .B1(n20020), .B2(n20046), .A(n20019), .ZN(P1_U2923) );
  INV_X1 U22904 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U22905 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20021) );
  OAI21_X1 U22906 ( .B1(n20022), .B2(n20046), .A(n20021), .ZN(P1_U2924) );
  INV_X1 U22907 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20024) );
  AOI22_X1 U22908 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20023) );
  OAI21_X1 U22909 ( .B1(n20024), .B2(n20046), .A(n20023), .ZN(P1_U2925) );
  INV_X1 U22910 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20026) );
  AOI22_X1 U22911 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20025) );
  OAI21_X1 U22912 ( .B1(n20026), .B2(n20046), .A(n20025), .ZN(P1_U2926) );
  INV_X1 U22913 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20028) );
  AOI22_X1 U22914 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20027) );
  OAI21_X1 U22915 ( .B1(n20028), .B2(n20046), .A(n20027), .ZN(P1_U2927) );
  INV_X1 U22916 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20030) );
  AOI22_X1 U22917 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20865), .B1(n20043), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20029) );
  OAI21_X1 U22918 ( .B1(n20030), .B2(n20046), .A(n20029), .ZN(P1_U2928) );
  AOI22_X1 U22919 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U22920 ( .B1(n13665), .B2(n20046), .A(n20031), .ZN(P1_U2929) );
  AOI22_X1 U22921 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U22922 ( .B1(n12027), .B2(n20046), .A(n20032), .ZN(P1_U2930) );
  AOI22_X1 U22923 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U22924 ( .B1(n20034), .B2(n20046), .A(n20033), .ZN(P1_U2931) );
  AOI22_X1 U22925 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U22926 ( .B1(n20036), .B2(n20046), .A(n20035), .ZN(P1_U2932) );
  AOI22_X1 U22927 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U22928 ( .B1(n20038), .B2(n20046), .A(n20037), .ZN(P1_U2933) );
  AOI22_X1 U22929 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20039) );
  OAI21_X1 U22930 ( .B1(n20040), .B2(n20046), .A(n20039), .ZN(P1_U2934) );
  AOI22_X1 U22931 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20041) );
  OAI21_X1 U22932 ( .B1(n20042), .B2(n20046), .A(n20041), .ZN(P1_U2935) );
  AOI22_X1 U22933 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20044), .B1(n20043), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20045) );
  OAI21_X1 U22934 ( .B1(n20047), .B2(n20046), .A(n20045), .ZN(P1_U2936) );
  AOI22_X1 U22935 ( .A1(n20076), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20075), .ZN(n20049) );
  NAND2_X1 U22936 ( .A1(n20061), .A2(n20048), .ZN(n20063) );
  NAND2_X1 U22937 ( .A1(n20049), .A2(n20063), .ZN(P1_U2945) );
  AOI22_X1 U22938 ( .A1(n20076), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20075), .ZN(n20051) );
  NAND2_X1 U22939 ( .A1(n20061), .A2(n20050), .ZN(n20065) );
  NAND2_X1 U22940 ( .A1(n20051), .A2(n20065), .ZN(P1_U2946) );
  AOI22_X1 U22941 ( .A1(n20076), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20075), .ZN(n20053) );
  NAND2_X1 U22942 ( .A1(n20061), .A2(n20052), .ZN(n20067) );
  NAND2_X1 U22943 ( .A1(n20053), .A2(n20067), .ZN(P1_U2947) );
  AOI22_X1 U22944 ( .A1(n20076), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20075), .ZN(n20055) );
  NAND2_X1 U22945 ( .A1(n20061), .A2(n20054), .ZN(n20069) );
  NAND2_X1 U22946 ( .A1(n20055), .A2(n20069), .ZN(P1_U2948) );
  AOI22_X1 U22947 ( .A1(n20076), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20075), .ZN(n20057) );
  NAND2_X1 U22948 ( .A1(n20061), .A2(n20056), .ZN(n20071) );
  NAND2_X1 U22949 ( .A1(n20057), .A2(n20071), .ZN(P1_U2949) );
  AOI22_X1 U22950 ( .A1(n20076), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20075), .ZN(n20059) );
  NAND2_X1 U22951 ( .A1(n20061), .A2(n20058), .ZN(n20073) );
  NAND2_X1 U22952 ( .A1(n20059), .A2(n20073), .ZN(P1_U2950) );
  AOI22_X1 U22953 ( .A1(n20076), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20075), .ZN(n20062) );
  NAND2_X1 U22954 ( .A1(n20061), .A2(n20060), .ZN(n20077) );
  NAND2_X1 U22955 ( .A1(n20062), .A2(n20077), .ZN(P1_U2951) );
  AOI22_X1 U22956 ( .A1(n20076), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20075), .ZN(n20064) );
  NAND2_X1 U22957 ( .A1(n20064), .A2(n20063), .ZN(P1_U2960) );
  AOI22_X1 U22958 ( .A1(n20076), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20075), .ZN(n20066) );
  NAND2_X1 U22959 ( .A1(n20066), .A2(n20065), .ZN(P1_U2961) );
  AOI22_X1 U22960 ( .A1(n20076), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20075), .ZN(n20068) );
  NAND2_X1 U22961 ( .A1(n20068), .A2(n20067), .ZN(P1_U2962) );
  AOI22_X1 U22962 ( .A1(n20076), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20075), .ZN(n20070) );
  NAND2_X1 U22963 ( .A1(n20070), .A2(n20069), .ZN(P1_U2963) );
  AOI22_X1 U22964 ( .A1(n20076), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20075), .ZN(n20072) );
  NAND2_X1 U22965 ( .A1(n20072), .A2(n20071), .ZN(P1_U2964) );
  AOI22_X1 U22966 ( .A1(n20076), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20075), .ZN(n20074) );
  NAND2_X1 U22967 ( .A1(n20074), .A2(n20073), .ZN(P1_U2965) );
  AOI22_X1 U22968 ( .A1(n20076), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20075), .ZN(n20078) );
  NAND2_X1 U22969 ( .A1(n20078), .A2(n20077), .ZN(P1_U2966) );
  INV_X1 U22970 ( .A(n20079), .ZN(n20083) );
  INV_X1 U22971 ( .A(n20080), .ZN(n20081) );
  AOI21_X1 U22972 ( .B1(n20083), .B2(n20082), .A(n20081), .ZN(n20095) );
  OR2_X1 U22973 ( .A1(n20085), .A2(n20084), .ZN(n20086) );
  AOI22_X1 U22974 ( .A1(n20095), .A2(n20087), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20086), .ZN(n20090) );
  NAND2_X1 U22975 ( .A1(n12840), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20089) );
  OAI211_X1 U22976 ( .C1(n20091), .C2(n20106), .A(n20090), .B(n20089), .ZN(
        P1_U2999) );
  AOI22_X1 U22977 ( .A1(n20095), .A2(n20094), .B1(n20093), .B2(n20092), .ZN(
        n20100) );
  OAI22_X1 U22978 ( .A1(n20098), .A2(n20097), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20096), .ZN(n20099) );
  OAI211_X1 U22979 ( .C1(n20847), .C2(n20101), .A(n20100), .B(n20099), .ZN(
        P1_U3031) );
  NOR2_X1 U22980 ( .A1(n20103), .A2(n20102), .ZN(P1_U3032) );
  AOI22_X1 U22981 ( .A1(DATAI_16_), .A2(n20147), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9571), .ZN(n20655) );
  INV_X1 U22982 ( .A(n20721), .ZN(n20652) );
  NAND2_X1 U22983 ( .A1(n20149), .A2(n20109), .ZN(n20709) );
  INV_X1 U22984 ( .A(n20709), .ZN(n20643) );
  NOR3_X1 U22985 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20167) );
  NAND2_X1 U22986 ( .A1(n20601), .A2(n20167), .ZN(n20113) );
  INV_X1 U22987 ( .A(n20113), .ZN(n20150) );
  AOI22_X1 U22988 ( .A1(n20770), .A2(n20652), .B1(n20643), .B2(n20150), .ZN(
        n20122) );
  AND2_X1 U22989 ( .A1(n20418), .A2(n20481), .ZN(n20272) );
  AND2_X1 U22990 ( .A1(n20117), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20639) );
  INV_X1 U22991 ( .A(n20770), .ZN(n20110) );
  NAND3_X1 U22992 ( .A1(n20110), .A2(n20716), .A3(n20183), .ZN(n20111) );
  NAND2_X1 U22993 ( .A1(n20111), .A2(n20162), .ZN(n20116) );
  OR2_X1 U22994 ( .A1(n20415), .A2(n20112), .ZN(n20230) );
  OR2_X1 U22995 ( .A1(n20230), .A2(n20646), .ZN(n20119) );
  AOI22_X1 U22996 ( .A1(n20116), .A2(n20119), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20113), .ZN(n20114) );
  OAI211_X1 U22997 ( .C1(n20272), .C2(n20856), .A(n20484), .B(n20114), .ZN(
        n20153) );
  NOR2_X2 U22998 ( .A1(n20115), .A2(n20279), .ZN(n20642) );
  INV_X1 U22999 ( .A(n20116), .ZN(n20120) );
  NOR2_X1 U23000 ( .A1(n20117), .A2(n20856), .ZN(n20421) );
  INV_X1 U23001 ( .A(n20421), .ZN(n20487) );
  INV_X1 U23002 ( .A(n20272), .ZN(n20118) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20153), .B1(
        n20642), .B2(n20152), .ZN(n20121) );
  OAI211_X1 U23004 ( .C1(n20655), .C2(n20183), .A(n20122), .B(n20121), .ZN(
        P1_U3033) );
  AOI22_X1 U23005 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9571), .B1(DATAI_25_), 
        .B2(n20147), .ZN(n20728) );
  INV_X1 U23006 ( .A(n20728), .ZN(n20658) );
  NAND2_X1 U23007 ( .A1(n20149), .A2(n11757), .ZN(n20723) );
  INV_X1 U23008 ( .A(n20723), .ZN(n20657) );
  AOI22_X1 U23009 ( .A1(n20770), .A2(n20658), .B1(n20657), .B2(n20150), .ZN(
        n20125) );
  NOR2_X2 U23010 ( .A1(n20123), .A2(n20279), .ZN(n20656) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20153), .B1(
        n20656), .B2(n20152), .ZN(n20124) );
  OAI211_X1 U23012 ( .C1(n20661), .C2(n20183), .A(n20125), .B(n20124), .ZN(
        P1_U3034) );
  AOI22_X1 U23013 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9571), .B1(DATAI_26_), 
        .B2(n20147), .ZN(n20735) );
  INV_X1 U23014 ( .A(n20735), .ZN(n20664) );
  NAND2_X1 U23015 ( .A1(n20149), .A2(n20126), .ZN(n20730) );
  INV_X1 U23016 ( .A(n20730), .ZN(n20663) );
  AOI22_X1 U23017 ( .A1(n20770), .A2(n20664), .B1(n20663), .B2(n20150), .ZN(
        n20129) );
  NOR2_X2 U23018 ( .A1(n20127), .A2(n20279), .ZN(n20662) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20153), .B1(
        n20662), .B2(n20152), .ZN(n20128) );
  OAI211_X1 U23020 ( .C1(n20667), .C2(n20183), .A(n20129), .B(n20128), .ZN(
        P1_U3035) );
  AOI22_X1 U23021 ( .A1(DATAI_19_), .A2(n20147), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9571), .ZN(n20673) );
  INV_X1 U23022 ( .A(n20742), .ZN(n20670) );
  NAND2_X1 U23023 ( .A1(n20149), .A2(n20130), .ZN(n20737) );
  INV_X1 U23024 ( .A(n20737), .ZN(n20669) );
  AOI22_X1 U23025 ( .A1(n20770), .A2(n20670), .B1(n20669), .B2(n20150), .ZN(
        n20133) );
  NOR2_X2 U23026 ( .A1(n20131), .A2(n20279), .ZN(n20668) );
  AOI22_X1 U23027 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20153), .B1(
        n20668), .B2(n20152), .ZN(n20132) );
  OAI211_X1 U23028 ( .C1(n20673), .C2(n20183), .A(n20133), .B(n20132), .ZN(
        P1_U3036) );
  AOI22_X1 U23029 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9571), .B1(DATAI_20_), 
        .B2(n20147), .ZN(n20679) );
  INV_X1 U23030 ( .A(n20749), .ZN(n20676) );
  NAND2_X1 U23031 ( .A1(n20149), .A2(n20134), .ZN(n20744) );
  INV_X1 U23032 ( .A(n20744), .ZN(n20675) );
  AOI22_X1 U23033 ( .A1(n20770), .A2(n20676), .B1(n20675), .B2(n20150), .ZN(
        n20137) );
  NOR2_X2 U23034 ( .A1(n20135), .A2(n20279), .ZN(n20674) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20153), .B1(
        n20674), .B2(n20152), .ZN(n20136) );
  OAI211_X1 U23036 ( .C1(n20679), .C2(n20183), .A(n20137), .B(n20136), .ZN(
        P1_U3037) );
  AOI22_X1 U23037 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9571), .B1(DATAI_29_), 
        .B2(n20147), .ZN(n20756) );
  INV_X1 U23038 ( .A(n20756), .ZN(n20682) );
  NAND2_X1 U23039 ( .A1(n20149), .A2(n20138), .ZN(n20751) );
  INV_X1 U23040 ( .A(n20751), .ZN(n20681) );
  AOI22_X1 U23041 ( .A1(n20770), .A2(n20682), .B1(n20681), .B2(n20150), .ZN(
        n20141) );
  NOR2_X2 U23042 ( .A1(n20139), .A2(n20279), .ZN(n20680) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20153), .B1(
        n20680), .B2(n20152), .ZN(n20140) );
  OAI211_X1 U23044 ( .C1(n20685), .C2(n20183), .A(n20141), .B(n20140), .ZN(
        P1_U3038) );
  AOI22_X1 U23045 ( .A1(DATAI_22_), .A2(n9570), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9571), .ZN(n20691) );
  INV_X1 U23046 ( .A(n20763), .ZN(n20688) );
  NAND2_X1 U23047 ( .A1(n20149), .A2(n20142), .ZN(n20758) );
  INV_X1 U23048 ( .A(n20758), .ZN(n20687) );
  AOI22_X1 U23049 ( .A1(n20770), .A2(n20688), .B1(n20687), .B2(n20150), .ZN(
        n20145) );
  NOR2_X2 U23050 ( .A1(n20143), .A2(n20279), .ZN(n20686) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20153), .B1(
        n20686), .B2(n20152), .ZN(n20144) );
  OAI211_X1 U23052 ( .C1(n20691), .C2(n20183), .A(n20145), .B(n20144), .ZN(
        P1_U3039) );
  AOI22_X1 U23053 ( .A1(DATAI_31_), .A2(n20147), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9571), .ZN(n20775) );
  INV_X1 U23054 ( .A(n20775), .ZN(n20696) );
  NAND2_X1 U23055 ( .A1(n20149), .A2(n20148), .ZN(n20767) );
  INV_X1 U23056 ( .A(n20767), .ZN(n20695) );
  AOI22_X1 U23057 ( .A1(n20770), .A2(n20696), .B1(n20695), .B2(n20150), .ZN(
        n20155) );
  NOR2_X2 U23058 ( .A1(n20151), .A2(n20279), .ZN(n20693) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20153), .B1(
        n20693), .B2(n20152), .ZN(n20154) );
  OAI211_X1 U23060 ( .C1(n20701), .C2(n20183), .A(n20155), .B(n20154), .ZN(
        P1_U3040) );
  INV_X1 U23061 ( .A(n20167), .ZN(n20156) );
  NOR2_X1 U23062 ( .A1(n20601), .A2(n20156), .ZN(n20185) );
  OR2_X1 U23063 ( .A1(n20230), .A2(n20157), .ZN(n20159) );
  INV_X1 U23064 ( .A(n20185), .ZN(n20158) );
  NAND2_X1 U23065 ( .A1(n20159), .A2(n20158), .ZN(n20163) );
  NAND2_X1 U23066 ( .A1(n20163), .A2(n20716), .ZN(n20161) );
  NAND2_X1 U23067 ( .A1(n20167), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20160) );
  NAND2_X1 U23068 ( .A1(n20161), .A2(n20160), .ZN(n20184) );
  AOI22_X1 U23069 ( .A1(n20643), .A2(n20185), .B1(n20642), .B2(n20184), .ZN(
        n20169) );
  NAND2_X1 U23070 ( .A1(n20227), .A2(n20377), .ZN(n20236) );
  INV_X1 U23071 ( .A(n20236), .ZN(n20165) );
  INV_X1 U23072 ( .A(n20162), .ZN(n20608) );
  INV_X1 U23073 ( .A(n20163), .ZN(n20164) );
  OAI21_X1 U23074 ( .B1(n20165), .B2(n20608), .A(n20164), .ZN(n20166) );
  OAI211_X1 U23075 ( .C1(n20377), .C2(n20167), .A(n20715), .B(n20166), .ZN(
        n20187) );
  INV_X1 U23076 ( .A(n20225), .ZN(n20180) );
  INV_X1 U23077 ( .A(n20655), .ZN(n20718) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20187), .B1(
        n20180), .B2(n20718), .ZN(n20168) );
  OAI211_X1 U23079 ( .C1(n20721), .C2(n20183), .A(n20169), .B(n20168), .ZN(
        P1_U3041) );
  AOI22_X1 U23080 ( .A1(n20657), .A2(n20185), .B1(n20656), .B2(n20184), .ZN(
        n20171) );
  INV_X1 U23081 ( .A(n20183), .ZN(n20186) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n20658), .ZN(n20170) );
  OAI211_X1 U23083 ( .C1(n20661), .C2(n20225), .A(n20171), .B(n20170), .ZN(
        P1_U3042) );
  AOI22_X1 U23084 ( .A1(n20663), .A2(n20185), .B1(n20662), .B2(n20184), .ZN(
        n20173) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n20664), .ZN(n20172) );
  OAI211_X1 U23086 ( .C1(n20667), .C2(n20225), .A(n20173), .B(n20172), .ZN(
        P1_U3043) );
  AOI22_X1 U23087 ( .A1(n20669), .A2(n20185), .B1(n20668), .B2(n20184), .ZN(
        n20175) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n20670), .ZN(n20174) );
  OAI211_X1 U23089 ( .C1(n20673), .C2(n20225), .A(n20175), .B(n20174), .ZN(
        P1_U3044) );
  AOI22_X1 U23090 ( .A1(n20675), .A2(n20185), .B1(n20674), .B2(n20184), .ZN(
        n20177) );
  INV_X1 U23091 ( .A(n20679), .ZN(n20746) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20187), .B1(
        n20180), .B2(n20746), .ZN(n20176) );
  OAI211_X1 U23093 ( .C1(n20749), .C2(n20183), .A(n20177), .B(n20176), .ZN(
        P1_U3045) );
  AOI22_X1 U23094 ( .A1(n20681), .A2(n20185), .B1(n20680), .B2(n20184), .ZN(
        n20179) );
  INV_X1 U23095 ( .A(n20685), .ZN(n20753) );
  AOI22_X1 U23096 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20187), .B1(
        n20180), .B2(n20753), .ZN(n20178) );
  OAI211_X1 U23097 ( .C1(n20756), .C2(n20183), .A(n20179), .B(n20178), .ZN(
        P1_U3046) );
  AOI22_X1 U23098 ( .A1(n20687), .A2(n20185), .B1(n20686), .B2(n20184), .ZN(
        n20182) );
  INV_X1 U23099 ( .A(n20691), .ZN(n20760) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20187), .B1(
        n20180), .B2(n20760), .ZN(n20181) );
  OAI211_X1 U23101 ( .C1(n20763), .C2(n20183), .A(n20182), .B(n20181), .ZN(
        P1_U3047) );
  AOI22_X1 U23102 ( .A1(n20695), .A2(n20185), .B1(n20693), .B2(n20184), .ZN(
        n20189) );
  AOI22_X1 U23103 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n20696), .ZN(n20188) );
  OAI211_X1 U23104 ( .C1(n20701), .C2(n20225), .A(n20189), .B(n20188), .ZN(
        P1_U3048) );
  INV_X1 U23105 ( .A(n20632), .ZN(n20190) );
  NAND3_X1 U23106 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20559), .A3(
        n20560), .ZN(n20239) );
  NOR2_X1 U23107 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20239), .ZN(
        n20193) );
  INV_X1 U23108 ( .A(n20193), .ZN(n20219) );
  OAI22_X1 U23109 ( .A1(n20263), .A2(n20655), .B1(n20709), .B2(n20219), .ZN(
        n20191) );
  INV_X1 U23110 ( .A(n20191), .ZN(n20200) );
  NAND2_X1 U23111 ( .A1(n20263), .A2(n20225), .ZN(n20192) );
  AOI21_X1 U23112 ( .B1(n20192), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20635), 
        .ZN(n20196) );
  OR2_X1 U23113 ( .A1(n20230), .A2(n14265), .ZN(n20197) );
  NOR2_X1 U23114 ( .A1(n20193), .A2(n20566), .ZN(n20194) );
  AOI21_X1 U23115 ( .B1(n20196), .B2(n20197), .A(n20194), .ZN(n20195) );
  OR2_X1 U23116 ( .A1(n20481), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20345) );
  NAND2_X1 U23117 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20345), .ZN(n20342) );
  NAND3_X1 U23118 ( .A1(n20484), .A2(n20195), .A3(n20342), .ZN(n20222) );
  INV_X1 U23119 ( .A(n20196), .ZN(n20198) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20222), .B1(
        n20642), .B2(n20221), .ZN(n20199) );
  OAI211_X1 U23121 ( .C1(n20721), .C2(n20225), .A(n20200), .B(n20199), .ZN(
        P1_U3049) );
  OAI22_X1 U23122 ( .A1(n20263), .A2(n20661), .B1(n20219), .B2(n20723), .ZN(
        n20201) );
  INV_X1 U23123 ( .A(n20201), .ZN(n20203) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20222), .B1(
        n20656), .B2(n20221), .ZN(n20202) );
  OAI211_X1 U23125 ( .C1(n20728), .C2(n20225), .A(n20203), .B(n20202), .ZN(
        P1_U3050) );
  OAI22_X1 U23126 ( .A1(n20263), .A2(n20667), .B1(n20219), .B2(n20730), .ZN(
        n20204) );
  INV_X1 U23127 ( .A(n20204), .ZN(n20206) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20222), .B1(
        n20662), .B2(n20221), .ZN(n20205) );
  OAI211_X1 U23129 ( .C1(n20735), .C2(n20225), .A(n20206), .B(n20205), .ZN(
        P1_U3051) );
  OAI22_X1 U23130 ( .A1(n20225), .A2(n20742), .B1(n20219), .B2(n20737), .ZN(
        n20207) );
  INV_X1 U23131 ( .A(n20207), .ZN(n20209) );
  AOI22_X1 U23132 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20222), .B1(
        n20668), .B2(n20221), .ZN(n20208) );
  OAI211_X1 U23133 ( .C1(n20673), .C2(n20263), .A(n20209), .B(n20208), .ZN(
        P1_U3052) );
  OAI22_X1 U23134 ( .A1(n20263), .A2(n20679), .B1(n20219), .B2(n20744), .ZN(
        n20210) );
  INV_X1 U23135 ( .A(n20210), .ZN(n20212) );
  AOI22_X1 U23136 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20222), .B1(
        n20674), .B2(n20221), .ZN(n20211) );
  OAI211_X1 U23137 ( .C1(n20749), .C2(n20225), .A(n20212), .B(n20211), .ZN(
        P1_U3053) );
  OAI22_X1 U23138 ( .A1(n20263), .A2(n20685), .B1(n20219), .B2(n20751), .ZN(
        n20213) );
  INV_X1 U23139 ( .A(n20213), .ZN(n20215) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20222), .B1(
        n20680), .B2(n20221), .ZN(n20214) );
  OAI211_X1 U23141 ( .C1(n20756), .C2(n20225), .A(n20215), .B(n20214), .ZN(
        P1_U3054) );
  OAI22_X1 U23142 ( .A1(n20263), .A2(n20691), .B1(n20219), .B2(n20758), .ZN(
        n20216) );
  INV_X1 U23143 ( .A(n20216), .ZN(n20218) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20222), .B1(
        n20686), .B2(n20221), .ZN(n20217) );
  OAI211_X1 U23145 ( .C1(n20763), .C2(n20225), .A(n20218), .B(n20217), .ZN(
        P1_U3055) );
  OAI22_X1 U23146 ( .A1(n20263), .A2(n20701), .B1(n20219), .B2(n20767), .ZN(
        n20220) );
  INV_X1 U23147 ( .A(n20220), .ZN(n20224) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20222), .B1(
        n20693), .B2(n20221), .ZN(n20223) );
  OAI211_X1 U23149 ( .C1(n20775), .C2(n20225), .A(n20224), .B(n20223), .ZN(
        P1_U3056) );
  INV_X1 U23150 ( .A(n20527), .ZN(n20226) );
  INV_X1 U23151 ( .A(n20228), .ZN(n20517) );
  NAND2_X1 U23152 ( .A1(n20517), .A2(n20559), .ZN(n20262) );
  OAI22_X1 U23153 ( .A1(n20263), .A2(n20721), .B1(n20709), .B2(n20262), .ZN(
        n20229) );
  INV_X1 U23154 ( .A(n20229), .ZN(n20243) );
  INV_X1 U23155 ( .A(n20230), .ZN(n20234) );
  NAND2_X1 U23156 ( .A1(n11916), .A2(n20231), .ZN(n20702) );
  INV_X1 U23157 ( .A(n20702), .ZN(n20233) );
  INV_X1 U23158 ( .A(n20262), .ZN(n20232) );
  AOI21_X1 U23159 ( .B1(n20234), .B2(n20233), .A(n20232), .ZN(n20241) );
  INV_X1 U23160 ( .A(n20713), .ZN(n20235) );
  INV_X1 U23161 ( .A(n20240), .ZN(n20237) );
  AOI22_X1 U23162 ( .A1(n20241), .A2(n20237), .B1(n20635), .B2(n20239), .ZN(
        n20238) );
  NAND2_X1 U23163 ( .A1(n20715), .A2(n20238), .ZN(n20266) );
  OAI22_X1 U23164 ( .A1(n20241), .A2(n20240), .B1(n20856), .B2(n20239), .ZN(
        n20265) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20266), .B1(
        n20642), .B2(n20265), .ZN(n20242) );
  OAI211_X1 U23166 ( .C1(n20655), .C2(n20276), .A(n20243), .B(n20242), .ZN(
        P1_U3057) );
  OAI22_X1 U23167 ( .A1(n20263), .A2(n20728), .B1(n20723), .B2(n20262), .ZN(
        n20244) );
  INV_X1 U23168 ( .A(n20244), .ZN(n20246) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20266), .B1(
        n20656), .B2(n20265), .ZN(n20245) );
  OAI211_X1 U23170 ( .C1(n20661), .C2(n20276), .A(n20246), .B(n20245), .ZN(
        P1_U3058) );
  OAI22_X1 U23171 ( .A1(n20276), .A2(n20667), .B1(n20730), .B2(n20262), .ZN(
        n20247) );
  INV_X1 U23172 ( .A(n20247), .ZN(n20249) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20266), .B1(
        n20662), .B2(n20265), .ZN(n20248) );
  OAI211_X1 U23174 ( .C1(n20735), .C2(n20263), .A(n20249), .B(n20248), .ZN(
        P1_U3059) );
  OAI22_X1 U23175 ( .A1(n20263), .A2(n20742), .B1(n20262), .B2(n20737), .ZN(
        n20250) );
  INV_X1 U23176 ( .A(n20250), .ZN(n20252) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20266), .B1(
        n20668), .B2(n20265), .ZN(n20251) );
  OAI211_X1 U23178 ( .C1(n20673), .C2(n20276), .A(n20252), .B(n20251), .ZN(
        P1_U3060) );
  OAI22_X1 U23179 ( .A1(n20276), .A2(n20679), .B1(n20744), .B2(n20262), .ZN(
        n20253) );
  INV_X1 U23180 ( .A(n20253), .ZN(n20255) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20266), .B1(
        n20674), .B2(n20265), .ZN(n20254) );
  OAI211_X1 U23182 ( .C1(n20749), .C2(n20263), .A(n20255), .B(n20254), .ZN(
        P1_U3061) );
  OAI22_X1 U23183 ( .A1(n20263), .A2(n20756), .B1(n20751), .B2(n20262), .ZN(
        n20256) );
  INV_X1 U23184 ( .A(n20256), .ZN(n20258) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20266), .B1(
        n20680), .B2(n20265), .ZN(n20257) );
  OAI211_X1 U23186 ( .C1(n20685), .C2(n20276), .A(n20258), .B(n20257), .ZN(
        P1_U3062) );
  OAI22_X1 U23187 ( .A1(n20263), .A2(n20763), .B1(n20758), .B2(n20262), .ZN(
        n20259) );
  INV_X1 U23188 ( .A(n20259), .ZN(n20261) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20266), .B1(
        n20686), .B2(n20265), .ZN(n20260) );
  OAI211_X1 U23190 ( .C1(n20691), .C2(n20276), .A(n20261), .B(n20260), .ZN(
        P1_U3063) );
  OAI22_X1 U23191 ( .A1(n20263), .A2(n20775), .B1(n20767), .B2(n20262), .ZN(
        n20264) );
  INV_X1 U23192 ( .A(n20264), .ZN(n20268) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20266), .B1(
        n20693), .B2(n20265), .ZN(n20267) );
  OAI211_X1 U23194 ( .C1(n20701), .C2(n20276), .A(n20268), .B(n20267), .ZN(
        P1_U3064) );
  NOR3_X1 U23195 ( .A1(n20560), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20317) );
  INV_X1 U23196 ( .A(n20317), .ZN(n20309) );
  NOR2_X1 U23197 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20309), .ZN(
        n20281) );
  INV_X1 U23198 ( .A(n20281), .ZN(n20303) );
  OR2_X1 U23199 ( .A1(n20564), .A2(n20270), .ZN(n20375) );
  NAND2_X1 U23200 ( .A1(n14265), .A2(n20716), .ZN(n20271) );
  OR2_X1 U23201 ( .A1(n20375), .A2(n20271), .ZN(n20274) );
  NAND2_X1 U23202 ( .A1(n20639), .A2(n20272), .ZN(n20273) );
  INV_X1 U23203 ( .A(n20642), .ZN(n20708) );
  OAI22_X1 U23204 ( .A1(n20709), .A2(n20303), .B1(n20302), .B2(n20708), .ZN(
        n20275) );
  INV_X1 U23205 ( .A(n20275), .ZN(n20283) );
  INV_X1 U23206 ( .A(n20339), .ZN(n20277) );
  OAI21_X1 U23207 ( .B1(n20305), .B2(n20277), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20278) );
  OAI21_X1 U23208 ( .B1(n20646), .B2(n20375), .A(n20278), .ZN(n20280) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20652), .ZN(n20282) );
  OAI211_X1 U23210 ( .C1(n20655), .C2(n20339), .A(n20283), .B(n20282), .ZN(
        P1_U3065) );
  INV_X1 U23211 ( .A(n20656), .ZN(n20722) );
  OAI22_X1 U23212 ( .A1(n20723), .A2(n20303), .B1(n20302), .B2(n20722), .ZN(
        n20284) );
  INV_X1 U23213 ( .A(n20284), .ZN(n20286) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20658), .ZN(n20285) );
  OAI211_X1 U23215 ( .C1(n20661), .C2(n20339), .A(n20286), .B(n20285), .ZN(
        P1_U3066) );
  INV_X1 U23216 ( .A(n20662), .ZN(n20729) );
  OAI22_X1 U23217 ( .A1(n20730), .A2(n20303), .B1(n20302), .B2(n20729), .ZN(
        n20287) );
  INV_X1 U23218 ( .A(n20287), .ZN(n20289) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20664), .ZN(n20288) );
  OAI211_X1 U23220 ( .C1(n20667), .C2(n20339), .A(n20289), .B(n20288), .ZN(
        P1_U3067) );
  INV_X1 U23221 ( .A(n20668), .ZN(n20736) );
  OAI22_X1 U23222 ( .A1(n20737), .A2(n20303), .B1(n20302), .B2(n20736), .ZN(
        n20290) );
  INV_X1 U23223 ( .A(n20290), .ZN(n20292) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20670), .ZN(n20291) );
  OAI211_X1 U23225 ( .C1(n20673), .C2(n20339), .A(n20292), .B(n20291), .ZN(
        P1_U3068) );
  INV_X1 U23226 ( .A(n20674), .ZN(n20743) );
  OAI22_X1 U23227 ( .A1(n20744), .A2(n20303), .B1(n20302), .B2(n20743), .ZN(
        n20293) );
  INV_X1 U23228 ( .A(n20293), .ZN(n20295) );
  AOI22_X1 U23229 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20676), .ZN(n20294) );
  OAI211_X1 U23230 ( .C1(n20679), .C2(n20339), .A(n20295), .B(n20294), .ZN(
        P1_U3069) );
  INV_X1 U23231 ( .A(n20680), .ZN(n20750) );
  OAI22_X1 U23232 ( .A1(n20751), .A2(n20303), .B1(n20302), .B2(n20750), .ZN(
        n20296) );
  INV_X1 U23233 ( .A(n20296), .ZN(n20298) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20682), .ZN(n20297) );
  OAI211_X1 U23235 ( .C1(n20685), .C2(n20339), .A(n20298), .B(n20297), .ZN(
        P1_U3070) );
  INV_X1 U23236 ( .A(n20686), .ZN(n20757) );
  OAI22_X1 U23237 ( .A1(n20758), .A2(n20303), .B1(n20302), .B2(n20757), .ZN(
        n20299) );
  INV_X1 U23238 ( .A(n20299), .ZN(n20301) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20688), .ZN(n20300) );
  OAI211_X1 U23240 ( .C1(n20691), .C2(n20339), .A(n20301), .B(n20300), .ZN(
        P1_U3071) );
  INV_X1 U23241 ( .A(n20693), .ZN(n20764) );
  OAI22_X1 U23242 ( .A1(n20767), .A2(n20303), .B1(n20302), .B2(n20764), .ZN(
        n20304) );
  INV_X1 U23243 ( .A(n20304), .ZN(n20308) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20306), .B1(
        n20305), .B2(n20696), .ZN(n20307) );
  OAI211_X1 U23245 ( .C1(n20701), .C2(n20339), .A(n20308), .B(n20307), .ZN(
        P1_U3072) );
  NOR2_X1 U23246 ( .A1(n20601), .A2(n20309), .ZN(n20334) );
  OR2_X1 U23247 ( .A1(n20375), .A2(n20157), .ZN(n20311) );
  INV_X1 U23248 ( .A(n20334), .ZN(n20310) );
  NAND2_X1 U23249 ( .A1(n20311), .A2(n20310), .ZN(n20314) );
  NAND2_X1 U23250 ( .A1(n20314), .A2(n20716), .ZN(n20313) );
  NAND2_X1 U23251 ( .A1(n20317), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20312) );
  NAND2_X1 U23252 ( .A1(n20313), .A2(n20312), .ZN(n20333) );
  AOI22_X1 U23253 ( .A1(n20643), .A2(n20334), .B1(n20642), .B2(n20333), .ZN(
        n20320) );
  NOR2_X1 U23254 ( .A1(n20385), .A2(n20635), .ZN(n20383) );
  INV_X1 U23255 ( .A(n20314), .ZN(n20315) );
  OAI21_X1 U23256 ( .B1(n20383), .B2(n20608), .A(n20315), .ZN(n20316) );
  OAI211_X1 U23257 ( .C1(n20377), .C2(n20317), .A(n20715), .B(n20316), .ZN(
        n20336) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20718), .ZN(n20319) );
  OAI211_X1 U23259 ( .C1(n20721), .C2(n20339), .A(n20320), .B(n20319), .ZN(
        P1_U3073) );
  AOI22_X1 U23260 ( .A1(n20657), .A2(n20334), .B1(n20656), .B2(n20333), .ZN(
        n20322) );
  INV_X1 U23261 ( .A(n20661), .ZN(n20725) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20725), .ZN(n20321) );
  OAI211_X1 U23263 ( .C1(n20728), .C2(n20339), .A(n20322), .B(n20321), .ZN(
        P1_U3074) );
  AOI22_X1 U23264 ( .A1(n20663), .A2(n20334), .B1(n20662), .B2(n20333), .ZN(
        n20324) );
  INV_X1 U23265 ( .A(n20667), .ZN(n20732) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20732), .ZN(n20323) );
  OAI211_X1 U23267 ( .C1(n20735), .C2(n20339), .A(n20324), .B(n20323), .ZN(
        P1_U3075) );
  AOI22_X1 U23268 ( .A1(n20669), .A2(n20334), .B1(n20668), .B2(n20333), .ZN(
        n20326) );
  INV_X1 U23269 ( .A(n20673), .ZN(n20739) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20739), .ZN(n20325) );
  OAI211_X1 U23271 ( .C1(n20742), .C2(n20339), .A(n20326), .B(n20325), .ZN(
        P1_U3076) );
  AOI22_X1 U23272 ( .A1(n20675), .A2(n20334), .B1(n20674), .B2(n20333), .ZN(
        n20328) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20746), .ZN(n20327) );
  OAI211_X1 U23274 ( .C1(n20749), .C2(n20339), .A(n20328), .B(n20327), .ZN(
        P1_U3077) );
  AOI22_X1 U23275 ( .A1(n20681), .A2(n20334), .B1(n20680), .B2(n20333), .ZN(
        n20330) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20753), .ZN(n20329) );
  OAI211_X1 U23277 ( .C1(n20756), .C2(n20339), .A(n20330), .B(n20329), .ZN(
        P1_U3078) );
  AOI22_X1 U23278 ( .A1(n20687), .A2(n20334), .B1(n20686), .B2(n20333), .ZN(
        n20332) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20760), .ZN(n20331) );
  OAI211_X1 U23280 ( .C1(n20763), .C2(n20339), .A(n20332), .B(n20331), .ZN(
        P1_U3079) );
  AOI22_X1 U23281 ( .A1(n20695), .A2(n20334), .B1(n20693), .B2(n20333), .ZN(
        n20338) );
  INV_X1 U23282 ( .A(n20701), .ZN(n20769) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20769), .ZN(n20337) );
  OAI211_X1 U23284 ( .C1(n20775), .C2(n20339), .A(n20338), .B(n20337), .ZN(
        P1_U3080) );
  NAND2_X1 U23285 ( .A1(n20601), .A2(n10079), .ZN(n20368) );
  OAI22_X1 U23286 ( .A1(n20406), .A2(n20655), .B1(n20709), .B2(n20368), .ZN(
        n20340) );
  INV_X1 U23287 ( .A(n20340), .ZN(n20349) );
  AOI21_X1 U23288 ( .B1(n20406), .B2(n20369), .A(n20857), .ZN(n20341) );
  NOR2_X1 U23289 ( .A1(n20341), .A2(n20635), .ZN(n20344) );
  OR2_X1 U23290 ( .A1(n20375), .A2(n14265), .ZN(n20346) );
  AOI22_X1 U23291 ( .A1(n20344), .A2(n20346), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20368), .ZN(n20343) );
  NAND3_X1 U23292 ( .A1(n20650), .A2(n20343), .A3(n20342), .ZN(n20372) );
  INV_X1 U23293 ( .A(n20344), .ZN(n20347) );
  INV_X1 U23294 ( .A(n20639), .ZN(n20570) );
  OAI22_X1 U23295 ( .A1(n20347), .A2(n20346), .B1(n20345), .B2(n20570), .ZN(
        n20371) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20372), .B1(
        n20642), .B2(n20371), .ZN(n20348) );
  OAI211_X1 U23297 ( .C1(n20721), .C2(n20369), .A(n20349), .B(n20348), .ZN(
        P1_U3081) );
  OAI22_X1 U23298 ( .A1(n20369), .A2(n20728), .B1(n20723), .B2(n20368), .ZN(
        n20350) );
  INV_X1 U23299 ( .A(n20350), .ZN(n20352) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20372), .B1(
        n20656), .B2(n20371), .ZN(n20351) );
  OAI211_X1 U23301 ( .C1(n20661), .C2(n20406), .A(n20352), .B(n20351), .ZN(
        P1_U3082) );
  OAI22_X1 U23302 ( .A1(n20369), .A2(n20735), .B1(n20730), .B2(n20368), .ZN(
        n20353) );
  INV_X1 U23303 ( .A(n20353), .ZN(n20355) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20372), .B1(
        n20662), .B2(n20371), .ZN(n20354) );
  OAI211_X1 U23305 ( .C1(n20667), .C2(n20406), .A(n20355), .B(n20354), .ZN(
        P1_U3083) );
  OAI22_X1 U23306 ( .A1(n20406), .A2(n20673), .B1(n20737), .B2(n20368), .ZN(
        n20356) );
  INV_X1 U23307 ( .A(n20356), .ZN(n20358) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20372), .B1(
        n20668), .B2(n20371), .ZN(n20357) );
  OAI211_X1 U23309 ( .C1(n20742), .C2(n20369), .A(n20358), .B(n20357), .ZN(
        P1_U3084) );
  OAI22_X1 U23310 ( .A1(n20406), .A2(n20679), .B1(n20744), .B2(n20368), .ZN(
        n20359) );
  INV_X1 U23311 ( .A(n20359), .ZN(n20361) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20372), .B1(
        n20674), .B2(n20371), .ZN(n20360) );
  OAI211_X1 U23313 ( .C1(n20749), .C2(n20369), .A(n20361), .B(n20360), .ZN(
        P1_U3085) );
  OAI22_X1 U23314 ( .A1(n20369), .A2(n20756), .B1(n20751), .B2(n20368), .ZN(
        n20362) );
  INV_X1 U23315 ( .A(n20362), .ZN(n20364) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20372), .B1(
        n20680), .B2(n20371), .ZN(n20363) );
  OAI211_X1 U23317 ( .C1(n20685), .C2(n20406), .A(n20364), .B(n20363), .ZN(
        P1_U3086) );
  OAI22_X1 U23318 ( .A1(n20406), .A2(n20691), .B1(n20758), .B2(n20368), .ZN(
        n20365) );
  INV_X1 U23319 ( .A(n20365), .ZN(n20367) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20372), .B1(
        n20686), .B2(n20371), .ZN(n20366) );
  OAI211_X1 U23321 ( .C1(n20763), .C2(n20369), .A(n20367), .B(n20366), .ZN(
        P1_U3087) );
  OAI22_X1 U23322 ( .A1(n20369), .A2(n20775), .B1(n20767), .B2(n20368), .ZN(
        n20370) );
  INV_X1 U23323 ( .A(n20370), .ZN(n20374) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20372), .B1(
        n20693), .B2(n20371), .ZN(n20373) );
  OAI211_X1 U23325 ( .C1(n20701), .C2(n20406), .A(n20374), .B(n20373), .ZN(
        P1_U3088) );
  OR2_X1 U23326 ( .A1(n20375), .A2(n20702), .ZN(n20376) );
  INV_X1 U23327 ( .A(n20382), .ZN(n20378) );
  NAND2_X1 U23328 ( .A1(n20378), .A2(n20377), .ZN(n20380) );
  NAND2_X1 U23329 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n10079), .ZN(n20379) );
  OAI22_X1 U23330 ( .A1(n20709), .A2(n20408), .B1(n20407), .B2(n20708), .ZN(
        n20381) );
  INV_X1 U23331 ( .A(n20381), .ZN(n20387) );
  OAI21_X1 U23332 ( .B1(n20713), .B2(n20383), .A(n20382), .ZN(n20384) );
  OAI211_X1 U23333 ( .C1(n10079), .C2(n20716), .A(n20715), .B(n20384), .ZN(
        n20411) );
  NAND2_X1 U23334 ( .A1(n20385), .A2(n20527), .ZN(n20414) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20411), .B1(
        n20444), .B2(n20718), .ZN(n20386) );
  OAI211_X1 U23336 ( .C1(n20721), .C2(n20406), .A(n20387), .B(n20386), .ZN(
        P1_U3089) );
  OAI22_X1 U23337 ( .A1(n20723), .A2(n20408), .B1(n20407), .B2(n20722), .ZN(
        n20388) );
  INV_X1 U23338 ( .A(n20388), .ZN(n20390) );
  INV_X1 U23339 ( .A(n20406), .ZN(n20410) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20658), .ZN(n20389) );
  OAI211_X1 U23341 ( .C1(n20661), .C2(n20414), .A(n20390), .B(n20389), .ZN(
        P1_U3090) );
  OAI22_X1 U23342 ( .A1(n20730), .A2(n20408), .B1(n20407), .B2(n20729), .ZN(
        n20391) );
  INV_X1 U23343 ( .A(n20391), .ZN(n20393) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20664), .ZN(n20392) );
  OAI211_X1 U23345 ( .C1(n20667), .C2(n20414), .A(n20393), .B(n20392), .ZN(
        P1_U3091) );
  OAI22_X1 U23346 ( .A1(n20737), .A2(n20408), .B1(n20407), .B2(n20736), .ZN(
        n20394) );
  INV_X1 U23347 ( .A(n20394), .ZN(n20396) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20411), .B1(
        n20444), .B2(n20739), .ZN(n20395) );
  OAI211_X1 U23349 ( .C1(n20742), .C2(n20406), .A(n20396), .B(n20395), .ZN(
        P1_U3092) );
  OAI22_X1 U23350 ( .A1(n20744), .A2(n20408), .B1(n20407), .B2(n20743), .ZN(
        n20397) );
  INV_X1 U23351 ( .A(n20397), .ZN(n20399) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20676), .ZN(n20398) );
  OAI211_X1 U23353 ( .C1(n20679), .C2(n20414), .A(n20399), .B(n20398), .ZN(
        P1_U3093) );
  OAI22_X1 U23354 ( .A1(n20751), .A2(n20408), .B1(n20407), .B2(n20750), .ZN(
        n20400) );
  INV_X1 U23355 ( .A(n20400), .ZN(n20402) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20682), .ZN(n20401) );
  OAI211_X1 U23357 ( .C1(n20685), .C2(n20414), .A(n20402), .B(n20401), .ZN(
        P1_U3094) );
  OAI22_X1 U23358 ( .A1(n20758), .A2(n20408), .B1(n20407), .B2(n20757), .ZN(
        n20403) );
  INV_X1 U23359 ( .A(n20403), .ZN(n20405) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20411), .B1(
        n20444), .B2(n20760), .ZN(n20404) );
  OAI211_X1 U23361 ( .C1(n20763), .C2(n20406), .A(n20405), .B(n20404), .ZN(
        P1_U3095) );
  OAI22_X1 U23362 ( .A1(n20767), .A2(n20408), .B1(n20407), .B2(n20764), .ZN(
        n20409) );
  INV_X1 U23363 ( .A(n20409), .ZN(n20413) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20696), .ZN(n20412) );
  OAI211_X1 U23365 ( .C1(n20701), .C2(n20414), .A(n20413), .B(n20412), .ZN(
        P1_U3096) );
  NOR3_X1 U23366 ( .A1(n20559), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20455) );
  INV_X1 U23367 ( .A(n20455), .ZN(n20448) );
  NOR2_X1 U23368 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20448), .ZN(
        n20443) );
  NAND2_X1 U23369 ( .A1(n20415), .A2(n20564), .ZN(n20518) );
  OR2_X1 U23370 ( .A1(n20518), .A2(n20646), .ZN(n20417) );
  INV_X1 U23371 ( .A(n20443), .ZN(n20416) );
  AND2_X1 U23372 ( .A1(n20417), .A2(n20416), .ZN(n20425) );
  OR2_X1 U23373 ( .A1(n20425), .A2(n20635), .ZN(n20423) );
  INV_X1 U23374 ( .A(n20418), .ZN(n20419) );
  NAND2_X1 U23375 ( .A1(n20419), .A2(n20481), .ZN(n20569) );
  INV_X1 U23376 ( .A(n20569), .ZN(n20420) );
  NAND2_X1 U23377 ( .A1(n20421), .A2(n20420), .ZN(n20422) );
  NAND2_X1 U23378 ( .A1(n20423), .A2(n20422), .ZN(n20442) );
  AOI22_X1 U23379 ( .A1(n20643), .A2(n20443), .B1(n20642), .B2(n20442), .ZN(
        n20429) );
  INV_X1 U23380 ( .A(n20475), .ZN(n20424) );
  OAI21_X1 U23381 ( .B1(n20424), .B2(n20444), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20426) );
  NAND2_X1 U23382 ( .A1(n20426), .A2(n20425), .ZN(n20427) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20652), .ZN(n20428) );
  OAI211_X1 U23384 ( .C1(n20655), .C2(n20475), .A(n20429), .B(n20428), .ZN(
        P1_U3097) );
  AOI22_X1 U23385 ( .A1(n20657), .A2(n20443), .B1(n20656), .B2(n20442), .ZN(
        n20431) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20658), .ZN(n20430) );
  OAI211_X1 U23387 ( .C1(n20661), .C2(n20475), .A(n20431), .B(n20430), .ZN(
        P1_U3098) );
  AOI22_X1 U23388 ( .A1(n20663), .A2(n20443), .B1(n20662), .B2(n20442), .ZN(
        n20433) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20664), .ZN(n20432) );
  OAI211_X1 U23390 ( .C1(n20667), .C2(n20475), .A(n20433), .B(n20432), .ZN(
        P1_U3099) );
  AOI22_X1 U23391 ( .A1(n20669), .A2(n20443), .B1(n20668), .B2(n20442), .ZN(
        n20435) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20670), .ZN(n20434) );
  OAI211_X1 U23393 ( .C1(n20673), .C2(n20475), .A(n20435), .B(n20434), .ZN(
        P1_U3100) );
  AOI22_X1 U23394 ( .A1(n20675), .A2(n20443), .B1(n20674), .B2(n20442), .ZN(
        n20437) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20676), .ZN(n20436) );
  OAI211_X1 U23396 ( .C1(n20679), .C2(n20475), .A(n20437), .B(n20436), .ZN(
        P1_U3101) );
  AOI22_X1 U23397 ( .A1(n20681), .A2(n20443), .B1(n20680), .B2(n20442), .ZN(
        n20439) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20682), .ZN(n20438) );
  OAI211_X1 U23399 ( .C1(n20685), .C2(n20475), .A(n20439), .B(n20438), .ZN(
        P1_U3102) );
  AOI22_X1 U23400 ( .A1(n20687), .A2(n20443), .B1(n20686), .B2(n20442), .ZN(
        n20441) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20688), .ZN(n20440) );
  OAI211_X1 U23402 ( .C1(n20691), .C2(n20475), .A(n20441), .B(n20440), .ZN(
        P1_U3103) );
  AOI22_X1 U23403 ( .A1(n20695), .A2(n20443), .B1(n20693), .B2(n20442), .ZN(
        n20447) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20445), .B1(
        n20444), .B2(n20696), .ZN(n20446) );
  OAI211_X1 U23405 ( .C1(n20701), .C2(n20475), .A(n20447), .B(n20446), .ZN(
        P1_U3104) );
  NOR2_X1 U23406 ( .A1(n20601), .A2(n20448), .ZN(n20471) );
  OR2_X1 U23407 ( .A1(n20518), .A2(n20157), .ZN(n20450) );
  INV_X1 U23408 ( .A(n20471), .ZN(n20449) );
  AND2_X1 U23409 ( .A1(n20450), .A2(n20449), .ZN(n20453) );
  OR2_X1 U23410 ( .A1(n20453), .A2(n20635), .ZN(n20452) );
  NAND2_X1 U23411 ( .A1(n20455), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20451) );
  NAND2_X1 U23412 ( .A1(n20452), .A2(n20451), .ZN(n20470) );
  AOI22_X1 U23413 ( .A1(n20643), .A2(n20471), .B1(n20642), .B2(n20470), .ZN(
        n20457) );
  NOR2_X1 U23414 ( .A1(n20528), .A2(n20635), .ZN(n20524) );
  OAI21_X1 U23415 ( .B1(n20524), .B2(n20608), .A(n20453), .ZN(n20454) );
  OAI211_X1 U23416 ( .C1(n20716), .C2(n20455), .A(n20715), .B(n20454), .ZN(
        n20472) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20718), .ZN(n20456) );
  OAI211_X1 U23418 ( .C1(n20721), .C2(n20475), .A(n20457), .B(n20456), .ZN(
        P1_U3105) );
  AOI22_X1 U23419 ( .A1(n20657), .A2(n20471), .B1(n20656), .B2(n20470), .ZN(
        n20459) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20725), .ZN(n20458) );
  OAI211_X1 U23421 ( .C1(n20728), .C2(n20475), .A(n20459), .B(n20458), .ZN(
        P1_U3106) );
  AOI22_X1 U23422 ( .A1(n20663), .A2(n20471), .B1(n20662), .B2(n20470), .ZN(
        n20461) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20732), .ZN(n20460) );
  OAI211_X1 U23424 ( .C1(n20735), .C2(n20475), .A(n20461), .B(n20460), .ZN(
        P1_U3107) );
  AOI22_X1 U23425 ( .A1(n20669), .A2(n20471), .B1(n20668), .B2(n20470), .ZN(
        n20463) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20739), .ZN(n20462) );
  OAI211_X1 U23427 ( .C1(n20742), .C2(n20475), .A(n20463), .B(n20462), .ZN(
        P1_U3108) );
  AOI22_X1 U23428 ( .A1(n20675), .A2(n20471), .B1(n20674), .B2(n20470), .ZN(
        n20465) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20746), .ZN(n20464) );
  OAI211_X1 U23430 ( .C1(n20749), .C2(n20475), .A(n20465), .B(n20464), .ZN(
        P1_U3109) );
  AOI22_X1 U23431 ( .A1(n20681), .A2(n20471), .B1(n20680), .B2(n20470), .ZN(
        n20467) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20753), .ZN(n20466) );
  OAI211_X1 U23433 ( .C1(n20756), .C2(n20475), .A(n20467), .B(n20466), .ZN(
        P1_U3110) );
  AOI22_X1 U23434 ( .A1(n20687), .A2(n20471), .B1(n20686), .B2(n20470), .ZN(
        n20469) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20760), .ZN(n20468) );
  OAI211_X1 U23436 ( .C1(n20763), .C2(n20475), .A(n20469), .B(n20468), .ZN(
        P1_U3111) );
  AOI22_X1 U23437 ( .A1(n20695), .A2(n20471), .B1(n20693), .B2(n20470), .ZN(
        n20474) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20472), .B1(
        n20479), .B2(n20769), .ZN(n20473) );
  OAI211_X1 U23439 ( .C1(n20775), .C2(n20475), .A(n20474), .B(n20473), .ZN(
        P1_U3112) );
  NOR3_X1 U23440 ( .A1(n20559), .A2(n20476), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20526) );
  INV_X1 U23441 ( .A(n20526), .ZN(n20477) );
  NOR2_X1 U23442 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20477), .ZN(
        n20482) );
  INV_X1 U23443 ( .A(n20482), .ZN(n20510) );
  OAI22_X1 U23444 ( .A1(n20511), .A2(n20721), .B1(n20709), .B2(n20510), .ZN(
        n20478) );
  INV_X1 U23445 ( .A(n20478), .ZN(n20491) );
  OAI21_X1 U23446 ( .B1(n20544), .B2(n20479), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20480) );
  NAND2_X1 U23447 ( .A1(n20480), .A2(n20377), .ZN(n20489) );
  NOR2_X1 U23448 ( .A1(n20518), .A2(n14265), .ZN(n20486) );
  OR2_X1 U23449 ( .A1(n20481), .A2(n20559), .ZN(n20637) );
  NAND2_X1 U23450 ( .A1(n20637), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20649) );
  OAI21_X1 U23451 ( .B1(n20566), .B2(n20482), .A(n20649), .ZN(n20483) );
  INV_X1 U23452 ( .A(n20483), .ZN(n20485) );
  OAI211_X1 U23453 ( .C1(n20489), .C2(n20486), .A(n20485), .B(n20484), .ZN(
        n20514) );
  INV_X1 U23454 ( .A(n20486), .ZN(n20488) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20514), .B1(
        n20642), .B2(n20513), .ZN(n20490) );
  OAI211_X1 U23456 ( .C1(n20655), .C2(n20557), .A(n20491), .B(n20490), .ZN(
        P1_U3113) );
  OAI22_X1 U23457 ( .A1(n20511), .A2(n20728), .B1(n20723), .B2(n20510), .ZN(
        n20492) );
  INV_X1 U23458 ( .A(n20492), .ZN(n20494) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20514), .B1(
        n20656), .B2(n20513), .ZN(n20493) );
  OAI211_X1 U23460 ( .C1(n20661), .C2(n20557), .A(n20494), .B(n20493), .ZN(
        P1_U3114) );
  OAI22_X1 U23461 ( .A1(n20557), .A2(n20667), .B1(n20730), .B2(n20510), .ZN(
        n20495) );
  INV_X1 U23462 ( .A(n20495), .ZN(n20497) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20514), .B1(
        n20662), .B2(n20513), .ZN(n20496) );
  OAI211_X1 U23464 ( .C1(n20735), .C2(n20511), .A(n20497), .B(n20496), .ZN(
        P1_U3115) );
  OAI22_X1 U23465 ( .A1(n20511), .A2(n20742), .B1(n20737), .B2(n20510), .ZN(
        n20498) );
  INV_X1 U23466 ( .A(n20498), .ZN(n20500) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20514), .B1(
        n20668), .B2(n20513), .ZN(n20499) );
  OAI211_X1 U23468 ( .C1(n20673), .C2(n20557), .A(n20500), .B(n20499), .ZN(
        P1_U3116) );
  OAI22_X1 U23469 ( .A1(n20557), .A2(n20679), .B1(n20744), .B2(n20510), .ZN(
        n20501) );
  INV_X1 U23470 ( .A(n20501), .ZN(n20503) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20514), .B1(
        n20674), .B2(n20513), .ZN(n20502) );
  OAI211_X1 U23472 ( .C1(n20749), .C2(n20511), .A(n20503), .B(n20502), .ZN(
        P1_U3117) );
  OAI22_X1 U23473 ( .A1(n20557), .A2(n20685), .B1(n20751), .B2(n20510), .ZN(
        n20504) );
  INV_X1 U23474 ( .A(n20504), .ZN(n20506) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20514), .B1(
        n20680), .B2(n20513), .ZN(n20505) );
  OAI211_X1 U23476 ( .C1(n20756), .C2(n20511), .A(n20506), .B(n20505), .ZN(
        P1_U3118) );
  OAI22_X1 U23477 ( .A1(n20511), .A2(n20763), .B1(n20758), .B2(n20510), .ZN(
        n20507) );
  INV_X1 U23478 ( .A(n20507), .ZN(n20509) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20514), .B1(
        n20686), .B2(n20513), .ZN(n20508) );
  OAI211_X1 U23480 ( .C1(n20691), .C2(n20557), .A(n20509), .B(n20508), .ZN(
        P1_U3119) );
  OAI22_X1 U23481 ( .A1(n20511), .A2(n20775), .B1(n20767), .B2(n20510), .ZN(
        n20512) );
  INV_X1 U23482 ( .A(n20512), .ZN(n20516) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20514), .B1(
        n20693), .B2(n20513), .ZN(n20515) );
  OAI211_X1 U23484 ( .C1(n20701), .C2(n20557), .A(n20516), .B(n20515), .ZN(
        P1_U3120) );
  NAND2_X1 U23485 ( .A1(n20517), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20551) );
  OR2_X1 U23486 ( .A1(n20518), .A2(n20702), .ZN(n20519) );
  OR2_X1 U23487 ( .A1(n20523), .A2(n20635), .ZN(n20521) );
  NAND2_X1 U23488 ( .A1(n20526), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20520) );
  OAI22_X1 U23489 ( .A1(n20709), .A2(n20551), .B1(n20550), .B2(n20708), .ZN(
        n20522) );
  INV_X1 U23490 ( .A(n20522), .ZN(n20530) );
  OAI21_X1 U23491 ( .B1(n20713), .B2(n20524), .A(n20523), .ZN(n20525) );
  OAI211_X1 U23492 ( .C1(n20716), .C2(n20526), .A(n20715), .B(n20525), .ZN(
        n20554) );
  INV_X1 U23493 ( .A(n20599), .ZN(n20553) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20554), .B1(
        n20553), .B2(n20718), .ZN(n20529) );
  OAI211_X1 U23495 ( .C1(n20721), .C2(n20557), .A(n20530), .B(n20529), .ZN(
        P1_U3121) );
  OAI22_X1 U23496 ( .A1(n20723), .A2(n20551), .B1(n20550), .B2(n20722), .ZN(
        n20531) );
  INV_X1 U23497 ( .A(n20531), .ZN(n20533) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20554), .B1(
        n20544), .B2(n20658), .ZN(n20532) );
  OAI211_X1 U23499 ( .C1(n20661), .C2(n20599), .A(n20533), .B(n20532), .ZN(
        P1_U3122) );
  OAI22_X1 U23500 ( .A1(n20730), .A2(n20551), .B1(n20550), .B2(n20729), .ZN(
        n20534) );
  INV_X1 U23501 ( .A(n20534), .ZN(n20536) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20554), .B1(
        n20544), .B2(n20664), .ZN(n20535) );
  OAI211_X1 U23503 ( .C1(n20667), .C2(n20599), .A(n20536), .B(n20535), .ZN(
        P1_U3123) );
  OAI22_X1 U23504 ( .A1(n20737), .A2(n20551), .B1(n20550), .B2(n20736), .ZN(
        n20537) );
  INV_X1 U23505 ( .A(n20537), .ZN(n20539) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20554), .B1(
        n20553), .B2(n20739), .ZN(n20538) );
  OAI211_X1 U23507 ( .C1(n20742), .C2(n20557), .A(n20539), .B(n20538), .ZN(
        P1_U3124) );
  OAI22_X1 U23508 ( .A1(n20744), .A2(n20551), .B1(n20550), .B2(n20743), .ZN(
        n20540) );
  INV_X1 U23509 ( .A(n20540), .ZN(n20542) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20554), .B1(
        n20553), .B2(n20746), .ZN(n20541) );
  OAI211_X1 U23511 ( .C1(n20749), .C2(n20557), .A(n20542), .B(n20541), .ZN(
        P1_U3125) );
  OAI22_X1 U23512 ( .A1(n20751), .A2(n20551), .B1(n20550), .B2(n20750), .ZN(
        n20543) );
  INV_X1 U23513 ( .A(n20543), .ZN(n20546) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20554), .B1(
        n20544), .B2(n20682), .ZN(n20545) );
  OAI211_X1 U23515 ( .C1(n20685), .C2(n20599), .A(n20546), .B(n20545), .ZN(
        P1_U3126) );
  OAI22_X1 U23516 ( .A1(n20758), .A2(n20551), .B1(n20550), .B2(n20757), .ZN(
        n20547) );
  INV_X1 U23517 ( .A(n20547), .ZN(n20549) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20554), .B1(
        n20553), .B2(n20760), .ZN(n20548) );
  OAI211_X1 U23519 ( .C1(n20763), .C2(n20557), .A(n20549), .B(n20548), .ZN(
        P1_U3127) );
  OAI22_X1 U23520 ( .A1(n20767), .A2(n20551), .B1(n20550), .B2(n20764), .ZN(
        n20552) );
  INV_X1 U23521 ( .A(n20552), .ZN(n20556) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20554), .B1(
        n20553), .B2(n20769), .ZN(n20555) );
  OAI211_X1 U23523 ( .C1(n20775), .C2(n20557), .A(n20556), .B(n20555), .ZN(
        P1_U3128) );
  NOR3_X1 U23524 ( .A1(n20560), .A2(n20559), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20610) );
  INV_X1 U23525 ( .A(n20610), .ZN(n20600) );
  NOR2_X1 U23526 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20600), .ZN(
        n20567) );
  INV_X1 U23527 ( .A(n20567), .ZN(n20593) );
  OAI22_X1 U23528 ( .A1(n20631), .A2(n20655), .B1(n20709), .B2(n20593), .ZN(
        n20561) );
  INV_X1 U23529 ( .A(n20561), .ZN(n20574) );
  NAND2_X1 U23530 ( .A1(n20599), .A2(n20631), .ZN(n20562) );
  AOI21_X1 U23531 ( .B1(n20562), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20635), 
        .ZN(n20568) );
  OR2_X1 U23532 ( .A1(n20564), .A2(n20563), .ZN(n20703) );
  OR2_X1 U23533 ( .A1(n20703), .A2(n20646), .ZN(n20571) );
  AOI22_X1 U23534 ( .A1(n20568), .A2(n20571), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20569), .ZN(n20565) );
  OAI211_X1 U23535 ( .C1(n20567), .C2(n20566), .A(n20650), .B(n20565), .ZN(
        n20596) );
  INV_X1 U23536 ( .A(n20568), .ZN(n20572) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20596), .B1(
        n20642), .B2(n20595), .ZN(n20573) );
  OAI211_X1 U23538 ( .C1(n20721), .C2(n20599), .A(n20574), .B(n20573), .ZN(
        P1_U3129) );
  OAI22_X1 U23539 ( .A1(n20631), .A2(n20661), .B1(n20723), .B2(n20593), .ZN(
        n20575) );
  INV_X1 U23540 ( .A(n20575), .ZN(n20577) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20596), .B1(
        n20656), .B2(n20595), .ZN(n20576) );
  OAI211_X1 U23542 ( .C1(n20728), .C2(n20599), .A(n20577), .B(n20576), .ZN(
        P1_U3130) );
  OAI22_X1 U23543 ( .A1(n20631), .A2(n20667), .B1(n20730), .B2(n20593), .ZN(
        n20578) );
  INV_X1 U23544 ( .A(n20578), .ZN(n20580) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20596), .B1(
        n20662), .B2(n20595), .ZN(n20579) );
  OAI211_X1 U23546 ( .C1(n20735), .C2(n20599), .A(n20580), .B(n20579), .ZN(
        P1_U3131) );
  OAI22_X1 U23547 ( .A1(n20631), .A2(n20673), .B1(n20737), .B2(n20593), .ZN(
        n20581) );
  INV_X1 U23548 ( .A(n20581), .ZN(n20583) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20596), .B1(
        n20668), .B2(n20595), .ZN(n20582) );
  OAI211_X1 U23550 ( .C1(n20742), .C2(n20599), .A(n20583), .B(n20582), .ZN(
        P1_U3132) );
  OAI22_X1 U23551 ( .A1(n20631), .A2(n20679), .B1(n20744), .B2(n20593), .ZN(
        n20584) );
  INV_X1 U23552 ( .A(n20584), .ZN(n20586) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20596), .B1(
        n20674), .B2(n20595), .ZN(n20585) );
  OAI211_X1 U23554 ( .C1(n20749), .C2(n20599), .A(n20586), .B(n20585), .ZN(
        P1_U3133) );
  OAI22_X1 U23555 ( .A1(n20631), .A2(n20685), .B1(n20751), .B2(n20593), .ZN(
        n20587) );
  INV_X1 U23556 ( .A(n20587), .ZN(n20589) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20596), .B1(
        n20680), .B2(n20595), .ZN(n20588) );
  OAI211_X1 U23558 ( .C1(n20756), .C2(n20599), .A(n20589), .B(n20588), .ZN(
        P1_U3134) );
  OAI22_X1 U23559 ( .A1(n20631), .A2(n20691), .B1(n20758), .B2(n20593), .ZN(
        n20590) );
  INV_X1 U23560 ( .A(n20590), .ZN(n20592) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20596), .B1(
        n20686), .B2(n20595), .ZN(n20591) );
  OAI211_X1 U23562 ( .C1(n20763), .C2(n20599), .A(n20592), .B(n20591), .ZN(
        P1_U3135) );
  OAI22_X1 U23563 ( .A1(n20631), .A2(n20701), .B1(n20767), .B2(n20593), .ZN(
        n20594) );
  INV_X1 U23564 ( .A(n20594), .ZN(n20598) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20596), .B1(
        n20693), .B2(n20595), .ZN(n20597) );
  OAI211_X1 U23566 ( .C1(n20775), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        P1_U3136) );
  NOR2_X1 U23567 ( .A1(n20601), .A2(n20600), .ZN(n20627) );
  OR2_X1 U23568 ( .A1(n20703), .A2(n20157), .ZN(n20603) );
  INV_X1 U23569 ( .A(n20627), .ZN(n20602) );
  NAND2_X1 U23570 ( .A1(n20603), .A2(n20602), .ZN(n20606) );
  NAND2_X1 U23571 ( .A1(n20606), .A2(n20377), .ZN(n20605) );
  NAND2_X1 U23572 ( .A1(n20610), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20604) );
  NAND2_X1 U23573 ( .A1(n20605), .A2(n20604), .ZN(n20626) );
  AOI22_X1 U23574 ( .A1(n20643), .A2(n20627), .B1(n20642), .B2(n20626), .ZN(
        n20613) );
  NOR2_X1 U23575 ( .A1(n20633), .A2(n20635), .ZN(n20712) );
  INV_X1 U23576 ( .A(n20606), .ZN(n20607) );
  OAI21_X1 U23577 ( .B1(n20712), .B2(n20608), .A(n20607), .ZN(n20609) );
  OAI211_X1 U23578 ( .C1(n20716), .C2(n20610), .A(n20715), .B(n20609), .ZN(
        n20628) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20718), .ZN(n20612) );
  OAI211_X1 U23580 ( .C1(n20721), .C2(n20631), .A(n20613), .B(n20612), .ZN(
        P1_U3137) );
  AOI22_X1 U23581 ( .A1(n20657), .A2(n20627), .B1(n20656), .B2(n20626), .ZN(
        n20615) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20725), .ZN(n20614) );
  OAI211_X1 U23583 ( .C1(n20728), .C2(n20631), .A(n20615), .B(n20614), .ZN(
        P1_U3138) );
  AOI22_X1 U23584 ( .A1(n20663), .A2(n20627), .B1(n20662), .B2(n20626), .ZN(
        n20617) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20732), .ZN(n20616) );
  OAI211_X1 U23586 ( .C1(n20735), .C2(n20631), .A(n20617), .B(n20616), .ZN(
        P1_U3139) );
  AOI22_X1 U23587 ( .A1(n20669), .A2(n20627), .B1(n20668), .B2(n20626), .ZN(
        n20619) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20739), .ZN(n20618) );
  OAI211_X1 U23589 ( .C1(n20742), .C2(n20631), .A(n20619), .B(n20618), .ZN(
        P1_U3140) );
  AOI22_X1 U23590 ( .A1(n20675), .A2(n20627), .B1(n20674), .B2(n20626), .ZN(
        n20621) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20746), .ZN(n20620) );
  OAI211_X1 U23592 ( .C1(n20749), .C2(n20631), .A(n20621), .B(n20620), .ZN(
        P1_U3141) );
  AOI22_X1 U23593 ( .A1(n20681), .A2(n20627), .B1(n20680), .B2(n20626), .ZN(
        n20623) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20753), .ZN(n20622) );
  OAI211_X1 U23595 ( .C1(n20756), .C2(n20631), .A(n20623), .B(n20622), .ZN(
        P1_U3142) );
  AOI22_X1 U23596 ( .A1(n20687), .A2(n20627), .B1(n20686), .B2(n20626), .ZN(
        n20625) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20760), .ZN(n20624) );
  OAI211_X1 U23598 ( .C1(n20763), .C2(n20631), .A(n20625), .B(n20624), .ZN(
        P1_U3143) );
  AOI22_X1 U23599 ( .A1(n20695), .A2(n20627), .B1(n20693), .B2(n20626), .ZN(
        n20630) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20628), .B1(
        n20697), .B2(n20769), .ZN(n20629) );
  OAI211_X1 U23601 ( .C1(n20775), .C2(n20631), .A(n20630), .B(n20629), .ZN(
        P1_U3144) );
  INV_X1 U23602 ( .A(n20717), .ZN(n20634) );
  NOR2_X1 U23603 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20634), .ZN(
        n20694) );
  OR2_X1 U23604 ( .A1(n14265), .A2(n20635), .ZN(n20636) );
  OR2_X1 U23605 ( .A1(n20703), .A2(n20636), .ZN(n20641) );
  INV_X1 U23606 ( .A(n20637), .ZN(n20638) );
  NAND2_X1 U23607 ( .A1(n20639), .A2(n20638), .ZN(n20640) );
  NAND2_X1 U23608 ( .A1(n20641), .A2(n20640), .ZN(n20692) );
  AOI22_X1 U23609 ( .A1(n20643), .A2(n20694), .B1(n20642), .B2(n20692), .ZN(
        n20654) );
  INV_X1 U23610 ( .A(n20703), .ZN(n20647) );
  INV_X1 U23611 ( .A(n20697), .ZN(n20644) );
  AOI21_X1 U23612 ( .B1(n20644), .B2(n20774), .A(n20857), .ZN(n20645) );
  AOI21_X1 U23613 ( .B1(n20647), .B2(n20646), .A(n20645), .ZN(n20648) );
  NOR2_X1 U23614 ( .A1(n20648), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20651) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20652), .ZN(n20653) );
  OAI211_X1 U23616 ( .C1(n20655), .C2(n20774), .A(n20654), .B(n20653), .ZN(
        P1_U3145) );
  AOI22_X1 U23617 ( .A1(n20657), .A2(n20694), .B1(n20656), .B2(n20692), .ZN(
        n20660) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20658), .ZN(n20659) );
  OAI211_X1 U23619 ( .C1(n20661), .C2(n20774), .A(n20660), .B(n20659), .ZN(
        P1_U3146) );
  AOI22_X1 U23620 ( .A1(n20663), .A2(n20694), .B1(n20662), .B2(n20692), .ZN(
        n20666) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20664), .ZN(n20665) );
  OAI211_X1 U23622 ( .C1(n20667), .C2(n20774), .A(n20666), .B(n20665), .ZN(
        P1_U3147) );
  AOI22_X1 U23623 ( .A1(n20669), .A2(n20694), .B1(n20668), .B2(n20692), .ZN(
        n20672) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20670), .ZN(n20671) );
  OAI211_X1 U23625 ( .C1(n20673), .C2(n20774), .A(n20672), .B(n20671), .ZN(
        P1_U3148) );
  AOI22_X1 U23626 ( .A1(n20675), .A2(n20694), .B1(n20674), .B2(n20692), .ZN(
        n20678) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20676), .ZN(n20677) );
  OAI211_X1 U23628 ( .C1(n20679), .C2(n20774), .A(n20678), .B(n20677), .ZN(
        P1_U3149) );
  AOI22_X1 U23629 ( .A1(n20681), .A2(n20694), .B1(n20680), .B2(n20692), .ZN(
        n20684) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20682), .ZN(n20683) );
  OAI211_X1 U23631 ( .C1(n20685), .C2(n20774), .A(n20684), .B(n20683), .ZN(
        P1_U3150) );
  AOI22_X1 U23632 ( .A1(n20687), .A2(n20694), .B1(n20686), .B2(n20692), .ZN(
        n20690) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20688), .ZN(n20689) );
  OAI211_X1 U23634 ( .C1(n20691), .C2(n20774), .A(n20690), .B(n20689), .ZN(
        P1_U3151) );
  AOI22_X1 U23635 ( .A1(n20695), .A2(n20694), .B1(n20693), .B2(n20692), .ZN(
        n20700) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20698), .B1(
        n20697), .B2(n20696), .ZN(n20699) );
  OAI211_X1 U23637 ( .C1(n20701), .C2(n20774), .A(n20700), .B(n20699), .ZN(
        P1_U3152) );
  OR2_X1 U23638 ( .A1(n20703), .A2(n20702), .ZN(n20704) );
  AND2_X1 U23639 ( .A1(n20704), .A2(n20766), .ZN(n20711) );
  INV_X1 U23640 ( .A(n20711), .ZN(n20705) );
  NAND2_X1 U23641 ( .A1(n20705), .A2(n20377), .ZN(n20707) );
  NAND2_X1 U23642 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20717), .ZN(n20706) );
  OAI22_X1 U23643 ( .A1(n20709), .A2(n20766), .B1(n20765), .B2(n20708), .ZN(
        n20710) );
  INV_X1 U23644 ( .A(n20710), .ZN(n20720) );
  OAI21_X1 U23645 ( .B1(n20713), .B2(n20712), .A(n20711), .ZN(n20714) );
  OAI211_X1 U23646 ( .C1(n20717), .C2(n20716), .A(n20715), .B(n20714), .ZN(
        n20771) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20718), .ZN(n20719) );
  OAI211_X1 U23648 ( .C1(n20721), .C2(n20774), .A(n20720), .B(n20719), .ZN(
        P1_U3153) );
  OAI22_X1 U23649 ( .A1(n20723), .A2(n20766), .B1(n20765), .B2(n20722), .ZN(
        n20724) );
  INV_X1 U23650 ( .A(n20724), .ZN(n20727) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20725), .ZN(n20726) );
  OAI211_X1 U23652 ( .C1(n20728), .C2(n20774), .A(n20727), .B(n20726), .ZN(
        P1_U3154) );
  OAI22_X1 U23653 ( .A1(n20730), .A2(n20766), .B1(n20765), .B2(n20729), .ZN(
        n20731) );
  INV_X1 U23654 ( .A(n20731), .ZN(n20734) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20732), .ZN(n20733) );
  OAI211_X1 U23656 ( .C1(n20735), .C2(n20774), .A(n20734), .B(n20733), .ZN(
        P1_U3155) );
  OAI22_X1 U23657 ( .A1(n20737), .A2(n20766), .B1(n20765), .B2(n20736), .ZN(
        n20738) );
  INV_X1 U23658 ( .A(n20738), .ZN(n20741) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20739), .ZN(n20740) );
  OAI211_X1 U23660 ( .C1(n20742), .C2(n20774), .A(n20741), .B(n20740), .ZN(
        P1_U3156) );
  OAI22_X1 U23661 ( .A1(n20744), .A2(n20766), .B1(n20765), .B2(n20743), .ZN(
        n20745) );
  INV_X1 U23662 ( .A(n20745), .ZN(n20748) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20746), .ZN(n20747) );
  OAI211_X1 U23664 ( .C1(n20749), .C2(n20774), .A(n20748), .B(n20747), .ZN(
        P1_U3157) );
  OAI22_X1 U23665 ( .A1(n20751), .A2(n20766), .B1(n20765), .B2(n20750), .ZN(
        n20752) );
  INV_X1 U23666 ( .A(n20752), .ZN(n20755) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20753), .ZN(n20754) );
  OAI211_X1 U23668 ( .C1(n20756), .C2(n20774), .A(n20755), .B(n20754), .ZN(
        P1_U3158) );
  OAI22_X1 U23669 ( .A1(n20758), .A2(n20766), .B1(n20765), .B2(n20757), .ZN(
        n20759) );
  INV_X1 U23670 ( .A(n20759), .ZN(n20762) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20760), .ZN(n20761) );
  OAI211_X1 U23672 ( .C1(n20763), .C2(n20774), .A(n20762), .B(n20761), .ZN(
        P1_U3159) );
  OAI22_X1 U23673 ( .A1(n20767), .A2(n20766), .B1(n20765), .B2(n20764), .ZN(
        n20768) );
  INV_X1 U23674 ( .A(n20768), .ZN(n20773) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20771), .B1(
        n20770), .B2(n20769), .ZN(n20772) );
  OAI211_X1 U23676 ( .C1(n20775), .C2(n20774), .A(n20773), .B(n20772), .ZN(
        P1_U3160) );
  NOR2_X1 U23677 ( .A1(n20777), .A2(n20776), .ZN(n20779) );
  OAI21_X1 U23678 ( .B1(n20779), .B2(n20856), .A(n20778), .ZN(P1_U3163) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20780), .ZN(
        P1_U3164) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20780), .ZN(
        P1_U3165) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20780), .ZN(
        P1_U3166) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20780), .ZN(
        P1_U3167) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20780), .ZN(
        P1_U3168) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20780), .ZN(
        P1_U3169) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20780), .ZN(
        P1_U3170) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20780), .ZN(
        P1_U3171) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20780), .ZN(
        P1_U3172) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20780), .ZN(
        P1_U3173) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20780), .ZN(
        P1_U3174) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20780), .ZN(
        P1_U3175) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20780), .ZN(
        P1_U3176) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20780), .ZN(
        P1_U3177) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20780), .ZN(
        P1_U3178) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20780), .ZN(
        P1_U3179) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20780), .ZN(
        P1_U3180) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20780), .ZN(
        P1_U3181) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20780), .ZN(
        P1_U3182) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20780), .ZN(
        P1_U3183) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20780), .ZN(
        P1_U3184) );
  AND2_X1 U23700 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20780), .ZN(
        P1_U3185) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20780), .ZN(P1_U3186) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20780), .ZN(P1_U3187) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20780), .ZN(P1_U3188) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20780), .ZN(P1_U3189) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20780), .ZN(P1_U3190) );
  AND2_X1 U23706 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20780), .ZN(P1_U3191) );
  AND2_X1 U23707 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20780), .ZN(P1_U3192) );
  AND2_X1 U23708 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20780), .ZN(P1_U3193) );
  AOI21_X1 U23709 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20781), .A(n20970), 
        .ZN(n20793) );
  NOR2_X1 U23710 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20783) );
  NOR2_X1 U23711 ( .A1(n20783), .A2(n20782), .ZN(n20784) );
  AOI211_X1 U23712 ( .C1(NA), .C2(n20970), .A(n20784), .B(n20790), .ZN(n20785)
         );
  OAI22_X1 U23713 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20793), .B1(n20868), 
        .B2(n20785), .ZN(P1_U3194) );
  NOR2_X1 U23714 ( .A1(n11754), .A2(n20794), .ZN(n20788) );
  OAI22_X1 U23715 ( .A1(n20788), .A2(n20787), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20786), .ZN(n20792) );
  OAI211_X1 U23716 ( .C1(NA), .C2(n20864), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20794), .ZN(n20789) );
  OAI211_X1 U23717 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20790), .A(HOLD), .B(
        n20789), .ZN(n20791) );
  OAI22_X1 U23718 ( .A1(n20793), .A2(n20792), .B1(n20970), .B2(n20791), .ZN(
        P1_U3196) );
  OR2_X1 U23719 ( .A1(n20869), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20839) );
  INV_X1 U23720 ( .A(n20835), .ZN(n20837) );
  AOI222_X1 U23721 ( .A1(n20833), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20837), .ZN(n20795) );
  INV_X1 U23722 ( .A(n20795), .ZN(P1_U3197) );
  AOI222_X1 U23723 ( .A1(n20837), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20833), .ZN(n20796) );
  INV_X1 U23724 ( .A(n20796), .ZN(P1_U3198) );
  OAI222_X1 U23725 ( .A1(n20835), .A2(n13620), .B1(n20797), .B2(n20868), .C1(
        n20799), .C2(n20839), .ZN(P1_U3199) );
  AOI22_X1 U23726 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20833), .ZN(n20798) );
  OAI21_X1 U23727 ( .B1(n20799), .B2(n20835), .A(n20798), .ZN(P1_U3200) );
  AOI22_X1 U23728 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20837), .ZN(n20800) );
  OAI21_X1 U23729 ( .B1(n20801), .B2(n20839), .A(n20800), .ZN(P1_U3201) );
  AOI222_X1 U23730 ( .A1(n20837), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20833), .ZN(n20802) );
  INV_X1 U23731 ( .A(n20802), .ZN(P1_U3202) );
  AOI222_X1 U23732 ( .A1(n20837), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20833), .ZN(n20803) );
  INV_X1 U23733 ( .A(n20803), .ZN(P1_U3203) );
  AOI222_X1 U23734 ( .A1(n20833), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20837), .ZN(n20804) );
  INV_X1 U23735 ( .A(n20804), .ZN(P1_U3204) );
  AOI222_X1 U23736 ( .A1(n20837), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20833), .ZN(n20805) );
  INV_X1 U23737 ( .A(n20805), .ZN(P1_U3205) );
  AOI222_X1 U23738 ( .A1(n20837), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20833), .ZN(n20806) );
  INV_X1 U23739 ( .A(n20806), .ZN(P1_U3206) );
  AOI222_X1 U23740 ( .A1(n20837), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20833), .ZN(n20807) );
  INV_X1 U23741 ( .A(n20807), .ZN(P1_U3207) );
  AOI222_X1 U23742 ( .A1(n20837), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20833), .ZN(n20808) );
  INV_X1 U23743 ( .A(n20808), .ZN(P1_U3208) );
  AOI22_X1 U23744 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20833), .ZN(n20809) );
  OAI21_X1 U23745 ( .B1(n20810), .B2(n20835), .A(n20809), .ZN(P1_U3209) );
  AOI22_X1 U23746 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20837), .ZN(n20811) );
  OAI21_X1 U23747 ( .B1(n20812), .B2(n20839), .A(n20811), .ZN(P1_U3210) );
  AOI222_X1 U23748 ( .A1(n20837), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20833), .ZN(n20813) );
  INV_X1 U23749 ( .A(n20813), .ZN(P1_U3211) );
  AOI222_X1 U23750 ( .A1(n20837), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20833), .ZN(n20814) );
  INV_X1 U23751 ( .A(n20814), .ZN(P1_U3212) );
  AOI222_X1 U23752 ( .A1(n20837), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20833), .ZN(n20815) );
  INV_X1 U23753 ( .A(n20815), .ZN(P1_U3213) );
  AOI222_X1 U23754 ( .A1(n20837), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20833), .ZN(n20816) );
  INV_X1 U23755 ( .A(n20816), .ZN(P1_U3214) );
  AOI22_X1 U23756 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20833), .ZN(n20817) );
  OAI21_X1 U23757 ( .B1(n20818), .B2(n20835), .A(n20817), .ZN(P1_U3215) );
  AOI22_X1 U23758 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20837), .ZN(n20819) );
  OAI21_X1 U23759 ( .B1(n20820), .B2(n20839), .A(n20819), .ZN(P1_U3216) );
  AOI222_X1 U23760 ( .A1(n20837), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20833), .ZN(n20821) );
  INV_X1 U23761 ( .A(n20821), .ZN(P1_U3217) );
  AOI22_X1 U23762 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20833), .ZN(n20822) );
  OAI21_X1 U23763 ( .B1(n20823), .B2(n20835), .A(n20822), .ZN(P1_U3218) );
  AOI22_X1 U23764 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20869), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20837), .ZN(n20824) );
  OAI21_X1 U23765 ( .B1(n20825), .B2(n20839), .A(n20824), .ZN(P1_U3219) );
  AOI222_X1 U23766 ( .A1(n20837), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20833), .ZN(n20826) );
  INV_X1 U23767 ( .A(n20826), .ZN(P1_U3220) );
  AOI222_X1 U23768 ( .A1(n20837), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20833), .ZN(n20827) );
  INV_X1 U23769 ( .A(n20827), .ZN(P1_U3221) );
  AOI22_X1 U23770 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20833), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20869), .ZN(n20828) );
  OAI21_X1 U23771 ( .B1(n20829), .B2(n20835), .A(n20828), .ZN(P1_U3222) );
  AOI22_X1 U23772 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20837), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20869), .ZN(n20830) );
  OAI21_X1 U23773 ( .B1(n20831), .B2(n20839), .A(n20830), .ZN(P1_U3223) );
  AOI222_X1 U23774 ( .A1(n20837), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20869), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20833), .ZN(n20832) );
  INV_X1 U23775 ( .A(n20832), .ZN(P1_U3224) );
  AOI22_X1 U23776 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20833), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20869), .ZN(n20834) );
  OAI21_X1 U23777 ( .B1(n20836), .B2(n20835), .A(n20834), .ZN(P1_U3225) );
  AOI22_X1 U23778 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20837), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20869), .ZN(n20838) );
  OAI21_X1 U23779 ( .B1(n20840), .B2(n20839), .A(n20838), .ZN(P1_U3226) );
  OAI22_X1 U23780 ( .A1(n20869), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20868), .ZN(n20841) );
  INV_X1 U23781 ( .A(n20841), .ZN(P1_U3458) );
  MUX2_X1 U23782 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(P1_BE_N_REG_2__SCAN_IN), .S(n20869), .Z(P1_U3459) );
  MUX2_X1 U23783 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(P1_BE_N_REG_1__SCAN_IN), .S(n20869), .Z(P1_U3460) );
  MUX2_X1 U23784 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(P1_BE_N_REG_0__SCAN_IN), .S(n20869), .Z(P1_U3461) );
  OAI21_X1 U23785 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20845), .A(n20843), 
        .ZN(n20842) );
  INV_X1 U23786 ( .A(n20842), .ZN(P1_U3464) );
  OAI21_X1 U23787 ( .B1(n20845), .B2(n20844), .A(n20843), .ZN(P1_U3465) );
  NAND2_X1 U23788 ( .A1(n20846), .A2(n20946), .ZN(n20852) );
  OAI21_X1 U23789 ( .B1(n20847), .B2(n20946), .A(n20853), .ZN(n20848) );
  OAI21_X1 U23790 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20853), .A(n20848), 
        .ZN(n20849) );
  OAI221_X1 U23791 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20851), .C1(n20850), .C2(n20852), .A(n20849), .ZN(P1_U3481) );
  OAI21_X1 U23792 ( .B1(n20853), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n20852), 
        .ZN(n20854) );
  INV_X1 U23793 ( .A(n20854), .ZN(P1_U3482) );
  AOI22_X1 U23794 ( .A1(n20868), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20855), 
        .B2(n20869), .ZN(P1_U3483) );
  AOI21_X1 U23795 ( .B1(n11773), .B2(n20857), .A(n20856), .ZN(n20860) );
  AOI211_X1 U23796 ( .C1(n20861), .C2(n20860), .A(n20859), .B(n20858), .ZN(
        n20867) );
  AOI211_X1 U23797 ( .C1(n20865), .C2(n20864), .A(n20863), .B(n20862), .ZN(
        n20866) );
  MUX2_X1 U23798 ( .A(n20867), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20866), 
        .Z(P1_U3485) );
  OAI22_X1 U23799 ( .A1(n20869), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20868), .ZN(n20870) );
  INV_X1 U23800 ( .A(n20870), .ZN(P1_U3486) );
  INV_X1 U23801 ( .A(keyinput26), .ZN(n20872) );
  AOI22_X1 U23802 ( .A1(n20873), .A2(keyinput3), .B1(P1_BE_N_REG_3__SCAN_IN), 
        .B2(n20872), .ZN(n20871) );
  OAI221_X1 U23803 ( .B1(n20873), .B2(keyinput3), .C1(n20872), .C2(
        P1_BE_N_REG_3__SCAN_IN), .A(n20871), .ZN(n20885) );
  AOI22_X1 U23804 ( .A1(n20876), .A2(keyinput51), .B1(keyinput11), .B2(n20875), 
        .ZN(n20874) );
  OAI221_X1 U23805 ( .B1(n20876), .B2(keyinput51), .C1(n20875), .C2(keyinput11), .A(n20874), .ZN(n20884) );
  INV_X1 U23806 ( .A(READY11_REG_SCAN_IN), .ZN(n20879) );
  INV_X1 U23807 ( .A(keyinput48), .ZN(n20878) );
  AOI22_X1 U23808 ( .A1(n20879), .A2(keyinput16), .B1(P3_LWORD_REG_4__SCAN_IN), 
        .B2(n20878), .ZN(n20877) );
  OAI221_X1 U23809 ( .B1(n20879), .B2(keyinput16), .C1(n20878), .C2(
        P3_LWORD_REG_4__SCAN_IN), .A(n20877), .ZN(n20883) );
  INV_X1 U23810 ( .A(DATAI_31_), .ZN(n20881) );
  AOI22_X1 U23811 ( .A1(n10488), .A2(keyinput29), .B1(keyinput30), .B2(n20881), 
        .ZN(n20880) );
  OAI221_X1 U23812 ( .B1(n10488), .B2(keyinput29), .C1(n20881), .C2(keyinput30), .A(n20880), .ZN(n20882) );
  NOR4_X1 U23813 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n21032) );
  INV_X1 U23814 ( .A(keyinput5), .ZN(n20887) );
  AOI22_X1 U23815 ( .A1(n20888), .A2(keyinput15), .B1(
        P2_MEMORYFETCH_REG_SCAN_IN), .B2(n20887), .ZN(n20886) );
  OAI221_X1 U23816 ( .B1(n20888), .B2(keyinput15), .C1(n20887), .C2(
        P2_MEMORYFETCH_REG_SCAN_IN), .A(n20886), .ZN(n20900) );
  INV_X1 U23817 ( .A(keyinput61), .ZN(n20890) );
  AOI22_X1 U23818 ( .A1(n20891), .A2(keyinput49), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n20890), .ZN(n20889) );
  OAI221_X1 U23819 ( .B1(n20891), .B2(keyinput49), .C1(n20890), .C2(
        P3_ADDRESS_REG_28__SCAN_IN), .A(n20889), .ZN(n20899) );
  INV_X1 U23820 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23821 ( .A1(n20894), .A2(keyinput42), .B1(keyinput2), .B2(n20893), 
        .ZN(n20892) );
  OAI221_X1 U23822 ( .B1(n20894), .B2(keyinput42), .C1(n20893), .C2(keyinput2), 
        .A(n20892), .ZN(n20898) );
  INV_X1 U23823 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U23824 ( .A1(n12386), .A2(keyinput24), .B1(keyinput12), .B2(n20896), 
        .ZN(n20895) );
  OAI221_X1 U23825 ( .B1(n12386), .B2(keyinput24), .C1(n20896), .C2(keyinput12), .A(n20895), .ZN(n20897) );
  NOR4_X1 U23826 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n21031) );
  AOI22_X1 U23827 ( .A1(n20902), .A2(keyinput58), .B1(n14067), .B2(keyinput39), 
        .ZN(n20901) );
  OAI221_X1 U23828 ( .B1(n20902), .B2(keyinput58), .C1(n14067), .C2(keyinput39), .A(n20901), .ZN(n20914) );
  INV_X1 U23829 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n20904) );
  AOI22_X1 U23830 ( .A1(n20905), .A2(keyinput32), .B1(keyinput50), .B2(n20904), 
        .ZN(n20903) );
  OAI221_X1 U23831 ( .B1(n20905), .B2(keyinput32), .C1(n20904), .C2(keyinput50), .A(n20903), .ZN(n20913) );
  INV_X1 U23832 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n20908) );
  INV_X1 U23833 ( .A(keyinput37), .ZN(n20907) );
  AOI22_X1 U23834 ( .A1(n20908), .A2(keyinput19), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n20907), .ZN(n20906) );
  OAI221_X1 U23835 ( .B1(n20908), .B2(keyinput19), .C1(n20907), .C2(
        P3_ADDRESS_REG_10__SCAN_IN), .A(n20906), .ZN(n20912) );
  AOI22_X1 U23836 ( .A1(n20910), .A2(keyinput53), .B1(n11236), .B2(keyinput41), 
        .ZN(n20909) );
  OAI221_X1 U23837 ( .B1(n20910), .B2(keyinput53), .C1(n11236), .C2(keyinput41), .A(n20909), .ZN(n20911) );
  NOR4_X1 U23838 ( .A1(n20914), .A2(n20913), .A3(n20912), .A4(n20911), .ZN(
        n20938) );
  XOR2_X1 U23839 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B(keyinput4), .Z(
        n20918) );
  XOR2_X1 U23840 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput55), .Z(
        n20917) );
  NOR3_X1 U23841 ( .A1(n20918), .A2(n20917), .A3(n20916), .ZN(n20923) );
  XOR2_X1 U23842 ( .A(keyinput38), .B(n20919), .Z(n20922) );
  XNOR2_X1 U23843 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B(keyinput9), .ZN(
        n20921) );
  XNOR2_X1 U23844 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput34), 
        .ZN(n20920) );
  NAND4_X1 U23845 ( .A1(n20923), .A2(n20922), .A3(n20921), .A4(n20920), .ZN(
        n20932) );
  INV_X1 U23846 ( .A(DATAI_4_), .ZN(n20926) );
  AOI22_X1 U23847 ( .A1(n20926), .A2(keyinput14), .B1(keyinput56), .B2(n20925), 
        .ZN(n20924) );
  OAI221_X1 U23848 ( .B1(n20926), .B2(keyinput14), .C1(n20925), .C2(keyinput56), .A(n20924), .ZN(n20931) );
  INV_X1 U23849 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n20928) );
  AOI22_X1 U23850 ( .A1(n20929), .A2(keyinput33), .B1(keyinput13), .B2(n20928), 
        .ZN(n20927) );
  OAI221_X1 U23851 ( .B1(n20929), .B2(keyinput33), .C1(n20928), .C2(keyinput13), .A(n20927), .ZN(n20930) );
  NOR3_X1 U23852 ( .A1(n20932), .A2(n20931), .A3(n20930), .ZN(n20937) );
  XOR2_X1 U23853 ( .A(keyinput52), .B(n20933), .Z(n20936) );
  XOR2_X1 U23854 ( .A(keyinput28), .B(n20934), .Z(n20935) );
  NAND4_X1 U23855 ( .A1(n20938), .A2(n20937), .A3(n20936), .A4(n20935), .ZN(
        n20964) );
  INV_X1 U23856 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n20940) );
  OAI22_X1 U23857 ( .A1(n20941), .A2(keyinput40), .B1(n20940), .B2(keyinput20), 
        .ZN(n20939) );
  AOI221_X1 U23858 ( .B1(n20941), .B2(keyinput40), .C1(keyinput20), .C2(n20940), .A(n20939), .ZN(n20962) );
  INV_X1 U23859 ( .A(keyinput63), .ZN(n20943) );
  OAI22_X1 U23860 ( .A1(keyinput22), .A2(n20944), .B1(n20943), .B2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20942) );
  AOI221_X1 U23861 ( .B1(n20944), .B2(keyinput22), .C1(n20943), .C2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A(n20942), .ZN(n20961) );
  INV_X1 U23862 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20947) );
  AOI22_X1 U23863 ( .A1(n20947), .A2(keyinput7), .B1(keyinput21), .B2(n20946), 
        .ZN(n20945) );
  OAI221_X1 U23864 ( .B1(n20947), .B2(keyinput7), .C1(n20946), .C2(keyinput21), 
        .A(n20945), .ZN(n20959) );
  AOI22_X1 U23865 ( .A1(n20950), .A2(keyinput17), .B1(n20949), .B2(keyinput27), 
        .ZN(n20948) );
  OAI221_X1 U23866 ( .B1(n20950), .B2(keyinput17), .C1(n20949), .C2(keyinput27), .A(n20948), .ZN(n20958) );
  AOI22_X1 U23867 ( .A1(n20953), .A2(keyinput46), .B1(keyinput35), .B2(n20952), 
        .ZN(n20951) );
  OAI221_X1 U23868 ( .B1(n20953), .B2(keyinput46), .C1(n20952), .C2(keyinput35), .A(n20951), .ZN(n20957) );
  AOI22_X1 U23869 ( .A1(n20955), .A2(keyinput60), .B1(n10885), .B2(keyinput31), 
        .ZN(n20954) );
  OAI221_X1 U23870 ( .B1(n20955), .B2(keyinput60), .C1(n10885), .C2(keyinput31), .A(n20954), .ZN(n20956) );
  NOR4_X1 U23871 ( .A1(n20959), .A2(n20958), .A3(n20957), .A4(n20956), .ZN(
        n20960) );
  NAND3_X1 U23872 ( .A1(n20962), .A2(n20961), .A3(n20960), .ZN(n20963) );
  NOR2_X1 U23873 ( .A1(n20964), .A2(n20963), .ZN(n20998) );
  INV_X1 U23874 ( .A(keyinput36), .ZN(n20966) );
  AOI22_X1 U23875 ( .A1(n20967), .A2(keyinput43), .B1(P3_DATAO_REG_12__SCAN_IN), .B2(n20966), .ZN(n20965) );
  OAI221_X1 U23876 ( .B1(n20967), .B2(keyinput43), .C1(n20966), .C2(
        P3_DATAO_REG_12__SCAN_IN), .A(n20965), .ZN(n20980) );
  AOI22_X1 U23877 ( .A1(n20970), .A2(keyinput10), .B1(keyinput8), .B2(n20969), 
        .ZN(n20968) );
  OAI221_X1 U23878 ( .B1(n20970), .B2(keyinput10), .C1(n20969), .C2(keyinput8), 
        .A(n20968), .ZN(n20979) );
  INV_X1 U23879 ( .A(keyinput54), .ZN(n20972) );
  AOI22_X1 U23880 ( .A1(n20973), .A2(keyinput62), .B1(
        P3_DATAWIDTH_REG_11__SCAN_IN), .B2(n20972), .ZN(n20971) );
  OAI221_X1 U23881 ( .B1(n20973), .B2(keyinput62), .C1(n20972), .C2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A(n20971), .ZN(n20978) );
  INV_X1 U23882 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U23883 ( .A1(n20976), .A2(keyinput18), .B1(n20975), .B2(keyinput6), 
        .ZN(n20974) );
  OAI221_X1 U23884 ( .B1(n20976), .B2(keyinput18), .C1(n20975), .C2(keyinput6), 
        .A(n20974), .ZN(n20977) );
  NOR4_X1 U23885 ( .A1(n20980), .A2(n20979), .A3(n20978), .A4(n20977), .ZN(
        n20997) );
  INV_X1 U23886 ( .A(keyinput57), .ZN(n20982) );
  AOI22_X1 U23887 ( .A1(n20983), .A2(keyinput25), .B1(
        P3_DATAWIDTH_REG_2__SCAN_IN), .B2(n20982), .ZN(n20981) );
  OAI221_X1 U23888 ( .B1(n20983), .B2(keyinput25), .C1(n20982), .C2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A(n20981), .ZN(n20995) );
  INV_X1 U23889 ( .A(keyinput45), .ZN(n20985) );
  AOI22_X1 U23890 ( .A1(n20986), .A2(keyinput44), .B1(
        P2_DATAWIDTH_REG_15__SCAN_IN), .B2(n20985), .ZN(n20984) );
  OAI221_X1 U23891 ( .B1(n20986), .B2(keyinput44), .C1(n20985), .C2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A(n20984), .ZN(n20994) );
  AOI22_X1 U23892 ( .A1(n12327), .A2(keyinput1), .B1(n20988), .B2(keyinput23), 
        .ZN(n20987) );
  OAI221_X1 U23893 ( .B1(n12327), .B2(keyinput1), .C1(n20988), .C2(keyinput23), 
        .A(n20987), .ZN(n20993) );
  INV_X1 U23894 ( .A(keyinput0), .ZN(n20990) );
  AOI22_X1 U23895 ( .A1(n20991), .A2(keyinput59), .B1(
        P2_BYTEENABLE_REG_1__SCAN_IN), .B2(n20990), .ZN(n20989) );
  OAI221_X1 U23896 ( .B1(n20991), .B2(keyinput59), .C1(n20990), .C2(
        P2_BYTEENABLE_REG_1__SCAN_IN), .A(n20989), .ZN(n20992) );
  NOR4_X1 U23897 ( .A1(n20995), .A2(n20994), .A3(n20993), .A4(n20992), .ZN(
        n20996) );
  AND3_X1 U23898 ( .A1(n20998), .A2(n20997), .A3(n20996), .ZN(n21030) );
  NAND3_X1 U23899 ( .A1(keyinput62), .A2(keyinput18), .A3(keyinput6), .ZN(
        n21004) );
  NAND4_X1 U23900 ( .A1(keyinput25), .A2(keyinput57), .A3(keyinput45), .A4(
        keyinput44), .ZN(n21003) );
  NOR2_X1 U23901 ( .A1(keyinput10), .A2(keyinput8), .ZN(n21001) );
  INV_X1 U23902 ( .A(keyinput1), .ZN(n20999) );
  NOR4_X1 U23903 ( .A1(keyinput59), .A2(keyinput23), .A3(keyinput0), .A4(
        n20999), .ZN(n21000) );
  NAND4_X1 U23904 ( .A1(keyinput36), .A2(keyinput43), .A3(n21001), .A4(n21000), 
        .ZN(n21002) );
  NOR4_X1 U23905 ( .A1(keyinput54), .A2(n21004), .A3(n21003), .A4(n21002), 
        .ZN(n21028) );
  NAND2_X1 U23906 ( .A1(keyinput39), .A2(keyinput55), .ZN(n21011) );
  NOR2_X1 U23907 ( .A1(keyinput19), .A2(keyinput52), .ZN(n21009) );
  NAND3_X1 U23908 ( .A1(keyinput53), .A2(keyinput41), .A3(keyinput32), .ZN(
        n21007) );
  INV_X1 U23909 ( .A(keyinput56), .ZN(n21005) );
  NAND3_X1 U23910 ( .A1(keyinput9), .A2(keyinput28), .A3(n21005), .ZN(n21006)
         );
  NOR4_X1 U23911 ( .A1(keyinput50), .A2(keyinput14), .A3(n21007), .A4(n21006), 
        .ZN(n21008) );
  NAND4_X1 U23912 ( .A1(keyinput37), .A2(keyinput4), .A3(n21009), .A4(n21008), 
        .ZN(n21010) );
  NOR4_X1 U23913 ( .A1(keyinput58), .A2(keyinput38), .A3(n21011), .A4(n21010), 
        .ZN(n21027) );
  NAND3_X1 U23914 ( .A1(keyinput61), .A2(keyinput49), .A3(keyinput15), .ZN(
        n21017) );
  NAND4_X1 U23915 ( .A1(keyinput51), .A2(keyinput11), .A3(keyinput26), .A4(
        keyinput3), .ZN(n21016) );
  NOR3_X1 U23916 ( .A1(keyinput12), .A2(keyinput42), .A3(keyinput2), .ZN(
        n21014) );
  INV_X1 U23917 ( .A(keyinput16), .ZN(n21012) );
  NOR3_X1 U23918 ( .A1(keyinput29), .A2(keyinput48), .A3(n21012), .ZN(n21013)
         );
  NAND4_X1 U23919 ( .A1(keyinput24), .A2(n21014), .A3(keyinput30), .A4(n21013), 
        .ZN(n21015) );
  NOR4_X1 U23920 ( .A1(keyinput5), .A2(n21017), .A3(n21016), .A4(n21015), .ZN(
        n21026) );
  NOR2_X1 U23921 ( .A1(keyinput13), .A2(keyinput47), .ZN(n21018) );
  NAND3_X1 U23922 ( .A1(keyinput33), .A2(keyinput34), .A3(n21018), .ZN(n21024)
         );
  NAND3_X1 U23923 ( .A1(keyinput17), .A2(keyinput7), .A3(keyinput21), .ZN(
        n21023) );
  NOR2_X1 U23924 ( .A1(keyinput63), .A2(keyinput20), .ZN(n21021) );
  INV_X1 U23925 ( .A(keyinput35), .ZN(n21019) );
  NOR4_X1 U23926 ( .A1(keyinput60), .A2(keyinput31), .A3(keyinput46), .A4(
        n21019), .ZN(n21020) );
  NAND4_X1 U23927 ( .A1(keyinput22), .A2(keyinput40), .A3(n21021), .A4(n21020), 
        .ZN(n21022) );
  NOR4_X1 U23928 ( .A1(keyinput27), .A2(n21024), .A3(n21023), .A4(n21022), 
        .ZN(n21025) );
  NAND4_X1 U23929 ( .A1(n21028), .A2(n21027), .A3(n21026), .A4(n21025), .ZN(
        n21029) );
  NAND4_X1 U23930 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21051) );
  AOI21_X1 U23931 ( .B1(n21034), .B2(n21038), .A(n21033), .ZN(n21035) );
  OAI21_X1 U23932 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21036), .A(n21035), 
        .ZN(n21049) );
  AOI21_X1 U23933 ( .B1(n21038), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n21037), 
        .ZN(n21046) );
  AOI21_X1 U23934 ( .B1(n21041), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n10709), 
        .ZN(n21044) );
  NOR3_X1 U23935 ( .A1(n21041), .A2(n21040), .A3(n21039), .ZN(n21043) );
  MUX2_X1 U23936 ( .A(n21044), .B(n21043), .S(n10710), .Z(n21045) );
  OAI21_X1 U23937 ( .B1(n21046), .B2(n21045), .A(n21049), .ZN(n21047) );
  OAI21_X1 U23938 ( .B1(n21049), .B2(n21048), .A(n21047), .ZN(n21050) );
  XNOR2_X1 U23939 ( .A(n21051), .B(n21050), .ZN(P2_U3610) );
  CLKBUF_X1 U11028 ( .A(n11792), .Z(n11793) );
  INV_X1 U11069 ( .A(n11562), .ZN(n11201) );
  NOR2_X2 U11140 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10431) );
  CLKBUF_X1 U11142 ( .A(n10703), .Z(n10743) );
  OR2_X1 U11307 ( .A1(n9857), .A2(n10816), .ZN(n10892) );
  CLKBUF_X1 U11346 ( .A(n13938), .Z(n16245) );
  CLKBUF_X1 U12101 ( .A(n10726), .Z(n13125) );
  INV_X1 U12264 ( .A(n9651), .ZN(n17238) );
  CLKBUF_X1 U12298 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n18726) );
  CLKBUF_X1 U12382 ( .A(n16533), .Z(n16541) );
  CLKBUF_X1 U12630 ( .A(n17549), .Z(n17560) );
  CLKBUF_X1 U12946 ( .A(n20044), .Z(n20865) );
endmodule

