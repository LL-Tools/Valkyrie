

module b20_C_SARLock_k_128_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308;

  INV_X1 U4943 ( .A(n6037), .ZN(n6065) );
  CLKBUF_X1 U4944 ( .A(n6529), .Z(n8764) );
  CLKBUF_X2 U4945 ( .A(n5322), .Z(n5688) );
  CLKBUF_X2 U4946 ( .A(n5297), .Z(n5757) );
  INV_X1 U4947 ( .A(n4660), .ZN(n6643) );
  NOR2_X2 U4948 ( .A1(n9609), .A2(n7081), .ZN(n9587) );
  INV_X2 U4949 ( .A(n9272), .ZN(n9609) );
  INV_X1 U4950 ( .A(P1_U3086), .ZN(n4436) );
  INV_X1 U4951 ( .A(n4436), .ZN(n4437) );
  INV_X1 U4952 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5255) );
  AND2_X1 U4953 ( .A1(n4793), .A2(n4792), .ZN(n5918) );
  OR2_X1 U4954 ( .A1(n5296), .A2(n6706), .ZN(n5270) );
  OR2_X1 U4955 ( .A1(n7885), .A2(n7961), .ZN(n5817) );
  INV_X1 U4956 ( .A(n5276), .ZN(n5577) );
  CLKBUF_X3 U4957 ( .A(n5298), .Z(n4439) );
  INV_X1 U4958 ( .A(n5236), .ZN(n5667) );
  INV_X2 U4959 ( .A(n4439), .ZN(n5283) );
  NOR2_X1 U4960 ( .A1(n9772), .A2(n8087), .ZN(n9791) );
  NAND2_X1 U4961 ( .A1(n6791), .A2(n7041), .ZN(n6668) );
  INV_X1 U4962 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U4963 ( .A1(n6724), .A2(n5876), .ZN(n5276) );
  INV_X1 U4964 ( .A(n8896), .ZN(n8911) );
  OAI22_X1 U4965 ( .A1(n9246), .A2(n9031), .B1(n9030), .B2(n4672), .ZN(n9234)
         );
  INV_X1 U4966 ( .A(n9009), .ZN(n4567) );
  NAND2_X1 U4967 ( .A1(n8479), .A2(n8477), .ZN(n5297) );
  NOR2_X2 U4968 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n5054) );
  OAI21_X2 U4969 ( .B1(n7703), .B2(n8073), .A(n4506), .ZN(n4533) );
  INV_X1 U4970 ( .A(n5235), .ZN(n8477) );
  OAI21_X1 U4971 ( .B1(n6994), .B2(n7060), .A(n7059), .ZN(n7058) );
  NAND4_X2 U4972 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n8934)
         );
  NAND2_X2 U4973 ( .A1(n8474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5229) );
  NAND2_X4 U4974 ( .A1(n6432), .A2(n6484), .ZN(n4603) );
  INV_X1 U4975 ( .A(n6522), .ZN(n8852) );
  NAND2_X2 U4976 ( .A1(n6321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5993) );
  BUF_X4 U4977 ( .A(n5296), .Z(n4438) );
  NAND2_X1 U4978 ( .A1(n8477), .A2(n5234), .ZN(n5296) );
  AOI22_X2 U4979 ( .A1(n8206), .A2(n5914), .B1(n8193), .B2(n8414), .ZN(n8191)
         );
  NAND2_X2 U4980 ( .A1(n4784), .A2(n4783), .ZN(n8206) );
  OAI21_X2 U4981 ( .B1(n5573), .B2(n5572), .A(n5134), .ZN(n5588) );
  OAI21_X2 U4982 ( .B1(n5555), .B2(n5129), .A(n5128), .ZN(n5573) );
  XNOR2_X2 U4983 ( .A(n5278), .B(n5277), .ZN(n6719) );
  AOI211_X1 U4984 ( .C1(n9382), .C2(n9311), .A(n9310), .B(n9309), .ZN(n9395)
         );
  NAND2_X1 U4985 ( .A1(n5201), .A2(n5200), .ZN(n7885) );
  NAND2_X1 U4986 ( .A1(n9311), .A2(n9058), .ZN(n9070) );
  OAI21_X1 U4987 ( .B1(n5725), .B2(SI_29_), .A(n5728), .ZN(n5744) );
  NAND2_X1 U4988 ( .A1(n4866), .A2(n5181), .ZN(n5727) );
  AND2_X1 U4989 ( .A1(n9063), .A2(n8731), .ZN(n9185) );
  AND2_X1 U4990 ( .A1(n6390), .A2(n6389), .ZN(n9196) );
  NAND2_X1 U4991 ( .A1(n6371), .A2(n6370), .ZN(n9421) );
  NAND2_X1 U4992 ( .A1(n6348), .A2(n6347), .ZN(n9429) );
  INV_X1 U4993 ( .A(n8076), .ZN(n5889) );
  INV_X1 U4994 ( .A(n7073), .ZN(n8078) );
  INV_X1 U4995 ( .A(n8077), .ZN(n9862) );
  NAND4_X1 U4996 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n7281)
         );
  INV_X1 U4997 ( .A(n6046), .ZN(n7180) );
  INV_X4 U4999 ( .A(n6065), .ZN(n6486) );
  INV_X2 U5000 ( .A(n5297), .ZN(n5282) );
  INV_X4 U5001 ( .A(n6636), .ZN(n5929) );
  NAND2_X2 U5002 ( .A1(n6345), .A2(n8911), .ZN(n6540) );
  CLKBUF_X2 U5003 ( .A(n6080), .Z(n8761) );
  NAND2_X1 U5004 ( .A1(n6668), .A2(n6640), .ZN(n6238) );
  NAND2_X1 U5005 ( .A1(n6014), .A2(n6017), .ZN(n6791) );
  INV_X4 U5006 ( .A(n6643), .ZN(n6640) );
  CLKBUF_X2 U5007 ( .A(n5060), .Z(n4660) );
  NAND2_X4 U5008 ( .A1(n4903), .A2(n4904), .ZN(n5060) );
  AND2_X1 U5009 ( .A1(n4475), .A2(n5972), .ZN(n4744) );
  AND2_X1 U5010 ( .A1(n4716), .A2(n6066), .ZN(n6081) );
  INV_X2 U5011 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X1 U5012 ( .B1(n6591), .B2(n9867), .A(n6590), .ZN(n6625) );
  AND2_X1 U5013 ( .A1(n4712), .A2(n9079), .ZN(n9393) );
  OAI21_X1 U5014 ( .B1(n6601), .B2(n9867), .A(n6600), .ZN(n8160) );
  NOR2_X1 U5015 ( .A1(n8180), .A2(n4798), .ZN(n8169) );
  NAND2_X1 U5016 ( .A1(n4871), .A2(n4870), .ZN(n4869) );
  MUX2_X1 U5017 ( .A(n8749), .B(n8748), .S(n8770), .Z(n8754) );
  OAI211_X1 U5018 ( .C1(n6404), .C2(n4612), .A(n4610), .B(n8507), .ZN(n8581)
         );
  XNOR2_X1 U5019 ( .A(n5750), .B(n5749), .ZN(n8760) );
  NAND2_X1 U5020 ( .A1(n5736), .A2(n5735), .ZN(n8392) );
  NAND2_X1 U5021 ( .A1(n4963), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U5022 ( .A1(n6489), .A2(n6488), .ZN(n9311) );
  NOR2_X1 U5023 ( .A1(n4612), .A2(n8614), .ZN(n4611) );
  NAND2_X1 U5024 ( .A1(n4855), .A2(n4853), .ZN(n7969) );
  INV_X1 U5025 ( .A(n8505), .ZN(n4612) );
  NAND2_X1 U5026 ( .A1(n5177), .A2(n5176), .ZN(n5713) );
  OR2_X1 U5027 ( .A1(n9216), .A2(n9217), .ZN(n9213) );
  NAND2_X1 U5028 ( .A1(n6406), .A2(n6405), .ZN(n9332) );
  NAND2_X1 U5029 ( .A1(n5157), .A2(n5156), .ZN(n5662) );
  NAND2_X1 U5030 ( .A1(n4974), .A2(n4485), .ZN(n8493) );
  NAND2_X1 U5031 ( .A1(n5606), .A2(n5605), .ZN(n8426) );
  AND2_X1 U5032 ( .A1(n9228), .A2(n8776), .ZN(n9249) );
  NAND2_X1 U5033 ( .A1(n7814), .A2(n8706), .ZN(n7815) );
  NAND2_X1 U5034 ( .A1(n4723), .A2(n4721), .ZN(n7814) );
  AND2_X1 U5035 ( .A1(n4836), .A2(n4835), .ZN(n7892) );
  NAND2_X1 U5036 ( .A1(n6277), .A2(n6276), .ZN(n9024) );
  AOI21_X1 U5037 ( .B1(n4620), .B2(n4619), .A(n4462), .ZN(n6177) );
  NOR2_X1 U5038 ( .A1(n9756), .A2(n4675), .ZN(n8086) );
  OR2_X1 U5039 ( .A1(n9738), .A2(n10262), .ZN(n4678) );
  OAI21_X1 U5040 ( .B1(n9146), .B2(n6477), .A(n6450), .ZN(n9052) );
  NAND2_X1 U5041 ( .A1(n5431), .A2(n4888), .ZN(n4886) );
  INV_X2 U5042 ( .A(n9661), .ZN(n9439) );
  NAND2_X2 U5043 ( .A1(n7080), .A2(n9236), .ZN(n9272) );
  NAND2_X1 U5044 ( .A1(n6920), .A2(n7300), .ZN(n5295) );
  NOR2_X2 U5045 ( .A1(n9475), .A2(n6713), .ZN(n6714) );
  OR2_X1 U5046 ( .A1(n8080), .A2(n6992), .ZN(n6979) );
  INV_X1 U5047 ( .A(n7640), .ZN(n4657) );
  NAND2_X1 U5048 ( .A1(n5290), .A2(n5289), .ZN(n8080) );
  INV_X1 U5049 ( .A(n7258), .ZN(n8075) );
  OAI211_X1 U5050 ( .C1(n5473), .C2(n6647), .A(n5311), .B(n5310), .ZN(n9852)
         );
  NAND4_X1 U5051 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n8077)
         );
  INV_X2 U5052 ( .A(n5473), .ZN(n5751) );
  AND4_X2 U5053 ( .A1(n5268), .A2(n5269), .A3(n5267), .A4(n5270), .ZN(n5881)
         );
  INV_X2 U5054 ( .A(n6304), .ZN(n8765) );
  AND2_X1 U5055 ( .A1(n5276), .A2(n6643), .ZN(n5275) );
  BUF_X2 U5056 ( .A(n6889), .Z(n8766) );
  AND2_X2 U5057 ( .A1(n5983), .A2(n5982), .ZN(n6889) );
  AND2_X2 U5058 ( .A1(n5983), .A2(n7889), .ZN(n6529) );
  AND2_X2 U5059 ( .A1(n5981), .A2(n7889), .ZN(n6074) );
  NAND2_X2 U5060 ( .A1(n6572), .A2(n6917), .ZN(n6636) );
  NAND2_X1 U5061 ( .A1(n9674), .A2(n6769), .ZN(n4688) );
  NAND2_X1 U5062 ( .A1(n4773), .A2(n4771), .ZN(n6724) );
  INV_X2 U5063 ( .A(n6238), .ZN(n8759) );
  NAND2_X1 U5064 ( .A1(n6506), .A2(n6001), .ZN(n8896) );
  XNOR2_X1 U5065 ( .A(n5576), .B(n5575), .ZN(n8125) );
  NAND2_X1 U5066 ( .A1(n5872), .A2(n4457), .ZN(n7865) );
  OR2_X1 U5067 ( .A1(n9676), .A2(n9677), .ZN(n9674) );
  OAI21_X1 U5068 ( .B1(n6008), .B2(n6007), .A(n6006), .ZN(n7874) );
  NAND2_X2 U5069 ( .A1(n6640), .A2(P1_U3086), .ZN(n7778) );
  XNOR2_X1 U5070 ( .A(n6003), .B(n6002), .ZN(n6522) );
  XNOR2_X1 U5071 ( .A(n6009), .B(n5972), .ZN(n7868) );
  NAND2_X1 U5072 ( .A1(n4459), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U5073 ( .A1(n6008), .A2(n6007), .ZN(n6006) );
  NAND2_X1 U5074 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6003) );
  XNOR2_X1 U5075 ( .A(n5996), .B(n5995), .ZN(n8808) );
  OR2_X1 U5076 ( .A1(n5542), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5556) );
  OR2_X1 U5077 ( .A1(n5994), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U5078 ( .A(n5341), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6905) );
  AND2_X1 U5079 ( .A1(n4549), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5053) );
  INV_X1 U5080 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6007) );
  NOR2_X2 U5081 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6047) );
  INV_X1 U5082 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5995) );
  INV_X1 U5083 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5558) );
  INV_X1 U5084 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6002) );
  INV_X1 U5085 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5992) );
  INV_X1 U5086 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5999) );
  INV_X1 U5087 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10248) );
  NOR2_X2 U5088 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4717) );
  INV_X1 U5089 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5508) );
  INV_X1 U5090 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5493) );
  INV_X1 U5091 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4549) );
  INV_X4 U5092 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5093 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5188) );
  INV_X1 U5094 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9007) );
  INV_X2 U5095 ( .A(n7112), .ZN(n7295) );
  AOI21_X2 U5096 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8126), .A(n9822), .ZN(
        n8092) );
  OR2_X1 U5097 ( .A1(n5298), .A2(n6705), .ZN(n5269) );
  NOR2_X1 U5098 ( .A1(n8181), .A2(n8186), .ZN(n8180) );
  NAND2_X2 U5099 ( .A1(n5295), .A2(n5768), .ZN(n5769) );
  NAND2_X1 U5100 ( .A1(n5235), .A2(n5234), .ZN(n5298) );
  OAI21_X2 U5101 ( .B1(n7070), .B2(n5888), .A(n5887), .ZN(n7207) );
  NAND2_X2 U5102 ( .A1(n5886), .A2(n5885), .ZN(n7070) );
  INV_X1 U5103 ( .A(n4439), .ZN(n4440) );
  NAND2_X1 U5104 ( .A1(n5600), .A2(n5929), .ZN(n4655) );
  NAND2_X1 U5105 ( .A1(n4998), .A2(n4495), .ZN(n4997) );
  NAND2_X1 U5106 ( .A1(n4999), .A2(n7812), .ZN(n4998) );
  INV_X1 U5107 ( .A(n5000), .ZN(n4999) );
  INV_X1 U5108 ( .A(n5522), .ZN(n5117) );
  NOR2_X1 U5109 ( .A1(n5871), .A2(n4943), .ZN(n5197) );
  OR2_X1 U5110 ( .A1(n8230), .A2(n8229), .ZN(n4790) );
  INV_X1 U5111 ( .A(n6441), .ZN(n4986) );
  OR2_X1 U5112 ( .A1(n9311), .A2(n9058), .ZN(n8829) );
  NAND2_X1 U5113 ( .A1(n9002), .A2(n8896), .ZN(n8770) );
  INV_X1 U5114 ( .A(n5102), .ZN(n4889) );
  CLKBUF_X1 U5115 ( .A(n5284), .Z(n5236) );
  OR2_X1 U5116 ( .A1(n5911), .A2(n7906), .ZN(n5044) );
  AND2_X1 U5117 ( .A1(n5698), .A2(n5697), .ZN(n8171) );
  INV_X1 U5118 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U5119 ( .A1(n5021), .A2(n5028), .ZN(n8564) );
  INV_X1 U5120 ( .A(n8653), .ZN(n5025) );
  NAND2_X1 U5121 ( .A1(n8662), .A2(n4446), .ZN(n4598) );
  NAND2_X1 U5122 ( .A1(n8667), .A2(n4477), .ZN(n4532) );
  NAND2_X1 U5123 ( .A1(n5628), .A2(n5627), .ZN(n4652) );
  NAND2_X1 U5124 ( .A1(n5716), .A2(n5717), .ZN(n5721) );
  NAND2_X1 U5125 ( .A1(n4780), .A2(n8073), .ZN(n4779) );
  INV_X1 U5126 ( .A(n5895), .ZN(n4780) );
  OR2_X1 U5127 ( .A1(n9301), .A2(n8752), .ZN(n8833) );
  NAND2_X1 U5128 ( .A1(n5120), .A2(n5119), .ZN(n5123) );
  INV_X1 U5129 ( .A(SI_17_), .ZN(n5119) );
  INV_X1 U5130 ( .A(n4850), .ZN(n4849) );
  INV_X1 U5131 ( .A(n8034), .ZN(n4865) );
  OR2_X1 U5132 ( .A1(n8005), .A2(n8209), .ZN(n5819) );
  INV_X1 U5133 ( .A(n5798), .ZN(n4938) );
  OR2_X1 U5134 ( .A1(n8432), .A2(n7972), .ZN(n5825) );
  OR2_X1 U5135 ( .A1(n8439), .A2(n7906), .ZN(n5795) );
  NAND2_X1 U5136 ( .A1(n4945), .A2(n4944), .ZN(n4943) );
  INV_X1 U5137 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4944) );
  INV_X1 U5138 ( .A(n4946), .ZN(n4945) );
  INV_X2 U5139 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n10121) );
  OR2_X1 U5140 ( .A1(n5527), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5417) );
  NOR2_X1 U5141 ( .A1(n5353), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5364) );
  OR2_X1 U5142 ( .A1(n6113), .A2(n7425), .ZN(n6112) );
  OR2_X1 U5143 ( .A1(n8582), .A2(n4986), .ZN(n4985) );
  INV_X1 U5144 ( .A(n7022), .ZN(n7113) );
  AND2_X1 U5145 ( .A1(n8833), .A2(n8841), .ZN(n9059) );
  INV_X1 U5146 ( .A(n8922), .ZN(n9054) );
  NAND4_X1 U5147 ( .A1(n5038), .A2(n5039), .A3(n4744), .A4(n4481), .ZN(n6015)
         );
  INV_X1 U5148 ( .A(n5974), .ZN(n4745) );
  NAND2_X1 U5149 ( .A1(n5169), .A2(n5168), .ZN(n5687) );
  AND2_X1 U5150 ( .A1(n5176), .A2(n5175), .ZN(n5686) );
  INV_X1 U5151 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5989) );
  AND2_X1 U5152 ( .A1(n5152), .A2(n5151), .ZN(n5630) );
  NAND2_X1 U5153 ( .A1(n5137), .A2(n5136), .ZN(n5604) );
  OAI21_X1 U5154 ( .B1(n5588), .B2(n5585), .A(n5135), .ZN(n5137) );
  OR2_X1 U5155 ( .A1(n6198), .A2(n5989), .ZN(n5990) );
  NAND3_X1 U5156 ( .A1(n5114), .A2(n5115), .A3(n4463), .ZN(n4893) );
  AND2_X1 U5157 ( .A1(n4582), .A2(n5079), .ZN(n4583) );
  INV_X1 U5158 ( .A(n5074), .ZN(n4584) );
  INV_X1 U5159 ( .A(n5355), .ZN(n4585) );
  OAI21_X1 U5161 ( .B1(n4455), .B2(n4828), .A(n4827), .ZN(n4826) );
  AND2_X1 U5162 ( .A1(n7924), .A2(n7957), .ZN(n4828) );
  NAND2_X1 U5163 ( .A1(n4455), .A2(n7957), .ZN(n4827) );
  OR2_X1 U5164 ( .A1(n4847), .A2(n4478), .ZN(n4844) );
  INV_X1 U5165 ( .A(n4848), .ZN(n4847) );
  OAI21_X1 U5166 ( .B1(n4851), .B2(n4849), .A(n8001), .ZN(n4848) );
  NOR2_X1 U5167 ( .A1(n7760), .A2(n4832), .ZN(n4831) );
  NOR2_X1 U5168 ( .A1(n4833), .A2(n4834), .ZN(n4832) );
  AND2_X1 U5169 ( .A1(n5613), .A2(n5612), .ZN(n7912) );
  AND2_X2 U5170 ( .A1(n6701), .A2(n5188), .ZN(n5340) );
  AND2_X1 U5171 ( .A1(n4916), .A2(n4648), .ZN(n4915) );
  OAI21_X1 U5172 ( .B1(n5876), .B2(n6643), .A(n4770), .ZN(n5322) );
  NAND2_X1 U5173 ( .A1(n4767), .A2(n4771), .ZN(n4770) );
  OAI21_X1 U5174 ( .B1(n5198), .B2(P2_IR_REG_27__SCAN_IN), .A(n4768), .ZN(
        n4765) );
  AND2_X1 U5175 ( .A1(n4795), .A2(n4524), .ZN(n4792) );
  AOI21_X1 U5176 ( .B1(n4786), .B2(n4788), .A(n4502), .ZN(n4783) );
  INV_X1 U5177 ( .A(n8328), .ZN(n9860) );
  OR2_X1 U5178 ( .A1(n8216), .A2(n4938), .ZN(n4936) );
  OR2_X1 U5179 ( .A1(n8363), .A2(n8012), .ZN(n5827) );
  OR2_X1 U5180 ( .A1(n5909), .A2(n8284), .ZN(n5046) );
  AND2_X1 U5181 ( .A1(n5792), .A2(n5829), .ZN(n4931) );
  INV_X1 U5182 ( .A(n8331), .ZN(n9867) );
  AOI21_X1 U5183 ( .B1(n4911), .B2(n4914), .A(n4909), .ZN(n4908) );
  INV_X1 U5184 ( .A(n5788), .ZN(n4914) );
  INV_X1 U5185 ( .A(n6711), .ZN(n8118) );
  INV_X1 U5186 ( .A(n4976), .ZN(n4975) );
  OAI21_X1 U5187 ( .B1(n4468), .B2(n4977), .A(n6270), .ZN(n4976) );
  NAND2_X1 U5188 ( .A1(n7412), .A2(n6146), .ZN(n4618) );
  NOR2_X1 U5189 ( .A1(n6426), .A2(n6425), .ZN(n6444) );
  NAND2_X1 U5190 ( .A1(n4963), .A2(n6403), .ZN(n4614) );
  CLKBUF_X1 U5191 ( .A(n6521), .Z(n8900) );
  NAND2_X1 U5192 ( .A1(n4982), .A2(n4468), .ZN(n4974) );
  AOI21_X1 U5193 ( .B1(n4587), .B2(n4586), .A(n8823), .ZN(n8742) );
  INV_X1 U5194 ( .A(n4559), .ZN(n4558) );
  OAI21_X1 U5195 ( .B1(n8753), .B2(n4567), .A(n4560), .ZN(n4559) );
  NAND2_X1 U5196 ( .A1(n4567), .A2(n8770), .ZN(n4560) );
  INV_X1 U5197 ( .A(n8764), .ZN(n6480) );
  INV_X1 U5198 ( .A(n6074), .ZN(n6477) );
  OR2_X1 U5199 ( .A1(n9408), .A2(n9052), .ZN(n5008) );
  INV_X1 U5200 ( .A(n4740), .ZN(n4739) );
  OAI21_X1 U5201 ( .B1(n4742), .B2(n4741), .A(n9280), .ZN(n4740) );
  INV_X1 U5202 ( .A(n8876), .ZN(n4741) );
  AND2_X1 U5203 ( .A1(n8829), .A2(n9070), .ZN(n9088) );
  NOR2_X1 U5204 ( .A1(n4489), .A2(n9261), .ZN(n5030) );
  NAND2_X1 U5205 ( .A1(n6262), .A2(n6261), .ZN(n9375) );
  NAND2_X1 U5206 ( .A1(n5036), .A2(n5034), .ZN(n6996) );
  NAND2_X1 U5207 ( .A1(n6668), .A2(n5035), .ZN(n5034) );
  NAND2_X1 U5208 ( .A1(n4508), .A2(n4450), .ZN(n5035) );
  NAND2_X1 U5209 ( .A1(n7027), .A2(n8910), .ZN(n9278) );
  NAND2_X1 U5210 ( .A1(n4886), .A2(n4488), .ZN(n5471) );
  INV_X1 U5211 ( .A(n5469), .ZN(n4890) );
  NAND2_X1 U5212 ( .A1(n5064), .A2(n5303), .ZN(n5306) );
  AND4_X1 U5213 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5533), .ZN(n8060)
         );
  AND2_X1 U5214 ( .A1(n5761), .A2(n5240), .ZN(n7961) );
  NAND2_X1 U5215 ( .A1(n5448), .A2(n6636), .ZN(n4650) );
  NAND2_X1 U5216 ( .A1(n5447), .A2(n5929), .ZN(n4649) );
  AND2_X1 U5217 ( .A1(n5795), .A2(n5792), .ZN(n4538) );
  INV_X1 U5218 ( .A(n8685), .ZN(n4591) );
  NAND2_X1 U5219 ( .A1(n8684), .A2(n8687), .ZN(n4595) );
  INV_X1 U5220 ( .A(n8704), .ZN(n4574) );
  OR2_X1 U5221 ( .A1(n4579), .A2(n4572), .ZN(n4571) );
  NOR2_X1 U5222 ( .A1(n8709), .A2(n8868), .ZN(n4572) );
  NAND2_X1 U5223 ( .A1(n8878), .A2(n8874), .ZN(n4579) );
  OAI21_X1 U5224 ( .B1(n8720), .B2(n8880), .A(n8719), .ZN(n4600) );
  AND2_X1 U5225 ( .A1(n7658), .A2(n8125), .ZN(n6568) );
  NAND2_X1 U5226 ( .A1(n7114), .A2(n7171), .ZN(n4731) );
  NOR2_X1 U5227 ( .A1(n9370), .A2(n9267), .ZN(n4673) );
  NAND2_X1 U5228 ( .A1(n5490), .A2(SI_14_), .ZN(n4898) );
  NAND2_X1 U5229 ( .A1(n5054), .A2(n9007), .ZN(n4903) );
  INV_X1 U5230 ( .A(n8008), .ZN(n4856) );
  INV_X1 U5231 ( .A(n7932), .ZN(n4813) );
  NAND2_X1 U5232 ( .A1(n6909), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5233 ( .A1(n7240), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U5234 ( .A1(n9717), .A2(n4625), .ZN(n8137) );
  OR2_X1 U5235 ( .A1(n9713), .A2(n10256), .ZN(n4625) );
  OR2_X1 U5236 ( .A1(n9789), .A2(n4703), .ZN(n4702) );
  NOR2_X1 U5237 ( .A1(n9780), .A2(n5500), .ZN(n4703) );
  NOR2_X1 U5238 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5190) );
  NOR2_X1 U5239 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5189) );
  OR2_X1 U5240 ( .A1(n5691), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5705) );
  AND2_X1 U5241 ( .A1(n8048), .A2(n8183), .ZN(n5806) );
  OR2_X1 U5242 ( .A1(n8048), .A2(n8183), .ZN(n5807) );
  OR2_X1 U5243 ( .A1(n8439), .A2(n8277), .ZN(n5910) );
  NOR2_X1 U5244 ( .A1(n5199), .A2(n8473), .ZN(n4772) );
  AOI21_X1 U5245 ( .B1(n4796), .B2(n4798), .A(n4510), .ZN(n4795) );
  OR2_X1 U5246 ( .A1(n7981), .A2(n8194), .ZN(n5803) );
  AND2_X1 U5247 ( .A1(n8414), .A2(n8221), .ZN(n5821) );
  NAND2_X1 U5248 ( .A1(n5195), .A2(n4947), .ZN(n4946) );
  OR2_X1 U5249 ( .A1(n6164), .A2(n7586), .ZN(n4619) );
  INV_X1 U5250 ( .A(n9492), .ZN(n4606) );
  NOR2_X1 U5251 ( .A1(n9332), .A2(n4671), .ZN(n4670) );
  NOR2_X1 U5252 ( .A1(n4671), .A2(n8923), .ZN(n5017) );
  INV_X1 U5253 ( .A(n5018), .ZN(n5013) );
  AND2_X1 U5254 ( .A1(n8839), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U5255 ( .A1(n9249), .A2(n4737), .ZN(n4736) );
  INV_X1 U5256 ( .A(n8837), .ZN(n4737) );
  INV_X1 U5257 ( .A(n9249), .ZN(n4738) );
  AND2_X1 U5258 ( .A1(n4743), .A2(n8707), .ZN(n4742) );
  INV_X1 U5259 ( .A(n8798), .ZN(n4743) );
  INV_X1 U5260 ( .A(n4990), .ZN(n4989) );
  OAI21_X1 U5261 ( .B1(n8677), .B2(n4991), .A(n7528), .ZN(n4990) );
  INV_X1 U5262 ( .A(n7499), .ZN(n4991) );
  NOR2_X1 U5263 ( .A1(n7492), .A2(n9588), .ZN(n4674) );
  INV_X1 U5264 ( .A(n4467), .ZN(n4961) );
  OR2_X1 U5265 ( .A1(n9348), .A2(n9036), .ZN(n9061) );
  OR2_X1 U5266 ( .A1(n9267), .A2(n8714), .ZN(n8837) );
  OR2_X1 U5267 ( .A1(n9370), .A2(n8694), .ZN(n8877) );
  NOR2_X1 U5268 ( .A1(n4997), .A2(n8794), .ZN(n4995) );
  INV_X1 U5269 ( .A(n4997), .ZN(n4994) );
  OR2_X1 U5270 ( .A1(n7738), .A2(n9381), .ZN(n7769) );
  AND2_X1 U5271 ( .A1(n8896), .A2(n6522), .ZN(n7024) );
  AND2_X1 U5272 ( .A1(n5168), .A2(n5167), .ZN(n5673) );
  INV_X1 U5273 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5964) );
  NOR2_X1 U5274 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5969) );
  NAND2_X1 U5275 ( .A1(n4876), .A2(n4874), .ZN(n5645) );
  AOI21_X1 U5276 ( .B1(n4878), .B2(n4881), .A(n4875), .ZN(n4874) );
  INV_X1 U5277 ( .A(n5152), .ZN(n4875) );
  NOR2_X1 U5278 ( .A1(n5616), .A2(n4885), .ZN(n4884) );
  INV_X1 U5279 ( .A(n5139), .ZN(n4885) );
  AOI21_X1 U5280 ( .B1(n4884), .B2(n5140), .A(n4883), .ZN(n4882) );
  INV_X1 U5281 ( .A(n5145), .ZN(n4883) );
  NOR2_X1 U5282 ( .A1(n5540), .A2(n4892), .ZN(n4891) );
  INV_X1 U5283 ( .A(n5118), .ZN(n4892) );
  NAND2_X1 U5284 ( .A1(n4896), .A2(n4894), .ZN(n5113) );
  INV_X1 U5285 ( .A(n4897), .ZN(n4894) );
  INV_X1 U5286 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U5287 ( .A1(n4813), .A2(n7897), .ZN(n4812) );
  AOI21_X1 U5288 ( .B1(n4859), .B2(n4864), .A(n4858), .ZN(n4857) );
  INV_X1 U5289 ( .A(n7949), .ZN(n4858) );
  AND2_X1 U5290 ( .A1(n7744), .A2(n8073), .ZN(n4833) );
  OAI21_X1 U5291 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7743) );
  NAND2_X1 U5292 ( .A1(n4814), .A2(n4442), .ZN(n4819) );
  OAI21_X1 U5293 ( .B1(n4815), .B2(n7095), .A(n7260), .ZN(n4814) );
  NAND2_X1 U5294 ( .A1(n7194), .A2(n4442), .ZN(n4820) );
  NAND2_X1 U5295 ( .A1(n4837), .A2(n4838), .ZN(n7920) );
  AOI21_X1 U5296 ( .B1(n4839), .B2(n4845), .A(n4441), .ZN(n4838) );
  AOI211_X1 U5297 ( .C1(n8391), .C2(n8392), .A(n5855), .B(n5815), .ZN(n5856)
         );
  AND2_X1 U5298 ( .A1(n6701), .A2(n5309), .ZN(n5323) );
  INV_X1 U5299 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U5300 ( .A1(n4688), .A2(n4695), .ZN(n4700) );
  OR2_X1 U5301 ( .A1(n7159), .A2(n4699), .ZN(n4694) );
  NAND2_X1 U5302 ( .A1(n6770), .A2(n4692), .ZN(n4687) );
  NAND2_X1 U5303 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5304 ( .A1(n4688), .A2(n4492), .ZN(n4690) );
  NAND2_X1 U5305 ( .A1(n4624), .A2(n4623), .ZN(n9701) );
  INV_X1 U5306 ( .A(n9697), .ZN(n4623) );
  INV_X1 U5307 ( .A(n9698), .ZN(n4624) );
  NAND2_X1 U5308 ( .A1(n4683), .A2(n7233), .ZN(n4686) );
  INV_X1 U5309 ( .A(n7162), .ZN(n4683) );
  NAND2_X1 U5310 ( .A1(n9701), .A2(n4621), .ZN(n7231) );
  NAND2_X1 U5311 ( .A1(n4622), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5312 ( .A1(n4681), .A2(n4686), .ZN(n4685) );
  INV_X1 U5313 ( .A(n4682), .ZN(n4681) );
  INV_X1 U5314 ( .A(n4685), .ZN(n7243) );
  NAND2_X1 U5315 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  XNOR2_X1 U5316 ( .A(n8137), .B(n9730), .ZN(n9732) );
  NAND2_X1 U5317 ( .A1(n4678), .A2(n4472), .ZN(n4677) );
  AND2_X1 U5318 ( .A1(n4677), .A2(n4676), .ZN(n9756) );
  INV_X1 U5319 ( .A(n9757), .ZN(n4676) );
  NOR2_X1 U5320 ( .A1(n9791), .A2(n9790), .ZN(n9789) );
  XNOR2_X1 U5321 ( .A(n4702), .B(n4701), .ZN(n9807) );
  NOR2_X1 U5322 ( .A1(n9807), .A2(n9806), .ZN(n9805) );
  INV_X1 U5323 ( .A(n8173), .ZN(n8168) );
  NAND2_X1 U5324 ( .A1(n5221), .A2(n10120), .ZN(n5677) );
  INV_X1 U5325 ( .A(n5665), .ZN(n5221) );
  OR2_X1 U5326 ( .A1(n5648), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5665) );
  OR2_X1 U5327 ( .A1(n5634), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5648) );
  OR2_X1 U5328 ( .A1(n5580), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5591) );
  OR2_X1 U5329 ( .A1(n5514), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U5330 ( .A1(n4762), .A2(n4764), .ZN(n4759) );
  INV_X1 U5331 ( .A(n4763), .ZN(n4762) );
  OAI21_X1 U5332 ( .B1(n5769), .B2(n6979), .A(n5768), .ZN(n9851) );
  NAND2_X1 U5333 ( .A1(n4775), .A2(n4774), .ZN(n5896) );
  AND2_X1 U5334 ( .A1(n6636), .A2(n6573), .ZN(n6617) );
  AOI21_X1 U5335 ( .B1(n4935), .B2(n4938), .A(n4934), .ZN(n4933) );
  INV_X1 U5336 ( .A(n4935), .ZN(n4932) );
  OR2_X1 U5337 ( .A1(n8408), .A2(n8209), .ZN(n5045) );
  OR2_X1 U5338 ( .A1(n8005), .A2(n8071), .ZN(n5915) );
  AND2_X1 U5339 ( .A1(n4937), .A2(n5800), .ZN(n4935) );
  INV_X1 U5340 ( .A(n5821), .ZN(n4937) );
  AND2_X1 U5341 ( .A1(n5626), .A2(n5625), .ZN(n8208) );
  INV_X1 U5342 ( .A(n8071), .ZN(n8209) );
  OR2_X1 U5343 ( .A1(n8420), .A2(n8208), .ZN(n5800) );
  INV_X1 U5344 ( .A(n8218), .ZN(n4789) );
  INV_X1 U5345 ( .A(n4787), .ZN(n4786) );
  OAI21_X1 U5346 ( .B1(n4443), .B2(n4788), .A(n8217), .ZN(n4787) );
  AOI21_X1 U5347 ( .B1(n4924), .B2(n4926), .A(n4922), .ZN(n4921) );
  INV_X1 U5348 ( .A(n5822), .ZN(n4922) );
  NAND2_X1 U5349 ( .A1(n4785), .A2(n4790), .ZN(n8228) );
  NAND2_X1 U5350 ( .A1(n8243), .A2(n4443), .ZN(n4785) );
  NOR2_X1 U5351 ( .A1(n5797), .A2(n4928), .ZN(n4927) );
  INV_X1 U5352 ( .A(n5827), .ZN(n4928) );
  AND2_X1 U5353 ( .A1(n4482), .A2(n5793), .ZN(n4929) );
  NAND2_X1 U5354 ( .A1(n4754), .A2(n4755), .ZN(n8274) );
  INV_X1 U5355 ( .A(n4756), .ZN(n4755) );
  OAI21_X1 U5356 ( .B1(n5847), .B2(n4757), .A(n8275), .ZN(n4756) );
  OR2_X1 U5357 ( .A1(n8451), .A2(n8060), .ZN(n5829) );
  NAND2_X1 U5358 ( .A1(n4758), .A2(n5847), .ZN(n8285) );
  INV_X1 U5359 ( .A(n8287), .ZN(n4758) );
  OR2_X1 U5360 ( .A1(n8462), .A2(n7899), .ZN(n5788) );
  NAND2_X1 U5361 ( .A1(n5786), .A2(n5785), .ZN(n8307) );
  AOI21_X1 U5362 ( .B1(n7808), .B2(n5783), .A(n4499), .ZN(n4940) );
  AND2_X1 U5363 ( .A1(n6922), .A2(n5929), .ZN(n8328) );
  INV_X1 U5364 ( .A(n9861), .ZN(n8326) );
  NAND2_X1 U5365 ( .A1(n5924), .A2(n5923), .ZN(n8331) );
  OR2_X1 U5366 ( .A1(n5244), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5864) );
  AOI21_X1 U5367 ( .B1(n5937), .B2(n7871), .A(n7877), .ZN(n6658) );
  XNOR2_X1 U5368 ( .A(n7865), .B(P2_B_REG_SCAN_IN), .ZN(n5937) );
  INV_X1 U5369 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U5370 ( .A1(n5871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4803) );
  AND2_X1 U5371 ( .A1(n5420), .A2(n5434), .ZN(n8133) );
  XNOR2_X1 U5372 ( .A(n5405), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U5373 ( .A1(n4609), .A2(n4608), .ZN(n4607) );
  INV_X1 U5374 ( .A(n6094), .ZN(n6073) );
  NAND2_X1 U5375 ( .A1(n6399), .A2(n6400), .ZN(n4963) );
  AOI21_X1 U5376 ( .B1(n4445), .B2(n4986), .A(n4484), .ZN(n4984) );
  OR2_X1 U5377 ( .A1(n7032), .A2(n7031), .ZN(n6535) );
  AND2_X1 U5378 ( .A1(n8493), .A2(n6285), .ZN(n5020) );
  OAI21_X1 U5379 ( .B1(n8754), .B2(n4565), .A(n4562), .ZN(n4557) );
  NAND2_X1 U5380 ( .A1(n9059), .A2(n4567), .ZN(n4565) );
  INV_X1 U5381 ( .A(n4563), .ZN(n4562) );
  AOI21_X1 U5382 ( .B1(n4558), .B2(n4561), .A(n4509), .ZN(n4555) );
  NAND2_X1 U5383 ( .A1(n9059), .A2(n9009), .ZN(n4561) );
  AOI21_X1 U5384 ( .B1(n6877), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6876), .ZN(
        n6880) );
  AOI21_X1 U5385 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n8987), .A(n9518), .ZN(
        n8977) );
  AND2_X1 U5386 ( .A1(n9540), .A2(n8991), .ZN(n9555) );
  AOI21_X1 U5387 ( .B1(n9549), .B2(n9548), .A(n8979), .ZN(n9559) );
  INV_X1 U5388 ( .A(n4666), .ZN(n4665) );
  NAND2_X1 U5389 ( .A1(n9093), .A2(n4663), .ZN(n4662) );
  NOR2_X1 U5390 ( .A1(n8772), .A2(n4466), .ZN(n4663) );
  OR2_X1 U5391 ( .A1(n9143), .A2(n9318), .ZN(n9121) );
  NOR2_X1 U5392 ( .A1(n9053), .A2(n5010), .ZN(n5007) );
  AND2_X1 U5393 ( .A1(n8828), .A2(n9067), .ZN(n9127) );
  NAND2_X1 U5394 ( .A1(n7815), .A2(n4742), .ZN(n8836) );
  NAND2_X1 U5395 ( .A1(n4447), .A2(n4479), .ZN(n5000) );
  AOI21_X1 U5396 ( .B1(n4724), .B2(n4726), .A(n4722), .ZN(n4721) );
  INV_X1 U5397 ( .A(n4725), .ZN(n4724) );
  NAND2_X1 U5398 ( .A1(n7670), .A2(n8794), .ZN(n7733) );
  NAND2_X1 U5399 ( .A1(n7665), .A2(n7669), .ZN(n7732) );
  OR2_X1 U5400 ( .A1(n7530), .A2(n7486), .ZN(n8683) );
  NAND2_X1 U5401 ( .A1(n7550), .A2(n8677), .ZN(n7549) );
  NAND2_X1 U5402 ( .A1(n4720), .A2(n4719), .ZN(n7483) );
  INV_X1 U5403 ( .A(n8783), .ZN(n4719) );
  INV_X1 U5404 ( .A(n8667), .ZN(n4720) );
  INV_X1 U5405 ( .A(n9278), .ZN(n9215) );
  NAND2_X1 U5406 ( .A1(n7026), .A2(n7025), .ZN(n7115) );
  NOR2_X1 U5407 ( .A1(n9059), .A2(n4961), .ZN(n4960) );
  OAI21_X1 U5408 ( .B1(n9059), .B2(n4959), .A(n4958), .ZN(n4957) );
  NOR2_X1 U5409 ( .A1(n4961), .A2(n4465), .ZN(n4959) );
  NAND2_X1 U5410 ( .A1(n9059), .A2(n4467), .ZN(n4958) );
  NAND2_X1 U5411 ( .A1(n6474), .A2(n6473), .ZN(n9113) );
  AOI21_X1 U5412 ( .B1(n5004), .B2(n5006), .A(n4504), .ZN(n5002) );
  NAND2_X1 U5413 ( .A1(n5019), .A2(n9041), .ZN(n5018) );
  NOR2_X1 U5414 ( .A1(n9043), .A2(n5016), .ZN(n5015) );
  INV_X1 U5415 ( .A(n9039), .ZN(n5016) );
  NOR2_X1 U5416 ( .A1(n5019), .A2(n9041), .ZN(n9043) );
  NOR2_X1 U5417 ( .A1(n9429), .A2(n9032), .ZN(n9034) );
  AND2_X1 U5418 ( .A1(n5032), .A2(n5031), .ZN(n9246) );
  NAND2_X1 U5419 ( .A1(n9267), .A2(n9028), .ZN(n5031) );
  AND2_X1 U5420 ( .A1(n8837), .A2(n8718), .ZN(n9261) );
  OR2_X1 U5421 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  OR2_X1 U5422 ( .A1(n9021), .A2(n9020), .ZN(n5049) );
  AND2_X1 U5423 ( .A1(n8877), .A2(n8878), .ZN(n9280) );
  OR2_X1 U5424 ( .A1(n9276), .A2(n9280), .ZN(n5033) );
  OR2_X1 U5425 ( .A1(n8770), .A2(n8895), .ZN(n9652) );
  XNOR2_X1 U5426 ( .A(n6507), .B(n10032), .ZN(n7840) );
  MUX2_X1 U5427 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6016), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n6017) );
  XNOR2_X1 U5428 ( .A(n6013), .B(n6012), .ZN(n7041) );
  OAI21_X1 U5429 ( .B1(n6004), .B2(n5974), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6013) );
  XNOR2_X1 U5430 ( .A(n5687), .B(n5686), .ZN(n8487) );
  XNOR2_X1 U5431 ( .A(n6005), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U5432 ( .A1(n6006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U5433 ( .A1(n6004), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6008) );
  OAI21_X1 U5434 ( .B1(n5604), .B2(n5140), .A(n5139), .ZN(n5617) );
  INV_X1 U5435 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6318) );
  AND2_X1 U5436 ( .A1(n6286), .A2(n5990), .ZN(n6299) );
  NAND2_X1 U5437 ( .A1(n4893), .A2(n5118), .ZN(n5541) );
  NAND2_X1 U5438 ( .A1(n5251), .A2(n5110), .ZN(n5492) );
  NAND2_X1 U5439 ( .A1(n5249), .A2(n5248), .ZN(n5251) );
  AOI21_X1 U5440 ( .B1(n5430), .B2(n4888), .A(n4511), .ZN(n4887) );
  XNOR2_X1 U5441 ( .A(n5416), .B(n5415), .ZN(n6685) );
  NAND2_X1 U5442 ( .A1(n5388), .A2(n5387), .ZN(n5402) );
  AND2_X1 U5443 ( .A1(n5079), .A2(n5078), .ZN(n5355) );
  NAND2_X1 U5444 ( .A1(n5337), .A2(n5336), .ZN(n5339) );
  AND2_X1 U5445 ( .A1(n4633), .A2(n5069), .ZN(n5319) );
  OR2_X1 U5446 ( .A1(n6047), .A2(n6198), .ZN(n6083) );
  NAND2_X1 U5447 ( .A1(n5062), .A2(n5271), .ZN(n5274) );
  NAND2_X1 U5448 ( .A1(n5936), .A2(n5874), .ZN(n6814) );
  NAND2_X1 U5449 ( .A1(n5579), .A2(n5578), .ZN(n8363) );
  NOR2_X1 U5450 ( .A1(n4448), .A2(n8050), .ZN(n4822) );
  INV_X1 U5451 ( .A(n7957), .ZN(n4825) );
  NAND2_X1 U5452 ( .A1(n4826), .A2(n4829), .ZN(n4824) );
  NAND2_X1 U5453 ( .A1(n4455), .A2(n4830), .ZN(n4829) );
  INV_X1 U5454 ( .A(n7924), .ZN(n4830) );
  NAND2_X1 U5455 ( .A1(n5715), .A2(n5714), .ZN(n7966) );
  AND3_X1 U5456 ( .A1(n5595), .A2(n5594), .A3(n5593), .ZN(n7972) );
  OR2_X1 U5457 ( .A1(n7984), .A2(n8300), .ZN(n7903) );
  AND2_X1 U5458 ( .A1(n7094), .A2(n7093), .ZN(n7096) );
  INV_X1 U5459 ( .A(n8059), .ZN(n8042) );
  INV_X1 U5460 ( .A(n8221), .ZN(n8193) );
  AND4_X1 U5461 ( .A1(n5551), .A2(n5550), .A3(n5549), .A4(n5548), .ZN(n8284)
         );
  NAND2_X1 U5462 ( .A1(n6828), .A2(n9857), .ZN(n8047) );
  NAND2_X1 U5463 ( .A1(n5711), .A2(n5710), .ZN(n8068) );
  INV_X1 U5464 ( .A(n7912), .ZN(n8244) );
  INV_X1 U5465 ( .A(P2_U3893), .ZN(n9475) );
  XNOR2_X1 U5466 ( .A(n7231), .B(n7226), .ZN(n7235) );
  AOI21_X1 U5467 ( .B1(n8152), .B2(n6714), .A(n8151), .ZN(n4628) );
  INV_X1 U5468 ( .A(n8097), .ZN(n4548) );
  NAND2_X1 U5469 ( .A1(n5633), .A2(n5632), .ZN(n8213) );
  INV_X1 U5470 ( .A(n8467), .ZN(n8334) );
  OR2_X1 U5471 ( .A1(n7809), .A2(n7808), .ZN(n8384) );
  NAND2_X1 U5472 ( .A1(n5477), .A2(n5476), .ZN(n8382) );
  OR2_X1 U5473 ( .A1(n6888), .A2(n5473), .ZN(n5477) );
  NOR2_X1 U5474 ( .A1(n6589), .A2(n6588), .ZN(n6590) );
  OR2_X1 U5475 ( .A1(n7882), .A2(n9902), .ZN(n5934) );
  NAND2_X1 U5476 ( .A1(n5513), .A2(n5512), .ZN(n8457) );
  AOI21_X1 U5477 ( .B1(n6129), .B2(n4964), .A(n4969), .ZN(n4968) );
  INV_X1 U5478 ( .A(n8630), .ZN(n4969) );
  OAI22_X1 U5479 ( .A1(n8498), .A2(n6065), .B1(n8693), .B2(n6432), .ZN(n8495)
         );
  INV_X1 U5480 ( .A(n8806), .ZN(n8915) );
  OAI21_X1 U5481 ( .B1(n9161), .B2(n6477), .A(n6431), .ZN(n9048) );
  NAND2_X1 U5482 ( .A1(n6074), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U5483 ( .A1(n6889), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5984) );
  AOI21_X1 U5484 ( .B1(n6877), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6872), .ZN(
        n6875) );
  NAND2_X1 U5485 ( .A1(n9092), .A2(n9091), .ZN(n9309) );
  NAND2_X1 U5486 ( .A1(n6221), .A2(n6220), .ZN(n7730) );
  NOR2_X1 U5487 ( .A1(n9304), .A2(n4713), .ZN(n4712) );
  INV_X1 U5488 ( .A(n9078), .ZN(n4713) );
  NAND2_X1 U5489 ( .A1(n4541), .A2(n4540), .ZN(n5344) );
  NAND2_X1 U5490 ( .A1(n4658), .A2(n4656), .ZN(n5429) );
  NAND2_X1 U5491 ( .A1(n5843), .A2(n5929), .ZN(n4656) );
  INV_X1 U5492 ( .A(n8309), .ZN(n4642) );
  INV_X1 U5493 ( .A(n5485), .ZN(n4646) );
  NAND2_X1 U5494 ( .A1(n4537), .A2(n6636), .ZN(n4536) );
  NAND2_X1 U5495 ( .A1(n5571), .A2(n5929), .ZN(n4539) );
  OR2_X1 U5496 ( .A1(n4594), .A2(n8770), .ZN(n4593) );
  NOR2_X1 U5497 ( .A1(n8709), .A2(n4574), .ZN(n4573) );
  OAI21_X1 U5498 ( .B1(n4601), .B2(n8770), .A(n4599), .ZN(n8727) );
  NAND2_X1 U5499 ( .A1(n6579), .A2(n5929), .ZN(n4870) );
  NAND2_X1 U5500 ( .A1(n5817), .A2(n5247), .ZN(n4871) );
  NOR2_X1 U5501 ( .A1(n4588), .A2(n8741), .ZN(n8743) );
  NAND2_X1 U5502 ( .A1(n5713), .A2(n5712), .ZN(n4866) );
  AOI21_X1 U5503 ( .B1(n4882), .B2(n4880), .A(n4879), .ZN(n4878) );
  INV_X1 U5504 ( .A(n5630), .ZN(n4879) );
  INV_X1 U5505 ( .A(n4884), .ZN(n4880) );
  INV_X1 U5506 ( .A(n4882), .ZN(n4881) );
  INV_X1 U5507 ( .A(n5602), .ZN(n5138) );
  NOR2_X1 U5508 ( .A1(n5490), .A2(SI_14_), .ZN(n4897) );
  INV_X1 U5509 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4905) );
  AND2_X1 U5510 ( .A1(n4905), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U5511 ( .A1(n7658), .A2(n6917), .ZN(n4805) );
  NAND2_X1 U5512 ( .A1(n4808), .A2(n6918), .ZN(n4807) );
  INV_X1 U5513 ( .A(n7977), .ZN(n4840) );
  INV_X1 U5514 ( .A(n4639), .ZN(n4638) );
  OAI21_X1 U5515 ( .B1(n4640), .B2(n6636), .A(n5853), .ZN(n4639) );
  NAND2_X1 U5516 ( .A1(n4638), .A2(n4640), .ZN(n4637) );
  OAI21_X1 U5517 ( .B1(n5722), .B2(n7966), .A(n5042), .ZN(n5723) );
  OAI211_X1 U5518 ( .C1(n4682), .C2(n4680), .A(n4505), .B(n4679), .ZN(n8081)
         );
  NAND2_X1 U5519 ( .A1(n4686), .A2(n7242), .ZN(n4680) );
  AOI21_X1 U5520 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8130), .A(n9722), .ZN(
        n8084) );
  NAND2_X1 U5521 ( .A1(n9748), .A2(n8139), .ZN(n8141) );
  NOR2_X1 U5522 ( .A1(n9747), .A2(n7806), .ZN(n4675) );
  INV_X1 U5523 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U5524 ( .A1(n4918), .A2(n5448), .ZN(n4916) );
  OAI21_X1 U5525 ( .B1(n7596), .B2(n7640), .A(n9897), .ZN(n4782) );
  NAND2_X1 U5526 ( .A1(n9897), .A2(n4657), .ZN(n5843) );
  NAND2_X1 U5527 ( .A1(n4763), .A2(n4496), .ZN(n4761) );
  OAI21_X1 U5528 ( .B1(n7403), .B2(n5839), .A(n5838), .ZN(n7457) );
  NAND2_X1 U5529 ( .A1(n5329), .A2(n5770), .ZN(n5884) );
  AND2_X1 U5530 ( .A1(n4769), .A2(n4660), .ZN(n4768) );
  NAND2_X1 U5531 ( .A1(n5199), .A2(n8473), .ZN(n4769) );
  NAND2_X1 U5532 ( .A1(n7480), .A2(n4657), .ZN(n4777) );
  NAND2_X1 U5533 ( .A1(n4513), .A2(n4779), .ZN(n4774) );
  NAND2_X1 U5534 ( .A1(n9897), .A2(n7640), .ZN(n4776) );
  OR2_X1 U5535 ( .A1(n5919), .A2(n8171), .ZN(n5809) );
  INV_X1 U5536 ( .A(n5801), .ZN(n4934) );
  INV_X1 U5537 ( .A(n4925), .ZN(n4924) );
  OAI21_X1 U5538 ( .B1(n4927), .B2(n4926), .A(n5823), .ZN(n4925) );
  OR2_X1 U5539 ( .A1(n8426), .A2(n7912), .ZN(n5823) );
  INV_X1 U5540 ( .A(n5790), .ZN(n4909) );
  NOR2_X1 U5541 ( .A1(n4913), .A2(n4498), .ZN(n4911) );
  INV_X1 U5542 ( .A(n5789), .ZN(n4913) );
  INV_X1 U5543 ( .A(n5787), .ZN(n4912) );
  NAND2_X1 U5544 ( .A1(n7480), .A2(n7640), .ZN(n5842) );
  INV_X1 U5545 ( .A(n6568), .ZN(n6919) );
  OR2_X1 U5546 ( .A1(n5417), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5418) );
  INV_X1 U5547 ( .A(n4979), .ZN(n4977) );
  NOR2_X1 U5548 ( .A1(n4977), .A2(n4973), .ZN(n4972) );
  INV_X1 U5549 ( .A(n7854), .ZN(n4973) );
  AOI21_X1 U5550 ( .B1(n8603), .B2(n8604), .A(n4980), .ZN(n4979) );
  INV_X1 U5551 ( .A(n6258), .ZN(n4980) );
  NAND2_X1 U5552 ( .A1(n8743), .A2(n8813), .ZN(n4587) );
  NOR2_X1 U5553 ( .A1(n9106), .A2(n8820), .ZN(n4586) );
  NAND2_X1 U5554 ( .A1(n9009), .A2(n8758), .ZN(n4564) );
  AOI21_X1 U5555 ( .B1(n9510), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9505), .ZN(
        n9520) );
  NOR2_X1 U5556 ( .A1(n9301), .A2(n9311), .ZN(n4666) );
  AND2_X1 U5557 ( .A1(n9332), .A2(n8732), .ZN(n9060) );
  AND2_X1 U5558 ( .A1(n9200), .A2(n9062), .ZN(n4750) );
  AND2_X1 U5559 ( .A1(n7821), .A2(n9021), .ZN(n9008) );
  INV_X1 U5560 ( .A(n8867), .ZN(n4726) );
  OAI21_X1 U5561 ( .B1(n8794), .B2(n4726), .A(n8870), .ZN(n4725) );
  NAND2_X1 U5562 ( .A1(n4718), .A2(n7517), .ZN(n8863) );
  NAND2_X1 U5563 ( .A1(n8792), .A2(n8788), .ZN(n8860) );
  NAND2_X1 U5564 ( .A1(n8785), .A2(n4730), .ZN(n4729) );
  INV_X1 U5565 ( .A(n4731), .ZN(n4730) );
  OR2_X1 U5566 ( .A1(n9113), .A2(n9055), .ZN(n8830) );
  NOR2_X1 U5567 ( .A1(n5005), .A2(n4501), .ZN(n5004) );
  NOR2_X1 U5568 ( .A1(n5007), .A2(n5006), .ZN(n5005) );
  INV_X1 U5569 ( .A(n5008), .ZN(n5006) );
  NAND2_X1 U5570 ( .A1(n9008), .A2(n4673), .ZN(n9265) );
  NAND2_X1 U5571 ( .A1(n9008), .A2(n9291), .ZN(n9284) );
  NOR2_X1 U5572 ( .A1(n7353), .A2(n7358), .ZN(n7352) );
  AND2_X1 U5573 ( .A1(n5745), .A2(n5734), .ZN(n5743) );
  INV_X1 U5574 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5973) );
  INV_X1 U5575 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6012) );
  AND2_X1 U5576 ( .A1(n5162), .A2(n5161), .ZN(n5661) );
  INV_X1 U5577 ( .A(SI_20_), .ZN(n5585) );
  INV_X1 U5578 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5116) );
  AOI21_X1 U5579 ( .B1(n4583), .B2(n4585), .A(n5362), .ZN(n4581) );
  INV_X1 U5580 ( .A(n4766), .ZN(n4773) );
  AOI21_X1 U5581 ( .B1(n5198), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_27__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5582 ( .A1(n6963), .A2(n6962), .ZN(n4804) );
  AOI21_X1 U5583 ( .B1(n4863), .B2(n4458), .A(n4451), .ZN(n4862) );
  INV_X1 U5584 ( .A(n8125), .ZN(n8096) );
  NAND2_X1 U5585 ( .A1(n7940), .A2(n8193), .ZN(n4850) );
  OR2_X1 U5586 ( .A1(n7940), .A2(n8193), .ZN(n4851) );
  NAND2_X1 U5587 ( .A1(n8017), .A2(n8018), .ZN(n8016) );
  OR2_X1 U5588 ( .A1(n7744), .A2(n8073), .ZN(n4834) );
  AND2_X1 U5589 ( .A1(n4812), .A2(n4527), .ZN(n4810) );
  NOR2_X1 U5590 ( .A1(n5855), .A2(n6918), .ZN(n4872) );
  AND2_X1 U5591 ( .A1(n5761), .A2(n5760), .ZN(n7433) );
  AND4_X1 U5592 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n7258)
         );
  INV_X1 U5593 ( .A(n5881), .ZN(n6920) );
  NAND2_X1 U5594 ( .A1(n4440), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5286) );
  OR2_X1 U5595 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NAND2_X1 U5596 ( .A1(n6757), .A2(n6756), .ZN(n6760) );
  AND2_X1 U5597 ( .A1(n6760), .A2(n6759), .ZN(n6901) );
  NOR2_X1 U5598 ( .A1(n6901), .A2(n4627), .ZN(n7156) );
  NOR2_X1 U5599 ( .A1(n6905), .A2(n6758), .ZN(n4627) );
  OAI21_X1 U5600 ( .B1(n8135), .B2(n8134), .A(n4626), .ZN(n9719) );
  OR2_X1 U5601 ( .A1(n8132), .A2(n8133), .ZN(n4626) );
  OR3_X1 U5602 ( .A1(n5417), .A2(P2_IR_REG_9__SCAN_IN), .A3(n5256), .ZN(n5451)
         );
  NAND2_X1 U5603 ( .A1(n9731), .A2(n8138), .ZN(n9749) );
  NAND2_X1 U5604 ( .A1(n9749), .A2(n9750), .ZN(n9748) );
  NOR2_X1 U5605 ( .A1(n5451), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U5606 ( .A(n8141), .B(n9764), .ZN(n9766) );
  NOR2_X1 U5607 ( .A1(n9805), .A2(n8090), .ZN(n9824) );
  INV_X1 U5608 ( .A(n4702), .ZN(n8089) );
  INV_X1 U5609 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5185) );
  INV_X1 U5610 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5253) );
  INV_X1 U5611 ( .A(n9482), .ZN(n4711) );
  NAND2_X1 U5612 ( .A1(n4711), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5613 ( .A1(n8093), .A2(n4711), .ZN(n4709) );
  INV_X1 U5614 ( .A(n5677), .ZN(n5223) );
  AND2_X1 U5615 ( .A1(n5684), .A2(n5807), .ZN(n8173) );
  NAND2_X1 U5616 ( .A1(n5220), .A2(n5219), .ZN(n5634) );
  NAND2_X1 U5617 ( .A1(n5218), .A2(n5217), .ZN(n5607) );
  INV_X1 U5618 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U5619 ( .A1(n5216), .A2(n10263), .ZN(n5580) );
  INV_X1 U5620 ( .A(n5563), .ZN(n5216) );
  NAND2_X1 U5621 ( .A1(n5215), .A2(n5214), .ZN(n5546) );
  INV_X1 U5622 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5214) );
  INV_X1 U5623 ( .A(n5531), .ZN(n5215) );
  NAND2_X1 U5624 ( .A1(n5213), .A2(n5212), .ZN(n5514) );
  INV_X1 U5625 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U5626 ( .A1(n5211), .A2(n5210), .ZN(n5498) );
  INV_X1 U5627 ( .A(n5480), .ZN(n5211) );
  NAND2_X1 U5628 ( .A1(n5209), .A2(n5208), .ZN(n5456) );
  INV_X1 U5629 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5208) );
  OR2_X1 U5630 ( .A1(n5456), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U5631 ( .A1(n5207), .A2(n5206), .ZN(n5423) );
  INV_X1 U5632 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5206) );
  INV_X1 U5633 ( .A(n5408), .ZN(n5207) );
  NAND2_X1 U5634 ( .A1(n7609), .A2(n5779), .ZN(n7707) );
  NAND2_X1 U5635 ( .A1(n4782), .A2(n4781), .ZN(n7611) );
  AND4_X1 U5636 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n7598)
         );
  INV_X1 U5637 ( .A(n7650), .ZN(n7705) );
  OR2_X1 U5638 ( .A1(n5394), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5408) );
  AND2_X1 U5639 ( .A1(n7599), .A2(n5444), .ZN(n7462) );
  INV_X1 U5640 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5203) );
  INV_X1 U5641 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5202) );
  NOR2_X1 U5642 ( .A1(n5889), .A2(n9879), .ZN(n4753) );
  AND2_X1 U5643 ( .A1(n5771), .A2(n5767), .ZN(n7071) );
  NAND2_X1 U5644 ( .A1(n7071), .A2(n7069), .ZN(n7068) );
  AND2_X1 U5645 ( .A1(n6571), .A2(n6570), .ZN(n6622) );
  XNOR2_X1 U5646 ( .A(n7966), .B(n6598), .ZN(n7959) );
  NAND2_X1 U5647 ( .A1(n8243), .A2(n8242), .ZN(n8241) );
  AOI21_X1 U5648 ( .B1(n5780), .B2(n7610), .A(n4919), .ZN(n4918) );
  INV_X1 U5649 ( .A(n5831), .ZN(n4919) );
  OR2_X1 U5650 ( .A1(n6636), .A2(n6919), .ZN(n5957) );
  NAND2_X1 U5651 ( .A1(n7775), .A2(n9853), .ZN(n9902) );
  NAND2_X1 U5652 ( .A1(n4942), .A2(n5199), .ZN(n4941) );
  INV_X1 U5653 ( .A(n4943), .ZN(n4942) );
  NAND2_X1 U5654 ( .A1(n5868), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5869) );
  OR2_X1 U5655 ( .A1(n5871), .A2(n4946), .ZN(n5868) );
  INV_X1 U5656 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5764) );
  INV_X1 U5657 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U5658 ( .A1(n8473), .A2(n5309), .ZN(n4704) );
  INV_X1 U5659 ( .A(n5323), .ZN(n4706) );
  NAND2_X1 U5660 ( .A1(n5308), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5661 ( .A1(n4966), .A2(n6112), .ZN(n4970) );
  INV_X1 U5662 ( .A(n6100), .ZN(n4966) );
  INV_X1 U5663 ( .A(n6112), .ZN(n4964) );
  NAND2_X1 U5664 ( .A1(n4614), .A2(n6404), .ZN(n8504) );
  XNOR2_X1 U5665 ( .A(n6025), .B(n6497), .ZN(n6026) );
  NAND2_X1 U5666 ( .A1(n4603), .A2(n6996), .ZN(n6023) );
  NAND2_X1 U5667 ( .A1(n8581), .A2(n8582), .ZN(n8580) );
  NAND2_X1 U5668 ( .A1(n4462), .A2(n4617), .ZN(n4615) );
  NAND2_X1 U5669 ( .A1(n4620), .A2(n4494), .ZN(n4616) );
  NAND2_X1 U5670 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  AOI21_X1 U5671 ( .B1(n8936), .B2(n6499), .A(n6040), .ZN(n6942) );
  OAI21_X1 U5672 ( .B1(n8851), .B2(n6065), .A(n6039), .ZN(n6040) );
  AND2_X1 U5673 ( .A1(n6350), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6372) );
  INV_X1 U5674 ( .A(n6360), .ZN(n8535) );
  AND2_X1 U5675 ( .A1(n6101), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6118) );
  AND2_X1 U5676 ( .A1(n6118), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6136) );
  NOR4_X1 U5677 ( .A1(n8807), .A2(n8806), .A3(n8893), .A4(n8805), .ZN(n8849)
         );
  INV_X1 U5678 ( .A(n4460), .ZN(n6304) );
  AOI21_X1 U5679 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7139), .A(n7130), .ZN(
        n7133) );
  AOI21_X1 U5680 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9510), .A(n9502), .ZN(
        n9515) );
  AOI21_X1 U5681 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8987), .A(n9514), .ZN(
        n8988) );
  OR2_X1 U5682 ( .A1(n9544), .A2(n9543), .ZN(n9540) );
  INV_X1 U5683 ( .A(n8921), .ZN(n9055) );
  NAND2_X1 U5684 ( .A1(n9104), .A2(n9069), .ZN(n9089) );
  NOR2_X1 U5685 ( .A1(n4669), .A2(n9408), .ZN(n4667) );
  OAI21_X1 U5686 ( .B1(n9201), .B2(n4748), .A(n4746), .ZN(n9175) );
  INV_X1 U5687 ( .A(n4749), .ZN(n4748) );
  AOI21_X1 U5688 ( .B1(n4749), .B2(n4747), .A(n8733), .ZN(n4746) );
  NOR2_X1 U5689 ( .A1(n4751), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U5690 ( .A1(n9190), .A2(n9196), .ZN(n9191) );
  NAND2_X1 U5691 ( .A1(n9190), .A2(n4670), .ZN(n9169) );
  NAND2_X1 U5692 ( .A1(n5012), .A2(n5011), .ZN(n9168) );
  NAND2_X1 U5693 ( .A1(n4512), .A2(n4444), .ZN(n5011) );
  NAND2_X1 U5694 ( .A1(n9040), .A2(n4486), .ZN(n5012) );
  AND2_X1 U5695 ( .A1(n8773), .A2(n9155), .ZN(n9176) );
  NAND2_X1 U5696 ( .A1(n6372), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6391) );
  AOI21_X1 U5697 ( .B1(n4735), .B2(n4738), .A(n4734), .ZN(n4733) );
  INV_X1 U5698 ( .A(n8883), .ZN(n4734) );
  OR2_X1 U5699 ( .A1(n9358), .A2(n9030), .ZN(n9228) );
  OR2_X1 U5700 ( .A1(n6324), .A2(n8622), .ZN(n6349) );
  INV_X1 U5701 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U5702 ( .A1(n9260), .A2(n8837), .ZN(n9248) );
  NAND2_X1 U5703 ( .A1(n9248), .A2(n9249), .ZN(n9247) );
  NAND2_X1 U5704 ( .A1(n9262), .A2(n9261), .ZN(n9260) );
  INV_X1 U5705 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6289) );
  NOR2_X1 U5706 ( .A1(n6290), .A2(n6289), .ZN(n6302) );
  INV_X1 U5707 ( .A(n9024), .ZN(n9021) );
  NOR2_X1 U5708 ( .A1(n7769), .A2(n9375), .ZN(n7821) );
  OR2_X1 U5709 ( .A1(n6263), .A2(n8496), .ZN(n6278) );
  AND2_X1 U5710 ( .A1(n7575), .A2(n7544), .ZN(n7633) );
  AND2_X1 U5711 ( .A1(n7633), .A2(n9655), .ZN(n7676) );
  INV_X1 U5712 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6186) );
  OR2_X1 U5713 ( .A1(n7522), .A2(n8787), .ZN(n7668) );
  NAND2_X1 U5714 ( .A1(n4988), .A2(n4987), .ZN(n7568) );
  AOI21_X1 U5715 ( .B1(n4989), .B2(n4991), .A(n4497), .ZN(n4987) );
  NAND2_X1 U5716 ( .A1(n4674), .A2(n9646), .ZN(n7573) );
  NOR2_X1 U5717 ( .A1(n7573), .A2(n7687), .ZN(n7575) );
  INV_X1 U5718 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6154) );
  INV_X1 U5719 ( .A(n4674), .ZN(n7557) );
  NAND2_X1 U5720 ( .A1(n7276), .A2(n7275), .ZN(n7354) );
  OR2_X1 U5721 ( .A1(n7173), .A2(n8778), .ZN(n7276) );
  OR2_X1 U5722 ( .A1(n6345), .A2(n6541), .ZN(n7632) );
  INV_X1 U5723 ( .A(n8785), .ZN(n7026) );
  NAND2_X1 U5724 ( .A1(n8936), .A2(n7083), .ZN(n7082) );
  CLKBUF_X1 U5725 ( .A(n7023), .Z(n8785) );
  AND2_X1 U5726 ( .A1(n6944), .A2(n9638), .ZN(n7078) );
  NAND2_X1 U5727 ( .A1(n9059), .A2(n4465), .ZN(n4962) );
  AND2_X1 U5728 ( .A1(n9013), .A2(n9075), .ZN(n9298) );
  NAND2_X1 U5729 ( .A1(n6456), .A2(n6455), .ZN(n9318) );
  NAND2_X1 U5730 ( .A1(n6301), .A2(n6300), .ZN(n9267) );
  NAND2_X1 U5731 ( .A1(n4994), .A2(n4500), .ZN(n4993) );
  NAND2_X1 U5732 ( .A1(n6242), .A2(n6241), .ZN(n9381) );
  INV_X1 U5733 ( .A(n9286), .ZN(n9333) );
  OAI21_X1 U5734 ( .B1(n9610), .B2(P1_D_REG_0__SCAN_IN), .A(n6505), .ZN(n7077)
         );
  XNOR2_X1 U5735 ( .A(n5744), .B(n5743), .ZN(n8755) );
  NAND2_X1 U5736 ( .A1(n5980), .A2(n9453), .ZN(n5982) );
  XNOR2_X1 U5737 ( .A(n5713), .B(n5712), .ZN(n8484) );
  XNOR2_X1 U5738 ( .A(n5674), .B(n5673), .ZN(n7875) );
  NOR2_X1 U5739 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5970) );
  NAND2_X1 U5740 ( .A1(n4877), .A2(n4882), .ZN(n5631) );
  NAND2_X1 U5741 ( .A1(n5604), .A2(n4884), .ZN(n4877) );
  INV_X1 U5742 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5988) );
  INV_X1 U5743 ( .A(n5113), .ZN(n5507) );
  NAND2_X1 U5744 ( .A1(n5471), .A2(n5105), .ZN(n5249) );
  NAND2_X1 U5745 ( .A1(n5433), .A2(n5102), .ZN(n5450) );
  AND2_X1 U5746 ( .A1(n6182), .A2(n6181), .ZN(n6218) );
  XNOR2_X1 U5747 ( .A(n5404), .B(n5403), .ZN(n6680) );
  CLKBUF_X1 U5748 ( .A(n6132), .Z(n6133) );
  INV_X1 U5749 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4716) );
  OAI21_X1 U5750 ( .B1(n5339), .B2(n4585), .A(n4583), .ZN(n5363) );
  NAND2_X1 U5751 ( .A1(n5274), .A2(n5063), .ZN(n5303) );
  NAND2_X1 U5752 ( .A1(n5059), .A2(n5063), .ZN(n5272) );
  NAND2_X1 U5753 ( .A1(n5060), .A2(n5061), .ZN(n4554) );
  OR2_X1 U5754 ( .A1(n7925), .A2(n7924), .ZN(n7958) );
  NAND2_X1 U5755 ( .A1(n4811), .A2(n4812), .ZN(n7934) );
  NAND2_X1 U5756 ( .A1(n5437), .A2(n5436), .ZN(n7653) );
  NAND2_X1 U5757 ( .A1(n4861), .A2(n4862), .ZN(n7951) );
  NAND2_X1 U5758 ( .A1(n7994), .A2(n4863), .ZN(n4861) );
  AOI21_X1 U5759 ( .B1(n4507), .B2(n4857), .A(n4854), .ZN(n4853) );
  NOR2_X1 U5760 ( .A1(n7910), .A2(n8252), .ZN(n4854) );
  NAND2_X1 U5761 ( .A1(n7760), .A2(n8072), .ZN(n4835) );
  NAND2_X1 U5762 ( .A1(n4841), .A2(n4844), .ZN(n7976) );
  NAND2_X1 U5763 ( .A1(n4843), .A2(n4842), .ZN(n4841) );
  INV_X1 U5764 ( .A(n7942), .ZN(n4843) );
  NAND2_X1 U5765 ( .A1(n7195), .A2(n7194), .ZN(n7261) );
  NAND2_X1 U5766 ( .A1(n4846), .A2(n4850), .ZN(n8000) );
  NAND2_X1 U5767 ( .A1(n7942), .A2(n4851), .ZN(n4846) );
  NAND2_X1 U5768 ( .A1(n5647), .A2(n5646), .ZN(n8005) );
  AND3_X1 U5769 ( .A1(n5584), .A2(n5583), .A3(n5582), .ZN(n8012) );
  NAND2_X1 U5770 ( .A1(n4852), .A2(n4857), .ZN(n8009) );
  OR2_X1 U5771 ( .A1(n7994), .A2(n4860), .ZN(n4852) );
  OR2_X1 U5772 ( .A1(n6924), .A2(n6826), .ZN(n8059) );
  INV_X1 U5773 ( .A(n9852), .ZN(n6935) );
  AOI21_X1 U5774 ( .B1(n7994), .B2(n7993), .A(n4458), .ZN(n8035) );
  NAND2_X1 U5775 ( .A1(n4819), .A2(n4820), .ZN(n4817) );
  NAND2_X1 U5776 ( .A1(n4816), .A2(n4819), .ZN(n7263) );
  OR2_X1 U5777 ( .A1(n7096), .A2(n4820), .ZN(n4816) );
  AOI21_X1 U5778 ( .B1(n8185), .B2(n5288), .A(n5670), .ZN(n8194) );
  NAND2_X1 U5779 ( .A1(n4811), .A2(n4809), .ZN(n8053) );
  AND2_X1 U5780 ( .A1(n4810), .A2(n8054), .ZN(n4809) );
  AND2_X1 U5781 ( .A1(n4811), .A2(n4810), .ZN(n8055) );
  NAND2_X1 U5782 ( .A1(n6824), .A2(n6823), .ZN(n8062) );
  XNOR2_X1 U5783 ( .A(n5243), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6572) );
  INV_X1 U5784 ( .A(n7433), .ZN(n8154) );
  INV_X1 U5785 ( .A(n8171), .ZN(n8069) );
  NAND2_X1 U5786 ( .A1(n5654), .A2(n5653), .ZN(n8071) );
  INV_X1 U5787 ( .A(n8208), .ZN(n8233) );
  CLKBUF_X1 U5788 ( .A(n6920), .Z(n8079) );
  NOR2_X2 U5789 ( .A1(n5325), .A2(n5340), .ZN(n9684) );
  NAND2_X1 U5790 ( .A1(n4700), .A2(n4692), .ZN(n4691) );
  XNOR2_X1 U5791 ( .A(n7156), .B(n4697), .ZN(n7158) );
  NAND2_X1 U5792 ( .A1(n4696), .A2(n4689), .ZN(n9693) );
  OAI211_X1 U5793 ( .C1(n4688), .C2(n4693), .A(n4690), .B(n4452), .ZN(n4689)
         );
  NAND2_X1 U5794 ( .A1(n4686), .A2(n7240), .ZN(n7163) );
  OAI22_X1 U5795 ( .A1(n7232), .A2(n7233), .B1(n7235), .B2(n7234), .ZN(n7236)
         );
  NAND2_X1 U5796 ( .A1(n4684), .A2(n7242), .ZN(n7337) );
  INV_X1 U5797 ( .A(n4678), .ZN(n9742) );
  INV_X1 U5798 ( .A(n4677), .ZN(n9758) );
  NOR2_X1 U5799 ( .A1(n4707), .A2(n9481), .ZN(n9483) );
  NOR2_X1 U5800 ( .A1(n9841), .A2(n4708), .ZN(n4707) );
  OR2_X1 U5801 ( .A1(n8093), .A2(n4711), .ZN(n4708) );
  INV_X1 U5802 ( .A(n8149), .ZN(n4632) );
  AND2_X1 U5803 ( .A1(n5690), .A2(n5689), .ZN(n8163) );
  INV_X1 U5804 ( .A(n6599), .ZN(n6600) );
  OAI22_X1 U5805 ( .A1(n6598), .A2(n9861), .B1(n9860), .B2(n8183), .ZN(n6599)
         );
  OR2_X1 U5806 ( .A1(n9909), .A2(n9853), .ZN(n8333) );
  INV_X1 U5807 ( .A(n7653), .ZN(n9910) );
  NAND2_X1 U5808 ( .A1(n5422), .A2(n5421), .ZN(n9906) );
  INV_X1 U5809 ( .A(n8318), .ZN(n9871) );
  AND3_X2 U5810 ( .A1(n5280), .A2(n5281), .A3(n5279), .ZN(n7002) );
  NAND2_X1 U5811 ( .A1(n8318), .A2(n6627), .ZN(n8339) );
  INV_X1 U5812 ( .A(n8176), .ZN(n8304) );
  OR2_X1 U5813 ( .A1(n6628), .A2(n8333), .ZN(n8176) );
  INV_X1 U5814 ( .A(n8163), .ZN(n5919) );
  INV_X1 U5815 ( .A(n8005), .ZN(n8408) );
  NAND2_X1 U5816 ( .A1(n4936), .A2(n4935), .ZN(n8198) );
  INV_X1 U5817 ( .A(n8213), .ZN(n8414) );
  NAND2_X1 U5818 ( .A1(n4936), .A2(n5800), .ZN(n8204) );
  NAND2_X1 U5819 ( .A1(n5619), .A2(n5618), .ZN(n8420) );
  OAI21_X1 U5820 ( .B1(n8243), .B2(n4788), .A(n4786), .ZN(n8220) );
  NAND2_X1 U5821 ( .A1(n4923), .A2(n5824), .ZN(n8227) );
  NAND2_X1 U5822 ( .A1(n5796), .A2(n4927), .ZN(n4923) );
  NAND2_X1 U5823 ( .A1(n5590), .A2(n5589), .ZN(n8432) );
  NAND2_X1 U5824 ( .A1(n5562), .A2(n5561), .ZN(n8439) );
  AND2_X1 U5825 ( .A1(n4930), .A2(n5793), .ZN(n8263) );
  NAND2_X1 U5826 ( .A1(n5545), .A2(n5544), .ZN(n8445) );
  NAND2_X1 U5827 ( .A1(n8285), .A2(n5908), .ZN(n8276) );
  NAND2_X1 U5828 ( .A1(n5791), .A2(n5829), .ZN(n8273) );
  NAND2_X1 U5829 ( .A1(n5530), .A2(n5529), .ZN(n8451) );
  NAND2_X1 U5830 ( .A1(n4910), .A2(n5788), .ZN(n8297) );
  NAND2_X1 U5831 ( .A1(n8307), .A2(n5787), .ZN(n4910) );
  NAND2_X1 U5832 ( .A1(n5497), .A2(n5496), .ZN(n8462) );
  NAND2_X1 U5833 ( .A1(n5260), .A2(n5259), .ZN(n8467) );
  OR2_X1 U5834 ( .A1(n6977), .A2(n5473), .ZN(n5260) );
  NAND2_X1 U5835 ( .A1(n8384), .A2(n5783), .ZN(n8323) );
  OAI21_X1 U5836 ( .B1(n5864), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U5837 ( .A1(n4802), .A2(n4801), .ZN(n5872) );
  NAND2_X1 U5838 ( .A1(n4947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4801) );
  NAND2_X1 U5839 ( .A1(n4803), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n4802) );
  AND2_X1 U5840 ( .A1(P2_U3151), .A2(n6640), .ZN(n8489) );
  INV_X1 U5841 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7776) );
  INV_X1 U5842 ( .A(n6572), .ZN(n7775) );
  INV_X1 U5843 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10029) );
  INV_X1 U5844 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7584) );
  INV_X1 U5845 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10138) );
  INV_X1 U5846 ( .A(n9813), .ZN(n8126) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10282) );
  INV_X1 U5848 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6686) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10071) );
  OR2_X1 U5850 ( .A1(n6021), .A2(n6635), .ZN(n6665) );
  NAND2_X1 U5851 ( .A1(n4607), .A2(n6197), .ZN(n9491) );
  XNOR2_X1 U5852 ( .A(n4620), .B(n6164), .ZN(n7587) );
  OR2_X1 U5853 ( .A1(n6457), .A2(n6445), .ZN(n9146) );
  AND2_X1 U5854 ( .A1(n8574), .A2(n8572), .ZN(n6313) );
  AND2_X1 U5855 ( .A1(n7252), .A2(n7250), .ZN(n6096) );
  NAND2_X1 U5856 ( .A1(n6334), .A2(n6333), .ZN(n9348) );
  OAI21_X1 U5857 ( .B1(n4982), .B2(n8604), .A(n4530), .ZN(n8602) );
  NAND2_X1 U5858 ( .A1(n7853), .A2(n6237), .ZN(n4978) );
  INV_X1 U5859 ( .A(n4614), .ZN(n4613) );
  OAI211_X1 U5860 ( .C1(n6238), .C2(n6647), .A(n6050), .B(n6049), .ZN(n7112)
         );
  OR2_X1 U5861 ( .A1(n6668), .A2(n6048), .ZN(n6049) );
  AND2_X1 U5862 ( .A1(n6329), .A2(n6328), .ZN(n8620) );
  AND2_X1 U5863 ( .A1(n6544), .A2(n6945), .ZN(n9501) );
  NAND2_X1 U5864 ( .A1(n4983), .A2(n4984), .ZN(n8643) );
  NAND2_X1 U5865 ( .A1(n6537), .A2(n6536), .ZN(n9489) );
  NAND2_X1 U5866 ( .A1(n5026), .A2(n5028), .ZN(n8654) );
  NAND2_X1 U5867 ( .A1(n4556), .A2(n4555), .ZN(n4566) );
  NAND2_X1 U5868 ( .A1(n8754), .A2(n4558), .ZN(n4556) );
  OR2_X1 U5869 ( .A1(n9123), .A2(n6477), .ZN(n6463) );
  NAND2_X1 U5870 ( .A1(n6412), .A2(n6411), .ZN(n9045) );
  CLKBUF_X2 U5871 ( .A(P1_U3973), .Z(n8935) );
  AOI21_X1 U5872 ( .B1(n6802), .B2(P1_REG1_REG_4__SCAN_IN), .A(n8968), .ZN(
        n6805) );
  AOI21_X1 U5873 ( .B1(n6802), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6790), .ZN(
        n6794) );
  AOI21_X1 U5874 ( .B1(n6838), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6837), .ZN(
        n6864) );
  AOI21_X1 U5875 ( .B1(n6838), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6832), .ZN(
        n6861) );
  AOI21_X1 U5876 ( .B1(n6852), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6849), .ZN(
        n6841) );
  AOI21_X1 U5877 ( .B1(n6852), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6846), .ZN(
        n6836) );
  AOI21_X1 U5878 ( .B1(n7012), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7011), .ZN(
        n7015) );
  AOI21_X1 U5879 ( .B1(n7012), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7006), .ZN(
        n7010) );
  AOI21_X1 U5880 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7139), .A(n7138), .ZN(
        n7143) );
  NOR2_X1 U5881 ( .A1(n9529), .A2(n8978), .ZN(n9549) );
  AND2_X1 U5882 ( .A1(n9554), .A2(n8994), .ZN(n9573) );
  NOR2_X1 U5883 ( .A1(n9010), .A2(n9286), .ZN(n9295) );
  NAND2_X1 U5884 ( .A1(n8772), .A2(n4466), .ZN(n4661) );
  NAND2_X1 U5885 ( .A1(n4954), .A2(n9606), .ZN(n4951) );
  NAND2_X1 U5886 ( .A1(n4957), .A2(n4962), .ZN(n4954) );
  NOR2_X1 U5887 ( .A1(n4955), .A2(n9294), .ZN(n4949) );
  INV_X1 U5888 ( .A(n4960), .ZN(n4956) );
  INV_X1 U5889 ( .A(n9318), .ZN(n9126) );
  NAND2_X1 U5890 ( .A1(n5003), .A2(n5008), .ZN(n9120) );
  NAND2_X1 U5891 ( .A1(n9049), .A2(n5007), .ZN(n5003) );
  NAND2_X1 U5892 ( .A1(n8836), .A2(n8876), .ZN(n9281) );
  NAND2_X1 U5893 ( .A1(n7815), .A2(n8707), .ZN(n7816) );
  NAND2_X1 U5894 ( .A1(n7732), .A2(n4469), .ZN(n4996) );
  NAND2_X1 U5895 ( .A1(n7733), .A2(n8867), .ZN(n7765) );
  NAND2_X1 U5896 ( .A1(n7732), .A2(n7731), .ZN(n7764) );
  NAND2_X1 U5897 ( .A1(n7549), .A2(n7499), .ZN(n7529) );
  NAND2_X1 U5898 ( .A1(n7483), .A2(n8856), .ZN(n7518) );
  INV_X1 U5899 ( .A(n9587), .ZN(n9602) );
  NAND2_X1 U5900 ( .A1(n7115), .A2(n7114), .ZN(n7172) );
  INV_X1 U5901 ( .A(n9241), .ZN(n9596) );
  OR2_X1 U5902 ( .A1(n9652), .A2(n6526), .ZN(n9236) );
  NAND2_X1 U5903 ( .A1(n4602), .A2(n6135), .ZN(n9588) );
  OR2_X1 U5904 ( .A1(n6679), .A2(n6238), .ZN(n4602) );
  OR2_X1 U5905 ( .A1(n7121), .A2(n7077), .ZN(n9665) );
  INV_X1 U5906 ( .A(n9113), .ZN(n9404) );
  NAND2_X1 U5907 ( .A1(n9049), .A2(n5009), .ZN(n9135) );
  NAND2_X1 U5908 ( .A1(n5014), .A2(n5018), .ZN(n9184) );
  NAND2_X1 U5909 ( .A1(n9040), .A2(n5015), .ZN(n5014) );
  AND2_X1 U5910 ( .A1(n5033), .A2(n4456), .ZN(n9259) );
  INV_X1 U5911 ( .A(n8670), .ZN(n8668) );
  INV_X1 U5912 ( .A(n6996), .ZN(n8850) );
  OR2_X1 U5913 ( .A1(n5979), .A2(n6198), .ZN(n5977) );
  INV_X1 U5914 ( .A(n5982), .ZN(n7889) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10111) );
  OR2_X1 U5916 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  INV_X1 U5917 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10193) );
  INV_X1 U5918 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10201) );
  AND2_X1 U5919 ( .A1(n6286), .A2(n4473), .ZN(n6319) );
  INV_X1 U5920 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U5921 ( .A1(n4886), .A2(n4887), .ZN(n5470) );
  AND2_X1 U5922 ( .A1(n6151), .A2(n6165), .ZN(n6877) );
  OAI21_X1 U5923 ( .B1(n5388), .B2(n5387), .A(n5402), .ZN(n6679) );
  NAND2_X1 U5924 ( .A1(n5355), .A2(n5356), .ZN(n5358) );
  NAND2_X1 U5925 ( .A1(n5339), .A2(n5074), .ZN(n5356) );
  NAND2_X1 U5926 ( .A1(n4551), .A2(n4550), .ZN(n5320) );
  NAND2_X1 U5927 ( .A1(n4824), .A2(n8052), .ZN(n4823) );
  NAND2_X1 U5928 ( .A1(n4631), .A2(n9839), .ZN(n4630) );
  XNOR2_X1 U5929 ( .A(n8150), .B(n4632), .ZN(n4631) );
  AOI21_X1 U5930 ( .B1(n9927), .B2(P2_REG1_REG_29__SCAN_IN), .A(n5047), .ZN(
        n6580) );
  AND2_X1 U5931 ( .A1(n6585), .A2(n6584), .ZN(n6593) );
  INV_X1 U5932 ( .A(n8346), .ZN(n4543) );
  INV_X1 U5933 ( .A(n8400), .ZN(n4545) );
  OR2_X1 U5934 ( .A1(n9398), .A2(n9372), .ZN(n4534) );
  NAND2_X1 U5935 ( .A1(n4715), .A2(n4493), .ZN(P1_U3519) );
  OR2_X1 U5936 ( .A1(n9393), .A2(n9661), .ZN(n4715) );
  OR2_X1 U5937 ( .A1(n9439), .A2(n10044), .ZN(n4714) );
  OR2_X1 U5938 ( .A1(n9398), .A2(n9449), .ZN(n4535) );
  AND2_X1 U5939 ( .A1(n7916), .A2(n8194), .ZN(n4441) );
  NAND2_X1 U5940 ( .A1(n4790), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U5941 ( .A1(n7259), .A2(n7258), .ZN(n4442) );
  AND2_X1 U5942 ( .A1(n4791), .A2(n8242), .ZN(n4443) );
  INV_X1 U5943 ( .A(n7159), .ZN(n4697) );
  OR2_X1 U5944 ( .A1(n9196), .A2(n9044), .ZN(n4444) );
  AND2_X1 U5945 ( .A1(n8556), .A2(n4985), .ZN(n4445) );
  INV_X1 U5946 ( .A(n8868), .ZN(n4722) );
  AND4_X1 U5947 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8770), .ZN(n4446)
         );
  OR2_X1 U5948 ( .A1(n9381), .A2(n8925), .ZN(n4447) );
  INV_X1 U5949 ( .A(n9062), .ZN(n4747) );
  NAND2_X1 U5950 ( .A1(n4963), .A2(n6404), .ZN(n8613) );
  INV_X1 U5951 ( .A(n4461), .ZN(n4640) );
  NAND2_X1 U5952 ( .A1(n4983), .A2(n4483), .ZN(n8645) );
  AND2_X1 U5953 ( .A1(n4826), .A2(n4487), .ZN(n4448) );
  INV_X1 U5954 ( .A(n4798), .ZN(n4797) );
  NOR2_X1 U5955 ( .A1(n7981), .A2(n4799), .ZN(n4798) );
  INV_X1 U5956 ( .A(n9408), .ZN(n9144) );
  NAND2_X1 U5957 ( .A1(n6443), .A2(n6442), .ZN(n9408) );
  AND2_X1 U5958 ( .A1(n4694), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5959 ( .A1(n6643), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4450) );
  AND2_X1 U5960 ( .A1(n7907), .A2(n7906), .ZN(n4451) );
  AND2_X1 U5961 ( .A1(n4687), .A2(n4449), .ZN(n4452) );
  AND2_X1 U5962 ( .A1(n4673), .A2(n4672), .ZN(n4453) );
  AND2_X1 U5963 ( .A1(n4813), .A2(n8018), .ZN(n4454) );
  AND2_X1 U5964 ( .A1(n5683), .A2(n5682), .ZN(n8183) );
  INV_X1 U5965 ( .A(n8194), .ZN(n4799) );
  NAND2_X1 U5966 ( .A1(n5940), .A2(n5939), .ZN(n4806) );
  XNOR2_X1 U5967 ( .A(n7960), .B(n7959), .ZN(n4455) );
  INV_X1 U5968 ( .A(n4603), .ZN(n6397) );
  NAND2_X1 U5969 ( .A1(n9370), .A2(n9027), .ZN(n4456) );
  OAI211_X1 U5970 ( .C1(n4807), .C2(n4806), .A(n6919), .B(n4805), .ZN(n6966)
         );
  OR2_X1 U5971 ( .A1(n5871), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n4457) );
  AND2_X1 U5972 ( .A1(n7905), .A2(n8284), .ZN(n4458) );
  OR2_X1 U5973 ( .A1(n6273), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4459) );
  INV_X1 U5974 ( .A(n6966), .ZN(n7504) );
  INV_X2 U5975 ( .A(n7504), .ZN(n7960) );
  AND2_X1 U5976 ( .A1(n5982), .A2(n5981), .ZN(n4460) );
  OR2_X1 U5977 ( .A1(n8392), .A2(n5742), .ZN(n4461) );
  AND2_X1 U5978 ( .A1(n6164), .A2(n7586), .ZN(n4462) );
  OR2_X1 U5979 ( .A1(n5117), .A2(SI_16_), .ZN(n4463) );
  AND2_X1 U5980 ( .A1(n9190), .A2(n4668), .ZN(n4464) );
  OR2_X1 U5981 ( .A1(n9311), .A2(n9077), .ZN(n4465) );
  OR2_X1 U5982 ( .A1(n4665), .A2(n9009), .ZN(n4466) );
  OR2_X1 U5983 ( .A1(n9099), .A2(n9058), .ZN(n4467) );
  NAND2_X1 U5984 ( .A1(n5664), .A2(n5663), .ZN(n7981) );
  AND2_X1 U5985 ( .A1(n8603), .A2(n4981), .ZN(n4468) );
  NAND2_X1 U5986 ( .A1(n6504), .A2(n6010), .ZN(n6021) );
  AND2_X1 U5987 ( .A1(n4447), .A2(n7731), .ZN(n4469) );
  OR2_X1 U5988 ( .A1(n6521), .A2(n8911), .ZN(n4470) );
  XNOR2_X1 U5989 ( .A(n5977), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5981) );
  AND4_X1 U5990 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(n7640)
         );
  AND2_X1 U5991 ( .A1(n5832), .A2(n7706), .ZN(n5780) );
  NAND2_X1 U5992 ( .A1(n8757), .A2(n8756), .ZN(n9009) );
  OR2_X1 U5993 ( .A1(n9906), .A2(n7650), .ZN(n4471) );
  OR2_X1 U5994 ( .A1(n9730), .A2(n8084), .ZN(n4472) );
  NAND2_X1 U5995 ( .A1(n8580), .A2(n6441), .ZN(n8555) );
  INV_X1 U5996 ( .A(n5824), .ZN(n4926) );
  XNOR2_X1 U5997 ( .A(n5869), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5936) );
  INV_X1 U5998 ( .A(n5936), .ZN(n7877) );
  AND2_X1 U5999 ( .A1(n5991), .A2(n5990), .ZN(n4473) );
  INV_X1 U6000 ( .A(n4860), .ZN(n4859) );
  NAND2_X1 U6001 ( .A1(n4862), .A2(n4529), .ZN(n4860) );
  AND2_X1 U6002 ( .A1(n9040), .A2(n9039), .ZN(n4474) );
  NAND2_X1 U6003 ( .A1(n6323), .A2(n6322), .ZN(n9358) );
  INV_X1 U6004 ( .A(n9358), .ZN(n4672) );
  AND4_X1 U6005 ( .A1(n6002), .A2(n5995), .A3(n5999), .A4(n10032), .ZN(n4475)
         );
  AND4_X1 U6006 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5558), .ZN(n4476)
         );
  AND2_X1 U6007 ( .A1(n5823), .A2(n5822), .ZN(n8230) );
  AND3_X1 U6008 ( .A1(n8666), .A2(n8856), .A3(n8758), .ZN(n4477) );
  AND2_X1 U6009 ( .A1(n5803), .A2(n5804), .ZN(n8186) );
  INV_X1 U6010 ( .A(n8186), .ZN(n4800) );
  AND2_X1 U6011 ( .A1(n7915), .A2(n8209), .ZN(n4478) );
  AND2_X1 U6012 ( .A1(n5407), .A2(n5406), .ZN(n9897) );
  INV_X1 U6013 ( .A(n9897), .ZN(n7480) );
  AND4_X1 U6014 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n7463)
         );
  INV_X1 U6015 ( .A(n7463), .ZN(n4764) );
  NAND2_X1 U6016 ( .A1(n6423), .A2(n6422), .ZN(n9329) );
  INV_X1 U6017 ( .A(n5487), .ZN(n4643) );
  AND2_X1 U6018 ( .A1(n9381), .A2(n8925), .ZN(n4479) );
  AND2_X1 U6019 ( .A1(n4471), .A2(n8073), .ZN(n4480) );
  AND2_X1 U6020 ( .A1(n4745), .A2(n6012), .ZN(n4481) );
  AND2_X1 U6021 ( .A1(n5795), .A2(n5794), .ZN(n4482) );
  AND2_X1 U6022 ( .A1(n4984), .A2(n6468), .ZN(n4483) );
  AND2_X1 U6023 ( .A1(n6454), .A2(n6453), .ZN(n4484) );
  NAND2_X1 U6024 ( .A1(n6288), .A2(n6287), .ZN(n9370) );
  AND2_X1 U6025 ( .A1(n4979), .A2(n6271), .ZN(n4485) );
  INV_X1 U6026 ( .A(n4864), .ZN(n4863) );
  OAI21_X1 U6027 ( .B1(n7993), .B2(n4458), .A(n4865), .ZN(n4864) );
  AND2_X1 U6028 ( .A1(n5015), .A2(n4444), .ZN(n4486) );
  AND2_X1 U6029 ( .A1(n5246), .A2(n5864), .ZN(n6917) );
  INV_X1 U6030 ( .A(n6917), .ZN(n4808) );
  OR2_X1 U6031 ( .A1(n4455), .A2(n4825), .ZN(n4487) );
  INV_X1 U6032 ( .A(n7780), .ZN(n4648) );
  INV_X1 U6033 ( .A(n4553), .ZN(n5271) );
  OAI211_X1 U6034 ( .C1(n5060), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4554), .ZN(n4553) );
  AND2_X1 U6035 ( .A1(n4890), .A2(n4887), .ZN(n4488) );
  AND2_X1 U6036 ( .A1(n9280), .A2(n4456), .ZN(n4489) );
  AND2_X1 U6037 ( .A1(n4613), .A2(n6404), .ZN(n4490) );
  NOR2_X1 U6038 ( .A1(n5449), .A2(n4889), .ZN(n4888) );
  AND2_X1 U6039 ( .A1(n8504), .A2(n8505), .ZN(n4491) );
  AND2_X1 U6040 ( .A1(n4695), .A2(n4697), .ZN(n4492) );
  AND2_X1 U6041 ( .A1(n9394), .A2(n4714), .ZN(n4493) );
  AND2_X1 U6042 ( .A1(n4619), .A2(n4617), .ZN(n4494) );
  INV_X1 U6043 ( .A(n4845), .ZN(n4842) );
  OR2_X1 U6044 ( .A1(n4478), .A2(n4849), .ZN(n4845) );
  INV_X1 U6045 ( .A(n5010), .ZN(n5009) );
  NAND2_X1 U6046 ( .A1(n9375), .A2(n8924), .ZN(n4495) );
  INV_X1 U6047 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6048 ( .A1(n5890), .A2(n4764), .ZN(n4496) );
  AND2_X1 U6049 ( .A1(n8772), .A2(n8771), .ZN(n8893) );
  NOR2_X1 U6050 ( .A1(n7530), .A2(n8930), .ZN(n4497) );
  OR2_X1 U6051 ( .A1(n9196), .A2(n8923), .ZN(n9063) );
  AND2_X1 U6052 ( .A1(n4912), .A2(n5788), .ZN(n4498) );
  INV_X1 U6053 ( .A(n4669), .ZN(n4668) );
  NAND2_X1 U6054 ( .A1(n4670), .A2(n9165), .ZN(n4669) );
  AND2_X1 U6055 ( .A1(n8467), .A2(n5784), .ZN(n4499) );
  NAND2_X1 U6056 ( .A1(n4469), .A2(n7812), .ZN(n4500) );
  INV_X1 U6057 ( .A(n5766), .ZN(n8391) );
  NAND2_X1 U6058 ( .A1(n5753), .A2(n5752), .ZN(n5766) );
  NOR2_X1 U6059 ( .A1(n9126), .A2(n9054), .ZN(n4501) );
  XNOR2_X1 U6060 ( .A(n5725), .B(SI_29_), .ZN(n7888) );
  NOR2_X1 U6061 ( .A1(n8420), .A2(n8233), .ZN(n4502) );
  NAND3_X1 U6062 ( .A1(n5038), .A2(n5039), .A3(n4475), .ZN(n4503) );
  AND2_X1 U6063 ( .A1(n9126), .A2(n9054), .ZN(n4504) );
  OR2_X1 U6064 ( .A1(n7338), .A2(n7604), .ZN(n4505) );
  INV_X1 U6065 ( .A(n7194), .ZN(n4815) );
  NAND2_X1 U6066 ( .A1(n5896), .A2(n9910), .ZN(n4506) );
  AND2_X1 U6067 ( .A1(n4860), .A2(n4856), .ZN(n4507) );
  OR2_X1 U6068 ( .A1(n6652), .A2(n6643), .ZN(n4508) );
  INV_X1 U6069 ( .A(n8398), .ZN(n8048) );
  AND2_X1 U6070 ( .A1(n5676), .A2(n5675), .ZN(n8398) );
  NAND2_X1 U6071 ( .A1(n8772), .A2(n9076), .ZN(n4509) );
  AND2_X1 U6072 ( .A1(n8398), .A2(n8183), .ZN(n4510) );
  NOR2_X1 U6073 ( .A1(n5103), .A2(SI_11_), .ZN(n4511) );
  INV_X1 U6074 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U6075 ( .A1(n4699), .A2(n7159), .ZN(n4693) );
  OR2_X1 U6076 ( .A1(n5017), .A2(n5013), .ZN(n4512) );
  INV_X1 U6077 ( .A(n6770), .ZN(n4695) );
  NAND2_X1 U6078 ( .A1(n4480), .A2(n4776), .ZN(n4513) );
  AND2_X1 U6079 ( .A1(n4857), .A2(n4856), .ZN(n4514) );
  AND2_X1 U6080 ( .A1(n8783), .A2(n8856), .ZN(n4515) );
  AND3_X1 U6081 ( .A1(n4650), .A2(n4649), .A3(n4648), .ZN(n4516) );
  AND2_X1 U6082 ( .A1(n5110), .A2(n4898), .ZN(n4517) );
  AND2_X1 U6083 ( .A1(n4779), .A2(n4777), .ZN(n4518) );
  NOR2_X1 U6084 ( .A1(n4897), .A2(n4895), .ZN(n4519) );
  AOI21_X1 U6085 ( .B1(n8186), .B2(n4797), .A(n5917), .ZN(n4796) );
  NOR2_X1 U6086 ( .A1(n6014), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5979) );
  AND2_X1 U6087 ( .A1(n7829), .A2(n4606), .ZN(n4520) );
  INV_X1 U6088 ( .A(n5908), .ZN(n4757) );
  AND2_X1 U6089 ( .A1(n4629), .A2(n4628), .ZN(n4521) );
  AND2_X1 U6090 ( .A1(n6487), .A2(n6472), .ZN(n4522) );
  AND2_X1 U6091 ( .A1(n4473), .A2(n6318), .ZN(n4523) );
  OR2_X1 U6092 ( .A1(n8445), .A2(n8284), .ZN(n5792) );
  NAND2_X1 U6093 ( .A1(n6046), .A2(n7295), .ZN(n8859) );
  NAND2_X1 U6094 ( .A1(n8163), .A2(n8171), .ZN(n4524) );
  AND2_X1 U6095 ( .A1(n4844), .A2(n4840), .ZN(n4839) );
  AND2_X1 U6096 ( .A1(n8763), .A2(n8762), .ZN(n9389) );
  INV_X2 U6097 ( .A(n4438), .ZN(n5288) );
  INV_X1 U6098 ( .A(n9196), .ZN(n4671) );
  XNOR2_X1 U6099 ( .A(n5354), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7159) );
  AND3_X1 U6100 ( .A1(n4607), .A2(n6197), .A3(n4606), .ZN(n7828) );
  INV_X1 U6101 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4906) );
  AND2_X1 U6102 ( .A1(n9008), .A2(n4453), .ZN(n4525) );
  INV_X1 U6103 ( .A(n9747), .ZN(n8129) );
  NAND2_X1 U6104 ( .A1(n4996), .A2(n5000), .ZN(n7813) );
  AND2_X1 U6105 ( .A1(n5390), .A2(n5417), .ZN(n7233) );
  INV_X1 U6106 ( .A(n7233), .ZN(n7226) );
  AND2_X1 U6107 ( .A1(n4982), .A2(n4981), .ZN(n4526) );
  INV_X1 U6108 ( .A(n8614), .ZN(n6403) );
  NAND2_X1 U6109 ( .A1(n4971), .A2(n4975), .ZN(n8492) );
  INV_X1 U6110 ( .A(n6285), .ZN(n5027) );
  INV_X1 U6111 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6112 ( .A1(n7898), .A2(n7899), .ZN(n4527) );
  NAND2_X2 U6113 ( .A1(n6628), .A2(n9857), .ZN(n8318) );
  INV_X1 U6114 ( .A(n9797), .ZN(n4701) );
  NOR2_X1 U6115 ( .A1(n9609), .A2(n7184), .ZN(n9606) );
  INV_X1 U6116 ( .A(n9606), .ZN(n9294) );
  NAND2_X1 U6117 ( .A1(n7474), .A2(n7473), .ZN(n7647) );
  AND2_X1 U6118 ( .A1(n7251), .A2(n6100), .ZN(n4528) );
  INV_X1 U6119 ( .A(n8378), .ZN(n9927) );
  INV_X2 U6120 ( .A(n9917), .ZN(n9915) );
  INV_X1 U6121 ( .A(n9780), .ZN(n8127) );
  XNOR2_X1 U6122 ( .A(n7743), .B(n8073), .ZN(n7745) );
  AND2_X1 U6123 ( .A1(n5891), .A2(n5890), .ZN(n7404) );
  OR2_X1 U6124 ( .A1(n7908), .A2(n8265), .ZN(n4529) );
  AOI21_X1 U6125 ( .B1(n7743), .B2(n4834), .A(n4833), .ZN(n7758) );
  AND2_X1 U6126 ( .A1(n8603), .A2(n4978), .ZN(n4530) );
  INV_X1 U6127 ( .A(n7853), .ZN(n4981) );
  OR2_X1 U6128 ( .A1(n8318), .A2(n6629), .ZN(n4531) );
  INV_X1 U6129 ( .A(SI_15_), .ZN(n4895) );
  INV_X1 U6130 ( .A(n4806), .ZN(n6916) );
  NAND2_X1 U6131 ( .A1(n7096), .A2(n7095), .ZN(n7195) );
  NAND2_X1 U6132 ( .A1(n4804), .A2(n6965), .ZN(n6967) );
  XNOR2_X1 U6133 ( .A(n5365), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7161) );
  INV_X1 U6134 ( .A(n7161), .ZN(n4622) );
  XNOR2_X1 U6135 ( .A(n5765), .B(n5764), .ZN(n7658) );
  AND2_X2 U6136 ( .A1(n6791), .A2(n6666), .ZN(n9012) );
  NAND3_X1 U6137 ( .A1(n8681), .A2(n4598), .A3(n4532), .ZN(n4597) );
  INV_X1 U6138 ( .A(n8721), .ZN(n4601) );
  NOR2_X1 U6139 ( .A1(n8716), .A2(n8715), .ZN(n8720) );
  AOI21_X1 U6140 ( .B1(n4557), .B2(n4569), .A(n8893), .ZN(n4568) );
  AOI21_X1 U6141 ( .B1(n8705), .B2(n4573), .A(n4571), .ZN(n4578) );
  OAI21_X1 U6142 ( .B1(n4576), .B2(n8770), .A(n4575), .ZN(n8712) );
  AOI211_X1 U6143 ( .C1(n8738), .C2(n8737), .A(n8736), .B(n9153), .ZN(n4588)
         );
  NAND2_X1 U6144 ( .A1(n7457), .A2(n7462), .ZN(n7600) );
  NAND2_X1 U6145 ( .A1(n5775), .A2(n5834), .ZN(n7403) );
  OAI21_X1 U6146 ( .B1(n8187), .B2(n5805), .A(n5804), .ZN(n8174) );
  NAND2_X1 U6147 ( .A1(n4930), .A2(n4929), .ZN(n8262) );
  NAND2_X1 U6148 ( .A1(n6594), .A2(n5808), .ZN(n5810) );
  INV_X1 U6149 ( .A(n5241), .ZN(n4752) );
  NAND2_X1 U6150 ( .A1(n4778), .A2(n5895), .ZN(n7703) );
  NAND2_X1 U6151 ( .A1(n5893), .A2(n5892), .ZN(n7459) );
  NAND2_X1 U6152 ( .A1(n7779), .A2(n5897), .ZN(n7803) );
  INV_X1 U6153 ( .A(n4533), .ZN(n7781) );
  NAND2_X1 U6154 ( .A1(n5912), .A2(n5044), .ZN(n8250) );
  OAI21_X2 U6155 ( .B1(n8325), .B2(n5904), .A(n5903), .ZN(n8299) );
  NAND2_X1 U6156 ( .A1(n5907), .A2(n5906), .ZN(n8287) );
  OAI22_X1 U6157 ( .A1(n7207), .A2(n4753), .B1(n8076), .B2(n7211), .ZN(n7305)
         );
  NAND2_X1 U6158 ( .A1(n9312), .A2(n4534), .ZN(P1_U3550) );
  NAND2_X1 U6159 ( .A1(n9397), .A2(n4535), .ZN(P1_U3518) );
  AOI21_X2 U6160 ( .B1(n7668), .B2(n7667), .A(n7666), .ZN(n7670) );
  NAND2_X1 U6161 ( .A1(n4539), .A2(n4536), .ZN(n5598) );
  OAI21_X1 U6162 ( .B1(n5570), .B2(n5569), .A(n4538), .ZN(n4537) );
  NAND2_X1 U6163 ( .A1(n4651), .A2(n4516), .ZN(n4647) );
  NAND2_X1 U6164 ( .A1(n4645), .A2(n7802), .ZN(n4644) );
  OAI21_X1 U6165 ( .B1(n5055), .B2(SI_2_), .A(n5065), .ZN(n5304) );
  AOI21_X1 U6166 ( .B1(n4655), .B2(n4654), .A(n5629), .ZN(n4653) );
  NAND2_X1 U6167 ( .A1(n5330), .A2(n5929), .ZN(n4540) );
  NAND2_X1 U6168 ( .A1(n4542), .A2(n6636), .ZN(n4541) );
  NAND2_X1 U6169 ( .A1(n5771), .A2(n5770), .ZN(n4542) );
  AOI21_X1 U6170 ( .B1(n5601), .B2(n6636), .A(n4926), .ZN(n4654) );
  NOR2_X1 U6171 ( .A1(n9532), .A2(n8990), .ZN(n9544) );
  NAND2_X1 U6172 ( .A1(n4647), .A2(n4646), .ZN(n4645) );
  AOI21_X1 U6173 ( .B1(n5724), .B2(n4638), .A(n4636), .ZN(n4634) );
  XNOR2_X2 U6174 ( .A(n6068), .B(P1_IR_REG_3__SCAN_IN), .ZN(n8950) );
  AOI21_X1 U6175 ( .B1(n4644), .B2(n5488), .A(n4641), .ZN(n5489) );
  NAND2_X1 U6176 ( .A1(n5463), .A2(n5462), .ZN(n4651) );
  NAND3_X1 U6177 ( .A1(n5340), .A2(n5525), .A3(n5191), .ZN(n5241) );
  NAND2_X1 U6178 ( .A1(n4544), .A2(n4543), .ZN(P2_U3485) );
  INV_X1 U6179 ( .A(n8347), .ZN(n4544) );
  NAND2_X1 U6180 ( .A1(n4546), .A2(n4545), .ZN(P2_U3453) );
  INV_X1 U6181 ( .A(n8401), .ZN(n4546) );
  NAND2_X1 U6182 ( .A1(n4547), .A2(n9740), .ZN(n4629) );
  XNOR2_X1 U6183 ( .A(n8095), .B(n4548), .ZN(n4547) );
  NAND2_X1 U6184 ( .A1(n5900), .A2(n5899), .ZN(n8325) );
  NAND2_X1 U6185 ( .A1(n6729), .A2(n6730), .ZN(n6765) );
  NAND2_X1 U6186 ( .A1(n4760), .A2(n4759), .ZN(n7461) );
  NAND2_X1 U6187 ( .A1(n4630), .A2(n4521), .ZN(P2_U3201) );
  NAND2_X1 U6188 ( .A1(n5163), .A2(n5162), .ZN(n5674) );
  NAND2_X1 U6189 ( .A1(n4637), .A2(n5857), .ZN(n4636) );
  XNOR2_X2 U6190 ( .A(n6083), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7052) );
  INV_X1 U6191 ( .A(n4869), .ZN(n4659) );
  NAND2_X1 U6192 ( .A1(n5306), .A2(n5065), .ZN(n4552) );
  INV_X1 U6193 ( .A(n5716), .ZN(n4868) );
  NAND2_X1 U6194 ( .A1(n4552), .A2(n5319), .ZN(n5321) );
  INV_X1 U6195 ( .A(n5319), .ZN(n4550) );
  INV_X1 U6196 ( .A(n4552), .ZN(n4551) );
  OAI21_X1 U6197 ( .B1(n8753), .B2(n9009), .A(n4564), .ZN(n4563) );
  NAND2_X1 U6198 ( .A1(n4568), .A2(n4566), .ZN(n8908) );
  AND2_X1 U6199 ( .A1(n8915), .A2(n8843), .ZN(n4569) );
  OR2_X1 U6200 ( .A1(n8710), .A2(n9024), .ZN(n4570) );
  NAND2_X1 U6201 ( .A1(n4570), .A2(n8877), .ZN(n4577) );
  NAND2_X1 U6202 ( .A1(n8711), .A2(n8770), .ZN(n4575) );
  NOR2_X1 U6203 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U6204 ( .A1(n4581), .A2(n4580), .ZN(n5385) );
  NAND2_X1 U6205 ( .A1(n5339), .A2(n4583), .ZN(n4580) );
  NAND2_X1 U6206 ( .A1(n5355), .A2(n4584), .ZN(n4582) );
  NAND2_X1 U6207 ( .A1(n4593), .A2(n4589), .ZN(n8699) );
  NAND2_X1 U6208 ( .A1(n4590), .A2(n8770), .ZN(n4589) );
  NAND2_X1 U6209 ( .A1(n4592), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U6210 ( .A1(n4597), .A2(n8686), .ZN(n4592) );
  AOI21_X1 U6211 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(n4594) );
  AND2_X1 U6212 ( .A1(n8682), .A2(n8683), .ZN(n4596) );
  NAND4_X1 U6213 ( .A1(n4600), .A2(n8770), .A3(n8774), .A4(n8883), .ZN(n4599)
         );
  NAND2_X1 U6214 ( .A1(n4603), .A2(n7083), .ZN(n6035) );
  NAND2_X1 U6215 ( .A1(n4603), .A2(n7112), .ZN(n6051) );
  NAND2_X1 U6216 ( .A1(n8645), .A2(n6472), .ZN(n6557) );
  NAND2_X1 U6217 ( .A1(n7830), .A2(n7829), .ZN(n4605) );
  NAND3_X1 U6218 ( .A1(n4607), .A2(n4520), .A3(n6197), .ZN(n4604) );
  NAND3_X1 U6219 ( .A1(n4605), .A2(n7854), .A3(n4604), .ZN(n4982) );
  AND2_X1 U6220 ( .A1(n4605), .A2(n4604), .ZN(n7827) );
  INV_X1 U6221 ( .A(n6195), .ZN(n4608) );
  INV_X1 U6222 ( .A(n6196), .ZN(n4609) );
  OAI21_X2 U6223 ( .B1(n7414), .B2(n6147), .A(n4618), .ZN(n4620) );
  NAND2_X1 U6224 ( .A1(n4616), .A2(n4615), .ZN(n7715) );
  INV_X1 U6225 ( .A(n6176), .ZN(n4617) );
  NAND2_X1 U6226 ( .A1(n6286), .A2(n4523), .ZN(n6321) );
  NOR2_X4 U6227 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6701) );
  NAND2_X1 U6228 ( .A1(n5321), .A2(n5069), .ZN(n5337) );
  NAND2_X1 U6229 ( .A1(n5068), .A2(n5067), .ZN(n4633) );
  NAND3_X1 U6230 ( .A1(n5723), .A2(n5853), .A3(n5929), .ZN(n4635) );
  NAND2_X1 U6231 ( .A1(n4635), .A2(n4634), .ZN(n4873) );
  NOR2_X1 U6232 ( .A1(n4643), .A2(n4642), .ZN(n4641) );
  OAI211_X1 U6233 ( .C1(n4653), .C2(n4652), .A(n5643), .B(n8197), .ZN(n5658)
         );
  NAND3_X1 U6234 ( .A1(n5842), .A2(n5778), .A3(n6636), .ZN(n4658) );
  NOR3_X2 U6235 ( .A1(n5704), .A2(n5703), .A3(n4659), .ZN(n5716) );
  MUX2_X1 U6236 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5060), .Z(n5066) );
  MUX2_X1 U6237 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4660), .Z(n5070) );
  MUX2_X1 U6238 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5060), .Z(n5075) );
  MUX2_X1 U6239 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4660), .Z(n5089) );
  MUX2_X1 U6240 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4660), .Z(n5080) );
  MUX2_X1 U6241 ( .A(n10071), .B(n5081), .S(n4660), .Z(n5083) );
  MUX2_X1 U6242 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4660), .Z(n5099) );
  MUX2_X1 U6243 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4660), .Z(n5103) );
  OR2_X1 U6244 ( .A1(n9093), .A2(n9389), .ZN(n4664) );
  NAND2_X1 U6245 ( .A1(n9093), .A2(n4666), .ZN(n9080) );
  NAND2_X1 U6246 ( .A1(n9093), .A2(n9099), .ZN(n9094) );
  NAND3_X1 U6247 ( .A1(n4664), .A2(n4662), .A3(n4661), .ZN(n9010) );
  NAND2_X1 U6248 ( .A1(n9190), .A2(n4667), .ZN(n9143) );
  NAND3_X1 U6249 ( .A1(n9240), .A2(n4453), .A3(n9008), .ZN(n9239) );
  NAND2_X1 U6250 ( .A1(n7241), .A2(n7242), .ZN(n4679) );
  NAND2_X1 U6251 ( .A1(n4685), .A2(n7240), .ZN(n4684) );
  NAND3_X1 U6252 ( .A1(n4691), .A2(n4694), .A3(n4690), .ZN(n7160) );
  NAND2_X1 U6253 ( .A1(n4698), .A2(n4697), .ZN(n4696) );
  MUX2_X1 U6254 ( .A(n6762), .B(P2_REG2_REG_2__SCAN_IN), .S(n6763), .Z(n6730)
         );
  AND3_X2 U6255 ( .A1(n4706), .A2(n4705), .A3(n4704), .ZN(n6763) );
  OAI21_X1 U6256 ( .B1(n9843), .B2(n4710), .A(n4709), .ZN(n9481) );
  NOR2_X1 U6257 ( .A1(n9843), .A2(n9842), .ZN(n9841) );
  NAND2_X1 U6258 ( .A1(n9079), .A2(n9078), .ZN(n9305) );
  NAND4_X2 U6259 ( .A1(n6081), .A2(n6047), .A3(n4717), .A4(n5963), .ZN(n6132)
         );
  NAND3_X1 U6260 ( .A1(n6081), .A2(n6047), .A3(n4717), .ZN(n6114) );
  AOI21_X1 U6261 ( .B1(n8667), .B2(n8856), .A(n4515), .ZN(n4718) );
  NAND2_X1 U6262 ( .A1(n8863), .A2(n8860), .ZN(n7522) );
  NAND2_X1 U6263 ( .A1(n7670), .A2(n4724), .ZN(n4723) );
  INV_X1 U6264 ( .A(n4727), .ZN(n4728) );
  OAI21_X1 U6265 ( .B1(n4731), .B2(n7025), .A(n8859), .ZN(n4727) );
  NAND2_X1 U6266 ( .A1(n4728), .A2(n4729), .ZN(n7173) );
  NAND2_X1 U6267 ( .A1(n9260), .A2(n4735), .ZN(n4732) );
  NAND2_X1 U6268 ( .A1(n4732), .A2(n4733), .ZN(n9216) );
  OAI21_X2 U6269 ( .B1(n7815), .B2(n4741), .A(n4739), .ZN(n9279) );
  INV_X1 U6270 ( .A(n6015), .ZN(n5976) );
  NAND3_X1 U6271 ( .A1(n5038), .A2(n5039), .A3(n4744), .ZN(n6004) );
  OAI21_X1 U6272 ( .B1(n9201), .B2(n9200), .A(n9062), .ZN(n9186) );
  INV_X1 U6273 ( .A(n9185), .ZN(n4751) );
  NAND2_X1 U6274 ( .A1(n5881), .A2(n7002), .ZN(n5768) );
  INV_X2 U6275 ( .A(n7002), .ZN(n7300) );
  NAND2_X2 U6276 ( .A1(n4752), .A2(n4476), .ZN(n5871) );
  NAND2_X1 U6277 ( .A1(n8287), .A2(n5908), .ZN(n4754) );
  NAND2_X1 U6278 ( .A1(n5891), .A2(n4761), .ZN(n4760) );
  OAI21_X1 U6279 ( .B1(n5890), .B2(n4764), .A(n9892), .ZN(n4763) );
  NAND2_X1 U6280 ( .A1(n5198), .A2(n4772), .ZN(n4771) );
  INV_X1 U6281 ( .A(n4765), .ZN(n4767) );
  NAND2_X1 U6282 ( .A1(n7596), .A2(n4518), .ZN(n4775) );
  NAND2_X1 U6283 ( .A1(n7596), .A2(n7640), .ZN(n4781) );
  NAND3_X1 U6284 ( .A1(n4782), .A2(n4781), .A3(n4471), .ZN(n4778) );
  NAND2_X1 U6285 ( .A1(n8243), .A2(n4786), .ZN(n4784) );
  INV_X1 U6286 ( .A(n8230), .ZN(n4791) );
  INV_X1 U6287 ( .A(n8181), .ZN(n4794) );
  NAND2_X1 U6288 ( .A1(n4793), .A2(n4795), .ZN(n6597) );
  NAND2_X1 U6289 ( .A1(n4794), .A2(n4796), .ZN(n4793) );
  OR2_X1 U6290 ( .A1(n5297), .A2(n10128), .ZN(n5268) );
  NAND2_X1 U6291 ( .A1(n5053), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U6292 ( .A1(n4873), .A2(n4872), .ZN(n5862) );
  NAND3_X1 U6293 ( .A1(n4804), .A2(n6965), .A3(n6969), .ZN(n7094) );
  NAND2_X1 U6294 ( .A1(n8017), .A2(n4454), .ZN(n4811) );
  NAND2_X1 U6295 ( .A1(n7096), .A2(n4819), .ZN(n4818) );
  NAND3_X1 U6296 ( .A1(n4818), .A2(n4817), .A3(n7262), .ZN(n7368) );
  NAND2_X1 U6297 ( .A1(n7925), .A2(n4822), .ZN(n4821) );
  OAI211_X1 U6298 ( .C1(n7925), .C2(n4823), .A(n4821), .B(n7967), .ZN(P2_U3160) );
  OAI21_X1 U6299 ( .B1(n7743), .B2(n4833), .A(n4831), .ZN(n4836) );
  INV_X1 U6300 ( .A(n4836), .ZN(n7759) );
  NAND2_X1 U6301 ( .A1(n7942), .A2(n4839), .ZN(n4837) );
  NAND2_X1 U6302 ( .A1(n7994), .A2(n4514), .ZN(n4855) );
  XNOR2_X2 U6303 ( .A(n5727), .B(n5726), .ZN(n5725) );
  NAND2_X1 U6304 ( .A1(n4868), .A2(n4867), .ZN(n5720) );
  NAND2_X1 U6305 ( .A1(n4869), .A2(n5717), .ZN(n4867) );
  NAND2_X1 U6306 ( .A1(n5604), .A2(n4878), .ZN(n4876) );
  NAND2_X1 U6307 ( .A1(n5101), .A2(n5100), .ZN(n5433) );
  NAND2_X1 U6308 ( .A1(n4893), .A2(n4891), .ZN(n5124) );
  NAND2_X1 U6309 ( .A1(n5115), .A2(n5114), .ZN(n5524) );
  NAND2_X1 U6310 ( .A1(n5251), .A2(n4517), .ZN(n4896) );
  NAND2_X1 U6311 ( .A1(n4896), .A2(n4519), .ZN(n5112) );
  NAND3_X1 U6312 ( .A1(n4899), .A2(n4902), .A3(n4901), .ZN(n5057) );
  NAND3_X1 U6313 ( .A1(n4904), .A2(n4906), .A3(n4903), .ZN(n4899) );
  NAND2_X1 U6314 ( .A1(n5053), .A2(n4900), .ZN(n4901) );
  NAND3_X1 U6315 ( .A1(n5054), .A2(n9007), .A3(n4905), .ZN(n4902) );
  INV_X1 U6316 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6317 ( .A1(n8307), .A2(n4911), .ZN(n4907) );
  NAND2_X1 U6318 ( .A1(n4907), .A2(n4908), .ZN(n8283) );
  OAI21_X1 U6319 ( .B1(n7609), .B2(n5448), .A(n4918), .ZN(n7785) );
  NAND2_X1 U6320 ( .A1(n4917), .A2(n4915), .ZN(n5782) );
  NAND2_X1 U6321 ( .A1(n7609), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U6322 ( .A1(n5796), .A2(n4924), .ZN(n4920) );
  NAND2_X1 U6323 ( .A1(n4920), .A2(n4921), .ZN(n8216) );
  NAND2_X1 U6324 ( .A1(n5796), .A2(n5827), .ZN(n8239) );
  OAI21_X2 U6325 ( .B1(n8174), .B2(n5806), .A(n5807), .ZN(n6594) );
  NAND2_X1 U6326 ( .A1(n5791), .A2(n4931), .ZN(n4930) );
  OAI21_X1 U6327 ( .B1(n5799), .B2(n4932), .A(n4933), .ZN(n5802) );
  NAND2_X1 U6328 ( .A1(n8078), .A2(n6935), .ZN(n5329) );
  INV_X1 U6329 ( .A(n5884), .ZN(n9859) );
  NAND2_X1 U6330 ( .A1(n9851), .A2(n9859), .ZN(n9850) );
  NAND2_X1 U6331 ( .A1(n4939), .A2(n4940), .ZN(n5786) );
  NAND2_X1 U6332 ( .A1(n7809), .A2(n5783), .ZN(n4939) );
  NOR2_X2 U6333 ( .A1(n5871), .A2(n4941), .ZN(n5227) );
  OR2_X1 U6334 ( .A1(n4962), .A2(n9087), .ZN(n4953) );
  NAND2_X1 U6335 ( .A1(n9087), .A2(n4960), .ZN(n4952) );
  NAND3_X1 U6336 ( .A1(n4950), .A2(n4948), .A3(n9086), .ZN(P1_U3356) );
  NAND2_X1 U6337 ( .A1(n9087), .A2(n4949), .ZN(n4948) );
  OR2_X1 U6338 ( .A1(n9087), .A2(n4951), .ZN(n4950) );
  NAND3_X1 U6339 ( .A1(n4953), .A2(n4952), .A3(n4957), .ZN(n9392) );
  AND2_X1 U6340 ( .A1(n4957), .A2(n4956), .ZN(n4955) );
  NAND2_X1 U6341 ( .A1(n6402), .A2(n6401), .ZN(n6404) );
  NAND2_X1 U6342 ( .A1(n4965), .A2(n7251), .ZN(n4967) );
  AND2_X1 U6343 ( .A1(n6129), .A2(n4970), .ZN(n4965) );
  NAND2_X1 U6344 ( .A1(n4968), .A2(n4967), .ZN(n7414) );
  NAND2_X1 U6345 ( .A1(n7827), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U6346 ( .A1(n8581), .A2(n4445), .ZN(n4983) );
  NAND2_X1 U6347 ( .A1(n7550), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U6348 ( .A1(n7665), .A2(n4995), .ZN(n4992) );
  NAND2_X1 U6349 ( .A1(n4992), .A2(n4993), .ZN(n9022) );
  NAND2_X1 U6350 ( .A1(n9049), .A2(n5004), .ZN(n5001) );
  NAND2_X1 U6351 ( .A1(n5001), .A2(n5002), .ZN(n9103) );
  NOR2_X1 U6352 ( .A1(n9165), .A2(n9050), .ZN(n5010) );
  INV_X1 U6353 ( .A(n9421), .ZN(n5019) );
  NAND2_X1 U6354 ( .A1(n5020), .A2(n6272), .ZN(n5028) );
  OAI211_X1 U6355 ( .C1(n6285), .C2(n6272), .A(n5022), .B(n5025), .ZN(n5021)
         );
  NAND2_X1 U6356 ( .A1(n5024), .A2(n5027), .ZN(n5022) );
  NAND2_X1 U6357 ( .A1(n5023), .A2(n5027), .ZN(n5026) );
  NAND2_X1 U6358 ( .A1(n6272), .A2(n8493), .ZN(n5023) );
  INV_X1 U6359 ( .A(n8493), .ZN(n5024) );
  NAND2_X1 U6360 ( .A1(n8564), .A2(n8565), .ZN(n8563) );
  NAND2_X1 U6361 ( .A1(n6558), .A2(n6559), .ZN(n6560) );
  NAND2_X1 U6362 ( .A1(n8645), .A2(n4522), .ZN(n6559) );
  NAND2_X1 U6363 ( .A1(n9276), .A2(n4456), .ZN(n5029) );
  NAND2_X1 U6364 ( .A1(n5029), .A2(n5030), .ZN(n5032) );
  INV_X1 U6365 ( .A(n5033), .ZN(n9275) );
  INV_X1 U6366 ( .A(n5032), .ZN(n9258) );
  NAND3_X1 U6367 ( .A1(n6791), .A2(n7041), .A3(n8943), .ZN(n5036) );
  AND2_X2 U6368 ( .A1(n6668), .A2(n6643), .ZN(n6080) );
  INV_X1 U6369 ( .A(n5968), .ZN(n5037) );
  NAND2_X1 U6370 ( .A1(n5039), .A2(n5038), .ZN(n5994) );
  AND2_X2 U6371 ( .A1(n5971), .A2(n5037), .ZN(n5038) );
  INV_X2 U6372 ( .A(n6132), .ZN(n5039) );
  NOR2_X1 U6373 ( .A1(n6132), .A2(n5968), .ZN(n6259) );
  NAND2_X1 U6374 ( .A1(n6625), .A2(n9915), .ZN(n6612) );
  NAND2_X1 U6375 ( .A1(n6625), .A2(n9929), .ZN(n6592) );
  XNOR2_X1 U6376 ( .A(n6966), .B(n9852), .ZN(n6964) );
  XNOR2_X1 U6377 ( .A(n6966), .B(n7002), .ZN(n6931) );
  INV_X1 U6378 ( .A(n6724), .ZN(n6711) );
  OAI21_X2 U6379 ( .B1(n7986), .B2(n7904), .A(n7903), .ZN(n7994) );
  AOI21_X2 U6380 ( .B1(n5933), .B2(n8331), .A(n5932), .ZN(n7887) );
  AND2_X1 U6381 ( .A1(n6060), .A2(n6059), .ZN(n7059) );
  NAND2_X1 U6382 ( .A1(n4460), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5986) );
  XNOR2_X1 U6383 ( .A(n7022), .B(n8850), .ZN(n7023) );
  INV_X1 U6384 ( .A(n5981), .ZN(n5983) );
  OAI22_X2 U6385 ( .A1(n8028), .A2(n8027), .B1(n7914), .B2(n8233), .ZN(n7942)
         );
  AOI21_X2 U6386 ( .B1(n7600), .B2(n5777), .A(n5776), .ZN(n7609) );
  AND2_X1 U6387 ( .A1(n9917), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5040) );
  AND2_X1 U6388 ( .A1(n6612), .A2(n6611), .ZN(n5041) );
  CLKBUF_X1 U6389 ( .A(n6677), .Z(n8483) );
  AND2_X1 U6390 ( .A1(n5721), .A2(n5817), .ZN(n5042) );
  AND2_X1 U6391 ( .A1(n8462), .A2(n8327), .ZN(n5043) );
  NOR2_X1 U6392 ( .A1(n6579), .A2(n8352), .ZN(n5047) );
  NOR2_X1 U6393 ( .A1(n6579), .A2(n8413), .ZN(n5048) );
  INV_X1 U6394 ( .A(n8352), .ZN(n6603) );
  INV_X1 U6395 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6396 ( .A1(n9915), .A2(n9907), .ZN(n8413) );
  INV_X1 U6397 ( .A(n8413), .ZN(n6608) );
  AND2_X1 U6398 ( .A1(n5858), .A2(n5857), .ZN(n5050) );
  INV_X1 U6399 ( .A(n6829), .ZN(n6992) );
  AND2_X1 U6400 ( .A1(n6630), .A2(n4531), .ZN(n5051) );
  INV_X1 U6401 ( .A(n9093), .ZN(n9112) );
  AND2_X1 U6402 ( .A1(n6550), .A2(n8634), .ZN(n5052) );
  AND2_X1 U6403 ( .A1(n5829), .A2(n5828), .ZN(n8288) );
  INV_X1 U6404 ( .A(n7462), .ZN(n5892) );
  INV_X1 U6405 ( .A(n7610), .ZN(n5779) );
  NAND2_X1 U6406 ( .A1(n6523), .A2(n6538), .ZN(n9493) );
  INV_X1 U6407 ( .A(n9493), .ZN(n8634) );
  INV_X1 U6408 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6409 ( .A1(n5766), .A2(n4640), .ZN(n5858) );
  INV_X1 U6410 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6629) );
  AND2_X1 U6411 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  INV_X1 U6412 ( .A(n7658), .ZN(n6918) );
  INV_X1 U6413 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5195) );
  INV_X1 U6414 ( .A(n6098), .ZN(n6099) );
  AND4_X1 U6415 ( .A1(n5970), .A2(n5969), .A3(n5989), .A4(n10248), .ZN(n5971)
         );
  INV_X1 U6416 ( .A(n5591), .ZN(n5218) );
  INV_X1 U6417 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U6418 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  NAND2_X1 U6419 ( .A1(n6097), .A2(n6099), .ZN(n6100) );
  INV_X1 U6420 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U6421 ( .A1(n6345), .A2(n8808), .ZN(n6521) );
  INV_X1 U6422 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10054) );
  INV_X1 U6423 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5972) );
  INV_X1 U6424 ( .A(SI_22_), .ZN(n5141) );
  INV_X1 U6425 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5125) );
  INV_X1 U6426 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5094) );
  INV_X1 U6427 ( .A(n7373), .ZN(n7370) );
  INV_X1 U6428 ( .A(n8068), .ZN(n6598) );
  INV_X1 U6429 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5199) );
  INV_X1 U6430 ( .A(n5620), .ZN(n5220) );
  OR2_X1 U6431 ( .A1(n5478), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5480) );
  OR2_X1 U6432 ( .A1(n5423), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5438) );
  NOR2_X1 U6433 ( .A1(n8171), .A2(n9860), .ZN(n6588) );
  NAND2_X1 U6434 ( .A1(n6038), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U6435 ( .A1(n6038), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6039) );
  INV_X1 U6436 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10162) );
  OR2_X1 U6437 ( .A1(n6391), .A2(n10171), .ZN(n6426) );
  OR2_X1 U6438 ( .A1(n6278), .A2(n10090), .ZN(n6290) );
  AND2_X1 U6439 ( .A1(n6222), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U6440 ( .A1(n9348), .A2(n9038), .ZN(n9039) );
  NAND2_X1 U6441 ( .A1(n7180), .A2(n7112), .ZN(n7171) );
  NAND2_X1 U6442 ( .A1(n5106), .A2(SI_13_), .ZN(n5110) );
  AND2_X1 U6443 ( .A1(n5935), .A2(n5873), .ZN(n5874) );
  OR2_X1 U6444 ( .A1(n7900), .A2(n7935), .ZN(n7901) );
  INV_X1 U6445 ( .A(n8329), .ZN(n8022) );
  OR2_X1 U6446 ( .A1(n6924), .A2(n6923), .ZN(n8045) );
  OR2_X1 U6447 ( .A1(P2_U3150), .A2(n6699), .ZN(n6908) );
  AND2_X1 U6448 ( .A1(n5817), .A2(n5816), .ZN(n5925) );
  NAND2_X1 U6449 ( .A1(n5223), .A2(n5222), .ZN(n5691) );
  OR2_X1 U6450 ( .A1(n5607), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5620) );
  OR2_X1 U6451 ( .A1(n5546), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5563) );
  INV_X1 U6452 ( .A(n5842), .ZN(n5776) );
  NAND2_X1 U6453 ( .A1(n6624), .A2(n6660), .ZN(n9857) );
  AND2_X1 U6454 ( .A1(n7658), .A2(n8096), .ZN(n9853) );
  AND2_X1 U6455 ( .A1(n5819), .A2(n5818), .ZN(n8200) );
  NAND2_X1 U6456 ( .A1(n6825), .A2(n5929), .ZN(n9861) );
  AND2_X1 U6457 ( .A1(n6809), .A2(n8333), .ZN(n6812) );
  INV_X1 U6458 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8496) );
  AND2_X1 U6459 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6101) );
  NAND2_X1 U6460 ( .A1(n6243), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6263) );
  NOR2_X1 U6461 ( .A1(n6202), .A2(n10162), .ZN(n6222) );
  INV_X1 U6462 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8622) );
  AND2_X1 U6463 ( .A1(n6444), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6457) );
  NOR2_X1 U6464 ( .A1(n6349), .A2(n8529), .ZN(n6350) );
  INV_X1 U6465 ( .A(n9060), .ZN(n9155) );
  NOR2_X1 U6466 ( .A1(n6155), .A2(n6154), .ZN(n6169) );
  NAND2_X1 U6467 ( .A1(n7275), .A2(n8855), .ZN(n8778) );
  NAND2_X1 U6468 ( .A1(n7171), .A2(n8859), .ZN(n8779) );
  AND2_X1 U6469 ( .A1(n5156), .A2(n5155), .ZN(n5644) );
  AND2_X1 U6470 ( .A1(n5110), .A2(n5109), .ZN(n5248) );
  INV_X1 U6471 ( .A(n5430), .ZN(n5100) );
  INV_X1 U6472 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5865) );
  AND4_X1 U6473 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n7747)
         );
  INV_X1 U6474 ( .A(n9696), .ZN(n9832) );
  INV_X1 U6475 ( .A(n9699), .ZN(n9839) );
  AND2_X1 U6476 ( .A1(n7600), .A2(n7458), .ZN(n7465) );
  INV_X1 U6477 ( .A(n8339), .ZN(n8260) );
  INV_X1 U6478 ( .A(n9857), .ZN(n8303) );
  NAND2_X1 U6479 ( .A1(n6622), .A2(n6621), .ZN(n6628) );
  AND2_X1 U6480 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  INV_X1 U6481 ( .A(n7981), .ZN(n8403) );
  NAND2_X1 U6482 ( .A1(n7775), .A2(n4808), .ZN(n9909) );
  INV_X1 U6483 ( .A(n9909), .ZN(n9907) );
  NAND2_X1 U6484 ( .A1(n7615), .A2(n9902), .ZN(n9914) );
  AND2_X1 U6485 ( .A1(n5953), .A2(n5952), .ZN(n6648) );
  XNOR2_X1 U6486 ( .A(n5435), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9713) );
  AND2_X1 U6487 ( .A1(n6665), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6670) );
  OR2_X1 U6488 ( .A1(n6187), .A2(n6186), .ZN(n6202) );
  INV_X1 U6489 ( .A(n9501), .ZN(n8656) );
  NAND2_X1 U6490 ( .A1(n6527), .A2(n9236), .ZN(n9497) );
  OR2_X1 U6491 ( .A1(n6562), .A2(n6477), .ZN(n6483) );
  INV_X1 U6492 ( .A(n9541), .ZN(n9570) );
  INV_X1 U6493 ( .A(n9565), .ZN(n9577) );
  INV_X1 U6494 ( .A(n6345), .ZN(n9002) );
  INV_X1 U6495 ( .A(n9236), .ZN(n9598) );
  NOR2_X1 U6496 ( .A1(n9665), .A2(n9384), .ZN(n9361) );
  INV_X1 U6497 ( .A(n9367), .ZN(n9354) );
  INV_X1 U6498 ( .A(n9065), .ZN(n9137) );
  INV_X1 U6499 ( .A(n9654), .ZN(n9382) );
  AND2_X1 U6500 ( .A1(n7626), .A2(n9652), .ZN(n9384) );
  NOR2_X1 U6501 ( .A1(n9661), .A2(n9384), .ZN(n9437) );
  INV_X1 U6502 ( .A(n9384), .ZN(n9650) );
  NAND2_X1 U6503 ( .A1(n6504), .A2(n6503), .ZN(n9610) );
  NOR2_X1 U6504 ( .A1(n6183), .A2(n6218), .ZN(n7012) );
  AND2_X1 U6505 ( .A1(n6107), .A2(n6087), .ZN(n6802) );
  XNOR2_X1 U6506 ( .A(n5866), .B(n5865), .ZN(n6815) );
  INV_X1 U6507 ( .A(n8047), .ZN(n8065) );
  INV_X1 U6508 ( .A(n8012), .ZN(n8265) );
  OR2_X1 U6509 ( .A1(n9668), .A2(n6711), .ZN(n9699) );
  OR2_X1 U6510 ( .A1(n9668), .A2(n8118), .ZN(n9845) );
  NAND2_X1 U6511 ( .A1(n9929), .A2(n9907), .ZN(n8352) );
  AND2_X1 U6512 ( .A1(n6622), .A2(n6577), .ZN(n8378) );
  NAND2_X1 U6513 ( .A1(n9929), .A2(n9914), .ZN(n8381) );
  INV_X1 U6514 ( .A(n9927), .ZN(n9929) );
  NOR2_X1 U6515 ( .A1(n5048), .A2(n5040), .ZN(n5961) );
  NAND2_X1 U6516 ( .A1(n9915), .A2(n9914), .ZN(n8470) );
  AND2_X1 U6517 ( .A1(n5960), .A2(n5959), .ZN(n9917) );
  INV_X1 U6518 ( .A(n9963), .ZN(n6663) );
  AND2_X1 U6519 ( .A1(n5875), .A2(n6815), .ZN(n6660) );
  INV_X1 U6520 ( .A(n5935), .ZN(n7871) );
  INV_X1 U6521 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7349) );
  INV_X1 U6522 ( .A(n9713), .ZN(n8130) );
  NAND2_X1 U6523 ( .A1(n6559), .A2(n6552), .ZN(n6553) );
  INV_X1 U6524 ( .A(n7730), .ZN(n7862) );
  INV_X1 U6525 ( .A(n9329), .ZN(n9165) );
  INV_X1 U6526 ( .A(n9497), .ZN(n8651) );
  NAND2_X1 U6527 ( .A1(n6483), .A2(n6482), .ZN(n8921) );
  NAND2_X1 U6528 ( .A1(n6463), .A2(n6462), .ZN(n8922) );
  OR2_X1 U6529 ( .A1(n6306), .A2(n6305), .ZN(n9028) );
  INV_X1 U6530 ( .A(n9547), .ZN(n9585) );
  NAND2_X1 U6531 ( .A1(n9667), .A2(n9382), .ZN(n9367) );
  INV_X2 U6532 ( .A(n9665), .ZN(n9667) );
  NAND2_X1 U6533 ( .A1(n9439), .A2(n9382), .ZN(n9444) );
  INV_X1 U6534 ( .A(n9437), .ZN(n9449) );
  OR2_X1 U6535 ( .A1(n7121), .A2(n7120), .ZN(n9661) );
  AND2_X1 U6536 ( .A1(n6508), .A2(n6021), .ZN(n9638) );
  INV_X1 U6537 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7872) );
  INV_X1 U6538 ( .A(n9462), .ZN(n9466) );
  AND2_X1 U6539 ( .A1(n6639), .A2(n6815), .ZN(P2_U3893) );
  NAND2_X1 U6540 ( .A1(n6593), .A2(n6592), .ZN(P2_U3487) );
  NOR2_X1 U6541 ( .A1(n6665), .A2(n4437), .ZN(P1_U3973) );
  MUX2_X1 U6542 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5060), .Z(n5055) );
  NAND2_X1 U6543 ( .A1(n5055), .A2(SI_2_), .ZN(n5065) );
  INV_X1 U6544 ( .A(n5304), .ZN(n5064) );
  INV_X1 U6545 ( .A(SI_1_), .ZN(n5056) );
  NAND2_X1 U6546 ( .A1(n5057), .A2(n5056), .ZN(n5059) );
  NAND2_X1 U6547 ( .A1(n5058), .A2(SI_1_), .ZN(n5063) );
  INV_X1 U6548 ( .A(n5272), .ZN(n5062) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10265) );
  INV_X1 U6550 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6551 ( .A1(n5066), .A2(SI_3_), .ZN(n5069) );
  INV_X1 U6552 ( .A(n5066), .ZN(n5068) );
  INV_X1 U6553 ( .A(SI_3_), .ZN(n5067) );
  NAND2_X1 U6554 ( .A1(n5070), .A2(SI_4_), .ZN(n5074) );
  INV_X1 U6555 ( .A(n5070), .ZN(n5072) );
  INV_X1 U6556 ( .A(SI_4_), .ZN(n5071) );
  NAND2_X1 U6557 ( .A1(n5072), .A2(n5071), .ZN(n5073) );
  AND2_X1 U6558 ( .A1(n5074), .A2(n5073), .ZN(n5336) );
  NAND2_X1 U6559 ( .A1(n5075), .A2(SI_5_), .ZN(n5079) );
  INV_X1 U6560 ( .A(n5075), .ZN(n5077) );
  INV_X1 U6561 ( .A(SI_5_), .ZN(n5076) );
  NAND2_X1 U6562 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  NAND2_X1 U6563 ( .A1(n5080), .A2(SI_6_), .ZN(n5384) );
  OAI21_X1 U6564 ( .B1(n5080), .B2(SI_6_), .A(n5384), .ZN(n5362) );
  INV_X1 U6565 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5081) );
  INV_X1 U6566 ( .A(SI_7_), .ZN(n5082) );
  NAND2_X1 U6567 ( .A1(n5083), .A2(n5082), .ZN(n5386) );
  INV_X1 U6568 ( .A(n5386), .ZN(n5088) );
  XNOR2_X1 U6569 ( .A(n5089), .B(SI_8_), .ZN(n5403) );
  INV_X1 U6570 ( .A(n5403), .ZN(n5085) );
  INV_X1 U6571 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6572 ( .A1(n5084), .A2(SI_7_), .ZN(n5401) );
  OAI211_X1 U6573 ( .C1(n5088), .C2(n5384), .A(n5085), .B(n5401), .ZN(n5086)
         );
  INV_X1 U6574 ( .A(n5086), .ZN(n5087) );
  OAI21_X1 U6575 ( .B1(n5385), .B2(n5088), .A(n5087), .ZN(n5093) );
  INV_X1 U6576 ( .A(n5089), .ZN(n5091) );
  INV_X1 U6577 ( .A(SI_8_), .ZN(n5090) );
  NAND2_X1 U6578 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  NAND2_X1 U6579 ( .A1(n5093), .A2(n5092), .ZN(n5416) );
  MUX2_X1 U6580 ( .A(n6686), .B(n5094), .S(n6640), .Z(n5096) );
  XNOR2_X1 U6581 ( .A(n5096), .B(SI_9_), .ZN(n5415) );
  NAND2_X1 U6582 ( .A1(n5416), .A2(n5415), .ZN(n5098) );
  INV_X1 U6583 ( .A(SI_9_), .ZN(n5095) );
  NAND2_X1 U6584 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  NAND2_X1 U6585 ( .A1(n5098), .A2(n5097), .ZN(n5431) );
  INV_X1 U6586 ( .A(n5431), .ZN(n5101) );
  NAND2_X1 U6587 ( .A1(n5099), .A2(SI_10_), .ZN(n5102) );
  OAI21_X1 U6588 ( .B1(n5099), .B2(SI_10_), .A(n5102), .ZN(n5430) );
  XNOR2_X1 U6589 ( .A(n5103), .B(SI_11_), .ZN(n5449) );
  MUX2_X1 U6590 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6640), .Z(n5104) );
  NAND2_X1 U6591 ( .A1(n5104), .A2(SI_12_), .ZN(n5105) );
  OAI21_X1 U6592 ( .B1(n5104), .B2(SI_12_), .A(n5105), .ZN(n5469) );
  MUX2_X1 U6593 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6640), .Z(n5106) );
  INV_X1 U6594 ( .A(n5106), .ZN(n5108) );
  INV_X1 U6595 ( .A(SI_13_), .ZN(n5107) );
  NAND2_X1 U6596 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  MUX2_X1 U6597 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6640), .Z(n5490) );
  MUX2_X1 U6598 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6640), .Z(n5505) );
  INV_X1 U6599 ( .A(n5505), .ZN(n5111) );
  NAND2_X1 U6600 ( .A1(n5112), .A2(n5111), .ZN(n5115) );
  NAND2_X1 U6601 ( .A1(n5113), .A2(n4895), .ZN(n5114) );
  MUX2_X1 U6602 ( .A(n10282), .B(n5116), .S(n6640), .Z(n5522) );
  NAND2_X1 U6603 ( .A1(n5117), .A2(SI_16_), .ZN(n5118) );
  MUX2_X1 U6604 ( .A(n7349), .B(n7347), .S(n6640), .Z(n5120) );
  INV_X1 U6605 ( .A(n5120), .ZN(n5121) );
  NAND2_X1 U6606 ( .A1(n5121), .A2(SI_17_), .ZN(n5122) );
  NAND2_X1 U6607 ( .A1(n5123), .A2(n5122), .ZN(n5540) );
  NAND2_X1 U6608 ( .A1(n5124), .A2(n5123), .ZN(n5555) );
  MUX2_X1 U6609 ( .A(n10138), .B(n5125), .S(n6640), .Z(n5126) );
  XNOR2_X1 U6610 ( .A(n5126), .B(SI_18_), .ZN(n5554) );
  INV_X1 U6611 ( .A(n5554), .ZN(n5129) );
  INV_X1 U6612 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6613 ( .A1(n5127), .A2(SI_18_), .ZN(n5128) );
  MUX2_X1 U6614 ( .A(n7584), .B(n10201), .S(n6640), .Z(n5131) );
  INV_X1 U6615 ( .A(SI_19_), .ZN(n5130) );
  NAND2_X1 U6616 ( .A1(n5131), .A2(n5130), .ZN(n5134) );
  INV_X1 U6617 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6618 ( .A1(n5132), .A2(SI_19_), .ZN(n5133) );
  NAND2_X1 U6619 ( .A1(n5134), .A2(n5133), .ZN(n5572) );
  MUX2_X1 U6620 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6640), .Z(n5586) );
  INV_X1 U6621 ( .A(n5586), .ZN(n5135) );
  NAND2_X1 U6622 ( .A1(n5588), .A2(n5585), .ZN(n5136) );
  MUX2_X1 U6623 ( .A(n10029), .B(n10193), .S(n6640), .Z(n5602) );
  NOR2_X1 U6624 ( .A1(n5138), .A2(SI_21_), .ZN(n5140) );
  NAND2_X1 U6625 ( .A1(n5138), .A2(SI_21_), .ZN(n5139) );
  MUX2_X1 U6626 ( .A(n7776), .B(n10111), .S(n6640), .Z(n5142) );
  NAND2_X1 U6627 ( .A1(n5142), .A2(n5141), .ZN(n5145) );
  INV_X1 U6628 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6629 ( .A1(n5143), .A2(SI_22_), .ZN(n5144) );
  NAND2_X1 U6630 ( .A1(n5145), .A2(n5144), .ZN(n5616) );
  INV_X1 U6631 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5147) );
  INV_X1 U6632 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5146) );
  MUX2_X1 U6633 ( .A(n5147), .B(n5146), .S(n6640), .Z(n5149) );
  INV_X1 U6634 ( .A(SI_23_), .ZN(n5148) );
  NAND2_X1 U6635 ( .A1(n5149), .A2(n5148), .ZN(n5152) );
  INV_X1 U6636 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6637 ( .A1(n5150), .A2(SI_23_), .ZN(n5151) );
  INV_X1 U6638 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7864) );
  INV_X1 U6639 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7866) );
  MUX2_X1 U6640 ( .A(n7864), .B(n7866), .S(n6640), .Z(n5153) );
  NAND2_X1 U6641 ( .A1(n5153), .A2(n10245), .ZN(n5156) );
  INV_X1 U6642 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6643 ( .A1(n5154), .A2(SI_24_), .ZN(n5155) );
  NAND2_X1 U6644 ( .A1(n5645), .A2(n5644), .ZN(n5157) );
  INV_X1 U6645 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7870) );
  MUX2_X1 U6646 ( .A(n7870), .B(n7872), .S(n6640), .Z(n5159) );
  INV_X1 U6647 ( .A(SI_25_), .ZN(n5158) );
  NAND2_X1 U6648 ( .A1(n5159), .A2(n5158), .ZN(n5162) );
  INV_X1 U6649 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6650 ( .A1(n5160), .A2(SI_25_), .ZN(n5161) );
  NAND2_X1 U6651 ( .A1(n5662), .A2(n5661), .ZN(n5163) );
  INV_X1 U6652 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7876) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10183) );
  MUX2_X1 U6654 ( .A(n7876), .B(n10183), .S(n6640), .Z(n5165) );
  INV_X1 U6655 ( .A(SI_26_), .ZN(n5164) );
  NAND2_X1 U6656 ( .A1(n5165), .A2(n5164), .ZN(n5168) );
  INV_X1 U6657 ( .A(n5165), .ZN(n5166) );
  NAND2_X1 U6658 ( .A1(n5166), .A2(SI_26_), .ZN(n5167) );
  NAND2_X1 U6659 ( .A1(n5674), .A2(n5673), .ZN(n5169) );
  INV_X1 U6660 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5171) );
  INV_X1 U6661 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5170) );
  MUX2_X1 U6662 ( .A(n5171), .B(n5170), .S(n6640), .Z(n5173) );
  INV_X1 U6663 ( .A(SI_27_), .ZN(n5172) );
  NAND2_X1 U6664 ( .A1(n5173), .A2(n5172), .ZN(n5176) );
  INV_X1 U6665 ( .A(n5173), .ZN(n5174) );
  NAND2_X1 U6666 ( .A1(n5174), .A2(SI_27_), .ZN(n5175) );
  NAND2_X1 U6667 ( .A1(n5687), .A2(n5686), .ZN(n5177) );
  INV_X1 U6668 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5178) );
  MUX2_X1 U6669 ( .A(n10054), .B(n5178), .S(n6640), .Z(n5180) );
  XNOR2_X1 U6670 ( .A(n5180), .B(SI_28_), .ZN(n5712) );
  INV_X1 U6671 ( .A(SI_28_), .ZN(n5179) );
  NAND2_X1 U6672 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  INV_X1 U6673 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10095) );
  INV_X1 U6674 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5182) );
  MUX2_X1 U6675 ( .A(n10095), .B(n5182), .S(n6640), .Z(n5726) );
  NOR2_X2 U6676 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5183) );
  NAND4_X1 U6677 ( .A1(n5183), .A2(n10121), .A3(n5493), .A4(n5508), .ZN(n5187)
         );
  INV_X2 U6678 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5257) );
  NAND4_X1 U6679 ( .A1(n5255), .A2(n5257), .A3(n5185), .A4(n5184), .ZN(n5186)
         );
  NOR2_X2 U6680 ( .A1(n5187), .A2(n5186), .ZN(n5525) );
  NOR2_X1 U6681 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5194) );
  NOR2_X1 U6682 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5193) );
  NOR2_X1 U6683 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5192) );
  OR2_X2 U6684 ( .A1(n5227), .A2(n8473), .ZN(n5231) );
  XNOR2_X2 U6685 ( .A(n5231), .B(n5196), .ZN(n5876) );
  INV_X1 U6686 ( .A(n5197), .ZN(n5198) );
  NAND2_X1 U6687 ( .A1(n7888), .A2(n5751), .ZN(n5201) );
  NAND2_X1 U6688 ( .A1(n5688), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6689 ( .A1(n5203), .A2(n5202), .ZN(n5369) );
  INV_X1 U6690 ( .A(n5369), .ZN(n5205) );
  NOR2_X1 U6691 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5204) );
  NAND2_X1 U6692 ( .A1(n5205), .A2(n5204), .ZN(n5394) );
  INV_X1 U6693 ( .A(n5438), .ZN(n5209) );
  INV_X1 U6694 ( .A(n5498), .ZN(n5213) );
  INV_X1 U6695 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5219) );
  INV_X1 U6696 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10120) );
  INV_X1 U6697 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5222) );
  INV_X1 U6698 ( .A(n5705), .ZN(n5225) );
  INV_X1 U6699 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6700 ( .A1(n5225), .A2(n5224), .ZN(n7878) );
  NOR2_X1 U6701 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5226) );
  NAND2_X1 U6702 ( .A1(n5227), .A2(n5226), .ZN(n8474) );
  INV_X1 U6703 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5228) );
  XNOR2_X2 U6704 ( .A(n5229), .B(n5228), .ZN(n5235) );
  NAND2_X1 U6705 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5230) );
  NAND2_X1 U6706 ( .A1(n5231), .A2(n5230), .ZN(n5233) );
  XNOR2_X2 U6707 ( .A(n5233), .B(n5232), .ZN(n5234) );
  OR2_X1 U6708 ( .A1(n7878), .A2(n5296), .ZN(n5761) );
  INV_X1 U6709 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7880) );
  INV_X1 U6710 ( .A(n5234), .ZN(n8479) );
  NAND2_X1 U6711 ( .A1(n5283), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6712 ( .A1(n8479), .A2(n5235), .ZN(n5284) );
  NAND2_X1 U6713 ( .A1(n5667), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5237) );
  OAI211_X1 U6714 ( .C1(n7880), .C2(n5757), .A(n5238), .B(n5237), .ZN(n5239)
         );
  INV_X1 U6715 ( .A(n5239), .ZN(n5240) );
  BUF_X1 U6716 ( .A(n5241), .Z(n5542) );
  NAND2_X1 U6717 ( .A1(n5558), .A2(n5575), .ZN(n5242) );
  NOR2_X2 U6718 ( .A1(n5556), .A2(n5242), .ZN(n5762) );
  NAND2_X1 U6719 ( .A1(n5762), .A2(n5764), .ZN(n5244) );
  NAND2_X1 U6720 ( .A1(n5864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6721 ( .A1(n5244), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5245) );
  MUX2_X1 U6722 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5245), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5246) );
  NAND2_X1 U6723 ( .A1(n7961), .A2(n5929), .ZN(n5247) );
  INV_X1 U6724 ( .A(n7885), .ZN(n6579) );
  OR2_X1 U6725 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  NAND2_X1 U6726 ( .A1(n5251), .A2(n5250), .ZN(n6977) );
  INV_X2 U6727 ( .A(n5275), .ZN(n5473) );
  NAND2_X1 U6728 ( .A1(n5340), .A2(n5252), .ZN(n5353) );
  NAND2_X1 U6729 ( .A1(n5364), .A2(n5253), .ZN(n5527) );
  INV_X1 U6730 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6731 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NAND2_X1 U6732 ( .A1(n5474), .A2(n5257), .ZN(n5258) );
  NAND2_X1 U6733 ( .A1(n5258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5494) );
  XNOR2_X1 U6734 ( .A(n5494), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U6735 ( .A1(n5688), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5577), .B2(
        n9764), .ZN(n5259) );
  INV_X1 U6736 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10242) );
  OR2_X1 U6737 ( .A1(n4439), .A2(n10242), .ZN(n5265) );
  INV_X1 U6738 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10217) );
  OR2_X1 U6739 ( .A1(n5236), .A2(n10217), .ZN(n5264) );
  NAND2_X1 U6740 ( .A1(n5480), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5261) );
  AND2_X1 U6741 ( .A1(n5498), .A2(n5261), .ZN(n8332) );
  OR2_X1 U6742 ( .A1(n4438), .A2(n8332), .ZN(n5263) );
  NAND2_X1 U6743 ( .A1(n5282), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5262) );
  NAND4_X1 U6744 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n8313)
         );
  INV_X1 U6745 ( .A(n8313), .ZN(n5784) );
  MUX2_X1 U6746 ( .A(n8334), .B(n5784), .S(n5929), .Z(n5487) );
  AND2_X1 U6747 ( .A1(n8467), .A2(n8313), .ZN(n8308) );
  INV_X1 U6748 ( .A(n8308), .ZN(n5830) );
  INV_X1 U6749 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6706) );
  INV_X1 U6750 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6705) );
  INV_X1 U6751 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6752 ( .A1(n5284), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U6753 ( .A1(n5272), .A2(n4553), .ZN(n5273) );
  NAND2_X1 U6754 ( .A1(n5274), .A2(n5273), .ZN(n6652) );
  NAND2_X1 U6755 ( .A1(n5275), .A2(n6652), .ZN(n5281) );
  NAND2_X1 U6756 ( .A1(n5322), .A2(n4906), .ZN(n5280) );
  INV_X1 U6757 ( .A(n5276), .ZN(n5326) );
  INV_X1 U6758 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6759 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5277) );
  NAND2_X1 U6760 ( .A1(n5326), .A2(n6719), .ZN(n5279) );
  INV_X1 U6761 ( .A(n5768), .ZN(n5294) );
  NAND2_X1 U6762 ( .A1(n5282), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5287) );
  INV_X1 U6763 ( .A(n5284), .ZN(n5314) );
  NAND2_X1 U6764 ( .A1(n5314), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5285) );
  AND3_X1 U6765 ( .A1(n5287), .A2(n5286), .A3(n5285), .ZN(n5290) );
  NAND2_X1 U6766 ( .A1(n5288), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6767 ( .A1(n6643), .A2(SI_0_), .ZN(n5291) );
  XNOR2_X1 U6768 ( .A(n5291), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8491) );
  MUX2_X1 U6769 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8491), .S(n5276), .Z(n6829) );
  AND2_X1 U6770 ( .A1(n8080), .A2(n6992), .ZN(n5835) );
  OAI21_X1 U6771 ( .B1(n5835), .B2(n4808), .A(n6979), .ZN(n5292) );
  AOI21_X1 U6772 ( .B1(n5292), .B2(n5295), .A(n5294), .ZN(n5293) );
  MUX2_X1 U6773 ( .A(n5294), .B(n5293), .S(n6636), .Z(n5313) );
  NOR3_X1 U6774 ( .A1(n5769), .A2(n5835), .A3(n6636), .ZN(n5312) );
  NAND2_X1 U6775 ( .A1(n5314), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5302) );
  INV_X1 U6776 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9856) );
  OR2_X1 U6777 ( .A1(n4438), .A2(n9856), .ZN(n5301) );
  INV_X1 U6778 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6762) );
  OR2_X1 U6779 ( .A1(n5297), .A2(n6762), .ZN(n5300) );
  INV_X1 U6780 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6732) );
  OR2_X1 U6781 ( .A1(n4439), .A2(n6732), .ZN(n5299) );
  AND4_X2 U6782 ( .A1(n5302), .A2(n5301), .A3(n5300), .A4(n5299), .ZN(n7073)
         );
  INV_X1 U6783 ( .A(n5303), .ZN(n5305) );
  NAND2_X1 U6784 ( .A1(n5305), .A2(n5304), .ZN(n5307) );
  NAND2_X1 U6785 ( .A1(n5307), .A2(n5306), .ZN(n6647) );
  NAND2_X1 U6786 ( .A1(n5322), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5311) );
  INV_X2 U6787 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8473) );
  NOR2_X1 U6788 ( .A1(n6701), .A2(n8473), .ZN(n5308) );
  NAND2_X1 U6789 ( .A1(n5326), .A2(n6763), .ZN(n5310) );
  NAND2_X1 U6790 ( .A1(n7073), .A2(n9852), .ZN(n5770) );
  NOR3_X1 U6791 ( .A1(n5313), .A2(n5312), .A3(n5884), .ZN(n5345) );
  OR2_X1 U6792 ( .A1(n4438), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6793 ( .A1(n5314), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6794 ( .A1(n5282), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6795 ( .A1(n5283), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6796 ( .A1(n5321), .A2(n5320), .ZN(n6645) );
  NAND2_X1 U6797 ( .A1(n5322), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5328) );
  NOR2_X1 U6798 ( .A1(n5323), .A2(n8473), .ZN(n5324) );
  MUX2_X1 U6799 ( .A(n8473), .B(n5324), .S(P2_IR_REG_3__SCAN_IN), .Z(n5325) );
  NAND2_X1 U6800 ( .A1(n5326), .A2(n9684), .ZN(n5327) );
  OAI211_X1 U6801 ( .C1(n5473), .C2(n6645), .A(n5328), .B(n5327), .ZN(n6974)
         );
  NAND2_X1 U6802 ( .A1(n9862), .A2(n6974), .ZN(n5771) );
  INV_X1 U6803 ( .A(n6974), .ZN(n7271) );
  NAND2_X1 U6804 ( .A1(n8077), .A2(n7271), .ZN(n5767) );
  NAND2_X1 U6805 ( .A1(n5767), .A2(n5329), .ZN(n5330) );
  NAND2_X1 U6806 ( .A1(n5283), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6807 ( .A1(n5314), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6808 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5331) );
  AND2_X1 U6809 ( .A1(n5369), .A2(n5331), .ZN(n7099) );
  OR2_X1 U6810 ( .A1(n4438), .A2(n7099), .ZN(n5333) );
  NAND2_X1 U6811 ( .A1(n5282), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5332) );
  NAND4_X1 U6812 ( .A1(n5335), .A2(n5334), .A3(n5333), .A4(n5332), .ZN(n8076)
         );
  OR2_X1 U6813 ( .A1(n5337), .A2(n5336), .ZN(n5338) );
  NAND2_X1 U6814 ( .A1(n5339), .A2(n5338), .ZN(n6657) );
  NAND2_X1 U6815 ( .A1(n5688), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5343) );
  OR2_X1 U6816 ( .A1(n5340), .A2(n8473), .ZN(n5341) );
  NAND2_X1 U6817 ( .A1(n5577), .A2(n6905), .ZN(n5342) );
  OAI211_X1 U6818 ( .C1(n5473), .C2(n6657), .A(n5343), .B(n5342), .ZN(n7211)
         );
  NAND2_X1 U6819 ( .A1(n5889), .A2(n7211), .ZN(n5773) );
  INV_X1 U6820 ( .A(n7211), .ZN(n9879) );
  NAND2_X1 U6821 ( .A1(n8076), .A2(n9879), .ZN(n5772) );
  AND2_X1 U6822 ( .A1(n5773), .A2(n5772), .ZN(n7206) );
  OAI21_X1 U6823 ( .B1(n5345), .B2(n5344), .A(n7206), .ZN(n5378) );
  INV_X1 U6824 ( .A(n5767), .ZN(n5361) );
  NAND2_X1 U6825 ( .A1(n5283), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5352) );
  INV_X1 U6826 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5346) );
  OR2_X1 U6827 ( .A1(n5236), .A2(n5346), .ZN(n5351) );
  INV_X1 U6828 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5347) );
  XNOR2_X1 U6829 ( .A(n5369), .B(n5347), .ZN(n7310) );
  OR2_X1 U6830 ( .A1(n4438), .A2(n7310), .ZN(n5350) );
  INV_X1 U6831 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5348) );
  OR2_X1 U6832 ( .A1(n5757), .A2(n5348), .ZN(n5349) );
  NAND2_X1 U6833 ( .A1(n5353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5354) );
  AOI22_X1 U6834 ( .A1(n5688), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5577), .B2(
        n7159), .ZN(n5360) );
  OR2_X1 U6835 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6836 ( .A1(n5358), .A2(n5357), .ZN(n6654) );
  OR2_X1 U6837 ( .A1(n6654), .A2(n5473), .ZN(n5359) );
  NAND2_X1 U6838 ( .A1(n5360), .A2(n5359), .ZN(n7312) );
  NAND2_X1 U6839 ( .A1(n7258), .A2(n7312), .ZN(n5834) );
  OAI211_X1 U6840 ( .C1(n5378), .C2(n5361), .A(n5834), .B(n5773), .ZN(n5375)
         );
  XNOR2_X1 U6841 ( .A(n5363), .B(n5362), .ZN(n6675) );
  NAND2_X1 U6842 ( .A1(n6675), .A2(n5751), .ZN(n5367) );
  OR2_X1 U6843 ( .A1(n5364), .A2(n8473), .ZN(n5365) );
  AOI22_X1 U6844 ( .A1(n5688), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5577), .B2(
        n7161), .ZN(n5366) );
  NAND2_X1 U6845 ( .A1(n5367), .A2(n5366), .ZN(n9892) );
  NAND2_X1 U6846 ( .A1(n5283), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5374) );
  INV_X1 U6847 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5368) );
  OR2_X1 U6848 ( .A1(n5236), .A2(n5368), .ZN(n5373) );
  OAI21_X1 U6849 ( .B1(n5369), .B2(P2_REG3_REG_5__SCAN_IN), .A(
        P2_REG3_REG_6__SCAN_IN), .ZN(n5370) );
  AND2_X1 U6850 ( .A1(n5370), .A2(n5394), .ZN(n7264) );
  OR2_X1 U6851 ( .A1(n4438), .A2(n7264), .ZN(n5372) );
  INV_X1 U6852 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7407) );
  OR2_X1 U6853 ( .A1(n5297), .A2(n7407), .ZN(n5371) );
  OR2_X1 U6854 ( .A1(n9892), .A2(n7463), .ZN(n5838) );
  INV_X1 U6855 ( .A(n7312), .ZN(n9883) );
  NAND2_X1 U6856 ( .A1(n9883), .A2(n8075), .ZN(n5833) );
  NAND3_X1 U6857 ( .A1(n5375), .A2(n5838), .A3(n5833), .ZN(n5376) );
  AND2_X1 U6858 ( .A1(n9892), .A2(n7463), .ZN(n5839) );
  INV_X1 U6859 ( .A(n5839), .ZN(n5379) );
  NAND2_X1 U6860 ( .A1(n5376), .A2(n5379), .ZN(n5383) );
  INV_X1 U6861 ( .A(n5771), .ZN(n5377) );
  OAI211_X1 U6862 ( .C1(n5378), .C2(n5377), .A(n5833), .B(n5772), .ZN(n5380)
         );
  NAND3_X1 U6863 ( .A1(n5380), .A2(n5379), .A3(n5834), .ZN(n5381) );
  NAND2_X1 U6864 ( .A1(n5381), .A2(n5838), .ZN(n5382) );
  MUX2_X1 U6865 ( .A(n5383), .B(n5382), .S(n5929), .Z(n5414) );
  NAND2_X1 U6866 ( .A1(n5385), .A2(n5384), .ZN(n5388) );
  AND2_X1 U6867 ( .A1(n5386), .A2(n5401), .ZN(n5387) );
  OR2_X1 U6868 ( .A1(n6679), .A2(n5473), .ZN(n5392) );
  NAND2_X1 U6869 ( .A1(n5527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5389) );
  MUX2_X1 U6870 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5389), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5390) );
  AOI22_X1 U6871 ( .A1(n5688), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5577), .B2(
        n7233), .ZN(n5391) );
  NAND2_X1 U6872 ( .A1(n5392), .A2(n5391), .ZN(n9896) );
  NAND2_X1 U6873 ( .A1(n5283), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5400) );
  INV_X1 U6874 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5393) );
  OR2_X1 U6875 ( .A1(n5236), .A2(n5393), .ZN(n5399) );
  NAND2_X1 U6876 ( .A1(n5394), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5395) );
  AND2_X1 U6877 ( .A1(n5408), .A2(n5395), .ZN(n7468) );
  OR2_X1 U6878 ( .A1(n4438), .A2(n7468), .ZN(n5398) );
  INV_X1 U6879 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5396) );
  OR2_X1 U6880 ( .A1(n5757), .A2(n5396), .ZN(n5397) );
  OR2_X1 U6881 ( .A1(n9896), .A2(n7598), .ZN(n7599) );
  NAND2_X1 U6882 ( .A1(n9896), .A2(n7598), .ZN(n5444) );
  NAND2_X1 U6883 ( .A1(n5402), .A2(n5401), .ZN(n5404) );
  NAND2_X1 U6884 ( .A1(n6680), .A2(n5751), .ZN(n5407) );
  NAND2_X1 U6885 ( .A1(n5417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5405) );
  AOI22_X1 U6886 ( .A1(n5688), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5577), .B2(
        n7338), .ZN(n5406) );
  NAND2_X1 U6887 ( .A1(n5667), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5413) );
  INV_X1 U6888 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7230) );
  OR2_X1 U6889 ( .A1(n4439), .A2(n7230), .ZN(n5412) );
  NAND2_X1 U6890 ( .A1(n5408), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5409) );
  AND2_X1 U6891 ( .A1(n5423), .A2(n5409), .ZN(n7603) );
  OR2_X1 U6892 ( .A1(n4438), .A2(n7603), .ZN(n5411) );
  INV_X1 U6893 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7604) );
  OR2_X1 U6894 ( .A1(n5757), .A2(n7604), .ZN(n5410) );
  AND2_X1 U6895 ( .A1(n5843), .A2(n7599), .ZN(n5777) );
  OAI22_X1 U6896 ( .A1(n5414), .A2(n5892), .B1(n5929), .B2(n5777), .ZN(n5463)
         );
  NAND2_X1 U6897 ( .A1(n6685), .A2(n5751), .ZN(n5422) );
  NAND2_X1 U6898 ( .A1(n5418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5419) );
  OR2_X1 U6899 ( .A1(n5419), .A2(n10121), .ZN(n5420) );
  NAND2_X1 U6900 ( .A1(n5419), .A2(n10121), .ZN(n5434) );
  AOI22_X1 U6901 ( .A1(n5688), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5577), .B2(
        n8133), .ZN(n5421) );
  NAND2_X1 U6902 ( .A1(n5283), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6903 ( .A1(n5667), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6904 ( .A1(n5423), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5424) );
  AND2_X1 U6905 ( .A1(n5438), .A2(n5424), .ZN(n7616) );
  OR2_X1 U6906 ( .A1(n4438), .A2(n7616), .ZN(n5426) );
  NAND2_X1 U6907 ( .A1(n5282), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5425) );
  NAND4_X1 U6908 ( .A1(n5428), .A2(n5427), .A3(n5426), .A4(n5425), .ZN(n7650)
         );
  NAND2_X1 U6909 ( .A1(n9906), .A2(n7705), .ZN(n5778) );
  OR2_X1 U6910 ( .A1(n9906), .A2(n7705), .ZN(n7706) );
  NAND2_X1 U6911 ( .A1(n5429), .A2(n7706), .ZN(n5446) );
  INV_X1 U6912 ( .A(n5446), .ZN(n5462) );
  NAND2_X1 U6913 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  NAND2_X1 U6914 ( .A1(n5433), .A2(n5432), .ZN(n6690) );
  OR2_X1 U6915 ( .A1(n6690), .A2(n5473), .ZN(n5437) );
  NAND2_X1 U6916 ( .A1(n5434), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5435) );
  AOI22_X1 U6917 ( .A1(n5688), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5577), .B2(
        n9713), .ZN(n5436) );
  NAND2_X1 U6918 ( .A1(n5283), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6919 ( .A1(n5438), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5439) );
  AND2_X1 U6920 ( .A1(n5456), .A2(n5439), .ZN(n7710) );
  OR2_X1 U6921 ( .A1(n4438), .A2(n7710), .ZN(n5442) );
  INV_X1 U6922 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8083) );
  OR2_X1 U6923 ( .A1(n5757), .A2(n8083), .ZN(n5441) );
  NAND2_X1 U6924 ( .A1(n5667), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5440) );
  NAND4_X1 U6925 ( .A1(n5443), .A2(n5442), .A3(n5441), .A4(n5440), .ZN(n8073)
         );
  INV_X1 U6926 ( .A(n8073), .ZN(n7754) );
  OR2_X1 U6927 ( .A1(n7653), .A2(n7754), .ZN(n5832) );
  INV_X1 U6928 ( .A(n5780), .ZN(n5448) );
  AND2_X1 U6929 ( .A1(n5842), .A2(n5444), .ZN(n5445) );
  NAND2_X1 U6930 ( .A1(n7653), .A2(n7754), .ZN(n5831) );
  OAI211_X1 U6931 ( .C1(n5446), .C2(n5445), .A(n5778), .B(n5831), .ZN(n5447)
         );
  XNOR2_X1 U6932 ( .A(n5450), .B(n5449), .ZN(n6779) );
  NAND2_X1 U6933 ( .A1(n6779), .A2(n5751), .ZN(n5454) );
  NAND2_X1 U6934 ( .A1(n5451), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U6935 ( .A(n5452), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9730) );
  AOI22_X1 U6936 ( .A1(n5688), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5577), .B2(
        n9730), .ZN(n5453) );
  NAND2_X1 U6937 ( .A1(n5454), .A2(n5453), .ZN(n7795) );
  NAND2_X1 U6938 ( .A1(n5667), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5461) );
  INV_X1 U6939 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5455) );
  OR2_X1 U6940 ( .A1(n4439), .A2(n5455), .ZN(n5460) );
  NAND2_X1 U6941 ( .A1(n5456), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5457) );
  AND2_X1 U6942 ( .A1(n5478), .A2(n5457), .ZN(n7797) );
  OR2_X1 U6943 ( .A1(n4438), .A2(n7797), .ZN(n5459) );
  INV_X1 U6944 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10262) );
  OR2_X1 U6945 ( .A1(n5757), .A2(n10262), .ZN(n5458) );
  OR2_X1 U6946 ( .A1(n7795), .A2(n7747), .ZN(n5465) );
  NAND2_X1 U6947 ( .A1(n7795), .A2(n7747), .ZN(n5781) );
  NAND2_X1 U6948 ( .A1(n5465), .A2(n5781), .ZN(n7780) );
  INV_X1 U6949 ( .A(n5781), .ZN(n5464) );
  OAI21_X1 U6950 ( .B1(n5464), .B2(n5832), .A(n5465), .ZN(n5468) );
  INV_X1 U6951 ( .A(n5465), .ZN(n5466) );
  AOI21_X1 U6952 ( .B1(n5831), .B2(n5781), .A(n5466), .ZN(n5467) );
  MUX2_X1 U6953 ( .A(n5468), .B(n5467), .S(n6636), .Z(n5485) );
  NAND2_X1 U6954 ( .A1(n5470), .A2(n5469), .ZN(n5472) );
  NAND2_X1 U6955 ( .A1(n5472), .A2(n5471), .ZN(n6888) );
  OR2_X1 U6956 ( .A1(n5474), .A2(n8473), .ZN(n5475) );
  XNOR2_X1 U6957 ( .A(n5475), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U6958 ( .A1(n5688), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5577), .B2(
        n9747), .ZN(n5476) );
  INV_X1 U6959 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7806) );
  OR2_X1 U6960 ( .A1(n5757), .A2(n7806), .ZN(n5484) );
  NAND2_X1 U6961 ( .A1(n5478), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5479) );
  AND2_X1 U6962 ( .A1(n5480), .A2(n5479), .ZN(n7805) );
  OR2_X1 U6963 ( .A1(n4438), .A2(n7805), .ZN(n5483) );
  INV_X1 U6964 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8128) );
  OR2_X1 U6965 ( .A1(n4439), .A2(n8128), .ZN(n5482) );
  NAND2_X1 U6966 ( .A1(n5667), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5481) );
  NAND4_X1 U6967 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n8329)
         );
  XNOR2_X1 U6968 ( .A(n8382), .B(n8022), .ZN(n7808) );
  INV_X1 U6969 ( .A(n7808), .ZN(n7802) );
  OR2_X1 U6970 ( .A1(n8382), .A2(n8022), .ZN(n5783) );
  NAND2_X1 U6971 ( .A1(n8382), .A2(n8022), .ZN(n5486) );
  MUX2_X1 U6972 ( .A(n5783), .B(n5486), .S(n6636), .Z(n5488) );
  NAND2_X1 U6973 ( .A1(n8334), .A2(n5784), .ZN(n8309) );
  AOI21_X1 U6974 ( .B1(n4643), .B2(n5830), .A(n5489), .ZN(n5521) );
  XNOR2_X1 U6975 ( .A(n5490), .B(SI_14_), .ZN(n5491) );
  XNOR2_X1 U6976 ( .A(n5492), .B(n5491), .ZN(n7037) );
  NAND2_X1 U6977 ( .A1(n7037), .A2(n5751), .ZN(n5497) );
  NAND2_X1 U6978 ( .A1(n5494), .A2(n5493), .ZN(n5495) );
  NAND2_X1 U6979 ( .A1(n5495), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5509) );
  XNOR2_X1 U6980 ( .A(n5509), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U6981 ( .A1(n9780), .A2(n5577), .B1(n5688), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5496) );
  INV_X1 U6982 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10169) );
  OR2_X1 U6983 ( .A1(n5236), .A2(n10169), .ZN(n5504) );
  INV_X1 U6984 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10123) );
  OR2_X1 U6985 ( .A1(n4439), .A2(n10123), .ZN(n5503) );
  NAND2_X1 U6986 ( .A1(n5498), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5499) );
  AND2_X1 U6987 ( .A1(n5514), .A2(n5499), .ZN(n8316) );
  OR2_X1 U6988 ( .A1(n4438), .A2(n8316), .ZN(n5502) );
  INV_X1 U6989 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5500) );
  OR2_X1 U6990 ( .A1(n5757), .A2(n5500), .ZN(n5501) );
  NAND4_X1 U6991 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n8327)
         );
  INV_X1 U6992 ( .A(n8327), .ZN(n7899) );
  NAND2_X1 U6993 ( .A1(n8462), .A2(n7899), .ZN(n5787) );
  NAND2_X1 U6994 ( .A1(n5788), .A2(n5787), .ZN(n8311) );
  MUX2_X1 U6995 ( .A(n5788), .B(n5787), .S(n6636), .Z(n5520) );
  XNOR2_X1 U6996 ( .A(n5505), .B(SI_15_), .ZN(n5506) );
  XNOR2_X1 U6997 ( .A(n5507), .B(n5506), .ZN(n7147) );
  NAND2_X1 U6998 ( .A1(n7147), .A2(n5751), .ZN(n5513) );
  NAND2_X1 U6999 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  NAND2_X1 U7000 ( .A1(n5510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5511) );
  XNOR2_X1 U7001 ( .A(n5511), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U7002 ( .A1(n9797), .A2(n5577), .B1(n5688), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5512) );
  INV_X1 U7003 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10060) );
  OR2_X1 U7004 ( .A1(n4439), .A2(n10060), .ZN(n5519) );
  NAND2_X1 U7005 ( .A1(n5514), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5515) );
  AND2_X1 U7006 ( .A1(n5531), .A2(n5515), .ZN(n8056) );
  OR2_X1 U7007 ( .A1(n4438), .A2(n8056), .ZN(n5518) );
  INV_X1 U7008 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9806) );
  OR2_X1 U7009 ( .A1(n5757), .A2(n9806), .ZN(n5517) );
  NAND2_X1 U7010 ( .A1(n5667), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5516) );
  NAND4_X1 U7011 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .ZN(n8314)
         );
  XNOR2_X1 U7012 ( .A(n8457), .B(n8314), .ZN(n8296) );
  OAI211_X1 U7013 ( .C1(n5521), .C2(n8311), .A(n5520), .B(n8296), .ZN(n5539)
         );
  XNOR2_X1 U7014 ( .A(n5522), .B(SI_16_), .ZN(n5523) );
  XNOR2_X1 U7015 ( .A(n5524), .B(n5523), .ZN(n7202) );
  NAND2_X1 U7016 ( .A1(n7202), .A2(n5751), .ZN(n5530) );
  INV_X1 U7017 ( .A(n5525), .ZN(n5526) );
  OAI21_X1 U7018 ( .B1(n5527), .B2(n5526), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5528) );
  XNOR2_X1 U7019 ( .A(n5528), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U7020 ( .A1(n5688), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5577), .B2(
        n9813), .ZN(n5529) );
  NAND2_X1 U7021 ( .A1(n5667), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5536) );
  INV_X1 U7022 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10161) );
  OR2_X1 U7023 ( .A1(n4439), .A2(n10161), .ZN(n5535) );
  NAND2_X1 U7024 ( .A1(n5531), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5532) );
  AND2_X1 U7025 ( .A1(n5546), .A2(n5532), .ZN(n8292) );
  OR2_X1 U7026 ( .A1(n4438), .A2(n8292), .ZN(n5534) );
  INV_X1 U7027 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8291) );
  OR2_X1 U7028 ( .A1(n5757), .A2(n8291), .ZN(n5533) );
  NAND2_X1 U7029 ( .A1(n8451), .A2(n8060), .ZN(n5828) );
  INV_X1 U7030 ( .A(n8314), .ZN(n7935) );
  OR2_X1 U7031 ( .A1(n8457), .A2(n7935), .ZN(n5790) );
  AND2_X1 U7032 ( .A1(n5829), .A2(n5790), .ZN(n5537) );
  NAND2_X1 U7033 ( .A1(n8457), .A2(n7935), .ZN(n5789) );
  MUX2_X1 U7034 ( .A(n5537), .B(n5789), .S(n5929), .Z(n5538) );
  NAND3_X1 U7035 ( .A1(n5539), .A2(n5828), .A3(n5538), .ZN(n5552) );
  XNOR2_X1 U7036 ( .A(n5541), .B(n5540), .ZN(n7346) );
  NAND2_X1 U7037 ( .A1(n7346), .A2(n5751), .ZN(n5545) );
  NAND2_X1 U7038 ( .A1(n5542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5543) );
  XNOR2_X1 U7039 ( .A(n5543), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U7040 ( .A1(n5688), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5577), .B2(
        n9831), .ZN(n5544) );
  NAND2_X1 U7041 ( .A1(n5546), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7042 ( .A1(n5563), .A2(n5547), .ZN(n8280) );
  NAND2_X1 U7043 ( .A1(n5288), .A2(n8280), .ZN(n5551) );
  INV_X1 U7044 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8369) );
  OR2_X1 U7045 ( .A1(n4439), .A2(n8369), .ZN(n5550) );
  INV_X1 U7046 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8443) );
  OR2_X1 U7047 ( .A1(n5236), .A2(n8443), .ZN(n5549) );
  INV_X1 U7048 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9842) );
  OR2_X1 U7049 ( .A1(n5757), .A2(n9842), .ZN(n5548) );
  NAND2_X1 U7050 ( .A1(n8445), .A2(n8284), .ZN(n5793) );
  NAND2_X1 U7051 ( .A1(n5792), .A2(n5793), .ZN(n8275) );
  INV_X1 U7052 ( .A(n8275), .ZN(n8272) );
  NAND2_X1 U7053 ( .A1(n5552), .A2(n8272), .ZN(n5570) );
  INV_X1 U7054 ( .A(n5829), .ZN(n5553) );
  NOR2_X1 U7055 ( .A1(n5570), .A2(n5553), .ZN(n5571) );
  INV_X1 U7056 ( .A(n5828), .ZN(n5569) );
  XNOR2_X1 U7057 ( .A(n5555), .B(n5554), .ZN(n7400) );
  NAND2_X1 U7058 ( .A1(n7400), .A2(n5751), .ZN(n5562) );
  NAND2_X1 U7059 ( .A1(n5556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5559) );
  INV_X1 U7060 ( .A(n5559), .ZN(n5557) );
  NAND2_X1 U7061 ( .A1(n5557), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7062 ( .A1(n5559), .A2(n5558), .ZN(n5574) );
  AND2_X1 U7063 ( .A1(n5560), .A2(n5574), .ZN(n9477) );
  AOI22_X1 U7064 ( .A1(n5688), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5577), .B2(
        n9477), .ZN(n5561) );
  INV_X1 U7065 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U7066 ( .A1(n5563), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7067 ( .A1(n5580), .A2(n5564), .ZN(n8269) );
  NAND2_X1 U7068 ( .A1(n8269), .A2(n5288), .ZN(n5568) );
  NAND2_X1 U7069 ( .A1(n5667), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5566) );
  INV_X1 U7070 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10228) );
  OR2_X1 U7071 ( .A1(n4439), .A2(n10228), .ZN(n5565) );
  AND2_X1 U7072 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  OAI211_X1 U7073 ( .C1(n5757), .C2(n8268), .A(n5568), .B(n5567), .ZN(n8277)
         );
  INV_X1 U7074 ( .A(n8277), .ZN(n7906) );
  XNOR2_X1 U7075 ( .A(n5573), .B(n5572), .ZN(n7583) );
  NAND2_X1 U7076 ( .A1(n7583), .A2(n5751), .ZN(n5579) );
  NAND2_X1 U7077 ( .A1(n5574), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5576) );
  AOI22_X1 U7078 ( .A1(n5688), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8096), .B2(
        n5577), .ZN(n5578) );
  NAND2_X1 U7079 ( .A1(n5580), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7080 ( .A1(n5591), .A2(n5581), .ZN(n8256) );
  NAND2_X1 U7081 ( .A1(n8256), .A2(n5288), .ZN(n5584) );
  AOI22_X1 U7082 ( .A1(n5282), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n5667), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7083 ( .A1(n5283), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7084 ( .A1(n8363), .A2(n8012), .ZN(n5826) );
  NAND2_X1 U7085 ( .A1(n8439), .A2(n7906), .ZN(n5794) );
  NAND3_X1 U7086 ( .A1(n5598), .A2(n5826), .A3(n5794), .ZN(n5596) );
  XNOR2_X1 U7087 ( .A(n5586), .B(n5585), .ZN(n5587) );
  XNOR2_X1 U7088 ( .A(n5588), .B(n5587), .ZN(n7656) );
  NAND2_X1 U7089 ( .A1(n7656), .A2(n5751), .ZN(n5590) );
  NAND2_X1 U7090 ( .A1(n5688), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7091 ( .A1(n5591), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7092 ( .A1(n5607), .A2(n5592), .ZN(n8240) );
  NAND2_X1 U7093 ( .A1(n8240), .A2(n5288), .ZN(n5595) );
  AOI22_X1 U7094 ( .A1(n5283), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5667), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7095 ( .A1(n5282), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5593) );
  NAND3_X1 U7096 ( .A1(n5596), .A2(n5825), .A3(n5827), .ZN(n5601) );
  NAND2_X1 U7097 ( .A1(n5794), .A2(n5793), .ZN(n5597) );
  OAI211_X1 U7098 ( .C1(n5598), .C2(n5597), .A(n5795), .B(n5827), .ZN(n5599)
         );
  NAND2_X1 U7099 ( .A1(n5599), .A2(n5826), .ZN(n5600) );
  NAND2_X1 U7100 ( .A1(n8432), .A2(n7972), .ZN(n5824) );
  XNOR2_X1 U7101 ( .A(n5602), .B(SI_21_), .ZN(n5603) );
  XNOR2_X1 U7102 ( .A(n5604), .B(n5603), .ZN(n7701) );
  NAND2_X1 U7103 ( .A1(n7701), .A2(n5751), .ZN(n5606) );
  NAND2_X1 U7104 ( .A1(n5688), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7105 ( .A1(n5607), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7106 ( .A1(n5620), .A2(n5608), .ZN(n8236) );
  NAND2_X1 U7107 ( .A1(n8236), .A2(n5288), .ZN(n5613) );
  INV_X1 U7108 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U7109 ( .A1(n5667), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7110 ( .A1(n5283), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5609) );
  OAI211_X1 U7111 ( .C1(n8235), .C2(n5757), .A(n5610), .B(n5609), .ZN(n5611)
         );
  INV_X1 U7112 ( .A(n5611), .ZN(n5612) );
  NAND2_X1 U7113 ( .A1(n8426), .A2(n7912), .ZN(n5822) );
  NAND2_X1 U7114 ( .A1(n5822), .A2(n5824), .ZN(n5615) );
  NAND2_X1 U7115 ( .A1(n5823), .A2(n5825), .ZN(n5614) );
  MUX2_X1 U7116 ( .A(n5615), .B(n5614), .S(n5929), .Z(n5629) );
  XNOR2_X1 U7117 ( .A(n5617), .B(n5616), .ZN(n7774) );
  NAND2_X1 U7118 ( .A1(n7774), .A2(n5751), .ZN(n5619) );
  NAND2_X1 U7119 ( .A1(n5688), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7120 ( .A1(n5620), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7121 ( .A1(n5634), .A2(n5621), .ZN(n8224) );
  NAND2_X1 U7122 ( .A1(n8224), .A2(n5288), .ZN(n5626) );
  INV_X1 U7123 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U7124 ( .A1(n5282), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7125 ( .A1(n5667), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5622) );
  OAI211_X1 U7126 ( .C1(n4439), .C2(n10124), .A(n5623), .B(n5622), .ZN(n5624)
         );
  INV_X1 U7127 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7128 ( .A1(n8420), .A2(n8208), .ZN(n5798) );
  NAND2_X1 U7129 ( .A1(n5800), .A2(n5798), .ZN(n8217) );
  INV_X1 U7130 ( .A(n8217), .ZN(n5628) );
  MUX2_X1 U7131 ( .A(n5822), .B(n5823), .S(n6636), .Z(n5627) );
  XNOR2_X1 U7132 ( .A(n5631), .B(n5630), .ZN(n7839) );
  NAND2_X1 U7133 ( .A1(n7839), .A2(n5751), .ZN(n5633) );
  NAND2_X1 U7134 ( .A1(n5688), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7135 ( .A1(n5634), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7136 ( .A1(n5648), .A2(n5635), .ZN(n8212) );
  NAND2_X1 U7137 ( .A1(n8212), .A2(n5288), .ZN(n5640) );
  INV_X1 U7138 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U7139 ( .A1(n5667), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7140 ( .A1(n5283), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U7141 ( .C1(n8211), .C2(n5757), .A(n5637), .B(n5636), .ZN(n5638)
         );
  INV_X1 U7142 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U7143 ( .A1(n5640), .A2(n5639), .ZN(n8221) );
  NAND2_X1 U7144 ( .A1(n8213), .A2(n8193), .ZN(n8197) );
  INV_X1 U7145 ( .A(n5800), .ZN(n5641) );
  NOR2_X1 U7146 ( .A1(n5821), .A2(n5641), .ZN(n5642) );
  MUX2_X1 U7147 ( .A(n5798), .B(n5642), .S(n5929), .Z(n5643) );
  XNOR2_X1 U7148 ( .A(n5645), .B(n5644), .ZN(n7863) );
  NAND2_X1 U7149 ( .A1(n7863), .A2(n5751), .ZN(n5647) );
  NAND2_X1 U7150 ( .A1(n5688), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7151 ( .A1(n5648), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7152 ( .A1(n5665), .A2(n5649), .ZN(n8196) );
  NAND2_X1 U7153 ( .A1(n8196), .A2(n5288), .ZN(n5654) );
  INV_X1 U7154 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U7155 ( .A1(n5667), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7156 ( .A1(n5282), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5650) );
  OAI211_X1 U7157 ( .C1(n10153), .C2(n4439), .A(n5651), .B(n5650), .ZN(n5652)
         );
  INV_X1 U7158 ( .A(n5652), .ZN(n5653) );
  INV_X1 U7159 ( .A(n5819), .ZN(n5657) );
  NOR2_X1 U7160 ( .A1(n5657), .A2(n5821), .ZN(n5656) );
  NAND2_X1 U7161 ( .A1(n8005), .A2(n8209), .ZN(n5818) );
  INV_X1 U7162 ( .A(n5818), .ZN(n5655) );
  AOI21_X1 U7163 ( .B1(n5658), .B2(n5656), .A(n5655), .ZN(n5660) );
  AND2_X1 U7164 ( .A1(n5818), .A2(n8197), .ZN(n5801) );
  AOI21_X1 U7165 ( .B1(n5658), .B2(n5801), .A(n5657), .ZN(n5659) );
  MUX2_X1 U7166 ( .A(n5660), .B(n5659), .S(n5929), .Z(n5672) );
  XNOR2_X1 U7167 ( .A(n5662), .B(n5661), .ZN(n7869) );
  NAND2_X1 U7168 ( .A1(n7869), .A2(n5751), .ZN(n5664) );
  NAND2_X1 U7169 ( .A1(n5688), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7170 ( .A1(n5665), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7171 ( .A1(n5677), .A2(n5666), .ZN(n8185) );
  INV_X1 U7172 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U7173 ( .A1(n5667), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7174 ( .A1(n5283), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5668) );
  OAI211_X1 U7175 ( .C1(n10205), .C2(n5757), .A(n5669), .B(n5668), .ZN(n5670)
         );
  NAND2_X1 U7176 ( .A1(n7981), .A2(n8194), .ZN(n5804) );
  MUX2_X1 U7177 ( .A(n5803), .B(n5804), .S(n6636), .Z(n5671) );
  OAI21_X1 U7178 ( .B1(n5672), .B2(n4800), .A(n5671), .ZN(n5700) );
  NAND2_X1 U7179 ( .A1(n7875), .A2(n5751), .ZN(n5676) );
  NAND2_X1 U7180 ( .A1(n5688), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7181 ( .A1(n5677), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7182 ( .A1(n5691), .A2(n5678), .ZN(n8172) );
  NAND2_X1 U7183 ( .A1(n8172), .A2(n5288), .ZN(n5683) );
  INV_X1 U7184 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U7185 ( .A1(n5283), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7186 ( .A1(n5667), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5679) );
  OAI211_X1 U7187 ( .C1(n8175), .C2(n5757), .A(n5680), .B(n5679), .ZN(n5681)
         );
  INV_X1 U7188 ( .A(n5681), .ZN(n5682) );
  INV_X1 U7189 ( .A(n5806), .ZN(n5684) );
  INV_X1 U7190 ( .A(n5807), .ZN(n5685) );
  MUX2_X1 U7191 ( .A(n5806), .B(n5685), .S(n5929), .Z(n5699) );
  NAND2_X1 U7192 ( .A1(n8487), .A2(n5751), .ZN(n5690) );
  NAND2_X1 U7193 ( .A1(n5688), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7194 ( .A1(n5691), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7195 ( .A1(n5705), .A2(n5692), .ZN(n8161) );
  NAND2_X1 U7196 ( .A1(n8161), .A2(n5288), .ZN(n5698) );
  INV_X1 U7197 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7198 ( .A1(n5667), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7199 ( .A1(n5283), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U7200 ( .C1(n5695), .C2(n5757), .A(n5694), .B(n5693), .ZN(n5696)
         );
  INV_X1 U7201 ( .A(n5696), .ZN(n5697) );
  NAND2_X1 U7202 ( .A1(n5919), .A2(n8171), .ZN(n5808) );
  NAND2_X1 U7203 ( .A1(n5809), .A2(n5808), .ZN(n6595) );
  AOI211_X1 U7204 ( .C1(n5700), .C2(n8173), .A(n5699), .B(n6595), .ZN(n5704)
         );
  INV_X1 U7205 ( .A(n5808), .ZN(n5702) );
  INV_X1 U7206 ( .A(n5809), .ZN(n5701) );
  MUX2_X1 U7207 ( .A(n5702), .B(n5701), .S(n6636), .Z(n5703) );
  NAND2_X1 U7208 ( .A1(n5705), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7209 ( .A1(n7878), .A2(n5706), .ZN(n7962) );
  NAND2_X1 U7210 ( .A1(n7962), .A2(n5288), .ZN(n5711) );
  NAND2_X1 U7211 ( .A1(n5283), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5708) );
  INV_X1 U7212 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10190) );
  OR2_X1 U7213 ( .A1(n5236), .A2(n10190), .ZN(n5707) );
  OAI211_X1 U7214 ( .C1(n6629), .C2(n5757), .A(n5708), .B(n5707), .ZN(n5709)
         );
  INV_X1 U7215 ( .A(n5709), .ZN(n5710) );
  NAND2_X1 U7216 ( .A1(n8484), .A2(n5751), .ZN(n5715) );
  NAND2_X1 U7217 ( .A1(n5688), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5714) );
  MUX2_X1 U7218 ( .A(n8068), .B(n7966), .S(n6636), .Z(n5717) );
  NAND2_X1 U7219 ( .A1(n5721), .A2(n8068), .ZN(n5719) );
  NAND2_X1 U7220 ( .A1(n7885), .A2(n7961), .ZN(n5816) );
  INV_X1 U7221 ( .A(n5816), .ZN(n5718) );
  AOI21_X1 U7222 ( .B1(n5719), .B2(n5720), .A(n5718), .ZN(n5724) );
  INV_X1 U7223 ( .A(n5720), .ZN(n5722) );
  NAND2_X1 U7224 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  INV_X1 U7225 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5730) );
  INV_X1 U7226 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n5729) );
  MUX2_X1 U7227 ( .A(n5730), .B(n5729), .S(n6640), .Z(n5732) );
  INV_X1 U7228 ( .A(SI_30_), .ZN(n5731) );
  NAND2_X1 U7229 ( .A1(n5732), .A2(n5731), .ZN(n5745) );
  INV_X1 U7230 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7231 ( .A1(n5733), .A2(SI_30_), .ZN(n5734) );
  NAND2_X1 U7232 ( .A1(n8755), .A2(n5751), .ZN(n5736) );
  NAND2_X1 U7233 ( .A1(n5688), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5735) );
  INV_X1 U7234 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7235 ( .A1(n5283), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7236 ( .A1(n5667), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7237 ( .C1(n5739), .C2(n5757), .A(n5738), .B(n5737), .ZN(n5740)
         );
  INV_X1 U7238 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7239 ( .A1(n5761), .A2(n5741), .ZN(n8067) );
  INV_X1 U7240 ( .A(n8067), .ZN(n5742) );
  NAND2_X1 U7241 ( .A1(n8392), .A2(n5742), .ZN(n5853) );
  NAND2_X1 U7242 ( .A1(n5744), .A2(n5743), .ZN(n5746) );
  NAND2_X1 U7243 ( .A1(n5746), .A2(n5745), .ZN(n5750) );
  INV_X1 U7244 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5747) );
  MUX2_X1 U7245 ( .A(n5747), .B(n10073), .S(n6640), .Z(n5748) );
  XNOR2_X1 U7246 ( .A(n5748), .B(SI_31_), .ZN(n5749) );
  NAND2_X1 U7247 ( .A1(n8760), .A2(n5751), .ZN(n5753) );
  NAND2_X1 U7248 ( .A1(n5688), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5752) );
  INV_X1 U7249 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7250 ( .A1(n5667), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5756) );
  INV_X1 U7251 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5754) );
  OR2_X1 U7252 ( .A1(n4439), .A2(n5754), .ZN(n5755) );
  OAI211_X1 U7253 ( .C1(n5758), .C2(n5757), .A(n5756), .B(n5755), .ZN(n5759)
         );
  INV_X1 U7254 ( .A(n5759), .ZN(n5760) );
  NAND2_X1 U7255 ( .A1(n5766), .A2(n7433), .ZN(n5857) );
  NOR2_X1 U7256 ( .A1(n5766), .A2(n7433), .ZN(n5855) );
  INV_X1 U7257 ( .A(n5762), .ZN(n5763) );
  NAND2_X1 U7258 ( .A1(n5763), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7259 ( .A1(n9850), .A2(n5770), .ZN(n7069) );
  NAND2_X1 U7260 ( .A1(n7068), .A2(n5771), .ZN(n7205) );
  NAND2_X1 U7261 ( .A1(n7205), .A2(n5772), .ZN(n5774) );
  NAND2_X1 U7262 ( .A1(n5774), .A2(n5773), .ZN(n7304) );
  NAND2_X1 U7263 ( .A1(n7304), .A2(n5833), .ZN(n5775) );
  NAND2_X1 U7264 ( .A1(n7706), .A2(n5778), .ZN(n7610) );
  NAND2_X1 U7265 ( .A1(n5782), .A2(n5781), .ZN(n7809) );
  NAND2_X1 U7266 ( .A1(n8334), .A2(n8313), .ZN(n5785) );
  NAND2_X1 U7267 ( .A1(n8283), .A2(n5828), .ZN(n5791) );
  NAND2_X1 U7268 ( .A1(n8262), .A2(n5795), .ZN(n8255) );
  NAND2_X1 U7269 ( .A1(n8255), .A2(n5826), .ZN(n5796) );
  INV_X1 U7270 ( .A(n5825), .ZN(n5797) );
  INV_X1 U7271 ( .A(n8216), .ZN(n5799) );
  NAND2_X1 U7272 ( .A1(n5802), .A2(n5819), .ZN(n8187) );
  INV_X1 U7273 ( .A(n5803), .ZN(n5805) );
  NAND2_X1 U7274 ( .A1(n5810), .A2(n5809), .ZN(n6582) );
  NAND2_X1 U7275 ( .A1(n7966), .A2(n6598), .ZN(n5811) );
  NAND2_X1 U7276 ( .A1(n6582), .A2(n5811), .ZN(n5813) );
  OR2_X1 U7277 ( .A1(n7966), .A2(n6598), .ZN(n5812) );
  NAND2_X1 U7278 ( .A1(n5813), .A2(n5812), .ZN(n5926) );
  INV_X1 U7279 ( .A(n5817), .ZN(n5814) );
  OAI211_X1 U7280 ( .C1(n5926), .C2(n5814), .A(n5853), .B(n5816), .ZN(n5815)
         );
  INV_X1 U7281 ( .A(n8197), .ZN(n5820) );
  NOR2_X1 U7282 ( .A1(n5821), .A2(n5820), .ZN(n8205) );
  NAND2_X1 U7283 ( .A1(n5825), .A2(n5824), .ZN(n8242) );
  NAND2_X1 U7284 ( .A1(n5827), .A2(n5826), .ZN(n8254) );
  INV_X1 U7285 ( .A(n8254), .ZN(n8251) );
  INV_X1 U7286 ( .A(n8288), .ZN(n5847) );
  INV_X1 U7287 ( .A(n8296), .ZN(n8298) );
  NAND2_X1 U7288 ( .A1(n5830), .A2(n8309), .ZN(n8324) );
  NAND2_X1 U7289 ( .A1(n5832), .A2(n5831), .ZN(n7708) );
  INV_X1 U7290 ( .A(n5769), .ZN(n6980) );
  NAND4_X1 U7291 ( .A1(n9859), .A2(n6980), .A3(n7071), .A4(n4808), .ZN(n5837)
         );
  INV_X1 U7292 ( .A(n7206), .ZN(n7204) );
  NAND2_X1 U7293 ( .A1(n5834), .A2(n5833), .ZN(n7306) );
  INV_X1 U7294 ( .A(n5835), .ZN(n5836) );
  NAND2_X1 U7295 ( .A1(n6979), .A2(n5836), .ZN(n6896) );
  NOR4_X1 U7296 ( .A1(n5837), .A2(n7204), .A3(n7306), .A4(n6896), .ZN(n5841)
         );
  INV_X1 U7297 ( .A(n5838), .ZN(n5840) );
  NOR2_X1 U7298 ( .A1(n5840), .A2(n5839), .ZN(n7405) );
  NAND3_X1 U7299 ( .A1(n7462), .A2(n5841), .A3(n7405), .ZN(n5844) );
  NAND2_X1 U7300 ( .A1(n5843), .A2(n5842), .ZN(n7601) );
  NOR4_X1 U7301 ( .A1(n7708), .A2(n5844), .A3(n7610), .A4(n7601), .ZN(n5845)
         );
  NAND4_X1 U7302 ( .A1(n8324), .A2(n4648), .A3(n5845), .A4(n7802), .ZN(n5846)
         );
  NOR4_X1 U7303 ( .A1(n5847), .A2(n8298), .A3(n8311), .A4(n5846), .ZN(n5848)
         );
  NAND4_X1 U7304 ( .A1(n8251), .A2(n8272), .A3(n4482), .A4(n5848), .ZN(n5849)
         );
  NOR4_X1 U7305 ( .A1(n8217), .A2(n4791), .A3(n8242), .A4(n5849), .ZN(n5850)
         );
  NAND4_X1 U7306 ( .A1(n8186), .A2(n8200), .A3(n8205), .A4(n5850), .ZN(n5851)
         );
  NOR4_X1 U7307 ( .A1(n7959), .A2(n6595), .A3(n8168), .A4(n5851), .ZN(n5852)
         );
  NAND4_X1 U7308 ( .A1(n5925), .A2(n4461), .A3(n5853), .A4(n5852), .ZN(n5854)
         );
  OAI22_X1 U7309 ( .A1(n5856), .A2(n4808), .B1(n5855), .B2(n5854), .ZN(n5859)
         );
  NAND2_X1 U7310 ( .A1(n5859), .A2(n5050), .ZN(n5860) );
  NAND2_X1 U7311 ( .A1(n5860), .A2(n6918), .ZN(n5861) );
  NAND2_X1 U7312 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  XNOR2_X1 U7313 ( .A(n5863), .B(n8125), .ZN(n5880) );
  INV_X1 U7314 ( .A(n6815), .ZN(n5867) );
  NAND2_X1 U7315 ( .A1(n5867), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7843) );
  INV_X1 U7316 ( .A(n5957), .ZN(n6985) );
  NAND2_X1 U7317 ( .A1(n4457), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U7318 ( .A(n5870), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5935) );
  INV_X1 U7319 ( .A(n7865), .ZN(n5873) );
  AND2_X1 U7320 ( .A1(n6814), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7321 ( .A1(n6985), .A2(n6660), .ZN(n6821) );
  NOR3_X1 U7322 ( .A1(n6821), .A2(n6711), .A3(n5876), .ZN(n5878) );
  OAI21_X1 U7323 ( .B1(n7843), .B2(n6572), .A(P2_B_REG_SCAN_IN), .ZN(n5877) );
  OR2_X1 U7324 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  OAI21_X1 U7325 ( .B1(n5880), .B2(n7843), .A(n5879), .ZN(P2_U3296) );
  NAND2_X1 U7326 ( .A1(n8080), .A2(n6829), .ZN(n6981) );
  NAND2_X1 U7327 ( .A1(n5769), .A2(n6981), .ZN(n5883) );
  NAND2_X1 U7328 ( .A1(n5881), .A2(n7300), .ZN(n5882) );
  NAND2_X1 U7329 ( .A1(n5883), .A2(n5882), .ZN(n9858) );
  NAND2_X1 U7330 ( .A1(n9858), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U7331 ( .A1(n7073), .A2(n6935), .ZN(n5885) );
  NOR2_X1 U7332 ( .A1(n8077), .A2(n6974), .ZN(n5888) );
  NAND2_X1 U7333 ( .A1(n8077), .A2(n6974), .ZN(n5887) );
  NAND2_X1 U7334 ( .A1(n7305), .A2(n7306), .ZN(n5891) );
  NAND2_X1 U7335 ( .A1(n7258), .A2(n9883), .ZN(n5890) );
  INV_X1 U7336 ( .A(n7461), .ZN(n5893) );
  INV_X1 U7337 ( .A(n7598), .ZN(n8074) );
  OR2_X1 U7338 ( .A1(n9896), .A2(n8074), .ZN(n5894) );
  NAND2_X2 U7339 ( .A1(n7459), .A2(n5894), .ZN(n7596) );
  NAND2_X1 U7340 ( .A1(n9906), .A2(n7650), .ZN(n5895) );
  NAND2_X1 U7341 ( .A1(n7781), .A2(n7780), .ZN(n7779) );
  INV_X1 U7342 ( .A(n7747), .ZN(n8072) );
  NAND2_X1 U7343 ( .A1(n7795), .A2(n8072), .ZN(n5897) );
  OR2_X1 U7344 ( .A1(n8382), .A2(n8329), .ZN(n5898) );
  NAND2_X1 U7345 ( .A1(n7803), .A2(n5898), .ZN(n5900) );
  NAND2_X1 U7346 ( .A1(n8382), .A2(n8329), .ZN(n5899) );
  OR2_X1 U7347 ( .A1(n8308), .A2(n5043), .ZN(n5904) );
  OR2_X1 U7348 ( .A1(n8462), .A2(n8327), .ZN(n5901) );
  AND2_X1 U7349 ( .A1(n8309), .A2(n5901), .ZN(n5902) );
  OR2_X1 U7350 ( .A1(n5043), .A2(n5902), .ZN(n5903) );
  NAND2_X1 U7351 ( .A1(n8457), .A2(n8314), .ZN(n5905) );
  NAND2_X1 U7352 ( .A1(n8299), .A2(n5905), .ZN(n5907) );
  OR2_X1 U7353 ( .A1(n8457), .A2(n8314), .ZN(n5906) );
  INV_X1 U7354 ( .A(n8060), .ZN(n8300) );
  NAND2_X1 U7355 ( .A1(n8451), .A2(n8300), .ZN(n5908) );
  INV_X1 U7356 ( .A(n8445), .ZN(n5909) );
  NAND2_X1 U7357 ( .A1(n8274), .A2(n5046), .ZN(n8264) );
  NAND2_X1 U7358 ( .A1(n8264), .A2(n5910), .ZN(n5912) );
  INV_X1 U7359 ( .A(n8439), .ZN(n5911) );
  AOI22_X2 U7360 ( .A1(n8250), .A2(n8254), .B1(n8265), .B2(n8363), .ZN(n8243)
         );
  INV_X1 U7361 ( .A(n8432), .ZN(n5913) );
  NAND2_X1 U7362 ( .A1(n5913), .A2(n7972), .ZN(n8229) );
  NOR2_X1 U7363 ( .A1(n8426), .A2(n8244), .ZN(n8218) );
  NAND2_X1 U7364 ( .A1(n8213), .A2(n8221), .ZN(n5914) );
  NAND2_X1 U7365 ( .A1(n8191), .A2(n5915), .ZN(n5916) );
  NAND2_X1 U7366 ( .A1(n5916), .A2(n5045), .ZN(n8181) );
  NOR2_X1 U7367 ( .A1(n8398), .A2(n8183), .ZN(n5917) );
  INV_X1 U7368 ( .A(n8183), .ZN(n8070) );
  AOI21_X2 U7369 ( .B1(n8069), .B2(n5919), .A(n5918), .ZN(n6586) );
  NAND2_X1 U7370 ( .A1(n7966), .A2(n8068), .ZN(n5921) );
  NOR2_X1 U7371 ( .A1(n7966), .A2(n8068), .ZN(n5920) );
  AOI21_X1 U7372 ( .B1(n6586), .B2(n5921), .A(n5920), .ZN(n5922) );
  XNOR2_X1 U7373 ( .A(n5922), .B(n5925), .ZN(n5933) );
  NAND2_X1 U7374 ( .A1(n6572), .A2(n8096), .ZN(n5924) );
  NAND2_X1 U7375 ( .A1(n6917), .A2(n6918), .ZN(n5923) );
  XNOR2_X1 U7376 ( .A(n5926), .B(n5925), .ZN(n7882) );
  AOI21_X1 U7377 ( .B1(n7775), .B2(n6918), .A(n8096), .ZN(n5927) );
  NAND3_X1 U7378 ( .A1(n5957), .A2(n5927), .A3(n9909), .ZN(n7615) );
  INV_X1 U7379 ( .A(n5876), .ZN(n6713) );
  NAND2_X1 U7380 ( .A1(n6713), .A2(n6711), .ZN(n5928) );
  NAND2_X1 U7381 ( .A1(n5276), .A2(n5928), .ZN(n6825) );
  INV_X1 U7382 ( .A(n6825), .ZN(n6922) );
  AND2_X1 U7383 ( .A1(n5276), .A2(P2_B_REG_SCAN_IN), .ZN(n5930) );
  NOR2_X1 U7384 ( .A1(n9861), .A2(n5930), .ZN(n8153) );
  AOI22_X1 U7385 ( .A1(n8068), .A2(n8328), .B1(n8067), .B2(n8153), .ZN(n5931)
         );
  OAI21_X1 U7386 ( .B1(n7882), .B2(n7615), .A(n5931), .ZN(n5932) );
  NAND2_X1 U7387 ( .A1(n7887), .A2(n5934), .ZN(n6578) );
  INV_X1 U7388 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7389 ( .A1(n6658), .A2(n5938), .ZN(n5940) );
  NAND2_X1 U7390 ( .A1(n7877), .A2(n7865), .ZN(n5939) );
  NOR2_X1 U7391 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n5944) );
  NOR4_X1 U7392 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5943) );
  NOR4_X1 U7393 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5942) );
  NOR4_X1 U7394 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5941) );
  NAND4_X1 U7395 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n5950)
         );
  NOR4_X1 U7396 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5948) );
  NOR4_X1 U7397 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5947) );
  NOR4_X1 U7398 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5946) );
  NOR4_X1 U7399 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5945) );
  NAND4_X1 U7400 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n5949)
         );
  OAI21_X1 U7401 ( .B1(n5950), .B2(n5949), .A(n6658), .ZN(n6569) );
  INV_X1 U7402 ( .A(n6569), .ZN(n5956) );
  NOR2_X1 U7403 ( .A1(n6916), .A2(n5956), .ZN(n5954) );
  INV_X1 U7404 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7405 ( .A1(n6658), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7406 ( .A1(n7877), .A2(n7871), .ZN(n5952) );
  INV_X1 U7407 ( .A(n6648), .ZN(n6618) );
  AND2_X1 U7408 ( .A1(n5954), .A2(n6618), .ZN(n6822) );
  NAND2_X1 U7409 ( .A1(n6822), .A2(n6660), .ZN(n6924) );
  NOR2_X1 U7410 ( .A1(n7658), .A2(n8125), .ZN(n5955) );
  NAND3_X1 U7411 ( .A1(n4808), .A2(n6572), .A3(n5955), .ZN(n6819) );
  NAND3_X1 U7412 ( .A1(n6819), .A2(n6636), .A3(n9909), .ZN(n6809) );
  OR2_X1 U7413 ( .A1(n6924), .A2(n6812), .ZN(n5960) );
  NAND2_X1 U7414 ( .A1(n6916), .A2(n6648), .ZN(n6570) );
  NOR2_X1 U7415 ( .A1(n6570), .A2(n5956), .ZN(n6813) );
  NAND2_X1 U7416 ( .A1(n6813), .A2(n6660), .ZN(n6827) );
  AND2_X1 U7417 ( .A1(n5957), .A2(n6819), .ZN(n5958) );
  OR2_X1 U7418 ( .A1(n6827), .A2(n5958), .ZN(n5959) );
  NAND2_X1 U7419 ( .A1(n6578), .A2(n9915), .ZN(n5962) );
  NAND2_X1 U7420 ( .A1(n5962), .A2(n5961), .ZN(P2_U3456) );
  NOR2_X1 U7421 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5967) );
  NOR2_X1 U7422 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5966) );
  NOR2_X1 U7423 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5965) );
  NAND4_X1 U7424 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n5968)
         );
  INV_X2 U7425 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U7426 ( .A1(n6007), .A2(n5973), .ZN(n5974) );
  INV_X1 U7427 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7428 ( .A1(n5976), .A2(n5975), .ZN(n6014) );
  NAND2_X1 U7429 ( .A1(n6014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5978) );
  MUX2_X1 U7430 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5978), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5980) );
  INV_X1 U7431 ( .A(n5979), .ZN(n9453) );
  NAND2_X1 U7432 ( .A1(n6529), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5985) );
  NAND4_X2 U7433 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n7022)
         );
  NAND2_X1 U7434 ( .A1(n6259), .A2(n5988), .ZN(n6273) );
  OR2_X1 U7435 ( .A1(n6198), .A2(n10248), .ZN(n5991) );
  XNOR2_X2 U7436 ( .A(n5993), .B(n5992), .ZN(n6345) );
  NAND2_X1 U7437 ( .A1(n5994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7438 ( .A1(n6003), .A2(n6002), .ZN(n5998) );
  NAND2_X1 U7439 ( .A1(n5998), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7440 ( .A1(n6000), .A2(n5999), .ZN(n6506) );
  NAND2_X1 U7441 ( .A1(n8852), .A2(n8808), .ZN(n6541) );
  NAND2_X1 U7442 ( .A1(n4503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  NOR2_X1 U7443 ( .A1(n7874), .A2(n7868), .ZN(n6010) );
  AND2_X1 U7444 ( .A1(n7632), .A2(n6021), .ZN(n6011) );
  NAND2_X2 U7445 ( .A1(n4470), .A2(n6011), .ZN(n6432) );
  INV_X2 U7446 ( .A(n6432), .ZN(n6499) );
  NAND2_X1 U7447 ( .A1(n6015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7448 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6018) );
  XNOR2_X1 U7449 ( .A(n6018), .B(P1_IR_REG_1__SCAN_IN), .ZN(n8943) );
  INV_X1 U7450 ( .A(n6541), .ZN(n6019) );
  AND2_X2 U7451 ( .A1(n6021), .A2(n6019), .ZN(n6037) );
  AND2_X1 U7452 ( .A1(n6996), .A2(n6037), .ZN(n6020) );
  AOI21_X1 U7453 ( .B1(n7022), .B2(n6499), .A(n6020), .ZN(n6027) );
  NAND2_X1 U7454 ( .A1(n7022), .A2(n6037), .ZN(n6024) );
  AND2_X1 U7455 ( .A1(n6021), .A2(n6541), .ZN(n6022) );
  NAND2_X4 U7456 ( .A1(n6540), .A2(n6022), .ZN(n6484) );
  NAND2_X1 U7457 ( .A1(n6026), .A2(n6027), .ZN(n6041) );
  OAI21_X1 U7458 ( .B1(n6027), .B2(n6026), .A(n6041), .ZN(n6993) );
  NAND2_X1 U7459 ( .A1(n6529), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7460 ( .A1(n6889), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7461 ( .A1(n4460), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6028) );
  AND3_X1 U7462 ( .A1(n6030), .A2(n6029), .A3(n6028), .ZN(n6032) );
  NAND2_X1 U7463 ( .A1(n6074), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6031) );
  NAND2_X2 U7464 ( .A1(n6032), .A2(n6031), .ZN(n8936) );
  NAND2_X1 U7465 ( .A1(n4660), .A2(SI_0_), .ZN(n6033) );
  XNOR2_X1 U7466 ( .A(n6033), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U7467 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9469), .S(n6668), .Z(n7083) );
  INV_X1 U7468 ( .A(n6021), .ZN(n6038) );
  AOI21_X2 U7469 ( .B1(n8936), .B2(n6486), .A(n6036), .ZN(n6941) );
  OAI22_X1 U7470 ( .A1(n6941), .A2(n6942), .B1(n7083), .B2(n6484), .ZN(n6995)
         );
  NOR2_X1 U7471 ( .A1(n6993), .A2(n6995), .ZN(n6994) );
  INV_X1 U7472 ( .A(n6041), .ZN(n7060) );
  NAND2_X1 U7473 ( .A1(n6074), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7474 ( .A1(n6889), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7475 ( .A1(n6529), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7476 ( .A1(n4460), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6042) );
  NAND4_X1 U7477 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n6046)
         );
  NAND2_X1 U7478 ( .A1(n6046), .A2(n6037), .ZN(n6052) );
  NAND2_X1 U7479 ( .A1(n6080), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6050) );
  INV_X1 U7480 ( .A(n7052), .ZN(n6048) );
  NAND2_X1 U7481 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  XNOR2_X1 U7482 ( .A(n6053), .B(n6497), .ZN(n6055) );
  AND2_X1 U7483 ( .A1(n7112), .A2(n6037), .ZN(n6054) );
  AOI21_X1 U7484 ( .B1(n6046), .B2(n6499), .A(n6054), .ZN(n6056) );
  NAND2_X1 U7485 ( .A1(n6055), .A2(n6056), .ZN(n6060) );
  INV_X1 U7486 ( .A(n6055), .ZN(n6058) );
  INV_X1 U7487 ( .A(n6056), .ZN(n6057) );
  NAND2_X1 U7488 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  NAND2_X1 U7489 ( .A1(n7058), .A2(n6060), .ZN(n8515) );
  INV_X1 U7490 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7187) );
  NAND2_X1 U7491 ( .A1(n6074), .A2(n7187), .ZN(n6064) );
  NAND2_X1 U7492 ( .A1(n8766), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7493 ( .A1(n6529), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7494 ( .A1(n4460), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7495 ( .A1(n6080), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6070) );
  INV_X2 U7496 ( .A(n6668), .ZN(n6346) );
  INV_X1 U7497 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7498 ( .A1(n6083), .A2(n6066), .ZN(n6067) );
  NAND2_X1 U7499 ( .A1(n6067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7500 ( .A1(n6346), .A2(n8950), .ZN(n6069) );
  OAI211_X1 U7501 ( .C1(n6238), .C2(n6645), .A(n6070), .B(n6069), .ZN(n8518)
         );
  INV_X2 U7502 ( .A(n6397), .ZN(n6433) );
  AOI22_X1 U7503 ( .A1(n8934), .A2(n6486), .B1(n8518), .B2(n6433), .ZN(n6071)
         );
  XNOR2_X1 U7504 ( .A(n6071), .B(n6484), .ZN(n6095) );
  AND2_X1 U7505 ( .A1(n8518), .A2(n6486), .ZN(n6072) );
  AOI21_X1 U7506 ( .B1(n8934), .B2(n6499), .A(n6072), .ZN(n6094) );
  XNOR2_X1 U7507 ( .A(n6095), .B(n6073), .ZN(n8516) );
  NAND2_X1 U7508 ( .A1(n8515), .A2(n8516), .ZN(n8514) );
  NAND2_X1 U7509 ( .A1(n8764), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7510 ( .A1(n8765), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6078) );
  NOR2_X1 U7511 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6075) );
  NOR2_X1 U7512 ( .A1(n6101), .A2(n6075), .ZN(n9599) );
  NAND2_X1 U7513 ( .A1(n6074), .A2(n9599), .ZN(n6077) );
  NAND2_X1 U7514 ( .A1(n8766), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7515 ( .A1(n7281), .A2(n6486), .ZN(n6091) );
  NAND2_X1 U7516 ( .A1(n8761), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7517 ( .A1(n6081), .A2(n6198), .ZN(n6082) );
  AND2_X1 U7518 ( .A1(n6083), .A2(n6082), .ZN(n6085) );
  INV_X1 U7519 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7520 ( .A1(n6085), .A2(n6084), .ZN(n6107) );
  INV_X1 U7521 ( .A(n6085), .ZN(n6086) );
  NAND2_X1 U7522 ( .A1(n6086), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7523 ( .A1(n6346), .A2(n6802), .ZN(n6088) );
  OAI211_X1 U7524 ( .C1(n6238), .C2(n6657), .A(n6089), .B(n6088), .ZN(n7358)
         );
  NAND2_X1 U7525 ( .A1(n6433), .A2(n7358), .ZN(n6090) );
  NAND2_X1 U7526 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7527 ( .A(n6092), .B(n6484), .ZN(n6097) );
  AND2_X1 U7528 ( .A1(n7358), .A2(n6037), .ZN(n6093) );
  AOI21_X1 U7529 ( .B1(n7281), .B2(n6499), .A(n6093), .ZN(n6098) );
  XNOR2_X1 U7530 ( .A(n6097), .B(n6098), .ZN(n7252) );
  NAND2_X1 U7531 ( .A1(n6095), .A2(n6094), .ZN(n7250) );
  NAND2_X1 U7532 ( .A1(n8514), .A2(n6096), .ZN(n7251) );
  NAND2_X1 U7533 ( .A1(n6889), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7534 ( .A1(n6529), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6105) );
  NOR2_X1 U7535 ( .A1(n6101), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6102) );
  NOR2_X1 U7536 ( .A1(n6118), .A2(n6102), .ZN(n7430) );
  NAND2_X1 U7537 ( .A1(n6074), .A2(n7430), .ZN(n6104) );
  NAND2_X1 U7538 ( .A1(n4460), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6103) );
  NAND4_X1 U7539 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n8933)
         );
  OR2_X1 U7540 ( .A1(n6654), .A2(n6238), .ZN(n6110) );
  NAND2_X1 U7541 ( .A1(n6107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6108) );
  XNOR2_X1 U7542 ( .A(n6108), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7543 ( .A1(n8761), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6346), .B2(
        n6838), .ZN(n6109) );
  NAND2_X1 U7544 ( .A1(n6110), .A2(n6109), .ZN(n8670) );
  AOI22_X1 U7545 ( .A1(n8933), .A2(n6037), .B1(n8670), .B2(n6433), .ZN(n6111)
         );
  XOR2_X1 U7546 ( .A(n6484), .B(n6111), .Z(n6113) );
  INV_X1 U7547 ( .A(n8933), .ZN(n8671) );
  OAI22_X1 U7548 ( .A1(n8671), .A2(n6432), .B1(n8668), .B2(n6065), .ZN(n7425)
         );
  INV_X1 U7549 ( .A(n6113), .ZN(n7423) );
  INV_X1 U7550 ( .A(n7425), .ZN(n6127) );
  NAND2_X1 U7551 ( .A1(n6675), .A2(n8759), .ZN(n6117) );
  NAND2_X1 U7552 ( .A1(n6114), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U7553 ( .A(n6115), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U7554 ( .A1(n8761), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6346), .B2(
        n6865), .ZN(n6116) );
  NAND2_X1 U7555 ( .A1(n6117), .A2(n6116), .ZN(n8674) );
  NAND2_X1 U7556 ( .A1(n8674), .A2(n6433), .ZN(n6125) );
  NAND2_X1 U7557 ( .A1(n6889), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7558 ( .A1(n6529), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6122) );
  NOR2_X1 U7559 ( .A1(n6118), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6119) );
  NOR2_X1 U7560 ( .A1(n6136), .A2(n6119), .ZN(n8638) );
  NAND2_X1 U7561 ( .A1(n6074), .A2(n8638), .ZN(n6121) );
  NAND2_X1 U7562 ( .A1(n4460), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6120) );
  NAND4_X1 U7563 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n8932)
         );
  NAND2_X1 U7564 ( .A1(n8932), .A2(n6037), .ZN(n6124) );
  NAND2_X1 U7565 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  XNOR2_X1 U7566 ( .A(n6126), .B(n6497), .ZN(n6131) );
  AOI22_X1 U7567 ( .A1(n8674), .A2(n6486), .B1(n8932), .B2(n6499), .ZN(n6130)
         );
  OR2_X1 U7568 ( .A1(n6131), .A2(n6130), .ZN(n8631) );
  OAI21_X1 U7569 ( .B1(n7423), .B2(n6127), .A(n8631), .ZN(n6128) );
  NAND2_X1 U7570 ( .A1(n6131), .A2(n6130), .ZN(n8630) );
  NAND2_X1 U7571 ( .A1(n6133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6134) );
  XNOR2_X1 U7572 ( .A(n6134), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6852) );
  AOI22_X1 U7573 ( .A1(n8761), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6346), .B2(
        n6852), .ZN(n6135) );
  NAND2_X1 U7574 ( .A1(n9588), .A2(n6433), .ZN(n6142) );
  NAND2_X1 U7575 ( .A1(n8764), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7576 ( .A1(n8766), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7577 ( .A1(n6136), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6155) );
  OAI21_X1 U7578 ( .B1(n6136), .B2(P1_REG3_REG_7__SCAN_IN), .A(n6155), .ZN(
        n7419) );
  INV_X1 U7579 ( .A(n7419), .ZN(n9586) );
  NAND2_X1 U7580 ( .A1(n6074), .A2(n9586), .ZN(n6138) );
  NAND2_X1 U7581 ( .A1(n8765), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6137) );
  NAND4_X1 U7582 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n8931)
         );
  NAND2_X1 U7583 ( .A1(n8931), .A2(n6486), .ZN(n6141) );
  NAND2_X1 U7584 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  XNOR2_X1 U7585 ( .A(n6143), .B(n6484), .ZN(n7412) );
  NAND2_X1 U7586 ( .A1(n9588), .A2(n6486), .ZN(n6145) );
  NAND2_X1 U7587 ( .A1(n8931), .A2(n6499), .ZN(n6144) );
  NAND2_X1 U7588 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  NOR2_X1 U7589 ( .A1(n7412), .A2(n6146), .ZN(n6147) );
  INV_X1 U7590 ( .A(n6146), .ZN(n7411) );
  NAND2_X1 U7591 ( .A1(n6680), .A2(n8759), .ZN(n6153) );
  NOR2_X1 U7592 ( .A1(n6133), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6179) );
  NOR2_X1 U7593 ( .A1(n6179), .A2(n6198), .ZN(n6148) );
  NAND2_X1 U7594 ( .A1(n6148), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6151) );
  INV_X1 U7595 ( .A(n6148), .ZN(n6150) );
  INV_X1 U7596 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7597 ( .A1(n6150), .A2(n6149), .ZN(n6165) );
  AOI22_X1 U7598 ( .A1(n6080), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6346), .B2(
        n6877), .ZN(n6152) );
  NAND2_X1 U7599 ( .A1(n6153), .A2(n6152), .ZN(n7530) );
  NAND2_X1 U7600 ( .A1(n7530), .A2(n6433), .ZN(n6162) );
  NAND2_X1 U7601 ( .A1(n6889), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7602 ( .A1(n6529), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6159) );
  AND2_X1 U7603 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  NOR2_X1 U7604 ( .A1(n6169), .A2(n6156), .ZN(n7593) );
  NAND2_X1 U7605 ( .A1(n6074), .A2(n7593), .ZN(n6158) );
  NAND2_X1 U7606 ( .A1(n8765), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6157) );
  NAND4_X1 U7607 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n8930)
         );
  NAND2_X1 U7608 ( .A1(n8930), .A2(n6037), .ZN(n6161) );
  NAND2_X1 U7609 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  XNOR2_X1 U7610 ( .A(n6163), .B(n6484), .ZN(n6164) );
  INV_X1 U7611 ( .A(n7530), .ZN(n9646) );
  INV_X1 U7612 ( .A(n8930), .ZN(n7486) );
  OAI22_X1 U7613 ( .A1(n9646), .A2(n6065), .B1(n7486), .B2(n6432), .ZN(n7586)
         );
  NAND2_X1 U7614 ( .A1(n6685), .A2(n8759), .ZN(n6168) );
  NAND2_X1 U7615 ( .A1(n6165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U7616 ( .A(n6166), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U7617 ( .A1(n6080), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6346), .B2(
        n6954), .ZN(n6167) );
  NAND2_X1 U7618 ( .A1(n6168), .A2(n6167), .ZN(n7687) );
  NAND2_X1 U7619 ( .A1(n8766), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7620 ( .A1(n6529), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7621 ( .A1(n6169), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7622 ( .A1(n6169), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6170) );
  AND2_X1 U7623 ( .A1(n6187), .A2(n6170), .ZN(n7725) );
  NAND2_X1 U7624 ( .A1(n6074), .A2(n7725), .ZN(n6172) );
  NAND2_X1 U7625 ( .A1(n8765), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6171) );
  NAND4_X1 U7626 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n8929)
         );
  AOI22_X1 U7627 ( .A1(n7687), .A2(n6433), .B1(n6486), .B2(n8929), .ZN(n6175)
         );
  XNOR2_X1 U7628 ( .A(n6175), .B(n6484), .ZN(n6176) );
  INV_X1 U7629 ( .A(n7687), .ZN(n7728) );
  INV_X1 U7630 ( .A(n8929), .ZN(n7515) );
  OAI22_X1 U7631 ( .A1(n7728), .A2(n6065), .B1(n7515), .B2(n6432), .ZN(n7718)
         );
  NAND2_X1 U7632 ( .A1(n6177), .A2(n6176), .ZN(n7716) );
  OAI21_X1 U7633 ( .B1(n7715), .B2(n7718), .A(n7716), .ZN(n6196) );
  OR2_X1 U7634 ( .A1(n6690), .A2(n6238), .ZN(n6185) );
  NOR2_X1 U7635 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6178) );
  AND2_X1 U7636 ( .A1(n6179), .A2(n6178), .ZN(n6182) );
  NOR2_X1 U7637 ( .A1(n6182), .A2(n6198), .ZN(n6180) );
  MUX2_X1 U7638 ( .A(n6198), .B(n6180), .S(P1_IR_REG_10__SCAN_IN), .Z(n6183)
         );
  INV_X1 U7639 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6181) );
  AOI22_X1 U7640 ( .A1(n6080), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6346), .B2(
        n7012), .ZN(n6184) );
  NAND2_X1 U7641 ( .A1(n6185), .A2(n6184), .ZN(n9498) );
  NAND2_X1 U7642 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  NAND2_X1 U7643 ( .A1(n6202), .A2(n6188), .ZN(n9500) );
  INV_X1 U7644 ( .A(n9500), .ZN(n6189) );
  NAND2_X1 U7645 ( .A1(n6074), .A2(n6189), .ZN(n6193) );
  NAND2_X1 U7646 ( .A1(n8765), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7647 ( .A1(n8764), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7648 ( .A1(n8766), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6190) );
  NAND4_X1 U7649 ( .A1(n6193), .A2(n6192), .A3(n6191), .A4(n6190), .ZN(n8928)
         );
  AOI22_X1 U7650 ( .A1(n9498), .A2(n4603), .B1(n6486), .B2(n8928), .ZN(n6194)
         );
  XNOR2_X1 U7651 ( .A(n6194), .B(n6484), .ZN(n6195) );
  NAND2_X1 U7652 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  INV_X1 U7653 ( .A(n9498), .ZN(n7544) );
  INV_X1 U7654 ( .A(n8928), .ZN(n7521) );
  OAI22_X1 U7655 ( .A1(n7544), .A2(n6065), .B1(n7521), .B2(n6432), .ZN(n9492)
         );
  INV_X1 U7656 ( .A(n6197), .ZN(n7830) );
  NAND2_X1 U7657 ( .A1(n6779), .A2(n8759), .ZN(n6201) );
  OR2_X1 U7658 ( .A1(n6218), .A2(n6198), .ZN(n6199) );
  XNOR2_X1 U7659 ( .A(n6199), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7139) );
  AOI22_X1 U7660 ( .A1(n6080), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6346), .B2(
        n7139), .ZN(n6200) );
  NAND2_X1 U7661 ( .A1(n6201), .A2(n6200), .ZN(n7661) );
  NAND2_X1 U7662 ( .A1(n7661), .A2(n4603), .ZN(n6209) );
  NAND2_X1 U7663 ( .A1(n8764), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6207) );
  AND2_X1 U7664 ( .A1(n6202), .A2(n10162), .ZN(n6203) );
  NOR2_X1 U7665 ( .A1(n6222), .A2(n6203), .ZN(n7836) );
  NAND2_X1 U7666 ( .A1(n6074), .A2(n7836), .ZN(n6206) );
  NAND2_X1 U7667 ( .A1(n8765), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7668 ( .A1(n6889), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6204) );
  NAND4_X1 U7669 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n8927)
         );
  NAND2_X1 U7670 ( .A1(n8927), .A2(n6486), .ZN(n6208) );
  NAND2_X1 U7671 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  XNOR2_X1 U7672 ( .A(n6210), .B(n6497), .ZN(n6212) );
  AND2_X1 U7673 ( .A1(n8927), .A2(n6499), .ZN(n6211) );
  AOI21_X1 U7674 ( .B1(n7661), .B2(n6486), .A(n6211), .ZN(n6213) );
  NAND2_X1 U7675 ( .A1(n6212), .A2(n6213), .ZN(n7854) );
  INV_X1 U7676 ( .A(n6212), .ZN(n6215) );
  INV_X1 U7677 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7678 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  AND2_X1 U7679 ( .A1(n7854), .A2(n6216), .ZN(n7829) );
  OR2_X1 U7680 ( .A1(n6888), .A2(n6238), .ZN(n6221) );
  INV_X1 U7681 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7682 ( .A1(n6218), .A2(n6217), .ZN(n6239) );
  NAND2_X1 U7683 ( .A1(n6239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6219) );
  XNOR2_X1 U7684 ( .A(n6219), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8985) );
  AOI22_X1 U7685 ( .A1(n6080), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6346), .B2(
        n8985), .ZN(n6220) );
  NAND2_X1 U7686 ( .A1(n7730), .A2(n4603), .ZN(n6229) );
  NAND2_X1 U7687 ( .A1(n8766), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7688 ( .A1(n8764), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6226) );
  NOR2_X1 U7689 ( .A1(n6222), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6223) );
  OR2_X1 U7690 ( .A1(n6243), .A2(n6223), .ZN(n7694) );
  INV_X1 U7691 ( .A(n7694), .ZN(n7859) );
  NAND2_X1 U7692 ( .A1(n6074), .A2(n7859), .ZN(n6225) );
  NAND2_X1 U7693 ( .A1(n8765), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6224) );
  NAND4_X1 U7694 ( .A1(n6227), .A2(n6226), .A3(n6225), .A4(n6224), .ZN(n8926)
         );
  NAND2_X1 U7695 ( .A1(n8926), .A2(n6037), .ZN(n6228) );
  NAND2_X1 U7696 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  XNOR2_X1 U7697 ( .A(n6230), .B(n6497), .ZN(n6232) );
  AND2_X1 U7698 ( .A1(n8926), .A2(n6499), .ZN(n6231) );
  AOI21_X1 U7699 ( .B1(n7730), .B2(n6486), .A(n6231), .ZN(n6233) );
  NAND2_X1 U7700 ( .A1(n6232), .A2(n6233), .ZN(n6237) );
  INV_X1 U7701 ( .A(n6232), .ZN(n6235) );
  INV_X1 U7702 ( .A(n6233), .ZN(n6234) );
  NAND2_X1 U7703 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  NAND2_X1 U7704 ( .A1(n6237), .A2(n6236), .ZN(n7853) );
  INV_X1 U7705 ( .A(n6237), .ZN(n8604) );
  OR2_X1 U7706 ( .A1(n6977), .A2(n6238), .ZN(n6242) );
  OAI21_X1 U7707 ( .B1(n6239), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6240) );
  XNOR2_X1 U7708 ( .A(n6240), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9510) );
  AOI22_X1 U7709 ( .A1(n6080), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6346), .B2(
        n9510), .ZN(n6241) );
  NAND2_X1 U7710 ( .A1(n9381), .A2(n4603), .ZN(n6250) );
  NAND2_X1 U7711 ( .A1(n8766), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7712 ( .A1(n8764), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6247) );
  OR2_X1 U7713 ( .A1(n6243), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6244) );
  AND2_X1 U7714 ( .A1(n6263), .A2(n6244), .ZN(n8609) );
  NAND2_X1 U7715 ( .A1(n6074), .A2(n8609), .ZN(n6246) );
  NAND2_X1 U7716 ( .A1(n8765), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6245) );
  NAND4_X1 U7717 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n8925)
         );
  NAND2_X1 U7718 ( .A1(n8925), .A2(n6486), .ZN(n6249) );
  NAND2_X1 U7719 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  XNOR2_X1 U7720 ( .A(n6251), .B(n6497), .ZN(n6253) );
  AND2_X1 U7721 ( .A1(n8925), .A2(n6499), .ZN(n6252) );
  AOI21_X1 U7722 ( .B1(n9381), .B2(n6486), .A(n6252), .ZN(n6254) );
  NAND2_X1 U7723 ( .A1(n6253), .A2(n6254), .ZN(n6258) );
  INV_X1 U7724 ( .A(n6253), .ZN(n6256) );
  INV_X1 U7725 ( .A(n6254), .ZN(n6255) );
  NAND2_X1 U7726 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  AND2_X1 U7727 ( .A1(n6258), .A2(n6257), .ZN(n8603) );
  NAND2_X1 U7728 ( .A1(n7037), .A2(n8759), .ZN(n6262) );
  OR2_X1 U7729 ( .A1(n6259), .A2(n6198), .ZN(n6260) );
  XNOR2_X1 U7730 ( .A(n6260), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8987) );
  AOI22_X1 U7731 ( .A1(n6080), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6346), .B2(
        n8987), .ZN(n6261) );
  NAND2_X1 U7732 ( .A1(n8766), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7733 ( .A1(n8764), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7734 ( .A1(n6263), .A2(n8496), .ZN(n6264) );
  AND2_X1 U7735 ( .A1(n6278), .A2(n6264), .ZN(n8501) );
  NAND2_X1 U7736 ( .A1(n6074), .A2(n8501), .ZN(n6266) );
  NAND2_X1 U7737 ( .A1(n8765), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6265) );
  NAND4_X1 U7738 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n8924)
         );
  AOI22_X1 U7739 ( .A1(n9375), .A2(n4603), .B1(n6486), .B2(n8924), .ZN(n6269)
         );
  XNOR2_X1 U7740 ( .A(n6269), .B(n6484), .ZN(n6270) );
  INV_X1 U7741 ( .A(n9375), .ZN(n8498) );
  INV_X1 U7742 ( .A(n8924), .ZN(n8693) );
  NAND2_X1 U7743 ( .A1(n8492), .A2(n8495), .ZN(n6272) );
  INV_X1 U7744 ( .A(n6270), .ZN(n6271) );
  NAND2_X1 U7745 ( .A1(n7147), .A2(n8759), .ZN(n6277) );
  NAND2_X1 U7746 ( .A1(n6273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6274) );
  MUX2_X1 U7747 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6274), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6275) );
  NAND2_X1 U7748 ( .A1(n6275), .A2(n4459), .ZN(n8989) );
  INV_X1 U7749 ( .A(n8989), .ZN(n9537) );
  AOI22_X1 U7750 ( .A1(n6080), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6346), .B2(
        n9537), .ZN(n6276) );
  NAND2_X1 U7751 ( .A1(n6529), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7752 ( .A1(n8766), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7753 ( .A1(n6278), .A2(n10090), .ZN(n6279) );
  AND2_X1 U7754 ( .A1(n6290), .A2(n6279), .ZN(n8655) );
  NAND2_X1 U7755 ( .A1(n6074), .A2(n8655), .ZN(n6281) );
  NAND2_X1 U7756 ( .A1(n8765), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6280) );
  NAND4_X1 U7757 ( .A1(n6283), .A2(n6282), .A3(n6281), .A4(n6280), .ZN(n9023)
         );
  AOI22_X1 U7758 ( .A1(n9024), .A2(n4603), .B1(n6486), .B2(n9023), .ZN(n6284)
         );
  XNOR2_X1 U7759 ( .A(n6284), .B(n6484), .ZN(n6285) );
  INV_X1 U7760 ( .A(n9023), .ZN(n9020) );
  OAI22_X1 U7761 ( .A1(n9021), .A2(n6065), .B1(n9020), .B2(n6432), .ZN(n8653)
         );
  NAND2_X1 U7762 ( .A1(n7202), .A2(n8759), .ZN(n6288) );
  XNOR2_X1 U7763 ( .A(n6286), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U7764 ( .A1(n6080), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6346), .B2(
        n9550), .ZN(n6287) );
  NAND2_X1 U7765 ( .A1(n9370), .A2(n4603), .ZN(n6297) );
  AND2_X1 U7766 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  NOR2_X1 U7767 ( .A1(n6302), .A2(n6291), .ZN(n9288) );
  NAND2_X1 U7768 ( .A1(n9288), .A2(n6074), .ZN(n6295) );
  NAND2_X1 U7769 ( .A1(n8766), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7770 ( .A1(n8764), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7771 ( .A1(n8765), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6292) );
  NAND4_X1 U7772 ( .A1(n6295), .A2(n6294), .A3(n6293), .A4(n6292), .ZN(n9027)
         );
  NAND2_X1 U7773 ( .A1(n9027), .A2(n6037), .ZN(n6296) );
  NAND2_X1 U7774 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  XNOR2_X1 U7775 ( .A(n6298), .B(n6484), .ZN(n6310) );
  AOI22_X1 U7776 ( .A1(n9370), .A2(n6486), .B1(n6499), .B2(n9027), .ZN(n6311)
         );
  XNOR2_X1 U7777 ( .A(n6310), .B(n6311), .ZN(n8565) );
  NAND2_X1 U7778 ( .A1(n7346), .A2(n8759), .ZN(n6301) );
  XNOR2_X1 U7779 ( .A(n6299), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8993) );
  AOI22_X1 U7780 ( .A1(n6080), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6346), .B2(
        n8993), .ZN(n6300) );
  NAND2_X1 U7781 ( .A1(n9267), .A2(n4603), .ZN(n6308) );
  NAND2_X1 U7782 ( .A1(n6302), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6324) );
  OR2_X1 U7783 ( .A1(n6302), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7784 ( .A1(n6324), .A2(n6303), .ZN(n8576) );
  INV_X1 U7785 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8992) );
  OAI22_X1 U7786 ( .A1(n8576), .A2(n6477), .B1(n6304), .B2(n8992), .ZN(n6306)
         );
  INV_X1 U7787 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9364) );
  INV_X1 U7788 ( .A(n8766), .ZN(n6395) );
  INV_X1 U7789 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9441) );
  OAI22_X1 U7790 ( .A1(n6480), .A2(n9364), .B1(n6395), .B2(n9441), .ZN(n6305)
         );
  NAND2_X1 U7791 ( .A1(n9028), .A2(n6037), .ZN(n6307) );
  NAND2_X1 U7792 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  XNOR2_X1 U7793 ( .A(n6309), .B(n6484), .ZN(n6316) );
  AOI22_X1 U7794 ( .A1(n9267), .A2(n6037), .B1(n6499), .B2(n9028), .ZN(n6314)
         );
  XNOR2_X1 U7795 ( .A(n6316), .B(n6314), .ZN(n8574) );
  INV_X1 U7796 ( .A(n6310), .ZN(n6312) );
  NAND2_X1 U7797 ( .A1(n6312), .A2(n6311), .ZN(n8572) );
  NAND2_X1 U7798 ( .A1(n8563), .A2(n6313), .ZN(n8573) );
  INV_X1 U7799 ( .A(n6314), .ZN(n6315) );
  NAND2_X1 U7800 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  NAND2_X1 U7801 ( .A1(n8573), .A2(n6317), .ZN(n8523) );
  NAND2_X1 U7802 ( .A1(n7400), .A2(n8759), .ZN(n6323) );
  OR2_X1 U7803 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  AND2_X1 U7804 ( .A1(n6321), .A2(n6320), .ZN(n9578) );
  AOI22_X1 U7805 ( .A1(n6080), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6346), .B2(
        n9578), .ZN(n6322) );
  NAND2_X1 U7806 ( .A1(n9358), .A2(n6486), .ZN(n6329) );
  NAND2_X1 U7807 ( .A1(n6324), .A2(n8622), .ZN(n6325) );
  NAND2_X1 U7808 ( .A1(n6349), .A2(n6325), .ZN(n9252) );
  AOI22_X1 U7809 ( .A1(n8764), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8765), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7810 ( .A1(n8766), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6326) );
  OAI211_X1 U7811 ( .C1(n9252), .C2(n6477), .A(n6327), .B(n6326), .ZN(n9029)
         );
  NAND2_X1 U7812 ( .A1(n9029), .A2(n6499), .ZN(n6328) );
  NAND2_X1 U7813 ( .A1(n9358), .A2(n6433), .ZN(n6331) );
  NAND2_X1 U7814 ( .A1(n9029), .A2(n6486), .ZN(n6330) );
  NAND2_X1 U7815 ( .A1(n6331), .A2(n6330), .ZN(n6332) );
  XNOR2_X1 U7816 ( .A(n6332), .B(n6497), .ZN(n6360) );
  NAND2_X1 U7817 ( .A1(n7656), .A2(n8759), .ZN(n6334) );
  NAND2_X1 U7818 ( .A1(n8761), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7819 ( .A1(n9348), .A2(n6433), .ZN(n6341) );
  NOR2_X1 U7820 ( .A1(n6350), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6335) );
  OR2_X1 U7821 ( .A1(n6372), .A2(n6335), .ZN(n9221) );
  INV_X1 U7822 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10168) );
  NAND2_X1 U7823 ( .A1(n6529), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7824 ( .A1(n8765), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6336) );
  OAI211_X1 U7825 ( .C1(n6395), .C2(n10168), .A(n6337), .B(n6336), .ZN(n6338)
         );
  INV_X1 U7826 ( .A(n6338), .ZN(n6339) );
  OAI21_X1 U7827 ( .B1(n9221), .B2(n6477), .A(n6339), .ZN(n9038) );
  NAND2_X1 U7828 ( .A1(n9038), .A2(n6486), .ZN(n6340) );
  NAND2_X1 U7829 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  XNOR2_X1 U7830 ( .A(n6342), .B(n6484), .ZN(n6364) );
  NAND2_X1 U7831 ( .A1(n9348), .A2(n6486), .ZN(n6344) );
  NAND2_X1 U7832 ( .A1(n9038), .A2(n6499), .ZN(n6343) );
  NAND2_X1 U7833 ( .A1(n6344), .A2(n6343), .ZN(n6365) );
  NAND2_X1 U7834 ( .A1(n6364), .A2(n6365), .ZN(n8541) );
  NAND2_X1 U7835 ( .A1(n7583), .A2(n8759), .ZN(n6348) );
  AOI22_X1 U7836 ( .A1(n6080), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6346), .B2(
        n9002), .ZN(n6347) );
  NAND2_X1 U7837 ( .A1(n9429), .A2(n6433), .ZN(n6355) );
  AND2_X1 U7838 ( .A1(n6349), .A2(n8529), .ZN(n6351) );
  OR2_X1 U7839 ( .A1(n6351), .A2(n6350), .ZN(n9237) );
  AOI22_X1 U7840 ( .A1(n8764), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8766), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7841 ( .A1(n8765), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6352) );
  OAI211_X1 U7842 ( .C1(n9237), .C2(n6477), .A(n6353), .B(n6352), .ZN(n9032)
         );
  NAND2_X1 U7843 ( .A1(n9032), .A2(n6037), .ZN(n6354) );
  NAND2_X1 U7844 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  XNOR2_X1 U7845 ( .A(n6356), .B(n6484), .ZN(n8525) );
  NAND2_X1 U7846 ( .A1(n9429), .A2(n6037), .ZN(n6358) );
  NAND2_X1 U7847 ( .A1(n9032), .A2(n6499), .ZN(n6357) );
  NAND2_X1 U7848 ( .A1(n6358), .A2(n6357), .ZN(n8524) );
  NAND2_X1 U7849 ( .A1(n8525), .A2(n8524), .ZN(n8540) );
  OAI211_X1 U7850 ( .C1(n8620), .C2(n6360), .A(n8541), .B(n8540), .ZN(n6359)
         );
  NOR2_X1 U7851 ( .A1(n8523), .A2(n6359), .ZN(n6384) );
  INV_X1 U7852 ( .A(n8541), .ZN(n6369) );
  INV_X1 U7853 ( .A(n8525), .ZN(n6363) );
  INV_X1 U7854 ( .A(n8620), .ZN(n8536) );
  OAI21_X1 U7855 ( .B1(n8535), .B2(n8536), .A(n8524), .ZN(n6362) );
  NOR3_X1 U7856 ( .A1(n8535), .A2(n8524), .A3(n8536), .ZN(n6361) );
  AOI21_X1 U7857 ( .B1(n6363), .B2(n6362), .A(n6361), .ZN(n6368) );
  INV_X1 U7858 ( .A(n6364), .ZN(n6367) );
  INV_X1 U7859 ( .A(n6365), .ZN(n6366) );
  NAND2_X1 U7860 ( .A1(n6367), .A2(n6366), .ZN(n8542) );
  OAI21_X1 U7861 ( .B1(n6369), .B2(n6368), .A(n8542), .ZN(n6383) );
  NAND2_X1 U7862 ( .A1(n7701), .A2(n8759), .ZN(n6371) );
  NAND2_X1 U7863 ( .A1(n6080), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U7864 ( .A1(n9421), .A2(n6433), .ZN(n6380) );
  OR2_X1 U7865 ( .A1(n6372), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6373) );
  AND2_X1 U7866 ( .A1(n6391), .A2(n6373), .ZN(n9206) );
  NAND2_X1 U7867 ( .A1(n9206), .A2(n6074), .ZN(n6378) );
  INV_X1 U7868 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U7869 ( .A1(n8764), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U7870 ( .A1(n8765), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6374) );
  OAI211_X1 U7871 ( .C1(n6395), .C2(n10075), .A(n6375), .B(n6374), .ZN(n6376)
         );
  INV_X1 U7872 ( .A(n6376), .ZN(n6377) );
  NAND2_X1 U7873 ( .A1(n6378), .A2(n6377), .ZN(n9042) );
  NAND2_X1 U7874 ( .A1(n9042), .A2(n6486), .ZN(n6379) );
  NAND2_X1 U7875 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  XNOR2_X1 U7876 ( .A(n6381), .B(n6484), .ZN(n6385) );
  AND2_X1 U7877 ( .A1(n9042), .A2(n6499), .ZN(n6382) );
  AOI21_X1 U7878 ( .B1(n9421), .B2(n6486), .A(n6382), .ZN(n6386) );
  XNOR2_X1 U7879 ( .A(n6385), .B(n6386), .ZN(n8543) );
  OAI21_X2 U7880 ( .B1(n6384), .B2(n6383), .A(n8543), .ZN(n8545) );
  INV_X1 U7881 ( .A(n6385), .ZN(n6387) );
  NAND2_X1 U7882 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U7883 ( .A1(n8545), .A2(n6388), .ZN(n6402) );
  INV_X1 U7884 ( .A(n6402), .ZN(n6399) );
  NAND2_X1 U7885 ( .A1(n7774), .A2(n8759), .ZN(n6390) );
  NAND2_X1 U7886 ( .A1(n8761), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6389) );
  INV_X1 U7887 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U7888 ( .A1(n6391), .A2(n10171), .ZN(n6392) );
  AND2_X1 U7889 ( .A1(n6426), .A2(n6392), .ZN(n9193) );
  INV_X1 U7890 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U7891 ( .A1(n6529), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U7892 ( .A1(n8765), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6393) );
  OAI211_X1 U7893 ( .C1(n6395), .C2(n10096), .A(n6394), .B(n6393), .ZN(n6396)
         );
  AOI21_X1 U7894 ( .B1(n9193), .B2(n6074), .A(n6396), .ZN(n9044) );
  OAI22_X1 U7895 ( .A1(n9196), .A2(n6397), .B1(n9044), .B2(n6065), .ZN(n6398)
         );
  XNOR2_X1 U7896 ( .A(n6398), .B(n6484), .ZN(n6400) );
  INV_X1 U7897 ( .A(n6400), .ZN(n6401) );
  OAI22_X1 U7898 ( .A1(n9196), .A2(n6065), .B1(n9044), .B2(n6432), .ZN(n8614)
         );
  NAND2_X1 U7899 ( .A1(n7839), .A2(n8759), .ZN(n6406) );
  NAND2_X1 U7900 ( .A1(n6080), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7901 ( .A1(n9332), .A2(n6433), .ZN(n6414) );
  XNOR2_X1 U7902 ( .A(n6426), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U7903 ( .A1(n9171), .A2(n6074), .ZN(n6412) );
  INV_X1 U7904 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U7905 ( .A1(n8766), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U7906 ( .A1(n8765), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6407) );
  OAI211_X1 U7907 ( .C1(n6480), .C2(n6409), .A(n6408), .B(n6407), .ZN(n6410)
         );
  INV_X1 U7908 ( .A(n6410), .ZN(n6411) );
  NAND2_X1 U7909 ( .A1(n9045), .A2(n6037), .ZN(n6413) );
  NAND2_X1 U7910 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  XNOR2_X1 U7911 ( .A(n6415), .B(n6484), .ZN(n6418) );
  NAND2_X1 U7912 ( .A1(n9332), .A2(n6037), .ZN(n6417) );
  NAND2_X1 U7913 ( .A1(n9045), .A2(n6499), .ZN(n6416) );
  NAND2_X1 U7914 ( .A1(n6417), .A2(n6416), .ZN(n6419) );
  NAND2_X1 U7915 ( .A1(n6418), .A2(n6419), .ZN(n8505) );
  INV_X1 U7916 ( .A(n6418), .ZN(n6421) );
  INV_X1 U7917 ( .A(n6419), .ZN(n6420) );
  NAND2_X1 U7918 ( .A1(n6421), .A2(n6420), .ZN(n8507) );
  NAND2_X1 U7919 ( .A1(n7863), .A2(n8759), .ZN(n6423) );
  NAND2_X1 U7920 ( .A1(n6080), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6422) );
  INV_X1 U7921 ( .A(n6426), .ZN(n6424) );
  AOI21_X1 U7922 ( .B1(n6424), .B2(P1_REG3_REG_23__SCAN_IN), .A(
        P1_REG3_REG_24__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U7923 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n6425) );
  OR2_X1 U7924 ( .A1(n6427), .A2(n6444), .ZN(n9161) );
  INV_X1 U7925 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U7926 ( .A1(n6889), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U7927 ( .A1(n8765), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6428) );
  OAI211_X1 U7928 ( .C1(n6480), .C2(n9330), .A(n6429), .B(n6428), .ZN(n6430)
         );
  INV_X1 U7929 ( .A(n6430), .ZN(n6431) );
  INV_X1 U7930 ( .A(n9048), .ZN(n9050) );
  OAI22_X1 U7931 ( .A1(n9165), .A2(n6065), .B1(n9050), .B2(n6432), .ZN(n6438)
         );
  NAND2_X1 U7932 ( .A1(n9329), .A2(n6433), .ZN(n6435) );
  NAND2_X1 U7933 ( .A1(n9048), .A2(n6486), .ZN(n6434) );
  NAND2_X1 U7934 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  XNOR2_X1 U7935 ( .A(n6436), .B(n6484), .ZN(n6437) );
  XOR2_X1 U7936 ( .A(n6438), .B(n6437), .Z(n8582) );
  INV_X1 U7937 ( .A(n6437), .ZN(n6440) );
  INV_X1 U7938 ( .A(n6438), .ZN(n6439) );
  NAND2_X1 U7939 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U7940 ( .A1(n7869), .A2(n8759), .ZN(n6443) );
  NAND2_X1 U7941 ( .A1(n8761), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6442) );
  NOR2_X1 U7942 ( .A1(n6444), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6445) );
  INV_X1 U7943 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7944 ( .A1(n8766), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U7945 ( .A1(n8765), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6446) );
  OAI211_X1 U7946 ( .C1(n6480), .C2(n6448), .A(n6447), .B(n6446), .ZN(n6449)
         );
  INV_X1 U7947 ( .A(n6449), .ZN(n6450) );
  AND2_X1 U7948 ( .A1(n9052), .A2(n6499), .ZN(n6451) );
  AOI21_X1 U7949 ( .B1(n9408), .B2(n6486), .A(n6451), .ZN(n6453) );
  AOI22_X1 U7950 ( .A1(n9408), .A2(n4603), .B1(n6486), .B2(n9052), .ZN(n6452)
         );
  XNOR2_X1 U7951 ( .A(n6452), .B(n6484), .ZN(n6454) );
  XOR2_X1 U7952 ( .A(n6453), .B(n6454), .Z(n8556) );
  NAND2_X1 U7953 ( .A1(n7875), .A2(n8759), .ZN(n6456) );
  NAND2_X1 U7954 ( .A1(n8761), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U7955 ( .A1(n6457), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6475) );
  OR2_X1 U7956 ( .A1(n6457), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U7957 ( .A1(n6475), .A2(n6458), .ZN(n9123) );
  INV_X1 U7958 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U7959 ( .A1(n6889), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U7960 ( .A1(n8765), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6459) );
  OAI211_X1 U7961 ( .C1(n6480), .C2(n10182), .A(n6460), .B(n6459), .ZN(n6461)
         );
  INV_X1 U7962 ( .A(n6461), .ZN(n6462) );
  AND2_X1 U7963 ( .A1(n8922), .A2(n6499), .ZN(n6464) );
  AOI21_X1 U7964 ( .B1(n9318), .B2(n6486), .A(n6464), .ZN(n6469) );
  NAND2_X1 U7965 ( .A1(n9318), .A2(n4603), .ZN(n6466) );
  NAND2_X1 U7966 ( .A1(n8922), .A2(n6037), .ZN(n6465) );
  NAND2_X1 U7967 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  XNOR2_X1 U7968 ( .A(n6467), .B(n6484), .ZN(n6471) );
  XOR2_X1 U7969 ( .A(n6469), .B(n6471), .Z(n8644) );
  INV_X1 U7970 ( .A(n8644), .ZN(n6468) );
  INV_X1 U7971 ( .A(n6469), .ZN(n6470) );
  NAND2_X1 U7972 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  NAND2_X1 U7973 ( .A1(n8487), .A2(n8759), .ZN(n6474) );
  NAND2_X1 U7974 ( .A1(n8761), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6473) );
  INV_X1 U7975 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10154) );
  NAND2_X1 U7976 ( .A1(n6475), .A2(n10154), .ZN(n6476) );
  NOR2_X1 U7977 ( .A1(n10154), .A2(n6475), .ZN(n6528) );
  INV_X1 U7978 ( .A(n6528), .ZN(n6490) );
  NAND2_X1 U7979 ( .A1(n6476), .A2(n6490), .ZN(n6562) );
  INV_X1 U7980 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U7981 ( .A1(n8766), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7982 ( .A1(n8765), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6478) );
  OAI211_X1 U7983 ( .C1(n6480), .C2(n9315), .A(n6479), .B(n6478), .ZN(n6481)
         );
  INV_X1 U7984 ( .A(n6481), .ZN(n6482) );
  AOI22_X1 U7985 ( .A1(n9113), .A2(n4603), .B1(n6486), .B2(n8921), .ZN(n6485)
         );
  XNOR2_X1 U7986 ( .A(n6485), .B(n6484), .ZN(n6547) );
  AOI22_X1 U7987 ( .A1(n9113), .A2(n6486), .B1(n6499), .B2(n8921), .ZN(n6546)
         );
  XNOR2_X1 U7988 ( .A(n6547), .B(n6546), .ZN(n6556) );
  INV_X1 U7989 ( .A(n6556), .ZN(n6487) );
  NAND2_X1 U7990 ( .A1(n8484), .A2(n8759), .ZN(n6489) );
  NAND2_X1 U7991 ( .A1(n8761), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7992 ( .A1(n9311), .A2(n4603), .ZN(n6496) );
  NAND2_X1 U7993 ( .A1(n6889), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7994 ( .A1(n8764), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6493) );
  XNOR2_X1 U7995 ( .A(P1_REG3_REG_28__SCAN_IN), .B(n6490), .ZN(n9096) );
  NAND2_X1 U7996 ( .A1(n6074), .A2(n9096), .ZN(n6492) );
  NAND2_X1 U7997 ( .A1(n8765), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6491) );
  NAND4_X1 U7998 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n9077)
         );
  NAND2_X1 U7999 ( .A1(n9077), .A2(n6037), .ZN(n6495) );
  NAND2_X1 U8000 ( .A1(n6496), .A2(n6495), .ZN(n6498) );
  XNOR2_X1 U8001 ( .A(n6498), .B(n6497), .ZN(n6501) );
  AOI22_X1 U8002 ( .A1(n9311), .A2(n6486), .B1(n6499), .B2(n9077), .ZN(n6500)
         );
  XNOR2_X1 U8003 ( .A(n6501), .B(n6500), .ZN(n6551) );
  INV_X1 U8004 ( .A(n6551), .ZN(n6524) );
  NAND2_X1 U8005 ( .A1(n7874), .A2(P1_B_REG_SCAN_IN), .ZN(n6502) );
  MUX2_X1 U8006 ( .A(P1_B_REG_SCAN_IN), .B(n6502), .S(n7868), .Z(n6503) );
  INV_X1 U8007 ( .A(n6504), .ZN(n9468) );
  NAND2_X1 U8008 ( .A1(n9468), .A2(n7868), .ZN(n6505) );
  NAND2_X1 U8009 ( .A1(n6506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6507) );
  AND2_X1 U8010 ( .A1(n7840), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6508) );
  INV_X1 U8011 ( .A(n9638), .ZN(n9612) );
  OR2_X1 U8012 ( .A1(n7077), .A2(n9612), .ZN(n9636) );
  NAND2_X1 U8013 ( .A1(n9468), .A2(n7874), .ZN(n6509) );
  OAI21_X1 U8014 ( .B1(n9610), .B2(P1_D_REG_1__SCAN_IN), .A(n6509), .ZN(n7032)
         );
  NOR4_X1 U8015 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6513) );
  NOR4_X1 U8016 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6512) );
  NOR4_X1 U8017 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6511) );
  NOR4_X1 U8018 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6510) );
  NAND4_X1 U8019 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(n6519)
         );
  NOR2_X1 U8020 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .ZN(
        n6517) );
  NOR4_X1 U8021 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6516) );
  NOR4_X1 U8022 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6515) );
  NOR4_X1 U8023 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6514) );
  NAND4_X1 U8024 ( .A1(n6517), .A2(n6516), .A3(n6515), .A4(n6514), .ZN(n6518)
         );
  NOR2_X1 U8025 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NOR2_X1 U8026 ( .A1(n9610), .A2(n6520), .ZN(n7031) );
  NOR2_X1 U8027 ( .A1(n9636), .A2(n6535), .ZN(n6523) );
  NAND2_X1 U8028 ( .A1(n8900), .A2(n7024), .ZN(n9654) );
  NAND2_X1 U8029 ( .A1(n8911), .A2(n8852), .ZN(n8845) );
  AND2_X1 U8030 ( .A1(n9654), .A2(n8845), .ZN(n6538) );
  NAND2_X1 U8031 ( .A1(n6524), .A2(n8634), .ZN(n6555) );
  INV_X1 U8032 ( .A(n9636), .ZN(n6536) );
  INV_X1 U8033 ( .A(n6535), .ZN(n7079) );
  INV_X1 U8034 ( .A(n8808), .ZN(n8895) );
  NAND2_X1 U8035 ( .A1(n7024), .A2(n8895), .ZN(n7081) );
  INV_X1 U8036 ( .A(n7081), .ZN(n6525) );
  NAND3_X1 U8037 ( .A1(n6536), .A2(n7079), .A3(n6525), .ZN(n6527) );
  NAND2_X1 U8038 ( .A1(n9638), .A2(n6522), .ZN(n6526) );
  OR2_X1 U8039 ( .A1(n6791), .A2(n8845), .ZN(n8508) );
  AND2_X1 U8040 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n6528), .ZN(n9082) );
  NAND2_X1 U8041 ( .A1(n6074), .A2(n9082), .ZN(n6533) );
  NAND2_X1 U8042 ( .A1(n6529), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8043 ( .A1(n8765), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8044 ( .A1(n8766), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6530) );
  NAND4_X1 U8045 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n8920)
         );
  INV_X1 U8046 ( .A(n8845), .ZN(n6666) );
  AND2_X1 U8047 ( .A1(n8920), .A2(n9012), .ZN(n6534) );
  AOI21_X1 U8048 ( .B1(n8921), .B2(n8595), .A(n6534), .ZN(n9091) );
  NOR2_X1 U8049 ( .A1(n6535), .A2(n8900), .ZN(n6537) );
  INV_X1 U8050 ( .A(n7077), .ZN(n7120) );
  NAND2_X1 U8051 ( .A1(n7079), .A2(n7120), .ZN(n6543) );
  NAND2_X1 U8052 ( .A1(n6543), .A2(n6538), .ZN(n6946) );
  NAND2_X1 U8053 ( .A1(n8900), .A2(n6666), .ZN(n6944) );
  NAND4_X1 U8054 ( .A1(n6946), .A2(n7840), .A3(n6021), .A4(n6944), .ZN(n6539)
         );
  NAND2_X1 U8055 ( .A1(n6539), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6544) );
  OR2_X1 U8056 ( .A1(n6540), .A2(n6541), .ZN(n7084) );
  OR2_X1 U8057 ( .A1(n7084), .A2(n9612), .ZN(n8899) );
  OAI21_X1 U8058 ( .B1(P1_U3086), .B2(n7081), .A(n8899), .ZN(n6542) );
  NAND2_X1 U8059 ( .A1(n6543), .A2(n6542), .ZN(n6945) );
  AOI22_X1 U8060 ( .A1(n8656), .A2(n9096), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        n4437), .ZN(n6545) );
  OAI21_X1 U8061 ( .B1(n9091), .B2(n9489), .A(n6545), .ZN(n6549) );
  NAND2_X1 U8062 ( .A1(n6547), .A2(n6546), .ZN(n6550) );
  NOR3_X1 U8063 ( .A1(n6551), .A2(n9493), .A3(n6550), .ZN(n6548) );
  AOI211_X1 U8064 ( .C1(n9311), .C2(n9497), .A(n6549), .B(n6548), .ZN(n6554)
         );
  AND2_X1 U8065 ( .A1(n6551), .A2(n5052), .ZN(n6552) );
  OAI211_X1 U8066 ( .C1(n6559), .C2(n6555), .A(n6554), .B(n6553), .ZN(P1_U3220) );
  NAND2_X1 U8067 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  NAND2_X1 U8068 ( .A1(n6560), .A2(n8634), .ZN(n6567) );
  AND2_X1 U8069 ( .A1(n9077), .A2(n9012), .ZN(n6561) );
  AOI21_X1 U8070 ( .B1(n8922), .B2(n8595), .A(n6561), .ZN(n9110) );
  NAND2_X1 U8071 ( .A1(n9113), .A2(n9497), .ZN(n6564) );
  INV_X1 U8072 ( .A(n6562), .ZN(n9114) );
  AOI22_X1 U8073 ( .A1(n9114), .A2(n8656), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6563) );
  OAI211_X1 U8074 ( .C1(n9110), .C2(n9489), .A(n6564), .B(n6563), .ZN(n6565)
         );
  INV_X1 U8075 ( .A(n6565), .ZN(n6566) );
  NAND2_X1 U8076 ( .A1(n6567), .A2(n6566), .ZN(P1_U3214) );
  OR2_X1 U8077 ( .A1(n6636), .A2(n6568), .ZN(n6816) );
  AND3_X1 U8078 ( .A1(n6660), .A2(n6569), .A3(n6816), .ZN(n6571) );
  OR2_X1 U8079 ( .A1(n9902), .A2(n6917), .ZN(n6623) );
  NAND2_X1 U8080 ( .A1(n6916), .A2(n6623), .ZN(n6574) );
  NAND3_X1 U8081 ( .A1(n6572), .A2(n6918), .A3(n8125), .ZN(n6573) );
  NAND2_X1 U8082 ( .A1(n6574), .A2(n6617), .ZN(n6576) );
  INV_X1 U8083 ( .A(n6617), .ZN(n6616) );
  NAND2_X1 U8084 ( .A1(n6618), .A2(n6616), .ZN(n6575) );
  NAND2_X1 U8085 ( .A1(n6578), .A2(n9929), .ZN(n6581) );
  NAND2_X1 U8086 ( .A1(n6581), .A2(n6580), .ZN(P2_U3488) );
  XOR2_X1 U8087 ( .A(n7959), .B(n6582), .Z(n6631) );
  INV_X1 U8088 ( .A(n7966), .ZN(n6613) );
  OAI22_X1 U8089 ( .A1(n6631), .A2(n8381), .B1(n6613), .B2(n8352), .ZN(n6583)
         );
  INV_X1 U8090 ( .A(n6583), .ZN(n6585) );
  NAND2_X1 U8091 ( .A1(n9927), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6584) );
  INV_X1 U8092 ( .A(n7959), .ZN(n6587) );
  XNOR2_X1 U8093 ( .A(n6587), .B(n6586), .ZN(n6591) );
  NOR2_X1 U8094 ( .A1(n9861), .A2(n7961), .ZN(n6589) );
  INV_X1 U8095 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6602) );
  XNOR2_X1 U8096 ( .A(n6594), .B(n6595), .ZN(n8165) );
  INV_X1 U8097 ( .A(n6595), .ZN(n6596) );
  XNOR2_X1 U8098 ( .A(n6597), .B(n6596), .ZN(n6601) );
  AOI21_X1 U8099 ( .B1(n9914), .B2(n8165), .A(n8160), .ZN(n6606) );
  MUX2_X1 U8100 ( .A(n6602), .B(n6606), .S(n8378), .Z(n6605) );
  NAND2_X1 U8101 ( .A1(n5919), .A2(n6603), .ZN(n6604) );
  NAND2_X1 U8102 ( .A1(n6605), .A2(n6604), .ZN(P2_U3486) );
  INV_X1 U8103 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6607) );
  MUX2_X1 U8104 ( .A(n6607), .B(n6606), .S(n9915), .Z(n6610) );
  NAND2_X1 U8105 ( .A1(n5919), .A2(n6608), .ZN(n6609) );
  NAND2_X1 U8106 ( .A1(n6610), .A2(n6609), .ZN(P2_U3454) );
  NAND2_X1 U8107 ( .A1(n9917), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6611) );
  OAI22_X1 U8108 ( .A1(n6631), .A2(n8470), .B1(n6613), .B2(n8413), .ZN(n6614)
         );
  INV_X1 U8109 ( .A(n6614), .ZN(n6615) );
  NAND2_X1 U8110 ( .A1(n5041), .A2(n6615), .ZN(P2_U3455) );
  NAND2_X1 U8111 ( .A1(n4806), .A2(n6616), .ZN(n6620) );
  NAND2_X1 U8112 ( .A1(n6618), .A2(n6617), .ZN(n6619) );
  AND2_X1 U8113 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  INV_X1 U8114 ( .A(n6623), .ZN(n6624) );
  NAND2_X1 U8115 ( .A1(n6625), .A2(n8318), .ZN(n6634) );
  AND2_X1 U8116 ( .A1(n6917), .A2(n9853), .ZN(n9869) );
  INV_X1 U8117 ( .A(n9869), .ZN(n6626) );
  NAND2_X1 U8118 ( .A1(n7615), .A2(n6626), .ZN(n6627) );
  AOI22_X1 U8119 ( .A1(n7966), .A2(n8304), .B1(n8303), .B2(n7962), .ZN(n6630)
         );
  OAI21_X1 U8120 ( .B1(n6631), .B2(n8339), .A(n5051), .ZN(n6632) );
  INV_X1 U8121 ( .A(n6632), .ZN(n6633) );
  NAND2_X1 U8122 ( .A1(n6634), .A2(n6633), .ZN(P2_U3205) );
  INV_X1 U8123 ( .A(n7840), .ZN(n6635) );
  NAND2_X1 U8124 ( .A1(n6636), .A2(n6814), .ZN(n6637) );
  NAND2_X1 U8125 ( .A1(n6637), .A2(n6815), .ZN(n6694) );
  NAND2_X1 U8126 ( .A1(n6694), .A2(n5276), .ZN(n6638) );
  NAND2_X1 U8127 ( .A1(n6638), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8128 ( .A1(n6814), .A2(P2_U3151), .ZN(n6639) );
  NOR2_X2 U8129 ( .A1(n6640), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9462) );
  AOI22_X1 U8130 ( .A1(n9462), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n7052), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6641) );
  OAI21_X1 U8131 ( .B1(n6647), .B2(n7778), .A(n6641), .ZN(P1_U3353) );
  AOI22_X1 U8132 ( .A1(n8950), .A2(P1_STATE_REG_SCAN_IN), .B1(n9462), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6642) );
  OAI21_X1 U8133 ( .B1(n6645), .B2(n7778), .A(n6642), .ZN(P1_U3352) );
  NAND2_X1 U8134 ( .A1(n6643), .A2(P2_U3151), .ZN(n6677) );
  INV_X2 U8135 ( .A(n8489), .ZN(n8480) );
  OAI222_X1 U8136 ( .A1(n8483), .A2(n6652), .B1(n6719), .B2(P2_U3151), .C1(
        n4906), .C2(n8480), .ZN(P2_U3294) );
  INV_X1 U8137 ( .A(n9684), .ZN(n6766) );
  INV_X1 U8138 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6644) );
  OAI222_X1 U8139 ( .A1(n8483), .A2(n6645), .B1(n6766), .B2(P2_U3151), .C1(
        n6644), .C2(n8480), .ZN(P2_U3292) );
  INV_X1 U8140 ( .A(n6763), .ZN(n6744) );
  INV_X1 U8141 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6646) );
  OAI222_X1 U8142 ( .A1(n8483), .A2(n6647), .B1(n6744), .B2(P2_U3151), .C1(
        n6646), .C2(n8480), .ZN(P2_U3293) );
  INV_X1 U8143 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6895) );
  INV_X1 U8144 ( .A(n6905), .ZN(n6909) );
  OAI222_X1 U8145 ( .A1(n8483), .A2(n6657), .B1(n8480), .B2(n6895), .C1(
        P2_U3151), .C2(n6909), .ZN(P2_U3291) );
  NAND2_X1 U8146 ( .A1(n6660), .A2(n6648), .ZN(n6649) );
  OAI21_X1 U8147 ( .B1(n6660), .B2(n5951), .A(n6649), .ZN(P2_U3377) );
  AOI22_X1 U8148 ( .A1(n6838), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9462), .ZN(n6650) );
  OAI21_X1 U8149 ( .B1(n6654), .B2(n7778), .A(n6650), .ZN(P1_U3350) );
  AOI22_X1 U8150 ( .A1(n9462), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n8943), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6651) );
  OAI21_X1 U8151 ( .B1(n6652), .B2(n7778), .A(n6651), .ZN(P1_U3354) );
  INV_X1 U8152 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6653) );
  OAI222_X1 U8153 ( .A1(n8483), .A2(n6654), .B1(n4697), .B2(P2_U3151), .C1(
        n6653), .C2(n8480), .ZN(P2_U3290) );
  NAND2_X1 U8154 ( .A1(n9612), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6655) );
  OAI21_X1 U8155 ( .B1(n9612), .B2(n7032), .A(n6655), .ZN(P1_U3440) );
  INV_X1 U8156 ( .A(n6802), .ZN(n8963) );
  INV_X1 U8157 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6656) );
  OAI222_X1 U8158 ( .A1(P1_U3086), .A2(n8963), .B1(n7778), .B2(n6657), .C1(
        n6656), .C2(n9466), .ZN(P1_U3351) );
  INV_X1 U8159 ( .A(n6658), .ZN(n6659) );
  NAND2_X1 U8160 ( .A1(n6660), .A2(n6659), .ZN(n9963) );
  AND4_X1 U8161 ( .A1(n6815), .A2(P2_STATE_REG_SCAN_IN), .A3(n7877), .A4(n7865), .ZN(n6661) );
  AOI21_X1 U8162 ( .B1(n9963), .B2(n5938), .A(n6661), .ZN(P2_U3376) );
  AND2_X1 U8163 ( .A1(n9963), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8164 ( .A1(n9963), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8165 ( .A1(n9963), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8166 ( .A1(n9963), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8167 ( .A1(n9963), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8168 ( .A1(n9963), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8169 ( .A1(n9963), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8170 ( .A1(n9963), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8171 ( .A1(n9963), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8172 ( .A1(n9963), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8173 ( .A1(n9963), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8174 ( .A1(n9963), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8175 ( .A1(n9963), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8176 ( .A1(n9963), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8177 ( .A1(n9963), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8178 ( .A1(n9963), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8179 ( .A1(n9963), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8180 ( .A1(n9963), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8181 ( .A1(n9963), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8182 ( .A1(n9963), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AOI22_X1 U8183 ( .A1(n6852), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9462), .ZN(n6662) );
  OAI21_X1 U8184 ( .B1(n6679), .B2(n7778), .A(n6662), .ZN(P1_U3348) );
  INV_X1 U8185 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U8186 ( .A1(n6663), .A2(n10175), .ZN(P2_U3251) );
  INV_X1 U8187 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U8188 ( .A1(n6663), .A2(n10158), .ZN(P2_U3240) );
  INV_X1 U8189 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10070) );
  NOR2_X1 U8190 ( .A1(n6663), .A2(n10070), .ZN(P2_U3234) );
  INV_X1 U8191 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U8192 ( .A1(n6663), .A2(n10055), .ZN(P2_U3243) );
  INV_X1 U8193 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U8194 ( .A1(n6663), .A2(n10061), .ZN(P2_U3244) );
  INV_X1 U8195 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U8196 ( .A1(n6663), .A2(n10198), .ZN(P2_U3237) );
  INV_X1 U8197 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U8198 ( .A1(n6663), .A2(n10092), .ZN(P2_U3238) );
  INV_X1 U8199 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U8200 ( .A1(n6663), .A2(n10106), .ZN(P2_U3245) );
  INV_X1 U8201 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10241) );
  NOR2_X1 U8202 ( .A1(n6663), .A2(n10241), .ZN(P2_U3250) );
  INV_X1 U8203 ( .A(n7041), .ZN(n9463) );
  INV_X1 U8204 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7090) );
  AOI21_X1 U8205 ( .B1(n9463), .B2(n7090), .A(n6791), .ZN(n7043) );
  OAI21_X1 U8206 ( .B1(n9463), .B2(P1_REG1_REG_0__SCAN_IN), .A(n7043), .ZN(
        n6664) );
  XOR2_X1 U8207 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6664), .Z(n6674) );
  NAND2_X1 U8208 ( .A1(n6666), .A2(n7840), .ZN(n6667) );
  AND2_X1 U8209 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  AND2_X1 U8210 ( .A1(n6670), .A2(n6669), .ZN(n6803) );
  INV_X1 U8211 ( .A(n6803), .ZN(n6673) );
  INV_X1 U8212 ( .A(n6669), .ZN(n6671) );
  AND2_X1 U8213 ( .A1(n6671), .A2(n6670), .ZN(n9547) );
  AOI22_X1 U8214 ( .A1(n9547), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n4437), .ZN(n6672) );
  OAI21_X1 U8215 ( .B1(n6674), .B2(n6673), .A(n6672), .ZN(P1_U3243) );
  INV_X1 U8216 ( .A(n6865), .ZN(n6676) );
  INV_X1 U8217 ( .A(n6675), .ZN(n6678) );
  INV_X1 U8218 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6692) );
  OAI222_X1 U8219 ( .A1(n4437), .A2(n6676), .B1(n7778), .B2(n6678), .C1(n9466), 
        .C2(n6692), .ZN(P1_U3349) );
  INV_X1 U8220 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10176) );
  OAI222_X1 U8221 ( .A1(n8480), .A2(n10176), .B1(n8483), .B2(n6678), .C1(
        P2_U3151), .C2(n4622), .ZN(P2_U3289) );
  OAI222_X1 U8222 ( .A1(n8483), .A2(n6679), .B1(n7226), .B2(P2_U3151), .C1(
        n10071), .C2(n8480), .ZN(P2_U3288) );
  INV_X1 U8223 ( .A(n6680), .ZN(n6683) );
  AOI22_X1 U8224 ( .A1(n6877), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9462), .ZN(n6681) );
  OAI21_X1 U8225 ( .B1(n6683), .B2(n7778), .A(n6681), .ZN(P1_U3347) );
  NAND2_X1 U8226 ( .A1(n7650), .A2(P2_U3893), .ZN(n6682) );
  OAI21_X1 U8227 ( .B1(P2_U3893), .B2(n5094), .A(n6682), .ZN(P2_U3500) );
  INV_X1 U8228 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6684) );
  INV_X1 U8229 ( .A(n7338), .ZN(n7239) );
  OAI222_X1 U8230 ( .A1(n8480), .A2(n6684), .B1(n8483), .B2(n6683), .C1(
        P2_U3151), .C2(n7239), .ZN(P2_U3287) );
  INV_X1 U8231 ( .A(n6685), .ZN(n6688) );
  INV_X1 U8232 ( .A(n8133), .ZN(n8105) );
  OAI222_X1 U8233 ( .A1(n8483), .A2(n6688), .B1(n8105), .B2(P2_U3151), .C1(
        n6686), .C2(n8480), .ZN(P2_U3286) );
  AOI22_X1 U8234 ( .A1(n7012), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9462), .ZN(n6687) );
  OAI21_X1 U8235 ( .B1(n6690), .B2(n7778), .A(n6687), .ZN(P1_U3345) );
  INV_X1 U8236 ( .A(n6954), .ZN(n6884) );
  OAI222_X1 U8237 ( .A1(n4437), .A2(n6884), .B1(n9466), .B2(n5094), .C1(n6688), 
        .C2(n7778), .ZN(P1_U3346) );
  INV_X1 U8238 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6689) );
  OAI222_X1 U8239 ( .A1(n8483), .A2(n6690), .B1(n8130), .B2(P2_U3151), .C1(
        n6689), .C2(n8480), .ZN(P2_U3285) );
  NAND2_X1 U8240 ( .A1(n4764), .A2(P2_U3893), .ZN(n6691) );
  OAI21_X1 U8241 ( .B1(P2_U3893), .B2(n6692), .A(n6691), .ZN(P2_U3497) );
  NOR2_X1 U8242 ( .A1(n8118), .A2(P2_U3151), .ZN(n8488) );
  NAND2_X1 U8243 ( .A1(n6694), .A2(n8488), .ZN(n6693) );
  MUX2_X1 U8244 ( .A(n6693), .B(n9475), .S(n6713), .Z(n9696) );
  NOR2_X1 U8245 ( .A1(n5876), .A2(P2_U3151), .ZN(n8485) );
  NAND2_X1 U8246 ( .A1(n8485), .A2(n6694), .ZN(n9668) );
  INV_X1 U8247 ( .A(n9845), .ZN(n9740) );
  INV_X1 U8248 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6700) );
  AND2_X1 U8249 ( .A1(n6700), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8250 ( .A1(n6701), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6727) );
  OAI21_X1 U8251 ( .B1(n6719), .B2(n6695), .A(n6727), .ZN(n6696) );
  INV_X1 U8252 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10128) );
  OR2_X1 U8253 ( .A1(n6696), .A2(n10128), .ZN(n6728) );
  NAND2_X1 U8254 ( .A1(n6696), .A2(n10128), .ZN(n6697) );
  NAND2_X1 U8255 ( .A1(n6728), .A2(n6697), .ZN(n6710) );
  INV_X1 U8256 ( .A(n6814), .ZN(n6698) );
  AND2_X1 U8257 ( .A1(n6698), .A2(n6815), .ZN(n6699) );
  INV_X1 U8258 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U8259 ( .A1(n6908), .A2(n9934), .ZN(n6709) );
  NAND2_X1 U8260 ( .A1(n6701), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8261 ( .A1(n6719), .A2(n6734), .ZN(n6704) );
  NAND2_X1 U8262 ( .A1(n6700), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6702) );
  OR2_X1 U8263 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  NAND2_X1 U8264 ( .A1(n6704), .A2(n6703), .ZN(n6733) );
  XNOR2_X1 U8265 ( .A(n6733), .B(n6705), .ZN(n6707) );
  OAI22_X1 U8266 ( .A1(n9699), .A2(n6707), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6706), .ZN(n6708) );
  AOI211_X1 U8267 ( .C1(n9740), .C2(n6710), .A(n6709), .B(n6708), .ZN(n6718)
         );
  INV_X1 U8268 ( .A(n6711), .ZN(n6745) );
  MUX2_X1 U8269 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6745), .Z(n6720) );
  XOR2_X1 U8270 ( .A(n6719), .B(n6720), .Z(n6716) );
  INV_X1 U8271 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6990) );
  INV_X1 U8272 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6712) );
  MUX2_X1 U8273 ( .A(n6990), .B(n6712), .S(n6745), .Z(n9669) );
  NAND2_X1 U8274 ( .A1(n9669), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U8275 ( .A1(n6716), .A2(n6715), .ZN(n6721) );
  OAI211_X1 U8276 ( .C1(n6716), .C2(n6715), .A(n6721), .B(n6714), .ZN(n6717)
         );
  OAI211_X1 U8277 ( .C1(n9696), .C2(n6719), .A(n6718), .B(n6717), .ZN(P2_U3183) );
  INV_X1 U8278 ( .A(n6719), .ZN(n6723) );
  INV_X1 U8279 ( .A(n6720), .ZN(n6722) );
  OAI21_X1 U8280 ( .B1(n6723), .B2(n6722), .A(n6721), .ZN(n6726) );
  MUX2_X1 U8281 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6724), .Z(n6746) );
  XNOR2_X1 U8282 ( .A(n6746), .B(n6763), .ZN(n6725) );
  NAND2_X1 U8283 ( .A1(n6726), .A2(n6725), .ZN(n6747) );
  OAI211_X1 U8284 ( .C1(n6726), .C2(n6725), .A(n6747), .B(n6714), .ZN(n6743)
         );
  INV_X1 U8285 ( .A(n6908), .ZN(n9830) );
  NAND2_X1 U8286 ( .A1(n6728), .A2(n6727), .ZN(n6729) );
  OAI21_X1 U8287 ( .B1(n6730), .B2(n6729), .A(n6765), .ZN(n6731) );
  NAND2_X1 U8288 ( .A1(n9740), .A2(n6731), .ZN(n6740) );
  MUX2_X1 U8289 ( .A(n6732), .B(P2_REG1_REG_2__SCAN_IN), .S(n6763), .Z(n6737)
         );
  NAND2_X1 U8290 ( .A1(n6733), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U8291 ( .A1(n6735), .A2(n6734), .ZN(n6736) );
  NAND2_X1 U8292 ( .A1(n6737), .A2(n6736), .ZN(n6754) );
  OAI21_X1 U8293 ( .B1(n6737), .B2(n6736), .A(n6754), .ZN(n6738) );
  NAND2_X1 U8294 ( .A1(n9839), .A2(n6738), .ZN(n6739) );
  OAI211_X1 U8295 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9856), .A(n6740), .B(n6739), .ZN(n6741) );
  AOI21_X1 U8296 ( .B1(n9830), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n6741), .ZN(
        n6742) );
  OAI211_X1 U8297 ( .C1(n9696), .C2(n6744), .A(n6743), .B(n6742), .ZN(P2_U3184) );
  MUX2_X1 U8298 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6745), .Z(n6749) );
  INV_X1 U8299 ( .A(n6749), .ZN(n6750) );
  INV_X1 U8300 ( .A(n6746), .ZN(n6748) );
  OAI21_X1 U8301 ( .B1(n6763), .B2(n6748), .A(n6747), .ZN(n9686) );
  XNOR2_X1 U8302 ( .A(n6749), .B(n6766), .ZN(n9687) );
  NOR2_X1 U8303 ( .A1(n9686), .A2(n9687), .ZN(n9685) );
  AOI21_X1 U8304 ( .B1(n9684), .B2(n6750), .A(n9685), .ZN(n6752) );
  MUX2_X1 U8305 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8118), .Z(n6902) );
  XNOR2_X1 U8306 ( .A(n6902), .B(n6905), .ZN(n6751) );
  NAND2_X1 U8307 ( .A1(n6752), .A2(n6751), .ZN(n6903) );
  OAI211_X1 U8308 ( .C1(n6752), .C2(n6751), .A(n6903), .B(n6714), .ZN(n6778)
         );
  NAND2_X1 U8309 ( .A1(n9830), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n6775) );
  OR2_X1 U8310 ( .A1(n6763), .A2(n6732), .ZN(n6753) );
  NAND2_X1 U8311 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  XNOR2_X1 U8312 ( .A(n6755), .B(n9684), .ZN(n9678) );
  NAND2_X1 U8313 ( .A1(n9678), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8314 ( .A1(n6755), .A2(n6766), .ZN(n6756) );
  INV_X1 U8315 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6758) );
  MUX2_X1 U8316 ( .A(n6758), .B(P2_REG1_REG_4__SCAN_IN), .S(n6905), .Z(n6759)
         );
  NOR2_X1 U8317 ( .A1(n6760), .A2(n6759), .ZN(n6761) );
  OAI21_X1 U8318 ( .B1(n6901), .B2(n6761), .A(n9839), .ZN(n6774) );
  OR2_X1 U8319 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  NAND2_X1 U8320 ( .A1(n6765), .A2(n6764), .ZN(n6767) );
  NAND2_X1 U8321 ( .A1(n6767), .A2(n6766), .ZN(n6769) );
  NAND2_X1 U8322 ( .A1(n6769), .A2(n6768), .ZN(n9676) );
  INV_X1 U8323 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9677) );
  INV_X1 U8324 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7209) );
  XNOR2_X1 U8325 ( .A(n6905), .B(n7209), .ZN(n6770) );
  NAND3_X1 U8326 ( .A1(n9674), .A2(n6770), .A3(n6769), .ZN(n6771) );
  NAND2_X1 U8327 ( .A1(n4700), .A2(n6771), .ZN(n6772) );
  NAND2_X1 U8328 ( .A1(n9740), .A2(n6772), .ZN(n6773) );
  NAND2_X1 U8329 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7097) );
  NAND4_X1 U8330 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n7097), .ZN(n6776)
         );
  AOI21_X1 U8331 ( .B1(n6905), .B2(n9832), .A(n6776), .ZN(n6777) );
  NAND2_X1 U8332 ( .A1(n6778), .A2(n6777), .ZN(P2_U3186) );
  INV_X1 U8333 ( .A(n6779), .ZN(n6871) );
  AOI22_X1 U8334 ( .A1(n7139), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9462), .ZN(n6780) );
  OAI21_X1 U8335 ( .B1(n6871), .B2(n7778), .A(n6780), .ZN(P1_U3344) );
  INV_X1 U8336 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8337 ( .A1(n6803), .A2(n6791), .ZN(n9565) );
  NAND2_X1 U8338 ( .A1(n9577), .A2(n6838), .ZN(n6781) );
  NAND2_X1 U8339 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7427) );
  OAI211_X1 U8340 ( .C1(n9585), .C2(n6782), .A(n6781), .B(n7427), .ZN(n6808)
         );
  INV_X1 U8341 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6783) );
  XNOR2_X1 U8342 ( .A(n7052), .B(n6783), .ZN(n7048) );
  INV_X1 U8343 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6784) );
  XNOR2_X1 U8344 ( .A(n8943), .B(n6784), .ZN(n8939) );
  AND2_X1 U8345 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8938) );
  NAND2_X1 U8346 ( .A1(n8939), .A2(n8938), .ZN(n8937) );
  NAND2_X1 U8347 ( .A1(n8943), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8348 ( .A1(n8937), .A2(n6785), .ZN(n7047) );
  NAND2_X1 U8349 ( .A1(n7048), .A2(n7047), .ZN(n7046) );
  NAND2_X1 U8350 ( .A1(n7052), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8351 ( .A1(n7046), .A2(n6786), .ZN(n8952) );
  INV_X1 U8352 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6787) );
  XNOR2_X1 U8353 ( .A(n8950), .B(n6787), .ZN(n8953) );
  NAND2_X1 U8354 ( .A1(n8952), .A2(n8953), .ZN(n8951) );
  NAND2_X1 U8355 ( .A1(n8950), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8356 ( .A1(n8951), .A2(n6788), .ZN(n8966) );
  INV_X1 U8357 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6789) );
  XNOR2_X1 U8358 ( .A(n6802), .B(n6789), .ZN(n8967) );
  NAND2_X1 U8359 ( .A1(n8966), .A2(n8967), .ZN(n8965) );
  INV_X1 U8360 ( .A(n8965), .ZN(n6790) );
  XNOR2_X1 U8361 ( .A(n6838), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6793) );
  NOR2_X1 U8362 ( .A1(n6794), .A2(n6793), .ZN(n6832) );
  INV_X1 U8363 ( .A(n6791), .ZN(n9459) );
  NAND2_X1 U8364 ( .A1(n9459), .A2(n9463), .ZN(n8898) );
  INV_X1 U8365 ( .A(n8898), .ZN(n6792) );
  NAND2_X1 U8366 ( .A1(n6803), .A2(n6792), .ZN(n9541) );
  AOI211_X1 U8367 ( .C1(n6794), .C2(n6793), .A(n6832), .B(n9541), .ZN(n6807)
         );
  INV_X1 U8368 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6795) );
  XNOR2_X1 U8369 ( .A(n7052), .B(n6795), .ZN(n7051) );
  INV_X1 U8370 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6796) );
  XNOR2_X1 U8371 ( .A(n8943), .B(n6796), .ZN(n8942) );
  AND2_X1 U8372 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8941) );
  NAND2_X1 U8373 ( .A1(n8942), .A2(n8941), .ZN(n8940) );
  NAND2_X1 U8374 ( .A1(n8943), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8375 ( .A1(n8940), .A2(n6797), .ZN(n7050) );
  NAND2_X1 U8376 ( .A1(n7051), .A2(n7050), .ZN(n7049) );
  NAND2_X1 U8377 ( .A1(n7052), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8378 ( .A1(n7049), .A2(n6798), .ZN(n8955) );
  INV_X1 U8379 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6799) );
  XNOR2_X1 U8380 ( .A(n8950), .B(n6799), .ZN(n8956) );
  NAND2_X1 U8381 ( .A1(n8955), .A2(n8956), .ZN(n8954) );
  NAND2_X1 U8382 ( .A1(n8950), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8383 ( .A1(n8954), .A2(n6800), .ZN(n8970) );
  INV_X1 U8384 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6801) );
  XNOR2_X1 U8385 ( .A(n6802), .B(n6801), .ZN(n8971) );
  AND2_X1 U8386 ( .A1(n8970), .A2(n8971), .ZN(n8968) );
  XNOR2_X1 U8387 ( .A(n6838), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6804) );
  NOR2_X1 U8388 ( .A1(n6805), .A2(n6804), .ZN(n6837) );
  NAND2_X1 U8389 ( .A1(n6803), .A2(n7041), .ZN(n9574) );
  AOI211_X1 U8390 ( .C1(n6805), .C2(n6804), .A(n6837), .B(n9574), .ZN(n6806)
         );
  OR3_X1 U8391 ( .A1(n6808), .A2(n6807), .A3(n6806), .ZN(P1_U3248) );
  INV_X1 U8392 ( .A(n6896), .ZN(n6986) );
  OR2_X1 U8393 ( .A1(n6924), .A2(n6819), .ZN(n6811) );
  OR2_X1 U8394 ( .A1(n6827), .A2(n6809), .ZN(n6810) );
  AND2_X2 U8395 ( .A1(n6811), .A2(n6810), .ZN(n8050) );
  OR2_X1 U8396 ( .A1(n6813), .A2(n6812), .ZN(n6818) );
  AND3_X1 U8397 ( .A1(n6816), .A2(n6815), .A3(n6814), .ZN(n6817) );
  OAI211_X1 U8398 ( .C1(n6822), .C2(n6819), .A(n6818), .B(n6817), .ZN(n6820)
         );
  NAND2_X1 U8399 ( .A1(n6820), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6824) );
  OR2_X1 U8400 ( .A1(n6822), .A2(n6821), .ZN(n6823) );
  INV_X1 U8401 ( .A(n8062), .ZN(n7989) );
  NAND2_X1 U8402 ( .A1(n7989), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8403 ( .A1(n6937), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U8404 ( .A1(n6825), .A2(n6985), .ZN(n6826) );
  OR2_X1 U8405 ( .A1(n6827), .A2(n9909), .ZN(n6828) );
  AOI22_X1 U8406 ( .A1(n8042), .A2(n8079), .B1(n8047), .B2(n6829), .ZN(n6830)
         );
  OAI211_X1 U8407 ( .C1(n6986), .C2(n8050), .A(n6831), .B(n6830), .ZN(P2_U3172) );
  INV_X1 U8408 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6833) );
  MUX2_X1 U8409 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6833), .S(n6865), .Z(n6834)
         );
  INV_X1 U8410 ( .A(n6834), .ZN(n6860) );
  NOR2_X1 U8411 ( .A1(n6861), .A2(n6860), .ZN(n6859) );
  AOI21_X1 U8412 ( .B1(n6865), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6859), .ZN(
        n6848) );
  XNOR2_X1 U8413 ( .A(n6852), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U8414 ( .A1(n6848), .A2(n6847), .ZN(n6846) );
  XNOR2_X1 U8415 ( .A(n6877), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6835) );
  NOR2_X1 U8416 ( .A1(n6836), .A2(n6835), .ZN(n6876) );
  AOI211_X1 U8417 ( .C1(n6836), .C2(n6835), .A(n9541), .B(n6876), .ZN(n6845)
         );
  INV_X1 U8418 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6839) );
  MUX2_X1 U8419 ( .A(n6839), .B(P1_REG1_REG_6__SCAN_IN), .S(n6865), .Z(n6863)
         );
  NOR2_X1 U8420 ( .A1(n6864), .A2(n6863), .ZN(n6862) );
  AOI21_X1 U8421 ( .B1(n6865), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6862), .ZN(
        n6851) );
  XNOR2_X1 U8422 ( .A(n6852), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U8423 ( .A1(n6851), .A2(n6850), .ZN(n6849) );
  XNOR2_X1 U8424 ( .A(n6877), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6840) );
  NOR2_X1 U8425 ( .A1(n6841), .A2(n6840), .ZN(n6872) );
  AOI211_X1 U8426 ( .C1(n6841), .C2(n6840), .A(n9574), .B(n6872), .ZN(n6844)
         );
  INV_X1 U8427 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U8428 ( .A1(n9577), .A2(n6877), .ZN(n6842) );
  NAND2_X1 U8429 ( .A1(n4437), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7589) );
  OAI211_X1 U8430 ( .C1(n9585), .C2(n10076), .A(n6842), .B(n7589), .ZN(n6843)
         );
  OR3_X1 U8431 ( .A1(n6845), .A2(n6844), .A3(n6843), .ZN(P1_U3251) );
  AOI211_X1 U8432 ( .C1(n6848), .C2(n6847), .A(n9541), .B(n6846), .ZN(n6858)
         );
  AOI211_X1 U8433 ( .C1(n6851), .C2(n6850), .A(n9574), .B(n6849), .ZN(n6857)
         );
  INV_X1 U8434 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8435 ( .A1(n9577), .A2(n6852), .ZN(n6854) );
  NAND2_X1 U8436 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(n4437), .ZN(n6853) );
  OAI211_X1 U8437 ( .C1(n9585), .C2(n6855), .A(n6854), .B(n6853), .ZN(n6856)
         );
  OR3_X1 U8438 ( .A1(n6858), .A2(n6857), .A3(n6856), .ZN(P1_U3250) );
  AOI211_X1 U8439 ( .C1(n6861), .C2(n6860), .A(n9541), .B(n6859), .ZN(n6870)
         );
  AOI211_X1 U8440 ( .C1(n6864), .C2(n6863), .A(n9574), .B(n6862), .ZN(n6869)
         );
  INV_X1 U8441 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U8442 ( .A1(n9577), .A2(n6865), .ZN(n6867) );
  NAND2_X1 U8443 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6866) );
  OAI211_X1 U8444 ( .C1(n9585), .C2(n10126), .A(n6867), .B(n6866), .ZN(n6868)
         );
  OR3_X1 U8445 ( .A1(n6870), .A2(n6869), .A3(n6868), .ZN(P1_U3249) );
  INV_X1 U8446 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10114) );
  INV_X1 U8447 ( .A(n9730), .ZN(n8136) );
  OAI222_X1 U8448 ( .A1(n8480), .A2(n10114), .B1(n8483), .B2(n6871), .C1(
        P2_U3151), .C2(n8136), .ZN(P2_U3284) );
  INV_X1 U8449 ( .A(n9574), .ZN(n9560) );
  INV_X1 U8450 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6873) );
  MUX2_X1 U8451 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6873), .S(n6954), .Z(n6874)
         );
  NAND2_X1 U8452 ( .A1(n6875), .A2(n6874), .ZN(n6953) );
  OAI21_X1 U8453 ( .B1(n6875), .B2(n6874), .A(n6953), .ZN(n6886) );
  INV_X1 U8454 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6878) );
  MUX2_X1 U8455 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6878), .S(n6954), .Z(n6879)
         );
  NAND2_X1 U8456 ( .A1(n6880), .A2(n6879), .ZN(n6949) );
  OAI21_X1 U8457 ( .B1(n6880), .B2(n6879), .A(n6949), .ZN(n6881) );
  NAND2_X1 U8458 ( .A1(n6881), .A2(n9570), .ZN(n6883) );
  AND2_X1 U8459 ( .A1(n4437), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7724) );
  AOI21_X1 U8460 ( .B1(n9547), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7724), .ZN(
        n6882) );
  OAI211_X1 U8461 ( .C1(n9565), .C2(n6884), .A(n6883), .B(n6882), .ZN(n6885)
         );
  AOI21_X1 U8462 ( .B1(n9560), .B2(n6886), .A(n6885), .ZN(n6887) );
  INV_X1 U8463 ( .A(n6887), .ZN(P1_U3252) );
  INV_X1 U8464 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10250) );
  OAI222_X1 U8465 ( .A1(n8483), .A2(n6888), .B1(n8129), .B2(P2_U3151), .C1(
        n10250), .C2(n8480), .ZN(P2_U3283) );
  NOR2_X1 U8466 ( .A1(n9547), .A2(n8935), .ZN(P1_U3085) );
  INV_X1 U8467 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10204) );
  INV_X1 U8468 ( .A(n8985), .ZN(n7135) );
  OAI222_X1 U8469 ( .A1(n9466), .A2(n10204), .B1(n7778), .B2(n6888), .C1(n7135), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U8470 ( .A1(n8764), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8471 ( .A1(n8765), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8472 ( .A1(n6889), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6890) );
  NAND3_X1 U8473 ( .A1(n6892), .A2(n6891), .A3(n6890), .ZN(n9013) );
  NAND2_X1 U8474 ( .A1(n9013), .A2(P1_U3973), .ZN(n6893) );
  OAI21_X1 U8475 ( .B1(n8935), .B2(n5747), .A(n6893), .ZN(P1_U3585) );
  NAND2_X1 U8476 ( .A1(n7281), .A2(P1_U3973), .ZN(n6894) );
  OAI21_X1 U8477 ( .B1(n8935), .B2(n6895), .A(n6894), .ZN(P1_U3558) );
  INV_X1 U8478 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8479 ( .B1(n8331), .B2(n9914), .A(n6896), .ZN(n6898) );
  NOR2_X1 U8480 ( .A1(n5881), .A2(n9861), .ZN(n6988) );
  INV_X1 U8481 ( .A(n6988), .ZN(n6897) );
  OAI211_X1 U8482 ( .C1(n9909), .C2(n6992), .A(n6898), .B(n6897), .ZN(n8388)
         );
  NAND2_X1 U8483 ( .A1(n8388), .A2(n9915), .ZN(n6899) );
  OAI21_X1 U8484 ( .B1(n6900), .B2(n9915), .A(n6899), .ZN(P2_U3390) );
  XOR2_X1 U8485 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7158), .Z(n6915) );
  INV_X1 U8486 ( .A(n6902), .ZN(n6904) );
  OAI21_X1 U8487 ( .B1(n6905), .B2(n6904), .A(n6903), .ZN(n6907) );
  MUX2_X1 U8488 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8118), .Z(n7151) );
  XNOR2_X1 U8489 ( .A(n7151), .B(n7159), .ZN(n6906) );
  NAND2_X1 U8490 ( .A1(n6907), .A2(n6906), .ZN(n7152) );
  OAI211_X1 U8491 ( .C1(n6907), .C2(n6906), .A(n7152), .B(n6714), .ZN(n6914)
         );
  INV_X1 U8492 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U8493 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7196) );
  OAI21_X1 U8494 ( .B1(n6908), .B2(n10156), .A(n7196), .ZN(n6912) );
  XNOR2_X1 U8495 ( .A(n7160), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n6910) );
  NOR2_X1 U8496 ( .A1(n6910), .A2(n9845), .ZN(n6911) );
  AOI211_X1 U8497 ( .C1(n9832), .C2(n7159), .A(n6912), .B(n6911), .ZN(n6913)
         );
  OAI211_X1 U8498 ( .C1(n6915), .C2(n9699), .A(n6914), .B(n6913), .ZN(P2_U3187) );
  XNOR2_X1 U8499 ( .A(n6931), .B(n8079), .ZN(n6929) );
  NAND2_X1 U8500 ( .A1(n7504), .A2(n6992), .ZN(n6921) );
  NAND2_X1 U8501 ( .A1(n6979), .A2(n6921), .ZN(n6930) );
  XOR2_X1 U8502 ( .A(n6929), .B(n6930), .Z(n6928) );
  NAND2_X1 U8503 ( .A1(n6922), .A2(n6985), .ZN(n6923) );
  INV_X1 U8504 ( .A(n8045), .ZN(n8057) );
  AOI22_X1 U8505 ( .A1(n8042), .A2(n8078), .B1(n8057), .B2(n8080), .ZN(n6925)
         );
  OAI21_X1 U8506 ( .B1(n8065), .B2(n7300), .A(n6925), .ZN(n6926) );
  AOI21_X1 U8507 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6937), .A(n6926), .ZN(
        n6927) );
  OAI21_X1 U8508 ( .B1(n6928), .B2(n8050), .A(n6927), .ZN(P2_U3162) );
  NAND2_X1 U8509 ( .A1(n6930), .A2(n6929), .ZN(n6933) );
  NAND2_X1 U8510 ( .A1(n6931), .A2(n5881), .ZN(n6932) );
  NAND2_X1 U8511 ( .A1(n6933), .A2(n6932), .ZN(n6963) );
  XNOR2_X1 U8512 ( .A(n6964), .B(n8078), .ZN(n6962) );
  XOR2_X1 U8513 ( .A(n6963), .B(n6962), .Z(n6939) );
  AOI22_X1 U8514 ( .A1(n8057), .A2(n8079), .B1(n8042), .B2(n8077), .ZN(n6934)
         );
  OAI21_X1 U8515 ( .B1(n6935), .B2(n8065), .A(n6934), .ZN(n6936) );
  AOI21_X1 U8516 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6937), .A(n6936), .ZN(
        n6938) );
  OAI21_X1 U8517 ( .B1(n6939), .B2(n8050), .A(n6938), .ZN(P2_U3177) );
  INV_X1 U8518 ( .A(n9764), .ZN(n8140) );
  INV_X1 U8519 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6940) );
  OAI222_X1 U8520 ( .A1(n8483), .A2(n6977), .B1(n8140), .B2(P2_U3151), .C1(
        n6940), .C2(n8480), .ZN(P2_U3282) );
  XNOR2_X1 U8521 ( .A(n6942), .B(n6941), .ZN(n7042) );
  INV_X1 U8522 ( .A(n9012), .ZN(n8548) );
  NAND2_X1 U8523 ( .A1(n7022), .A2(n9012), .ZN(n7215) );
  INV_X1 U8524 ( .A(n7215), .ZN(n6943) );
  INV_X1 U8525 ( .A(n9489), .ZN(n8636) );
  AOI22_X1 U8526 ( .A1(n6943), .A2(n8636), .B1(n7083), .B2(n9497), .ZN(n6948)
         );
  AND3_X1 U8527 ( .A1(n6946), .A2(n6945), .A3(n7078), .ZN(n7067) );
  INV_X1 U8528 ( .A(n7067), .ZN(n6998) );
  NAND2_X1 U8529 ( .A1(n6998), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6947) );
  OAI211_X1 U8530 ( .C1(n7042), .C2(n9493), .A(n6948), .B(n6947), .ZN(P1_U3232) );
  XNOR2_X1 U8531 ( .A(n7012), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6951) );
  OAI21_X1 U8532 ( .B1(n6954), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6949), .ZN(
        n6950) );
  NOR2_X1 U8533 ( .A1(n6950), .A2(n6951), .ZN(n7006) );
  AOI211_X1 U8534 ( .C1(n6951), .C2(n6950), .A(n9541), .B(n7006), .ZN(n6961)
         );
  INV_X1 U8535 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6952) );
  MUX2_X1 U8536 ( .A(n6952), .B(P1_REG1_REG_10__SCAN_IN), .S(n7012), .Z(n6956)
         );
  OAI21_X1 U8537 ( .B1(n6954), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6953), .ZN(
        n6955) );
  NOR2_X1 U8538 ( .A1(n6955), .A2(n6956), .ZN(n7011) );
  AOI211_X1 U8539 ( .C1(n6956), .C2(n6955), .A(n9574), .B(n7011), .ZN(n6960)
         );
  INV_X1 U8540 ( .A(n7012), .ZN(n6958) );
  NAND2_X1 U8541 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U8542 ( .A1(n9547), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n6957) );
  OAI211_X1 U8543 ( .C1(n9565), .C2(n6958), .A(n9488), .B(n6957), .ZN(n6959)
         );
  OR3_X1 U8544 ( .A1(n6961), .A2(n6960), .A3(n6959), .ZN(P1_U3253) );
  NAND2_X1 U8545 ( .A1(n6964), .A2(n7073), .ZN(n6965) );
  XNOR2_X1 U8546 ( .A(n7960), .B(n6974), .ZN(n7091) );
  XNOR2_X1 U8547 ( .A(n7091), .B(n9862), .ZN(n6968) );
  AOI21_X1 U8548 ( .B1(n6967), .B2(n6968), .A(n8050), .ZN(n6970) );
  INV_X1 U8549 ( .A(n6968), .ZN(n6969) );
  NAND2_X1 U8550 ( .A1(n6970), .A2(n7094), .ZN(n6976) );
  NAND2_X1 U8551 ( .A1(n8042), .A2(n8076), .ZN(n6971) );
  NAND2_X1 U8552 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9680) );
  OAI211_X1 U8553 ( .C1(n7073), .C2(n8045), .A(n6971), .B(n9680), .ZN(n6973)
         );
  NOR2_X1 U8554 ( .A1(n7989), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6972) );
  AOI211_X1 U8555 ( .C1(n6974), .C2(n8047), .A(n6973), .B(n6972), .ZN(n6975)
         );
  NAND2_X1 U8556 ( .A1(n6976), .A2(n6975), .ZN(P2_U3158) );
  INV_X1 U8557 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6978) );
  INV_X1 U8558 ( .A(n9510), .ZN(n8982) );
  OAI222_X1 U8559 ( .A1(n9466), .A2(n6978), .B1(n7778), .B2(n6977), .C1(n8982), 
        .C2(n4437), .ZN(P1_U3342) );
  INV_X1 U8560 ( .A(n9914), .ZN(n9887) );
  XNOR2_X1 U8561 ( .A(n6980), .B(n6979), .ZN(n7005) );
  XNOR2_X1 U8562 ( .A(n5769), .B(n6981), .ZN(n6982) );
  AOI222_X1 U8563 ( .A1(n8331), .A2(n6982), .B1(n8078), .B2(n8326), .C1(n8080), 
        .C2(n8328), .ZN(n7001) );
  OAI21_X1 U8564 ( .B1(n9887), .B2(n7005), .A(n7001), .ZN(n7302) );
  OAI22_X1 U8565 ( .A1(n8413), .A2(n7300), .B1(n5266), .B2(n9915), .ZN(n6983)
         );
  AOI21_X1 U8566 ( .B1(n7302), .B2(n9915), .A(n6983), .ZN(n6984) );
  INV_X1 U8567 ( .A(n6984), .ZN(P2_U3393) );
  INV_X1 U8568 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10057) );
  NOR3_X1 U8569 ( .A1(n6986), .A2(n6985), .A3(n9907), .ZN(n6987) );
  AOI211_X1 U8570 ( .C1(n8303), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6988), .B(
        n6987), .ZN(n6989) );
  MUX2_X1 U8571 ( .A(n6990), .B(n6989), .S(n8318), .Z(n6991) );
  OAI21_X1 U8572 ( .B1(n8176), .B2(n6992), .A(n6991), .ZN(P2_U3233) );
  AOI21_X1 U8573 ( .B1(n6995), .B2(n6993), .A(n6994), .ZN(n7000) );
  INV_X2 U8574 ( .A(n8508), .ZN(n8595) );
  AOI22_X1 U8575 ( .A1(n9012), .A2(n6046), .B1(n8936), .B2(n8595), .ZN(n7029)
         );
  OAI22_X1 U8576 ( .A1(n7029), .A2(n9489), .B1(n8850), .B2(n8651), .ZN(n6997)
         );
  AOI21_X1 U8577 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6998), .A(n6997), .ZN(
        n6999) );
  OAI21_X1 U8578 ( .B1(n7000), .B2(n9493), .A(n6999), .ZN(P1_U3222) );
  MUX2_X1 U8579 ( .A(n10128), .B(n7001), .S(n8318), .Z(n7004) );
  AOI22_X1 U8580 ( .A1(n8304), .A2(n7002), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8303), .ZN(n7003) );
  OAI211_X1 U8581 ( .C1(n7005), .C2(n8339), .A(n7004), .B(n7003), .ZN(P2_U3232) );
  INV_X1 U8582 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7007) );
  MUX2_X1 U8583 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7007), .S(n7139), .Z(n7008)
         );
  INV_X1 U8584 ( .A(n7008), .ZN(n7009) );
  NOR2_X1 U8585 ( .A1(n7010), .A2(n7009), .ZN(n7138) );
  AOI211_X1 U8586 ( .C1(n7010), .C2(n7009), .A(n9541), .B(n7138), .ZN(n7020)
         );
  INV_X1 U8587 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7013) );
  MUX2_X1 U8588 ( .A(n7013), .B(P1_REG1_REG_11__SCAN_IN), .S(n7139), .Z(n7014)
         );
  NOR2_X1 U8589 ( .A1(n7015), .A2(n7014), .ZN(n7130) );
  AOI211_X1 U8590 ( .C1(n7015), .C2(n7014), .A(n9574), .B(n7130), .ZN(n7019)
         );
  INV_X1 U8591 ( .A(n7139), .ZN(n7017) );
  NAND2_X1 U8592 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7833) );
  NAND2_X1 U8593 ( .A1(n9547), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n7016) );
  OAI211_X1 U8594 ( .C1(n9565), .C2(n7017), .A(n7833), .B(n7016), .ZN(n7018)
         );
  OR3_X1 U8595 ( .A1(n7020), .A2(n7019), .A3(n7018), .ZN(P1_U3254) );
  INV_X1 U8596 ( .A(n7024), .ZN(n7217) );
  NAND2_X1 U8597 ( .A1(n8900), .A2(n6540), .ZN(n7021) );
  NAND3_X1 U8598 ( .A1(n7084), .A2(n7217), .A3(n7021), .ZN(n7626) );
  NAND2_X1 U8599 ( .A1(n7082), .A2(n7023), .ZN(n7108) );
  OAI21_X1 U8600 ( .B1(n8785), .B2(n7082), .A(n7108), .ZN(n7324) );
  NAND2_X1 U8601 ( .A1(n7024), .A2(n8808), .ZN(n9286) );
  NOR2_X1 U8602 ( .A1(n6996), .A2(n7083), .ZN(n7110) );
  AOI211_X1 U8603 ( .C1(n7083), .C2(n6996), .A(n9286), .B(n7110), .ZN(n7328)
         );
  INV_X1 U8604 ( .A(n7083), .ZN(n8851) );
  NOR2_X1 U8605 ( .A1(n8936), .A2(n8851), .ZN(n7025) );
  OAI21_X1 U8606 ( .B1(n7026), .B2(n7025), .A(n7115), .ZN(n7028) );
  OR2_X1 U8607 ( .A1(n6345), .A2(n8896), .ZN(n7027) );
  OR2_X1 U8608 ( .A1(n6522), .A2(n8808), .ZN(n8910) );
  NAND2_X1 U8609 ( .A1(n7028), .A2(n9278), .ZN(n7030) );
  NAND2_X1 U8610 ( .A1(n7030), .A2(n7029), .ZN(n7325) );
  AOI211_X1 U8611 ( .C1(n9650), .C2(n7324), .A(n7328), .B(n7325), .ZN(n7129)
         );
  INV_X1 U8612 ( .A(n7031), .ZN(n7033) );
  AND2_X1 U8613 ( .A1(n7033), .A2(n7032), .ZN(n7034) );
  OAI211_X1 U8614 ( .C1(n8852), .C2(n9652), .A(n7034), .B(n7078), .ZN(n7121)
         );
  OAI22_X1 U8615 ( .A1(n9367), .A2(n8850), .B1(n9667), .B2(n6796), .ZN(n7035)
         );
  INV_X1 U8616 ( .A(n7035), .ZN(n7036) );
  OAI21_X1 U8617 ( .B1(n7129), .B2(n9665), .A(n7036), .ZN(P1_U3523) );
  INV_X1 U8618 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7038) );
  INV_X1 U8619 ( .A(n7037), .ZN(n7039) );
  INV_X1 U8620 ( .A(n8987), .ZN(n9524) );
  OAI222_X1 U8621 ( .A1(n9466), .A2(n7038), .B1(n7778), .B2(n7039), .C1(n4437), 
        .C2(n9524), .ZN(P1_U3341) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7040) );
  OAI222_X1 U8623 ( .A1(n8480), .A2(n7040), .B1(n8483), .B2(n7039), .C1(
        P2_U3151), .C2(n8127), .ZN(P2_U3281) );
  MUX2_X1 U8624 ( .A(n8938), .B(n7042), .S(n7041), .Z(n7045) );
  OAI21_X1 U8625 ( .B1(n7043), .B2(P1_IR_REG_0__SCAN_IN), .A(P1_U3973), .ZN(
        n7044) );
  AOI21_X1 U8626 ( .B1(n7045), .B2(n9459), .A(n7044), .ZN(n8960) );
  OAI211_X1 U8627 ( .C1(n7048), .C2(n7047), .A(n9570), .B(n7046), .ZN(n7056)
         );
  AOI22_X1 U8628 ( .A1(n9547), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n4437), .ZN(n7055) );
  OAI211_X1 U8629 ( .C1(n7051), .C2(n7050), .A(n9560), .B(n7049), .ZN(n7054)
         );
  NAND2_X1 U8630 ( .A1(n9577), .A2(n7052), .ZN(n7053) );
  NAND4_X1 U8631 ( .A1(n7056), .A2(n7055), .A3(n7054), .A4(n7053), .ZN(n7057)
         );
  OR2_X1 U8632 ( .A1(n8960), .A2(n7057), .ZN(P1_U3245) );
  INV_X1 U8633 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7066) );
  INV_X1 U8634 ( .A(n7058), .ZN(n7062) );
  NOR3_X1 U8635 ( .A1(n6994), .A2(n7060), .A3(n7059), .ZN(n7061) );
  OAI21_X1 U8636 ( .B1(n7062), .B2(n7061), .A(n8634), .ZN(n7065) );
  AOI22_X1 U8637 ( .A1(n9012), .A2(n8934), .B1(n7022), .B2(n8595), .ZN(n7116)
         );
  INV_X1 U8638 ( .A(n7116), .ZN(n7063) );
  AOI22_X1 U8639 ( .A1(n7063), .A2(n8636), .B1(n7112), .B2(n9497), .ZN(n7064)
         );
  OAI211_X1 U8640 ( .C1(n7067), .C2(n7066), .A(n7065), .B(n7064), .ZN(P1_U3237) );
  OAI21_X1 U8641 ( .B1(n7069), .B2(n7071), .A(n7068), .ZN(n7224) );
  XNOR2_X1 U8642 ( .A(n7070), .B(n7071), .ZN(n7072) );
  OAI222_X1 U8643 ( .A1(n9860), .A2(n7073), .B1(n9861), .B2(n5889), .C1(n9867), 
        .C2(n7072), .ZN(n7221) );
  AOI21_X1 U8644 ( .B1(n9914), .B2(n7224), .A(n7221), .ZN(n7274) );
  INV_X1 U8645 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7074) );
  OAI22_X1 U8646 ( .A1(n8413), .A2(n7271), .B1(n7074), .B2(n9915), .ZN(n7075)
         );
  INV_X1 U8647 ( .A(n7075), .ZN(n7076) );
  OAI21_X1 U8648 ( .B1(n7274), .B2(n9917), .A(n7076), .ZN(P2_U3399) );
  NAND3_X1 U8649 ( .A1(n7079), .A2(n7078), .A3(n7077), .ZN(n7080) );
  NAND2_X1 U8650 ( .A1(n9272), .A2(n6345), .ZN(n9241) );
  NOR2_X1 U8651 ( .A1(n9241), .A2(n9286), .ZN(n9182) );
  OAI21_X1 U8652 ( .B1(n9182), .B2(n9587), .A(n7083), .ZN(n7089) );
  INV_X1 U8653 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7086) );
  OAI21_X1 U8654 ( .B1(n8936), .B2(n7083), .A(n7082), .ZN(n8780) );
  INV_X1 U8655 ( .A(n8780), .ZN(n7214) );
  NAND3_X1 U8656 ( .A1(n7214), .A2(n7084), .A3(n7217), .ZN(n7085) );
  OAI211_X1 U8657 ( .C1(n9236), .C2(n7086), .A(n7085), .B(n7215), .ZN(n7087)
         );
  NAND2_X1 U8658 ( .A1(n7087), .A2(n9272), .ZN(n7088) );
  OAI211_X1 U8659 ( .C1(n7090), .C2(n9272), .A(n7089), .B(n7088), .ZN(P1_U3293) );
  INV_X1 U8660 ( .A(n7091), .ZN(n7092) );
  NAND2_X1 U8661 ( .A1(n7092), .A2(n8077), .ZN(n7093) );
  XNOR2_X1 U8662 ( .A(n7960), .B(n7211), .ZN(n7193) );
  XNOR2_X1 U8663 ( .A(n7193), .B(n8076), .ZN(n7095) );
  OAI21_X1 U8664 ( .B1(n7096), .B2(n7095), .A(n7195), .ZN(n7105) );
  INV_X1 U8665 ( .A(n8050), .ZN(n8052) );
  INV_X1 U8666 ( .A(n7097), .ZN(n7098) );
  AOI21_X1 U8667 ( .B1(n8057), .B2(n8077), .A(n7098), .ZN(n7103) );
  INV_X1 U8668 ( .A(n7099), .ZN(n7210) );
  NAND2_X1 U8669 ( .A1(n8062), .A2(n7210), .ZN(n7102) );
  NAND2_X1 U8670 ( .A1(n8047), .A2(n7211), .ZN(n7101) );
  NAND2_X1 U8671 ( .A1(n8042), .A2(n8075), .ZN(n7100) );
  NAND4_X1 U8672 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7104)
         );
  AOI21_X1 U8673 ( .B1(n7105), .B2(n8052), .A(n7104), .ZN(n7106) );
  INV_X1 U8674 ( .A(n7106), .ZN(P2_U3170) );
  NAND2_X1 U8675 ( .A1(n7113), .A2(n8850), .ZN(n7107) );
  NAND2_X1 U8676 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  NAND2_X1 U8677 ( .A1(n7109), .A2(n8779), .ZN(n7182) );
  OAI21_X1 U8678 ( .B1(n7109), .B2(n8779), .A(n7182), .ZN(n7297) );
  INV_X1 U8679 ( .A(n7110), .ZN(n7111) );
  NAND2_X1 U8680 ( .A1(n7110), .A2(n7295), .ZN(n7185) );
  INV_X1 U8681 ( .A(n7185), .ZN(n7186) );
  AOI211_X1 U8682 ( .C1(n7112), .C2(n7111), .A(n9286), .B(n7186), .ZN(n7292)
         );
  NAND2_X1 U8683 ( .A1(n7113), .A2(n6996), .ZN(n7114) );
  XNOR2_X1 U8684 ( .A(n7172), .B(n8779), .ZN(n7117) );
  OAI21_X1 U8685 ( .B1(n7117), .B2(n9215), .A(n7116), .ZN(n7291) );
  AOI211_X1 U8686 ( .C1(n9650), .C2(n7297), .A(n7292), .B(n7291), .ZN(n7125)
         );
  OAI22_X1 U8687 ( .A1(n9367), .A2(n7295), .B1(n9667), .B2(n6795), .ZN(n7118)
         );
  INV_X1 U8688 ( .A(n7118), .ZN(n7119) );
  OAI21_X1 U8689 ( .B1(n7125), .B2(n9665), .A(n7119), .ZN(P1_U3524) );
  INV_X1 U8690 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7122) );
  OAI22_X1 U8691 ( .A1(n9444), .A2(n7295), .B1(n9439), .B2(n7122), .ZN(n7123)
         );
  INV_X1 U8692 ( .A(n7123), .ZN(n7124) );
  OAI21_X1 U8693 ( .B1(n7125), .B2(n9661), .A(n7124), .ZN(P1_U3459) );
  INV_X1 U8694 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7126) );
  OAI22_X1 U8695 ( .A1(n9444), .A2(n8850), .B1(n9439), .B2(n7126), .ZN(n7127)
         );
  INV_X1 U8696 ( .A(n7127), .ZN(n7128) );
  OAI21_X1 U8697 ( .B1(n7129), .B2(n9661), .A(n7128), .ZN(P1_U3456) );
  INV_X1 U8698 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7131) );
  MUX2_X1 U8699 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7131), .S(n8985), .Z(n7132)
         );
  NAND2_X1 U8700 ( .A1(n7133), .A2(n7132), .ZN(n8976) );
  OAI21_X1 U8701 ( .B1(n7133), .B2(n7132), .A(n8976), .ZN(n7137) );
  NAND2_X1 U8702 ( .A1(n9547), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U8703 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7856) );
  OAI211_X1 U8704 ( .C1(n9565), .C2(n7135), .A(n7134), .B(n7856), .ZN(n7136)
         );
  AOI21_X1 U8705 ( .B1(n7137), .B2(n9560), .A(n7136), .ZN(n7146) );
  INV_X1 U8706 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7140) );
  MUX2_X1 U8707 ( .A(n7140), .B(P1_REG2_REG_12__SCAN_IN), .S(n8985), .Z(n7141)
         );
  INV_X1 U8708 ( .A(n7141), .ZN(n7142) );
  NAND2_X1 U8709 ( .A1(n7143), .A2(n7142), .ZN(n8984) );
  OAI21_X1 U8710 ( .B1(n7143), .B2(n7142), .A(n8984), .ZN(n7144) );
  NAND2_X1 U8711 ( .A1(n7144), .A2(n9570), .ZN(n7145) );
  NAND2_X1 U8712 ( .A1(n7146), .A2(n7145), .ZN(P1_U3255) );
  INV_X1 U8713 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7148) );
  INV_X1 U8714 ( .A(n7147), .ZN(n7149) );
  OAI222_X1 U8715 ( .A1(n9466), .A2(n7148), .B1(n7778), .B2(n7149), .C1(
        P1_U3086), .C2(n8989), .ZN(P1_U3340) );
  INV_X1 U8716 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7150) );
  OAI222_X1 U8717 ( .A1(n8480), .A2(n7150), .B1(n8483), .B2(n7149), .C1(
        P2_U3151), .C2(n4701), .ZN(P2_U3280) );
  MUX2_X1 U8718 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8118), .Z(n7227) );
  XOR2_X1 U8719 ( .A(n7233), .B(n7227), .Z(n7228) );
  MUX2_X1 U8720 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8118), .Z(n7154) );
  INV_X1 U8721 ( .A(n7154), .ZN(n7155) );
  INV_X1 U8722 ( .A(n7151), .ZN(n7153) );
  OAI21_X1 U8723 ( .B1(n7159), .B2(n7153), .A(n7152), .ZN(n9706) );
  XOR2_X1 U8724 ( .A(n7161), .B(n7154), .Z(n9707) );
  NOR2_X1 U8725 ( .A1(n9706), .A2(n9707), .ZN(n9705) );
  AOI21_X1 U8726 ( .B1(n7161), .B2(n7155), .A(n9705), .ZN(n7229) );
  XOR2_X1 U8727 ( .A(n7228), .B(n7229), .Z(n7170) );
  INV_X1 U8728 ( .A(n6714), .ZN(n9708) );
  INV_X1 U8729 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9922) );
  INV_X1 U8730 ( .A(n7156), .ZN(n7157) );
  AOI22_X1 U8731 ( .A1(n7158), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n4697), .B2(
        n7157), .ZN(n9698) );
  MUX2_X1 U8732 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9922), .S(n7161), .Z(n9697)
         );
  XOR2_X1 U8733 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7235), .Z(n7168) );
  MUX2_X1 U8734 ( .A(n7407), .B(P2_REG2_REG_6__SCAN_IN), .S(n7161), .Z(n9694)
         );
  NAND2_X1 U8735 ( .A1(n9693), .A2(n9694), .ZN(n9692) );
  OAI21_X1 U8736 ( .B1(n7161), .B2(n7407), .A(n9692), .ZN(n7162) );
  NAND2_X1 U8737 ( .A1(n7162), .A2(n7226), .ZN(n7240) );
  AOI21_X1 U8738 ( .B1(n5396), .B2(n7163), .A(n7243), .ZN(n7166) );
  INV_X1 U8739 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U8740 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10031), .ZN(n7375) );
  NOR2_X1 U8741 ( .A1(n9696), .A2(n7226), .ZN(n7164) );
  AOI211_X1 U8742 ( .C1(n9830), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7375), .B(
        n7164), .ZN(n7165) );
  OAI21_X1 U8743 ( .B1(n7166), .B2(n9845), .A(n7165), .ZN(n7167) );
  AOI21_X1 U8744 ( .B1(n7168), .B2(n9839), .A(n7167), .ZN(n7169) );
  OAI21_X1 U8745 ( .B1(n7170), .B2(n9708), .A(n7169), .ZN(P2_U3189) );
  INV_X1 U8746 ( .A(n8934), .ZN(n7278) );
  NAND2_X1 U8747 ( .A1(n7278), .A2(n8518), .ZN(n7275) );
  INV_X1 U8748 ( .A(n8518), .ZN(n9640) );
  NAND2_X1 U8749 ( .A1(n8934), .A2(n9640), .ZN(n8855) );
  NAND2_X1 U8750 ( .A1(n7173), .A2(n8778), .ZN(n7174) );
  NAND2_X1 U8751 ( .A1(n7276), .A2(n7174), .ZN(n7175) );
  NAND2_X1 U8752 ( .A1(n7175), .A2(n9278), .ZN(n7179) );
  NAND2_X1 U8753 ( .A1(n6046), .A2(n8595), .ZN(n7177) );
  NAND2_X1 U8754 ( .A1(n7281), .A2(n9012), .ZN(n7176) );
  NAND2_X1 U8755 ( .A1(n7177), .A2(n7176), .ZN(n8519) );
  INV_X1 U8756 ( .A(n8519), .ZN(n7178) );
  NAND2_X1 U8757 ( .A1(n7179), .A2(n7178), .ZN(n9641) );
  INV_X1 U8758 ( .A(n9641), .ZN(n7192) );
  NAND2_X1 U8759 ( .A1(n7180), .A2(n7295), .ZN(n7181) );
  NAND2_X1 U8760 ( .A1(n7182), .A2(n7181), .ZN(n7183) );
  NAND2_X1 U8761 ( .A1(n7183), .A2(n8778), .ZN(n7280) );
  OAI21_X1 U8762 ( .B1(n7183), .B2(n8778), .A(n7280), .ZN(n9643) );
  AND2_X1 U8763 ( .A1(n7626), .A2(n7632), .ZN(n7184) );
  OR2_X1 U8764 ( .A1(n7185), .A2(n8518), .ZN(n7353) );
  OAI211_X1 U8765 ( .C1(n7186), .C2(n9640), .A(n9333), .B(n7353), .ZN(n9639)
         );
  AOI22_X1 U8766 ( .A1(n9609), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9598), .B2(
        n7187), .ZN(n7189) );
  NAND2_X1 U8767 ( .A1(n9587), .A2(n8518), .ZN(n7188) );
  OAI211_X1 U8768 ( .C1(n9639), .C2(n9241), .A(n7189), .B(n7188), .ZN(n7190)
         );
  AOI21_X1 U8769 ( .B1(n9643), .B2(n9606), .A(n7190), .ZN(n7191) );
  OAI21_X1 U8770 ( .B1(n7192), .B2(n9609), .A(n7191), .ZN(P1_U3290) );
  NAND2_X1 U8771 ( .A1(n7193), .A2(n5889), .ZN(n7194) );
  XNOR2_X1 U8772 ( .A(n7312), .B(n7960), .ZN(n7259) );
  XNOR2_X1 U8773 ( .A(n7259), .B(n8075), .ZN(n7260) );
  XOR2_X1 U8774 ( .A(n7261), .B(n7260), .Z(n7201) );
  NAND2_X1 U8775 ( .A1(n8057), .A2(n8076), .ZN(n7197) );
  OAI211_X1 U8776 ( .C1(n7463), .C2(n8059), .A(n7197), .B(n7196), .ZN(n7199)
         );
  NOR2_X1 U8777 ( .A1(n7989), .A2(n7310), .ZN(n7198) );
  AOI211_X1 U8778 ( .C1(n7312), .C2(n8047), .A(n7199), .B(n7198), .ZN(n7200)
         );
  OAI21_X1 U8779 ( .B1(n7201), .B2(n8050), .A(n7200), .ZN(P2_U3167) );
  INV_X1 U8780 ( .A(n7202), .ZN(n7220) );
  AOI22_X1 U8781 ( .A1(n9550), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9462), .ZN(n7203) );
  OAI21_X1 U8782 ( .B1(n7220), .B2(n7778), .A(n7203), .ZN(P1_U3339) );
  XNOR2_X1 U8783 ( .A(n7205), .B(n7204), .ZN(n9877) );
  XNOR2_X1 U8784 ( .A(n7207), .B(n7206), .ZN(n7208) );
  AOI222_X1 U8785 ( .A1(n8331), .A2(n7208), .B1(n8077), .B2(n8328), .C1(n8075), 
        .C2(n8326), .ZN(n9878) );
  MUX2_X1 U8786 ( .A(n7209), .B(n9878), .S(n8318), .Z(n7213) );
  AOI22_X1 U8787 ( .A1(n8304), .A2(n7211), .B1(n8303), .B2(n7210), .ZN(n7212)
         );
  OAI211_X1 U8788 ( .C1(n8339), .C2(n9877), .A(n7213), .B(n7212), .ZN(P2_U3229) );
  INV_X1 U8789 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7219) );
  OAI21_X1 U8790 ( .B1(n9278), .B2(n9650), .A(n7214), .ZN(n7216) );
  OAI211_X1 U8791 ( .C1(n7217), .C2(n8851), .A(n7216), .B(n7215), .ZN(n9386)
         );
  NAND2_X1 U8792 ( .A1(n9386), .A2(n9439), .ZN(n7218) );
  OAI21_X1 U8793 ( .B1(n9439), .B2(n7219), .A(n7218), .ZN(P1_U3453) );
  OAI222_X1 U8794 ( .A1(n8483), .A2(n7220), .B1(n8126), .B2(P2_U3151), .C1(
        n10282), .C2(n8480), .ZN(P2_U3279) );
  OAI22_X1 U8795 ( .A1(n8176), .A2(n7271), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9857), .ZN(n7223) );
  MUX2_X1 U8796 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7221), .S(n8318), .Z(n7222)
         );
  AOI211_X1 U8797 ( .C1(n8260), .C2(n7224), .A(n7223), .B(n7222), .ZN(n7225)
         );
  INV_X1 U8798 ( .A(n7225), .ZN(P2_U3230) );
  MUX2_X1 U8799 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8118), .Z(n7333) );
  XNOR2_X1 U8800 ( .A(n7333), .B(n7338), .ZN(n7335) );
  OAI22_X1 U8801 ( .A1(n7229), .A2(n7228), .B1(n7227), .B2(n7226), .ZN(n7336)
         );
  XOR2_X1 U8802 ( .A(n7335), .B(n7336), .Z(n7249) );
  MUX2_X1 U8803 ( .A(n7230), .B(P2_REG1_REG_8__SCAN_IN), .S(n7338), .Z(n7237)
         );
  INV_X1 U8804 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7234) );
  INV_X1 U8805 ( .A(n7231), .ZN(n7232) );
  NAND2_X1 U8806 ( .A1(n7236), .A2(n7237), .ZN(n7332) );
  OAI21_X1 U8807 ( .B1(n7237), .B2(n7236), .A(n7332), .ZN(n7247) );
  NAND2_X1 U8808 ( .A1(n9830), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U8809 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7475) );
  OAI211_X1 U8810 ( .C1(n9696), .C2(n7239), .A(n7238), .B(n7475), .ZN(n7246)
         );
  INV_X1 U8811 ( .A(n7240), .ZN(n7241) );
  MUX2_X1 U8812 ( .A(n7604), .B(P2_REG2_REG_8__SCAN_IN), .S(n7338), .Z(n7242)
         );
  OR3_X1 U8813 ( .A1(n7243), .A2(n7242), .A3(n7241), .ZN(n7244) );
  AOI21_X1 U8814 ( .B1(n7337), .B2(n7244), .A(n9845), .ZN(n7245) );
  AOI211_X1 U8815 ( .C1(n7247), .C2(n9839), .A(n7246), .B(n7245), .ZN(n7248)
         );
  OAI21_X1 U8816 ( .B1(n7249), .B2(n9708), .A(n7248), .ZN(P2_U3190) );
  INV_X1 U8817 ( .A(n9599), .ZN(n7257) );
  AND2_X1 U8818 ( .A1(n8514), .A2(n7250), .ZN(n7253) );
  OAI211_X1 U8819 ( .C1(n7253), .C2(n7252), .A(n8634), .B(n7251), .ZN(n7256)
         );
  OAI22_X1 U8820 ( .A1(n8671), .A2(n8548), .B1(n7278), .B2(n8508), .ZN(n7355)
         );
  INV_X1 U8821 ( .A(n7358), .ZN(n9603) );
  NAND2_X1 U8822 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(n4437), .ZN(n8962) );
  OAI21_X1 U8823 ( .B1(n8651), .B2(n9603), .A(n8962), .ZN(n7254) );
  AOI21_X1 U8824 ( .B1(n7355), .B2(n8636), .A(n7254), .ZN(n7255) );
  OAI211_X1 U8825 ( .C1(n9501), .C2(n7257), .A(n7256), .B(n7255), .ZN(P1_U3230) );
  INV_X1 U8826 ( .A(n9892), .ZN(n7269) );
  XNOR2_X1 U8827 ( .A(n9892), .B(n7960), .ZN(n7365) );
  XNOR2_X1 U8828 ( .A(n7365), .B(n4764), .ZN(n7262) );
  OAI211_X1 U8829 ( .C1(n7263), .C2(n7262), .A(n7368), .B(n8052), .ZN(n7268)
         );
  INV_X1 U8830 ( .A(n7264), .ZN(n7408) );
  NAND2_X1 U8831 ( .A1(n8057), .A2(n8075), .ZN(n7265) );
  NAND2_X1 U8832 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9695) );
  OAI211_X1 U8833 ( .C1(n7598), .C2(n8059), .A(n7265), .B(n9695), .ZN(n7266)
         );
  AOI21_X1 U8834 ( .B1(n7408), .B2(n8062), .A(n7266), .ZN(n7267) );
  OAI211_X1 U8835 ( .C1(n7269), .C2(n8065), .A(n7268), .B(n7267), .ZN(P2_U3179) );
  INV_X1 U8836 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7270) );
  OAI22_X1 U8837 ( .A1(n8352), .A2(n7271), .B1(n8378), .B2(n7270), .ZN(n7272)
         );
  INV_X1 U8838 ( .A(n7272), .ZN(n7273) );
  OAI21_X1 U8839 ( .B1(n7274), .B2(n9927), .A(n7273), .ZN(P2_U3462) );
  NAND2_X1 U8840 ( .A1(n7281), .A2(n9603), .ZN(n8857) );
  NAND2_X1 U8841 ( .A1(n7354), .A2(n8857), .ZN(n8662) );
  INV_X1 U8842 ( .A(n7281), .ZN(n7282) );
  NAND2_X1 U8843 ( .A1(n7282), .A2(n7358), .ZN(n8664) );
  NAND2_X1 U8844 ( .A1(n8662), .A2(n8664), .ZN(n8667) );
  NAND2_X1 U8845 ( .A1(n8671), .A2(n8670), .ZN(n8663) );
  NAND2_X1 U8846 ( .A1(n8933), .A2(n8668), .ZN(n8856) );
  NAND2_X1 U8847 ( .A1(n8663), .A2(n8856), .ZN(n8783) );
  XNOR2_X1 U8848 ( .A(n8667), .B(n8783), .ZN(n7277) );
  AOI22_X1 U8849 ( .A1(n9012), .A2(n8932), .B1(n7281), .B2(n8595), .ZN(n7428)
         );
  OAI21_X1 U8850 ( .B1(n7277), .B2(n9215), .A(n7428), .ZN(n7316) );
  INV_X1 U8851 ( .A(n7316), .ZN(n7290) );
  NAND2_X1 U8852 ( .A1(n7278), .A2(n9640), .ZN(n7279) );
  NAND2_X1 U8853 ( .A1(n7280), .A2(n7279), .ZN(n7351) );
  XNOR2_X1 U8854 ( .A(n7281), .B(n9603), .ZN(n8784) );
  NAND2_X1 U8855 ( .A1(n7351), .A2(n8784), .ZN(n7350) );
  NAND2_X1 U8856 ( .A1(n7282), .A2(n9603), .ZN(n7283) );
  NAND2_X1 U8857 ( .A1(n7350), .A2(n7283), .ZN(n7284) );
  NAND2_X1 U8858 ( .A1(n7284), .A2(n8783), .ZN(n7436) );
  OAI21_X1 U8859 ( .B1(n7284), .B2(n8783), .A(n7436), .ZN(n7321) );
  OAI21_X1 U8860 ( .B1(n7352), .B2(n8668), .A(n9333), .ZN(n7285) );
  AND2_X1 U8861 ( .A1(n7352), .A2(n8668), .ZN(n7443) );
  NOR2_X1 U8862 ( .A1(n7285), .A2(n7443), .ZN(n7315) );
  NAND2_X1 U8863 ( .A1(n7315), .A2(n9596), .ZN(n7287) );
  AOI22_X1 U8864 ( .A1(n9609), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7430), .B2(
        n9598), .ZN(n7286) );
  OAI211_X1 U8865 ( .C1(n8668), .C2(n9602), .A(n7287), .B(n7286), .ZN(n7288)
         );
  AOI21_X1 U8866 ( .B1(n7321), .B2(n9606), .A(n7288), .ZN(n7289) );
  OAI21_X1 U8867 ( .B1(n7290), .B2(n9609), .A(n7289), .ZN(P1_U3288) );
  INV_X1 U8868 ( .A(n7291), .ZN(n7299) );
  NAND2_X1 U8869 ( .A1(n7292), .A2(n9596), .ZN(n7294) );
  AOI22_X1 U8870 ( .A1(n9609), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9598), .ZN(n7293) );
  OAI211_X1 U8871 ( .C1(n7295), .C2(n9602), .A(n7294), .B(n7293), .ZN(n7296)
         );
  AOI21_X1 U8872 ( .B1(n9606), .B2(n7297), .A(n7296), .ZN(n7298) );
  OAI21_X1 U8873 ( .B1(n9609), .B2(n7299), .A(n7298), .ZN(P1_U3291) );
  OAI22_X1 U8874 ( .A1(n8352), .A2(n7300), .B1(n8378), .B2(n6705), .ZN(n7301)
         );
  AOI21_X1 U8875 ( .B1(n7302), .B2(n8378), .A(n7301), .ZN(n7303) );
  INV_X1 U8876 ( .A(n7303), .ZN(P2_U3460) );
  XNOR2_X1 U8877 ( .A(n7304), .B(n7306), .ZN(n9884) );
  NAND2_X1 U8878 ( .A1(n8318), .A2(n9869), .ZN(n7881) );
  XNOR2_X1 U8879 ( .A(n7305), .B(n7306), .ZN(n7308) );
  OAI22_X1 U8880 ( .A1(n5889), .A2(n9860), .B1(n7463), .B2(n9861), .ZN(n7307)
         );
  AOI21_X1 U8881 ( .B1(n7308), .B2(n8331), .A(n7307), .ZN(n7309) );
  OAI21_X1 U8882 ( .B1(n9884), .B2(n7615), .A(n7309), .ZN(n9886) );
  NAND2_X1 U8883 ( .A1(n9886), .A2(n8318), .ZN(n7314) );
  OAI22_X1 U8884 ( .A1(n8318), .A2(n5348), .B1(n7310), .B2(n9857), .ZN(n7311)
         );
  AOI21_X1 U8885 ( .B1(n8304), .B2(n7312), .A(n7311), .ZN(n7313) );
  OAI211_X1 U8886 ( .C1(n9884), .C2(n7881), .A(n7314), .B(n7313), .ZN(P2_U3228) );
  NOR2_X1 U8887 ( .A1(n7316), .A2(n7315), .ZN(n7323) );
  INV_X1 U8888 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7317) );
  OAI22_X1 U8889 ( .A1(n9444), .A2(n8668), .B1(n9439), .B2(n7317), .ZN(n7318)
         );
  AOI21_X1 U8890 ( .B1(n7321), .B2(n9437), .A(n7318), .ZN(n7319) );
  OAI21_X1 U8891 ( .B1(n7323), .B2(n9661), .A(n7319), .ZN(P1_U3468) );
  INV_X1 U8892 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10139) );
  OAI22_X1 U8893 ( .A1(n9367), .A2(n8668), .B1(n9667), .B2(n10139), .ZN(n7320)
         );
  AOI21_X1 U8894 ( .B1(n7321), .B2(n9361), .A(n7320), .ZN(n7322) );
  OAI21_X1 U8895 ( .B1(n7323), .B2(n9665), .A(n7322), .ZN(P1_U3527) );
  INV_X1 U8896 ( .A(n7324), .ZN(n7331) );
  NAND2_X1 U8897 ( .A1(n7325), .A2(n9272), .ZN(n7330) );
  AOI22_X1 U8898 ( .A1(n9609), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9598), .ZN(n7326) );
  OAI21_X1 U8899 ( .B1(n9602), .B2(n8850), .A(n7326), .ZN(n7327) );
  AOI21_X1 U8900 ( .B1(n9596), .B2(n7328), .A(n7327), .ZN(n7329) );
  OAI211_X1 U8901 ( .C1(n7331), .C2(n9294), .A(n7330), .B(n7329), .ZN(P1_U3292) );
  OAI21_X1 U8902 ( .B1(n7338), .B2(n7230), .A(n7332), .ZN(n8131) );
  XOR2_X1 U8903 ( .A(n8133), .B(n8131), .Z(n8135) );
  XNOR2_X1 U8904 ( .A(n8135), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7345) );
  INV_X1 U8905 ( .A(n7333), .ZN(n7334) );
  AOI22_X1 U8906 ( .A1(n7336), .A2(n7335), .B1(n7338), .B2(n7334), .ZN(n8108)
         );
  MUX2_X1 U8907 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8118), .Z(n8106) );
  XOR2_X1 U8908 ( .A(n8133), .B(n8106), .Z(n8107) );
  XNOR2_X1 U8909 ( .A(n8108), .B(n8107), .ZN(n7343) );
  XNOR2_X1 U8910 ( .A(n8081), .B(n8133), .ZN(n8082) );
  INV_X1 U8911 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7617) );
  XNOR2_X1 U8912 ( .A(n8082), .B(n7617), .ZN(n7339) );
  NOR2_X1 U8913 ( .A1(n7339), .A2(n9845), .ZN(n7342) );
  NAND2_X1 U8914 ( .A1(n9830), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U8915 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7507) );
  OAI211_X1 U8916 ( .C1(n9696), .C2(n8105), .A(n7340), .B(n7507), .ZN(n7341)
         );
  AOI211_X1 U8917 ( .C1(n7343), .C2(n6714), .A(n7342), .B(n7341), .ZN(n7344)
         );
  OAI21_X1 U8918 ( .B1(n7345), .B2(n9699), .A(n7344), .ZN(P2_U3191) );
  INV_X1 U8919 ( .A(n7346), .ZN(n7348) );
  INV_X1 U8920 ( .A(n8993), .ZN(n9564) );
  OAI222_X1 U8921 ( .A1(n9466), .A2(n7347), .B1(n7778), .B2(n7348), .C1(n4437), 
        .C2(n9564), .ZN(P1_U3338) );
  INV_X1 U8922 ( .A(n9831), .ZN(n8146) );
  OAI222_X1 U8923 ( .A1(n8480), .A2(n7349), .B1(n8483), .B2(n7348), .C1(
        P2_U3151), .C2(n8146), .ZN(P2_U3278) );
  OAI21_X1 U8924 ( .B1(n7351), .B2(n8784), .A(n7350), .ZN(n9605) );
  AOI211_X1 U8925 ( .C1(n7358), .C2(n7353), .A(n9286), .B(n7352), .ZN(n9597)
         );
  XOR2_X1 U8926 ( .A(n8784), .B(n7354), .Z(n7356) );
  AOI21_X1 U8927 ( .B1(n7356), .B2(n9278), .A(n7355), .ZN(n9608) );
  INV_X1 U8928 ( .A(n9608), .ZN(n7357) );
  AOI211_X1 U8929 ( .C1(n9650), .C2(n9605), .A(n9597), .B(n7357), .ZN(n7363)
         );
  AOI22_X1 U8930 ( .A1(n9354), .A2(n7358), .B1(n9665), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7359) );
  OAI21_X1 U8931 ( .B1(n7363), .B2(n9665), .A(n7359), .ZN(P1_U3526) );
  INV_X1 U8932 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7360) );
  OAI22_X1 U8933 ( .A1(n9444), .A2(n9603), .B1(n9439), .B2(n7360), .ZN(n7361)
         );
  INV_X1 U8934 ( .A(n7361), .ZN(n7362) );
  OAI21_X1 U8935 ( .B1(n7363), .B2(n9661), .A(n7362), .ZN(P1_U3465) );
  NAND2_X1 U8936 ( .A1(n9475), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7364) );
  OAI21_X1 U8937 ( .B1(n7961), .B2(n9475), .A(n7364), .ZN(P2_U3520) );
  XNOR2_X1 U8938 ( .A(n9896), .B(n7917), .ZN(n7472) );
  XNOR2_X1 U8939 ( .A(n7472), .B(n7598), .ZN(n7373) );
  INV_X1 U8940 ( .A(n7365), .ZN(n7366) );
  NAND2_X1 U8941 ( .A1(n7366), .A2(n4764), .ZN(n7367) );
  NAND2_X1 U8942 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  INV_X1 U8943 ( .A(n7369), .ZN(n7371) );
  NAND2_X1 U8944 ( .A1(n7371), .A2(n7370), .ZN(n7474) );
  INV_X1 U8945 ( .A(n7474), .ZN(n7372) );
  AOI21_X1 U8946 ( .B1(n7373), .B2(n7369), .A(n7372), .ZN(n7379) );
  NOR2_X1 U8947 ( .A1(n8045), .A2(n7463), .ZN(n7374) );
  AOI211_X1 U8948 ( .C1(n8042), .C2(n4657), .A(n7375), .B(n7374), .ZN(n7376)
         );
  OAI21_X1 U8949 ( .B1(n7468), .B2(n7989), .A(n7376), .ZN(n7377) );
  AOI21_X1 U8950 ( .B1(n9896), .B2(n8047), .A(n7377), .ZN(n7378) );
  OAI21_X1 U8951 ( .B1(n7379), .B2(n8050), .A(n7378), .ZN(P2_U3153) );
  INV_X1 U8952 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9936) );
  NOR2_X1 U8953 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7380) );
  AOI21_X1 U8954 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7380), .ZN(n9941) );
  NOR2_X1 U8955 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7381) );
  AOI21_X1 U8956 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7381), .ZN(n9944) );
  NOR2_X1 U8957 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7382) );
  AOI21_X1 U8958 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7382), .ZN(n9947) );
  NOR2_X1 U8959 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7383) );
  AOI21_X1 U8960 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7383), .ZN(n9950) );
  NOR2_X1 U8961 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7384) );
  AOI21_X1 U8962 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7384), .ZN(n9953) );
  NOR2_X1 U8963 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7385) );
  AOI21_X1 U8964 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7385), .ZN(n9956) );
  NOR2_X1 U8965 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7386) );
  AOI21_X1 U8966 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7386), .ZN(n9959) );
  NOR2_X1 U8967 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7387) );
  AOI21_X1 U8968 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7387), .ZN(n9962) );
  NOR2_X1 U8969 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7388) );
  AOI21_X1 U8970 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7388), .ZN(n10293) );
  NOR2_X1 U8971 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7389) );
  AOI21_X1 U8972 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7389), .ZN(n10299) );
  NOR2_X1 U8973 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7390) );
  AOI21_X1 U8974 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7390), .ZN(n10296) );
  NOR2_X1 U8975 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7391) );
  AOI21_X1 U8976 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7391), .ZN(n10287) );
  NOR2_X1 U8977 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7392) );
  AOI21_X1 U8978 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7392), .ZN(n10290) );
  AND2_X1 U8979 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7393) );
  NOR2_X1 U8980 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7393), .ZN(n9931) );
  INV_X1 U8981 ( .A(n9931), .ZN(n9932) );
  NAND3_X1 U8982 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U8983 ( .A1(n9934), .A2(n9933), .ZN(n9930) );
  NAND2_X1 U8984 ( .A1(n9932), .A2(n9930), .ZN(n10302) );
  NAND2_X1 U8985 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7394) );
  OAI21_X1 U8986 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7394), .ZN(n10301) );
  NOR2_X1 U8987 ( .A1(n10302), .A2(n10301), .ZN(n10300) );
  AOI21_X1 U8988 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10300), .ZN(n10305) );
  NAND2_X1 U8989 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7395) );
  OAI21_X1 U8990 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7395), .ZN(n10304) );
  NOR2_X1 U8991 ( .A1(n10305), .A2(n10304), .ZN(n10303) );
  AOI21_X1 U8992 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10303), .ZN(n10308) );
  NOR2_X1 U8993 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7396) );
  AOI21_X1 U8994 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7396), .ZN(n10307) );
  NAND2_X1 U8995 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  OAI21_X1 U8996 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10306), .ZN(n10289) );
  NAND2_X1 U8997 ( .A1(n10290), .A2(n10289), .ZN(n10288) );
  OAI21_X1 U8998 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10288), .ZN(n10286) );
  NAND2_X1 U8999 ( .A1(n10287), .A2(n10286), .ZN(n10285) );
  OAI21_X1 U9000 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10285), .ZN(n10295) );
  NAND2_X1 U9001 ( .A1(n10296), .A2(n10295), .ZN(n10294) );
  OAI21_X1 U9002 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10294), .ZN(n10298) );
  NAND2_X1 U9003 ( .A1(n10299), .A2(n10298), .ZN(n10297) );
  OAI21_X1 U9004 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10297), .ZN(n10292) );
  NAND2_X1 U9005 ( .A1(n10293), .A2(n10292), .ZN(n10291) );
  OAI21_X1 U9006 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10291), .ZN(n9961) );
  NAND2_X1 U9007 ( .A1(n9962), .A2(n9961), .ZN(n9960) );
  OAI21_X1 U9008 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9960), .ZN(n9958) );
  NAND2_X1 U9009 ( .A1(n9959), .A2(n9958), .ZN(n9957) );
  OAI21_X1 U9010 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9957), .ZN(n9955) );
  NAND2_X1 U9011 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  OAI21_X1 U9012 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9954), .ZN(n9952) );
  NAND2_X1 U9013 ( .A1(n9953), .A2(n9952), .ZN(n9951) );
  OAI21_X1 U9014 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9951), .ZN(n9949) );
  NAND2_X1 U9015 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  OAI21_X1 U9016 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9948), .ZN(n9946) );
  NAND2_X1 U9017 ( .A1(n9947), .A2(n9946), .ZN(n9945) );
  OAI21_X1 U9018 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9945), .ZN(n9943) );
  NAND2_X1 U9019 ( .A1(n9944), .A2(n9943), .ZN(n9942) );
  OAI21_X1 U9020 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9942), .ZN(n9940) );
  NAND2_X1 U9021 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  OAI21_X1 U9022 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9939), .ZN(n9937) );
  NOR2_X1 U9023 ( .A1(n9936), .A2(n9937), .ZN(n7397) );
  NAND2_X1 U9024 ( .A1(n9936), .A2(n9937), .ZN(n9935) );
  OAI21_X1 U9025 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7397), .A(n9935), .ZN(
        n7399) );
  XNOR2_X1 U9026 ( .A(n9007), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7398) );
  XNOR2_X1 U9027 ( .A(n7399), .B(n7398), .ZN(ADD_1068_U4) );
  INV_X1 U9028 ( .A(n7400), .ZN(n7402) );
  AOI22_X1 U9029 ( .A1(n9578), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9462), .ZN(n7401) );
  OAI21_X1 U9030 ( .B1(n7402), .B2(n7778), .A(n7401), .ZN(P1_U3337) );
  INV_X1 U9031 ( .A(n9477), .ZN(n9479) );
  OAI222_X1 U9032 ( .A1(n8483), .A2(n7402), .B1(n9479), .B2(P2_U3151), .C1(
        n10138), .C2(n8480), .ZN(P2_U3277) );
  XOR2_X1 U9033 ( .A(n7403), .B(n7405), .Z(n9888) );
  XNOR2_X1 U9034 ( .A(n7404), .B(n7405), .ZN(n7406) );
  AOI222_X1 U9035 ( .A1(n8331), .A2(n7406), .B1(n8074), .B2(n8326), .C1(n8075), 
        .C2(n8328), .ZN(n9889) );
  MUX2_X1 U9036 ( .A(n7407), .B(n9889), .S(n8318), .Z(n7410) );
  AOI22_X1 U9037 ( .A1(n9892), .A2(n8304), .B1(n8303), .B2(n7408), .ZN(n7409)
         );
  OAI211_X1 U9038 ( .C1(n8339), .C2(n9888), .A(n7410), .B(n7409), .ZN(P2_U3227) );
  XNOR2_X1 U9039 ( .A(n7412), .B(n7411), .ZN(n7413) );
  XNOR2_X1 U9040 ( .A(n7414), .B(n7413), .ZN(n7421) );
  NAND2_X1 U9041 ( .A1(n8932), .A2(n8595), .ZN(n7416) );
  NAND2_X1 U9042 ( .A1(n8930), .A2(n9012), .ZN(n7415) );
  NAND2_X1 U9043 ( .A1(n7416), .A2(n7415), .ZN(n7555) );
  AOI22_X1 U9044 ( .A1(n7555), .A2(n8636), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7418) );
  NAND2_X1 U9045 ( .A1(n9588), .A2(n9497), .ZN(n7417) );
  OAI211_X1 U9046 ( .C1(n9501), .C2(n7419), .A(n7418), .B(n7417), .ZN(n7420)
         );
  AOI21_X1 U9047 ( .B1(n7421), .B2(n8634), .A(n7420), .ZN(n7422) );
  INV_X1 U9048 ( .A(n7422), .ZN(P1_U3213) );
  NAND2_X1 U9049 ( .A1(n4528), .A2(n7423), .ZN(n8627) );
  OAI21_X1 U9050 ( .B1(n4528), .B2(n7423), .A(n8627), .ZN(n7424) );
  NOR2_X1 U9051 ( .A1(n7424), .A2(n7425), .ZN(n8629) );
  AOI21_X1 U9052 ( .B1(n7425), .B2(n7424), .A(n8629), .ZN(n7432) );
  NAND2_X1 U9053 ( .A1(n9497), .A2(n8670), .ZN(n7426) );
  OAI211_X1 U9054 ( .C1(n7428), .C2(n9489), .A(n7427), .B(n7426), .ZN(n7429)
         );
  AOI21_X1 U9055 ( .B1(n7430), .B2(n8656), .A(n7429), .ZN(n7431) );
  OAI21_X1 U9056 ( .B1(n7432), .B2(n9493), .A(n7431), .ZN(P1_U3227) );
  INV_X1 U9057 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U9058 ( .A1(n8154), .A2(P2_U3893), .ZN(n7434) );
  OAI21_X1 U9059 ( .B1(P2_U3893), .B2(n10073), .A(n7434), .ZN(P2_U3522) );
  NAND2_X1 U9060 ( .A1(n8671), .A2(n8668), .ZN(n7435) );
  NAND2_X1 U9061 ( .A1(n7436), .A2(n7435), .ZN(n7437) );
  INV_X1 U9062 ( .A(n8674), .ZN(n8672) );
  NAND2_X1 U9063 ( .A1(n8672), .A2(n8932), .ZN(n8666) );
  INV_X1 U9064 ( .A(n8932), .ZN(n8673) );
  NAND2_X1 U9065 ( .A1(n8673), .A2(n8674), .ZN(n8665) );
  NAND2_X1 U9066 ( .A1(n8666), .A2(n8665), .ZN(n7439) );
  NAND2_X1 U9067 ( .A1(n7437), .A2(n7439), .ZN(n7498) );
  OAI21_X1 U9068 ( .B1(n7437), .B2(n7439), .A(n7498), .ZN(n7438) );
  INV_X1 U9069 ( .A(n7438), .ZN(n7456) );
  XNOR2_X1 U9070 ( .A(n7518), .B(n7439), .ZN(n7442) );
  NAND2_X1 U9071 ( .A1(n8933), .A2(n8595), .ZN(n7441) );
  NAND2_X1 U9072 ( .A1(n8931), .A2(n9012), .ZN(n7440) );
  NAND2_X1 U9073 ( .A1(n7441), .A2(n7440), .ZN(n8637) );
  AOI21_X1 U9074 ( .B1(n7442), .B2(n9278), .A(n8637), .ZN(n7450) );
  INV_X1 U9075 ( .A(n7443), .ZN(n7444) );
  NAND2_X1 U9076 ( .A1(n7443), .A2(n8672), .ZN(n7492) );
  INV_X1 U9077 ( .A(n7492), .ZN(n7558) );
  AOI21_X1 U9078 ( .B1(n8674), .B2(n7444), .A(n7558), .ZN(n7453) );
  AOI22_X1 U9079 ( .A1(n7453), .A2(n9333), .B1(n9382), .B2(n8674), .ZN(n7445)
         );
  OAI211_X1 U9080 ( .C1(n9384), .C2(n7456), .A(n7450), .B(n7445), .ZN(n7447)
         );
  NAND2_X1 U9081 ( .A1(n7447), .A2(n9667), .ZN(n7446) );
  OAI21_X1 U9082 ( .B1(n9667), .B2(n6839), .A(n7446), .ZN(P1_U3528) );
  INV_X1 U9083 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7449) );
  NAND2_X1 U9084 ( .A1(n7447), .A2(n9439), .ZN(n7448) );
  OAI21_X1 U9085 ( .B1(n9439), .B2(n7449), .A(n7448), .ZN(P1_U3471) );
  MUX2_X1 U9086 ( .A(n7450), .B(n6833), .S(n9609), .Z(n7455) );
  INV_X1 U9087 ( .A(n8638), .ZN(n7451) );
  OAI22_X1 U9088 ( .A1(n9602), .A2(n8672), .B1(n7451), .B2(n9236), .ZN(n7452)
         );
  AOI21_X1 U9089 ( .B1(n7453), .B2(n9182), .A(n7452), .ZN(n7454) );
  OAI211_X1 U9090 ( .C1(n7456), .C2(n9294), .A(n7455), .B(n7454), .ZN(P1_U3287) );
  OR2_X1 U9091 ( .A1(n7457), .A2(n7462), .ZN(n7458) );
  INV_X1 U9092 ( .A(n7465), .ZN(n9893) );
  INV_X1 U9093 ( .A(n7459), .ZN(n7460) );
  AOI21_X1 U9094 ( .B1(n7462), .B2(n7461), .A(n7460), .ZN(n7467) );
  INV_X1 U9095 ( .A(n7615), .ZN(n9864) );
  OAI22_X1 U9096 ( .A1(n7463), .A2(n9860), .B1(n7640), .B2(n9861), .ZN(n7464)
         );
  AOI21_X1 U9097 ( .B1(n7465), .B2(n9864), .A(n7464), .ZN(n7466) );
  OAI21_X1 U9098 ( .B1(n7467), .B2(n9867), .A(n7466), .ZN(n9894) );
  NAND2_X1 U9099 ( .A1(n9894), .A2(n8318), .ZN(n7471) );
  OAI22_X1 U9100 ( .A1(n8318), .A2(n5396), .B1(n7468), .B2(n9857), .ZN(n7469)
         );
  AOI21_X1 U9101 ( .B1(n9896), .B2(n8304), .A(n7469), .ZN(n7470) );
  OAI211_X1 U9102 ( .C1(n9893), .C2(n7881), .A(n7471), .B(n7470), .ZN(P2_U3226) );
  NAND2_X1 U9103 ( .A1(n7472), .A2(n7598), .ZN(n7473) );
  XNOR2_X1 U9104 ( .A(n9897), .B(n7960), .ZN(n7642) );
  XNOR2_X1 U9105 ( .A(n7647), .B(n7642), .ZN(n7503) );
  XNOR2_X1 U9106 ( .A(n7503), .B(n4657), .ZN(n7482) );
  INV_X1 U9107 ( .A(n7475), .ZN(n7477) );
  NOR2_X1 U9108 ( .A1(n8045), .A2(n7598), .ZN(n7476) );
  AOI211_X1 U9109 ( .C1(n8042), .C2(n7650), .A(n7477), .B(n7476), .ZN(n7478)
         );
  OAI21_X1 U9110 ( .B1(n7603), .B2(n7989), .A(n7478), .ZN(n7479) );
  AOI21_X1 U9111 ( .B1(n7480), .B2(n8047), .A(n7479), .ZN(n7481) );
  OAI21_X1 U9112 ( .B1(n7482), .B2(n8050), .A(n7481), .ZN(P2_U3161) );
  NAND3_X1 U9113 ( .A1(n7483), .A2(n8666), .A3(n8856), .ZN(n7484) );
  NAND2_X1 U9114 ( .A1(n7484), .A2(n8665), .ZN(n7552) );
  INV_X1 U9115 ( .A(n8931), .ZN(n7485) );
  OR2_X1 U9116 ( .A1(n9588), .A2(n7485), .ZN(n8682) );
  NAND2_X1 U9117 ( .A1(n9588), .A2(n7485), .ZN(n7514) );
  NAND2_X1 U9118 ( .A1(n8682), .A2(n7514), .ZN(n8677) );
  INV_X1 U9119 ( .A(n8677), .ZN(n7553) );
  NAND2_X1 U9120 ( .A1(n7552), .A2(n7553), .ZN(n7551) );
  NAND2_X1 U9121 ( .A1(n7530), .A2(n7486), .ZN(n8684) );
  NAND2_X1 U9122 ( .A1(n8683), .A2(n8684), .ZN(n7528) );
  INV_X1 U9123 ( .A(n7528), .ZN(n7487) );
  NAND3_X1 U9124 ( .A1(n7551), .A2(n7487), .A3(n7514), .ZN(n7569) );
  NAND2_X1 U9125 ( .A1(n7569), .A2(n9278), .ZN(n7491) );
  AOI21_X1 U9126 ( .B1(n7551), .B2(n7514), .A(n7487), .ZN(n7490) );
  NAND2_X1 U9127 ( .A1(n8931), .A2(n8595), .ZN(n7489) );
  NAND2_X1 U9128 ( .A1(n8929), .A2(n9012), .ZN(n7488) );
  AND2_X1 U9129 ( .A1(n7489), .A2(n7488), .ZN(n7590) );
  OAI21_X1 U9130 ( .B1(n7491), .B2(n7490), .A(n7590), .ZN(n9647) );
  AOI21_X1 U9131 ( .B1(n7593), .B2(n9598), .A(n9647), .ZN(n7502) );
  AOI21_X1 U9132 ( .B1(n7557), .B2(n7530), .A(n9286), .ZN(n7493) );
  NAND2_X1 U9133 ( .A1(n7493), .A2(n7573), .ZN(n9645) );
  INV_X1 U9134 ( .A(n9645), .ZN(n7496) );
  INV_X1 U9135 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7494) );
  OAI22_X1 U9136 ( .A1(n9646), .A2(n9602), .B1(n7494), .B2(n9272), .ZN(n7495)
         );
  AOI21_X1 U9137 ( .B1(n7496), .B2(n9596), .A(n7495), .ZN(n7501) );
  OR2_X1 U9138 ( .A1(n8932), .A2(n8674), .ZN(n7497) );
  NAND2_X1 U9139 ( .A1(n7498), .A2(n7497), .ZN(n7550) );
  OR2_X1 U9140 ( .A1(n9588), .A2(n8931), .ZN(n7499) );
  XNOR2_X1 U9141 ( .A(n7529), .B(n7528), .ZN(n9649) );
  NAND2_X1 U9142 ( .A1(n9649), .A2(n9606), .ZN(n7500) );
  OAI211_X1 U9143 ( .C1(n7502), .C2(n9609), .A(n7501), .B(n7500), .ZN(P1_U3285) );
  INV_X1 U9144 ( .A(n7642), .ZN(n7639) );
  AOI22_X1 U9145 ( .A1(n7503), .A2(n7640), .B1(n7647), .B2(n7639), .ZN(n7506)
         );
  XNOR2_X1 U9146 ( .A(n9906), .B(n7504), .ZN(n7643) );
  XNOR2_X1 U9147 ( .A(n7643), .B(n7705), .ZN(n7505) );
  XNOR2_X1 U9148 ( .A(n7506), .B(n7505), .ZN(n7513) );
  INV_X1 U9149 ( .A(n7507), .ZN(n7509) );
  NOR2_X1 U9150 ( .A1(n8045), .A2(n7640), .ZN(n7508) );
  AOI211_X1 U9151 ( .C1(n8042), .C2(n8073), .A(n7509), .B(n7508), .ZN(n7510)
         );
  OAI21_X1 U9152 ( .B1(n7616), .B2(n7989), .A(n7510), .ZN(n7511) );
  AOI21_X1 U9153 ( .B1(n9906), .B2(n8047), .A(n7511), .ZN(n7512) );
  OAI21_X1 U9154 ( .B1(n7513), .B2(n8050), .A(n7512), .ZN(P2_U3171) );
  AND2_X1 U9155 ( .A1(n8684), .A2(n7514), .ZN(n8686) );
  OR2_X1 U9156 ( .A1(n7687), .A2(n7515), .ZN(n8698) );
  NAND2_X1 U9157 ( .A1(n8683), .A2(n8698), .ZN(n8685) );
  OR2_X1 U9158 ( .A1(n8686), .A2(n8685), .ZN(n7516) );
  NAND2_X1 U9159 ( .A1(n7687), .A2(n7515), .ZN(n8687) );
  NAND2_X1 U9160 ( .A1(n7516), .A2(n8687), .ZN(n7519) );
  INV_X1 U9161 ( .A(n8665), .ZN(n8789) );
  NOR2_X1 U9162 ( .A1(n7519), .A2(n8789), .ZN(n7517) );
  INV_X1 U9163 ( .A(n7519), .ZN(n8792) );
  INV_X1 U9164 ( .A(n8666), .ZN(n8669) );
  INV_X1 U9165 ( .A(n8682), .ZN(n7520) );
  OR3_X1 U9166 ( .A1(n8685), .A2(n8669), .A3(n7520), .ZN(n8788) );
  OR2_X1 U9167 ( .A1(n9498), .A2(n7521), .ZN(n8861) );
  NAND2_X1 U9168 ( .A1(n9498), .A2(n7521), .ZN(n8688) );
  NAND2_X1 U9169 ( .A1(n8861), .A2(n8688), .ZN(n8787) );
  NAND2_X1 U9170 ( .A1(n7522), .A2(n8787), .ZN(n7523) );
  NAND2_X1 U9171 ( .A1(n7668), .A2(n7523), .ZN(n7527) );
  NAND2_X1 U9172 ( .A1(n8929), .A2(n8595), .ZN(n7525) );
  NAND2_X1 U9173 ( .A1(n8927), .A2(n9012), .ZN(n7524) );
  AND2_X1 U9174 ( .A1(n7525), .A2(n7524), .ZN(n9490) );
  INV_X1 U9175 ( .A(n9490), .ZN(n7526) );
  AOI21_X1 U9176 ( .B1(n7527), .B2(n9278), .A(n7526), .ZN(n7541) );
  NAND2_X1 U9177 ( .A1(n8698), .A2(n8687), .ZN(n7571) );
  NAND2_X1 U9178 ( .A1(n7568), .A2(n7571), .ZN(n7567) );
  OR2_X1 U9179 ( .A1(n7687), .A2(n8929), .ZN(n7531) );
  NAND2_X1 U9180 ( .A1(n7567), .A2(n7531), .ZN(n7532) );
  NAND2_X1 U9181 ( .A1(n7532), .A2(n8787), .ZN(n7622) );
  OAI21_X1 U9182 ( .B1(n7532), .B2(n8787), .A(n7622), .ZN(n7539) );
  NAND2_X1 U9183 ( .A1(n7539), .A2(n9606), .ZN(n7538) );
  INV_X1 U9184 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7533) );
  OAI22_X1 U9185 ( .A1(n9272), .A2(n7533), .B1(n9500), .B2(n9236), .ZN(n7536)
         );
  INV_X1 U9186 ( .A(n7633), .ZN(n7534) );
  OAI211_X1 U9187 ( .C1(n7544), .C2(n7575), .A(n7534), .B(n9333), .ZN(n7540)
         );
  NOR2_X1 U9188 ( .A1(n7540), .A2(n9241), .ZN(n7535) );
  AOI211_X1 U9189 ( .C1(n9587), .C2(n9498), .A(n7536), .B(n7535), .ZN(n7537)
         );
  OAI211_X1 U9190 ( .C1(n9609), .C2(n7541), .A(n7538), .B(n7537), .ZN(P1_U3283) );
  INV_X1 U9191 ( .A(n7539), .ZN(n7548) );
  INV_X1 U9192 ( .A(n9361), .ZN(n9372) );
  NAND2_X1 U9193 ( .A1(n7541), .A2(n7540), .ZN(n7546) );
  OAI22_X1 U9194 ( .A1(n7544), .A2(n9367), .B1(n9667), .B2(n6952), .ZN(n7542)
         );
  AOI21_X1 U9195 ( .B1(n7546), .B2(n9667), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9196 ( .B1(n7548), .B2(n9372), .A(n7543), .ZN(P1_U3532) );
  INV_X1 U9197 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10105) );
  OAI22_X1 U9198 ( .A1(n7544), .A2(n9444), .B1(n9439), .B2(n10105), .ZN(n7545)
         );
  AOI21_X1 U9199 ( .B1(n7546), .B2(n9439), .A(n7545), .ZN(n7547) );
  OAI21_X1 U9200 ( .B1(n7548), .B2(n9449), .A(n7547), .ZN(P1_U3483) );
  INV_X1 U9201 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7562) );
  OAI21_X1 U9202 ( .B1(n7550), .B2(n8677), .A(n7549), .ZN(n9592) );
  INV_X1 U9203 ( .A(n9592), .ZN(n7559) );
  OAI21_X1 U9204 ( .B1(n7553), .B2(n7552), .A(n7551), .ZN(n7556) );
  NOR2_X1 U9205 ( .A1(n7559), .A2(n7626), .ZN(n7554) );
  AOI211_X1 U9206 ( .C1(n9278), .C2(n7556), .A(n7555), .B(n7554), .ZN(n9595)
         );
  INV_X1 U9207 ( .A(n9588), .ZN(n7563) );
  OAI211_X1 U9208 ( .C1(n7558), .C2(n7563), .A(n9333), .B(n7557), .ZN(n9589)
         );
  OAI211_X1 U9209 ( .C1(n7559), .C2(n9652), .A(n9595), .B(n9589), .ZN(n7565)
         );
  NAND2_X1 U9210 ( .A1(n7565), .A2(n9667), .ZN(n7561) );
  NAND2_X1 U9211 ( .A1(n9354), .A2(n9588), .ZN(n7560) );
  OAI211_X1 U9212 ( .C1(n9667), .C2(n7562), .A(n7561), .B(n7560), .ZN(P1_U3529) );
  INV_X1 U9213 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10062) );
  OAI22_X1 U9214 ( .A1(n7563), .A2(n9444), .B1(n9439), .B2(n10062), .ZN(n7564)
         );
  AOI21_X1 U9215 ( .B1(n7565), .B2(n9439), .A(n7564), .ZN(n7566) );
  INV_X1 U9216 ( .A(n7566), .ZN(P1_U3474) );
  OAI21_X1 U9217 ( .B1(n7568), .B2(n7571), .A(n7567), .ZN(n7686) );
  INV_X1 U9218 ( .A(n7686), .ZN(n7582) );
  NAND2_X1 U9219 ( .A1(n7569), .A2(n8683), .ZN(n7570) );
  XOR2_X1 U9220 ( .A(n7571), .B(n7570), .Z(n7572) );
  NAND2_X1 U9221 ( .A1(n8930), .A2(n8595), .ZN(n7722) );
  OAI21_X1 U9222 ( .B1(n7572), .B2(n9215), .A(n7722), .ZN(n7684) );
  NAND2_X1 U9223 ( .A1(n7684), .A2(n9272), .ZN(n7581) );
  INV_X1 U9224 ( .A(n7573), .ZN(n7574) );
  OAI21_X1 U9225 ( .B1(n7574), .B2(n7728), .A(n9333), .ZN(n7576) );
  NAND2_X1 U9226 ( .A1(n8928), .A2(n9012), .ZN(n7721) );
  OAI21_X1 U9227 ( .B1(n7576), .B2(n7575), .A(n7721), .ZN(n7685) );
  NOR2_X1 U9228 ( .A1(n7728), .A2(n9602), .ZN(n7579) );
  INV_X1 U9229 ( .A(n7725), .ZN(n7577) );
  OAI22_X1 U9230 ( .A1(n9272), .A2(n6878), .B1(n7577), .B2(n9236), .ZN(n7578)
         );
  AOI211_X1 U9231 ( .C1(n7685), .C2(n9596), .A(n7579), .B(n7578), .ZN(n7580)
         );
  OAI211_X1 U9232 ( .C1(n7582), .C2(n9294), .A(n7581), .B(n7580), .ZN(P1_U3284) );
  INV_X1 U9233 ( .A(n7583), .ZN(n7585) );
  OAI222_X1 U9234 ( .A1(n8480), .A2(n7584), .B1(n8483), .B2(n7585), .C1(n8125), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9235 ( .A1(n9466), .A2(n10201), .B1(n7778), .B2(n7585), .C1(n4437), .C2(n6345), .ZN(P1_U3336) );
  XNOR2_X1 U9236 ( .A(n7587), .B(n7586), .ZN(n7588) );
  NAND2_X1 U9237 ( .A1(n7588), .A2(n8634), .ZN(n7595) );
  INV_X1 U9238 ( .A(n7589), .ZN(n7592) );
  NOR2_X1 U9239 ( .A1(n7590), .A2(n9489), .ZN(n7591) );
  AOI211_X1 U9240 ( .C1(n7593), .C2(n8656), .A(n7592), .B(n7591), .ZN(n7594)
         );
  OAI211_X1 U9241 ( .C1(n9646), .C2(n8651), .A(n7595), .B(n7594), .ZN(P1_U3221) );
  XOR2_X1 U9242 ( .A(n7596), .B(n7601), .Z(n7597) );
  OAI222_X1 U9243 ( .A1(n9861), .A2(n7705), .B1(n9860), .B2(n7598), .C1(n9867), 
        .C2(n7597), .ZN(n9898) );
  INV_X1 U9244 ( .A(n9898), .ZN(n7608) );
  NAND2_X1 U9245 ( .A1(n7600), .A2(n7599), .ZN(n7602) );
  XNOR2_X1 U9246 ( .A(n7602), .B(n7601), .ZN(n9900) );
  NOR2_X1 U9247 ( .A1(n9897), .A2(n8176), .ZN(n7606) );
  OAI22_X1 U9248 ( .A1(n8318), .A2(n7604), .B1(n7603), .B2(n9857), .ZN(n7605)
         );
  AOI211_X1 U9249 ( .C1(n9900), .C2(n8260), .A(n7606), .B(n7605), .ZN(n7607)
         );
  OAI21_X1 U9250 ( .B1(n7608), .B2(n9871), .A(n7607), .ZN(P2_U3225) );
  OAI21_X1 U9251 ( .B1(n7609), .B2(n5779), .A(n7707), .ZN(n9903) );
  XNOR2_X1 U9252 ( .A(n7611), .B(n7610), .ZN(n7612) );
  NAND2_X1 U9253 ( .A1(n7612), .A2(n8331), .ZN(n7614) );
  AOI22_X1 U9254 ( .A1(n4657), .A2(n8328), .B1(n8326), .B2(n8073), .ZN(n7613)
         );
  OAI211_X1 U9255 ( .C1(n7615), .C2(n9903), .A(n7614), .B(n7613), .ZN(n9904)
         );
  NAND2_X1 U9256 ( .A1(n9904), .A2(n8318), .ZN(n7620) );
  OAI22_X1 U9257 ( .A1(n8318), .A2(n7617), .B1(n7616), .B2(n9857), .ZN(n7618)
         );
  AOI21_X1 U9258 ( .B1(n9906), .B2(n8304), .A(n7618), .ZN(n7619) );
  OAI211_X1 U9259 ( .C1(n9903), .C2(n7881), .A(n7620), .B(n7619), .ZN(P2_U3224) );
  OR2_X1 U9260 ( .A1(n9498), .A2(n8928), .ZN(n7621) );
  NAND2_X1 U9261 ( .A1(n7622), .A2(n7621), .ZN(n7624) );
  INV_X1 U9262 ( .A(n8927), .ZN(n7623) );
  OR2_X1 U9263 ( .A1(n7661), .A2(n7623), .ZN(n8700) );
  NAND2_X1 U9264 ( .A1(n7661), .A2(n7623), .ZN(n8701) );
  NAND2_X1 U9265 ( .A1(n8700), .A2(n8701), .ZN(n8777) );
  NAND2_X1 U9266 ( .A1(n7624), .A2(n8777), .ZN(n7663) );
  OR2_X1 U9267 ( .A1(n7624), .A2(n8777), .ZN(n7625) );
  NAND2_X1 U9268 ( .A1(n7663), .A2(n7625), .ZN(n9658) );
  INV_X1 U9269 ( .A(n7626), .ZN(n7768) );
  NAND2_X1 U9270 ( .A1(n7668), .A2(n8688), .ZN(n7627) );
  XNOR2_X1 U9271 ( .A(n7627), .B(n8777), .ZN(n7630) );
  NAND2_X1 U9272 ( .A1(n8926), .A2(n9012), .ZN(n7629) );
  NAND2_X1 U9273 ( .A1(n8928), .A2(n8595), .ZN(n7628) );
  AND2_X1 U9274 ( .A1(n7629), .A2(n7628), .ZN(n7834) );
  OAI21_X1 U9275 ( .B1(n7630), .B2(n9215), .A(n7834), .ZN(n7631) );
  AOI21_X1 U9276 ( .B1(n9658), .B2(n7768), .A(n7631), .ZN(n9660) );
  NOR2_X1 U9277 ( .A1(n9609), .A2(n7632), .ZN(n9591) );
  INV_X1 U9278 ( .A(n7661), .ZN(n9655) );
  OAI21_X1 U9279 ( .B1(n7633), .B2(n9655), .A(n9333), .ZN(n7634) );
  OR2_X1 U9280 ( .A1(n7676), .A2(n7634), .ZN(n9653) );
  AOI22_X1 U9281 ( .A1(n9609), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7836), .B2(
        n9598), .ZN(n7636) );
  NAND2_X1 U9282 ( .A1(n7661), .A2(n9587), .ZN(n7635) );
  OAI211_X1 U9283 ( .C1(n9653), .C2(n9241), .A(n7636), .B(n7635), .ZN(n7637)
         );
  AOI21_X1 U9284 ( .B1(n9658), .B2(n9591), .A(n7637), .ZN(n7638) );
  OAI21_X1 U9285 ( .B1(n9660), .B2(n9609), .A(n7638), .ZN(P1_U3282) );
  OAI22_X1 U9286 ( .A1(n7642), .A2(n4657), .B1(n7643), .B2(n7650), .ZN(n7646)
         );
  OAI21_X1 U9287 ( .B1(n7639), .B2(n7640), .A(n7705), .ZN(n7644) );
  NOR2_X1 U9288 ( .A1(n7705), .A2(n7640), .ZN(n7641) );
  AOI22_X1 U9289 ( .A1(n7644), .A2(n7643), .B1(n7642), .B2(n7641), .ZN(n7645)
         );
  XNOR2_X1 U9290 ( .A(n9910), .B(n7917), .ZN(n7744) );
  XOR2_X1 U9291 ( .A(n7745), .B(n7744), .Z(n7655) );
  NAND2_X1 U9292 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9727) );
  INV_X1 U9293 ( .A(n9727), .ZN(n7649) );
  NOR2_X1 U9294 ( .A1(n8059), .A2(n7747), .ZN(n7648) );
  AOI211_X1 U9295 ( .C1(n8057), .C2(n7650), .A(n7649), .B(n7648), .ZN(n7651)
         );
  OAI21_X1 U9296 ( .B1(n7710), .B2(n7989), .A(n7651), .ZN(n7652) );
  AOI21_X1 U9297 ( .B1(n7653), .B2(n8047), .A(n7652), .ZN(n7654) );
  OAI21_X1 U9298 ( .B1(n7655), .B2(n8050), .A(n7654), .ZN(P2_U3157) );
  INV_X1 U9299 ( .A(n7656), .ZN(n7660) );
  INV_X1 U9300 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7657) );
  OAI222_X1 U9301 ( .A1(n6677), .A2(n7660), .B1(P2_U3151), .B2(n7658), .C1(
        n7657), .C2(n8480), .ZN(P2_U3275) );
  INV_X1 U9302 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7659) );
  OAI222_X1 U9303 ( .A1(P1_U3086), .A2(n8808), .B1(n7778), .B2(n7660), .C1(
        n7659), .C2(n9466), .ZN(P1_U3335) );
  OR2_X1 U9304 ( .A1(n7661), .A2(n8927), .ZN(n7662) );
  NAND2_X1 U9305 ( .A1(n7663), .A2(n7662), .ZN(n7665) );
  INV_X1 U9306 ( .A(n8926), .ZN(n7664) );
  OR2_X1 U9307 ( .A1(n7730), .A2(n7664), .ZN(n8704) );
  NAND2_X1 U9308 ( .A1(n7730), .A2(n7664), .ZN(n8867) );
  NAND2_X1 U9309 ( .A1(n8704), .A2(n8867), .ZN(n7669) );
  OAI21_X1 U9310 ( .B1(n7665), .B2(n7669), .A(n7732), .ZN(n7693) );
  INV_X1 U9311 ( .A(n7693), .ZN(n7683) );
  INV_X1 U9312 ( .A(n8688), .ZN(n8697) );
  NOR2_X1 U9313 ( .A1(n8777), .A2(n8697), .ZN(n7667) );
  INV_X1 U9314 ( .A(n8700), .ZN(n7666) );
  INV_X1 U9315 ( .A(n7669), .ZN(n8794) );
  OR2_X1 U9316 ( .A1(n7670), .A2(n8794), .ZN(n7671) );
  NAND2_X1 U9317 ( .A1(n7733), .A2(n7671), .ZN(n7675) );
  NAND2_X1 U9318 ( .A1(n8925), .A2(n9012), .ZN(n7673) );
  NAND2_X1 U9319 ( .A1(n8927), .A2(n8595), .ZN(n7672) );
  AND2_X1 U9320 ( .A1(n7673), .A2(n7672), .ZN(n7857) );
  INV_X1 U9321 ( .A(n7857), .ZN(n7674) );
  AOI21_X1 U9322 ( .B1(n7675), .B2(n9278), .A(n7674), .ZN(n7700) );
  NAND2_X1 U9323 ( .A1(n7676), .A2(n7862), .ZN(n7738) );
  OAI211_X1 U9324 ( .C1(n7676), .C2(n7862), .A(n9333), .B(n7738), .ZN(n7695)
         );
  NAND2_X1 U9325 ( .A1(n7700), .A2(n7695), .ZN(n7681) );
  INV_X1 U9326 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7677) );
  OAI22_X1 U9327 ( .A1(n7862), .A2(n9444), .B1(n9439), .B2(n7677), .ZN(n7678)
         );
  AOI21_X1 U9328 ( .B1(n7681), .B2(n9439), .A(n7678), .ZN(n7679) );
  OAI21_X1 U9329 ( .B1(n7683), .B2(n9449), .A(n7679), .ZN(P1_U3489) );
  OAI22_X1 U9330 ( .A1(n7862), .A2(n9367), .B1(n9667), .B2(n7131), .ZN(n7680)
         );
  AOI21_X1 U9331 ( .B1(n7681), .B2(n9667), .A(n7680), .ZN(n7682) );
  OAI21_X1 U9332 ( .B1(n7683), .B2(n9372), .A(n7682), .ZN(P1_U3534) );
  AOI211_X1 U9333 ( .C1(n9650), .C2(n7686), .A(n7685), .B(n7684), .ZN(n7692)
         );
  AOI22_X1 U9334 ( .A1(n7687), .A2(n9354), .B1(n9665), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7688) );
  OAI21_X1 U9335 ( .B1(n7692), .B2(n9665), .A(n7688), .ZN(P1_U3531) );
  INV_X1 U9336 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7689) );
  OAI22_X1 U9337 ( .A1(n7728), .A2(n9444), .B1(n9439), .B2(n7689), .ZN(n7690)
         );
  INV_X1 U9338 ( .A(n7690), .ZN(n7691) );
  OAI21_X1 U9339 ( .B1(n7692), .B2(n9661), .A(n7691), .ZN(P1_U3480) );
  NAND2_X1 U9340 ( .A1(n7693), .A2(n9606), .ZN(n7699) );
  OAI22_X1 U9341 ( .A1(n9272), .A2(n7140), .B1(n7694), .B2(n9236), .ZN(n7697)
         );
  NOR2_X1 U9342 ( .A1(n7695), .A2(n9241), .ZN(n7696) );
  AOI211_X1 U9343 ( .C1(n9587), .C2(n7730), .A(n7697), .B(n7696), .ZN(n7698)
         );
  OAI211_X1 U9344 ( .C1(n9609), .C2(n7700), .A(n7699), .B(n7698), .ZN(P1_U3281) );
  INV_X1 U9345 ( .A(n7701), .ZN(n7702) );
  OAI222_X1 U9346 ( .A1(n8483), .A2(n7702), .B1(P2_U3151), .B2(n4808), .C1(
        n10029), .C2(n8480), .ZN(P2_U3274) );
  OAI222_X1 U9347 ( .A1(n9466), .A2(n10193), .B1(n7778), .B2(n7702), .C1(n6522), .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U9348 ( .A(n7703), .B(n7708), .ZN(n7704) );
  OAI222_X1 U9349 ( .A1(n9860), .A2(n7705), .B1(n9861), .B2(n7747), .C1(n7704), 
        .C2(n9867), .ZN(n9911) );
  INV_X1 U9350 ( .A(n9911), .ZN(n7714) );
  NAND2_X1 U9351 ( .A1(n7707), .A2(n7706), .ZN(n7709) );
  XNOR2_X1 U9352 ( .A(n7709), .B(n7708), .ZN(n9913) );
  NOR2_X1 U9353 ( .A1(n9910), .A2(n8176), .ZN(n7712) );
  OAI22_X1 U9354 ( .A1(n8318), .A2(n8083), .B1(n7710), .B2(n9857), .ZN(n7711)
         );
  AOI211_X1 U9355 ( .C1(n9913), .C2(n8260), .A(n7712), .B(n7711), .ZN(n7713)
         );
  OAI21_X1 U9356 ( .B1(n7714), .B2(n9871), .A(n7713), .ZN(P2_U3223) );
  INV_X1 U9357 ( .A(n7715), .ZN(n7717) );
  NAND2_X1 U9358 ( .A1(n7717), .A2(n7716), .ZN(n7719) );
  XNOR2_X1 U9359 ( .A(n7719), .B(n7718), .ZN(n7720) );
  NAND2_X1 U9360 ( .A1(n7720), .A2(n8634), .ZN(n7727) );
  AOI21_X1 U9361 ( .B1(n7722), .B2(n7721), .A(n9489), .ZN(n7723) );
  AOI211_X1 U9362 ( .C1(n8656), .C2(n7725), .A(n7724), .B(n7723), .ZN(n7726)
         );
  OAI211_X1 U9363 ( .C1(n7728), .C2(n8651), .A(n7727), .B(n7726), .ZN(P1_U3231) );
  INV_X1 U9364 ( .A(n9381), .ZN(n8612) );
  NAND2_X1 U9365 ( .A1(n8612), .A2(n8925), .ZN(n8870) );
  INV_X1 U9366 ( .A(n8925), .ZN(n7729) );
  NAND2_X1 U9367 ( .A1(n9381), .A2(n7729), .ZN(n8868) );
  NAND2_X1 U9368 ( .A1(n8870), .A2(n8868), .ZN(n8796) );
  OR2_X1 U9369 ( .A1(n7730), .A2(n8926), .ZN(n7731) );
  XOR2_X1 U9370 ( .A(n8796), .B(n7764), .Z(n9385) );
  XNOR2_X1 U9371 ( .A(n7765), .B(n8796), .ZN(n7736) );
  NAND2_X1 U9372 ( .A1(n8924), .A2(n9012), .ZN(n7735) );
  NAND2_X1 U9373 ( .A1(n8926), .A2(n8595), .ZN(n7734) );
  AND2_X1 U9374 ( .A1(n7735), .A2(n7734), .ZN(n8607) );
  OAI21_X1 U9375 ( .B1(n7736), .B2(n9215), .A(n8607), .ZN(n9379) );
  INV_X1 U9376 ( .A(n7769), .ZN(n7737) );
  AOI211_X1 U9377 ( .C1(n9381), .C2(n7738), .A(n9286), .B(n7737), .ZN(n9380)
         );
  NAND2_X1 U9378 ( .A1(n9380), .A2(n9596), .ZN(n7740) );
  AOI22_X1 U9379 ( .A1(n9609), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8609), .B2(
        n9598), .ZN(n7739) );
  OAI211_X1 U9380 ( .C1(n8612), .C2(n9602), .A(n7740), .B(n7739), .ZN(n7741)
         );
  AOI21_X1 U9381 ( .B1(n9272), .B2(n9379), .A(n7741), .ZN(n7742) );
  OAI21_X1 U9382 ( .B1(n9385), .B2(n9294), .A(n7742), .ZN(P1_U3280) );
  XNOR2_X1 U9383 ( .A(n7780), .B(n7960), .ZN(n7760) );
  XNOR2_X1 U9384 ( .A(n8382), .B(n7960), .ZN(n7891) );
  XNOR2_X1 U9385 ( .A(n7891), .B(n8022), .ZN(n7746) );
  XNOR2_X1 U9386 ( .A(n7892), .B(n7746), .ZN(n7753) );
  NAND2_X1 U9387 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9761) );
  INV_X1 U9388 ( .A(n9761), .ZN(n7749) );
  NOR2_X1 U9389 ( .A1(n8045), .A2(n7747), .ZN(n7748) );
  AOI211_X1 U9390 ( .C1(n8042), .C2(n8313), .A(n7749), .B(n7748), .ZN(n7750)
         );
  OAI21_X1 U9391 ( .B1(n7805), .B2(n7989), .A(n7750), .ZN(n7751) );
  AOI21_X1 U9392 ( .B1(n8382), .B2(n8047), .A(n7751), .ZN(n7752) );
  OAI21_X1 U9393 ( .B1(n7753), .B2(n8050), .A(n7752), .ZN(P2_U3164) );
  NAND2_X1 U9394 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9744) );
  INV_X1 U9395 ( .A(n9744), .ZN(n7756) );
  NOR2_X1 U9396 ( .A1(n7754), .A2(n8045), .ZN(n7755) );
  AOI211_X1 U9397 ( .C1(n8042), .C2(n8329), .A(n7756), .B(n7755), .ZN(n7757)
         );
  OAI21_X1 U9398 ( .B1(n7797), .B2(n7989), .A(n7757), .ZN(n7762) );
  AOI211_X1 U9399 ( .C1(n7760), .C2(n7758), .A(n8050), .B(n7759), .ZN(n7761)
         );
  AOI211_X1 U9400 ( .C1(n7795), .C2(n8047), .A(n7762), .B(n7761), .ZN(n7763)
         );
  INV_X1 U9401 ( .A(n7763), .ZN(P2_U3176) );
  XNOR2_X1 U9402 ( .A(n9375), .B(n8924), .ZN(n8706) );
  XNOR2_X1 U9403 ( .A(n7813), .B(n8706), .ZN(n9373) );
  INV_X1 U9404 ( .A(n8706), .ZN(n8797) );
  XNOR2_X1 U9405 ( .A(n7814), .B(n8797), .ZN(n7766) );
  AOI22_X1 U9406 ( .A1(n9012), .A2(n9023), .B1(n8925), .B2(n8595), .ZN(n8497)
         );
  OAI21_X1 U9407 ( .B1(n7766), .B2(n9215), .A(n8497), .ZN(n7767) );
  AOI21_X1 U9408 ( .B1(n9373), .B2(n7768), .A(n7767), .ZN(n9377) );
  AOI211_X1 U9409 ( .C1(n9375), .C2(n7769), .A(n9286), .B(n7821), .ZN(n9374)
         );
  NAND2_X1 U9410 ( .A1(n9374), .A2(n9596), .ZN(n7771) );
  AOI22_X1 U9411 ( .A1(n9609), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8501), .B2(
        n9598), .ZN(n7770) );
  OAI211_X1 U9412 ( .C1(n8498), .C2(n9602), .A(n7771), .B(n7770), .ZN(n7772)
         );
  AOI21_X1 U9413 ( .B1(n9373), .B2(n9591), .A(n7772), .ZN(n7773) );
  OAI21_X1 U9414 ( .B1(n9377), .B2(n9609), .A(n7773), .ZN(P1_U3279) );
  INV_X1 U9415 ( .A(n7774), .ZN(n7777) );
  OAI222_X1 U9416 ( .A1(n8480), .A2(n7776), .B1(n8483), .B2(n7777), .C1(n7775), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9417 ( .A1(n9466), .A2(n10111), .B1(n7778), .B2(n7777), .C1(
        P1_U3086), .C2(n8896), .ZN(P1_U3333) );
  OAI211_X1 U9418 ( .C1(n7781), .C2(n7780), .A(n7779), .B(n8331), .ZN(n7783)
         );
  AOI22_X1 U9419 ( .A1(n8328), .A2(n8073), .B1(n8329), .B2(n8326), .ZN(n7782)
         );
  NAND2_X1 U9420 ( .A1(n7783), .A2(n7782), .ZN(n7793) );
  MUX2_X1 U9421 ( .A(n7793), .B(P2_REG0_REG_11__SCAN_IN), .S(n9917), .Z(n7784)
         );
  INV_X1 U9422 ( .A(n7784), .ZN(n7788) );
  XNOR2_X1 U9423 ( .A(n7785), .B(n4648), .ZN(n7799) );
  INV_X1 U9424 ( .A(n8470), .ZN(n7786) );
  AOI22_X1 U9425 ( .A1(n7799), .A2(n7786), .B1(n6608), .B2(n7795), .ZN(n7787)
         );
  NAND2_X1 U9426 ( .A1(n7788), .A2(n7787), .ZN(P2_U3423) );
  MUX2_X1 U9427 ( .A(n7793), .B(P2_REG1_REG_11__SCAN_IN), .S(n9927), .Z(n7789)
         );
  INV_X1 U9428 ( .A(n7789), .ZN(n7792) );
  INV_X1 U9429 ( .A(n8381), .ZN(n7790) );
  AOI22_X1 U9430 ( .A1(n7799), .A2(n7790), .B1(n6603), .B2(n7795), .ZN(n7791)
         );
  NAND2_X1 U9431 ( .A1(n7792), .A2(n7791), .ZN(P2_U3470) );
  MUX2_X1 U9432 ( .A(n7793), .B(P2_REG2_REG_11__SCAN_IN), .S(n9871), .Z(n7794)
         );
  INV_X1 U9433 ( .A(n7794), .ZN(n7801) );
  NAND2_X1 U9434 ( .A1(n7795), .A2(n8304), .ZN(n7796) );
  OAI21_X1 U9435 ( .B1(n7797), .B2(n9857), .A(n7796), .ZN(n7798) );
  AOI21_X1 U9436 ( .B1(n7799), .B2(n8260), .A(n7798), .ZN(n7800) );
  NAND2_X1 U9437 ( .A1(n7801), .A2(n7800), .ZN(P2_U3222) );
  XNOR2_X1 U9438 ( .A(n7803), .B(n7802), .ZN(n7804) );
  AOI222_X1 U9439 ( .A1(n8331), .A2(n7804), .B1(n8313), .B2(n8326), .C1(n8072), 
        .C2(n8328), .ZN(n8386) );
  OAI22_X1 U9440 ( .A1(n8318), .A2(n7806), .B1(n7805), .B2(n9857), .ZN(n7807)
         );
  AOI21_X1 U9441 ( .B1(n8382), .B2(n8304), .A(n7807), .ZN(n7811) );
  NAND2_X1 U9442 ( .A1(n7809), .A2(n7808), .ZN(n8383) );
  NAND3_X1 U9443 ( .A1(n8384), .A2(n8383), .A3(n8260), .ZN(n7810) );
  OAI211_X1 U9444 ( .C1(n8386), .C2(n9871), .A(n7811), .B(n7810), .ZN(P2_U3221) );
  OR2_X1 U9445 ( .A1(n9024), .A2(n9020), .ZN(n8876) );
  NAND2_X1 U9446 ( .A1(n9024), .A2(n9020), .ZN(n8708) );
  NAND2_X1 U9447 ( .A1(n8876), .A2(n8708), .ZN(n8798) );
  NAND2_X1 U9448 ( .A1(n8498), .A2(n8693), .ZN(n7812) );
  XOR2_X1 U9449 ( .A(n8798), .B(n9022), .Z(n7852) );
  NAND2_X1 U9450 ( .A1(n9375), .A2(n8693), .ZN(n8707) );
  AOI21_X1 U9451 ( .B1(n7816), .B2(n8798), .A(n9215), .ZN(n7820) );
  NAND2_X1 U9452 ( .A1(n8924), .A2(n8595), .ZN(n7818) );
  NAND2_X1 U9453 ( .A1(n9027), .A2(n9012), .ZN(n7817) );
  AND2_X1 U9454 ( .A1(n7818), .A2(n7817), .ZN(n8658) );
  INV_X1 U9455 ( .A(n8658), .ZN(n7819) );
  AOI21_X1 U9456 ( .B1(n7820), .B2(n8836), .A(n7819), .ZN(n7846) );
  INV_X1 U9457 ( .A(n7846), .ZN(n7825) );
  INV_X1 U9458 ( .A(n9008), .ZN(n9287) );
  OAI211_X1 U9459 ( .C1(n9021), .C2(n7821), .A(n9287), .B(n9333), .ZN(n7845)
         );
  AOI22_X1 U9460 ( .A1(n9609), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8655), .B2(
        n9598), .ZN(n7823) );
  NAND2_X1 U9461 ( .A1(n9024), .A2(n9587), .ZN(n7822) );
  OAI211_X1 U9462 ( .C1(n7845), .C2(n9241), .A(n7823), .B(n7822), .ZN(n7824)
         );
  AOI21_X1 U9463 ( .B1(n7825), .B2(n9272), .A(n7824), .ZN(n7826) );
  OAI21_X1 U9464 ( .B1(n7852), .B2(n9294), .A(n7826), .ZN(P1_U3278) );
  INV_X1 U9465 ( .A(n7827), .ZN(n7832) );
  NOR3_X1 U9466 ( .A1(n7828), .A2(n7830), .A3(n7829), .ZN(n7831) );
  OAI21_X1 U9467 ( .B1(n7832), .B2(n7831), .A(n8634), .ZN(n7838) );
  OAI21_X1 U9468 ( .B1(n7834), .B2(n9489), .A(n7833), .ZN(n7835) );
  AOI21_X1 U9469 ( .B1(n7836), .B2(n8656), .A(n7835), .ZN(n7837) );
  OAI211_X1 U9470 ( .C1(n9655), .C2(n8651), .A(n7838), .B(n7837), .ZN(P1_U3236) );
  INV_X1 U9471 ( .A(n7839), .ZN(n7844) );
  OR2_X1 U9472 ( .A1(n7840), .A2(P1_U3086), .ZN(n8912) );
  INV_X1 U9473 ( .A(n8912), .ZN(n8902) );
  AOI21_X1 U9474 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9462), .A(n8902), .ZN(
        n7841) );
  OAI21_X1 U9475 ( .B1(n7844), .B2(n7778), .A(n7841), .ZN(P1_U3332) );
  NAND2_X1 U9476 ( .A1(n8489), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7842) );
  OAI211_X1 U9477 ( .C1(n7844), .C2(n8483), .A(n7843), .B(n7842), .ZN(P2_U3272) );
  NAND2_X1 U9478 ( .A1(n7846), .A2(n7845), .ZN(n7849) );
  MUX2_X1 U9479 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n7849), .S(n9667), .Z(n7847)
         );
  AOI21_X1 U9480 ( .B1(n9354), .B2(n9024), .A(n7847), .ZN(n7848) );
  OAI21_X1 U9481 ( .B1(n7852), .B2(n9372), .A(n7848), .ZN(P1_U3537) );
  INV_X1 U9482 ( .A(n9444), .ZN(n9430) );
  MUX2_X1 U9483 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n7849), .S(n9439), .Z(n7850)
         );
  AOI21_X1 U9484 ( .B1(n9430), .B2(n9024), .A(n7850), .ZN(n7851) );
  OAI21_X1 U9485 ( .B1(n7852), .B2(n9449), .A(n7851), .ZN(P1_U3498) );
  AND3_X1 U9486 ( .A1(n7827), .A2(n7854), .A3(n7853), .ZN(n7855) );
  OAI21_X1 U9487 ( .B1(n4526), .B2(n7855), .A(n8634), .ZN(n7861) );
  OAI21_X1 U9488 ( .B1(n7857), .B2(n9489), .A(n7856), .ZN(n7858) );
  AOI21_X1 U9489 ( .B1(n7859), .B2(n8656), .A(n7858), .ZN(n7860) );
  OAI211_X1 U9490 ( .C1(n7862), .C2(n8651), .A(n7861), .B(n7860), .ZN(P1_U3224) );
  INV_X1 U9491 ( .A(n7863), .ZN(n7867) );
  OAI222_X1 U9492 ( .A1(n6677), .A2(n7867), .B1(P2_U3151), .B2(n7865), .C1(
        n7864), .C2(n8480), .ZN(P2_U3271) );
  OAI222_X1 U9493 ( .A1(n7868), .A2(n4437), .B1(n7778), .B2(n7867), .C1(n7866), 
        .C2(n9466), .ZN(P1_U3331) );
  INV_X1 U9494 ( .A(n7869), .ZN(n7873) );
  OAI222_X1 U9495 ( .A1(n6677), .A2(n7873), .B1(P2_U3151), .B2(n7871), .C1(
        n7870), .C2(n8480), .ZN(P2_U3270) );
  OAI222_X1 U9496 ( .A1(n7874), .A2(P1_U3086), .B1(n7778), .B2(n7873), .C1(
        n7872), .C2(n9466), .ZN(P1_U3330) );
  INV_X1 U9497 ( .A(n7875), .ZN(n9467) );
  OAI222_X1 U9498 ( .A1(n6677), .A2(n9467), .B1(P2_U3151), .B2(n7877), .C1(
        n7876), .C2(n8480), .ZN(P2_U3269) );
  INV_X1 U9499 ( .A(n7878), .ZN(n7879) );
  NAND2_X1 U9500 ( .A1(n7879), .A2(n8303), .ZN(n8155) );
  OAI21_X1 U9501 ( .B1(n8318), .B2(n7880), .A(n8155), .ZN(n7884) );
  NOR2_X1 U9502 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  AOI211_X1 U9503 ( .C1(n8304), .C2(n7885), .A(n7884), .B(n7883), .ZN(n7886)
         );
  OAI21_X1 U9504 ( .B1(n7887), .B2(n9871), .A(n7886), .ZN(P2_U3204) );
  INV_X1 U9505 ( .A(n7888), .ZN(n8482) );
  AOI22_X1 U9506 ( .A1(n7889), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9462), .ZN(n7890) );
  OAI21_X1 U9507 ( .B1(n8482), .B2(n7778), .A(n7890), .ZN(P1_U3326) );
  XNOR2_X1 U9508 ( .A(n8462), .B(n7960), .ZN(n7898) );
  INV_X1 U9509 ( .A(n7891), .ZN(n7895) );
  INV_X1 U9510 ( .A(n7892), .ZN(n7894) );
  AOI21_X1 U9511 ( .B1(n7892), .B2(n7891), .A(n8022), .ZN(n7893) );
  AOI21_X1 U9512 ( .B1(n7895), .B2(n7894), .A(n7893), .ZN(n8017) );
  XNOR2_X1 U9513 ( .A(n8467), .B(n7504), .ZN(n7896) );
  NOR2_X1 U9514 ( .A1(n7896), .A2(n8313), .ZN(n7897) );
  AOI21_X1 U9515 ( .B1(n7896), .B2(n8313), .A(n7897), .ZN(n8018) );
  INV_X1 U9516 ( .A(n7897), .ZN(n7931) );
  XNOR2_X1 U9517 ( .A(n7898), .B(n7899), .ZN(n7932) );
  XNOR2_X1 U9518 ( .A(n8457), .B(n7960), .ZN(n7900) );
  XNOR2_X1 U9519 ( .A(n7900), .B(n8314), .ZN(n8054) );
  NAND2_X1 U9520 ( .A1(n8053), .A2(n7901), .ZN(n7986) );
  XOR2_X1 U9521 ( .A(n7960), .B(n8451), .Z(n7984) );
  INV_X1 U9522 ( .A(n7984), .ZN(n7902) );
  NOR2_X1 U9523 ( .A1(n7902), .A2(n8060), .ZN(n7904) );
  XNOR2_X1 U9524 ( .A(n8445), .B(n7917), .ZN(n7905) );
  XOR2_X1 U9525 ( .A(n8284), .B(n7905), .Z(n7993) );
  XNOR2_X1 U9526 ( .A(n8439), .B(n7917), .ZN(n7907) );
  XNOR2_X1 U9527 ( .A(n7907), .B(n7906), .ZN(n8034) );
  XNOR2_X1 U9528 ( .A(n8363), .B(n7504), .ZN(n7908) );
  NAND2_X1 U9529 ( .A1(n7908), .A2(n8265), .ZN(n7949) );
  XNOR2_X1 U9530 ( .A(n8432), .B(n7917), .ZN(n7909) );
  XNOR2_X1 U9531 ( .A(n7909), .B(n7972), .ZN(n8008) );
  INV_X1 U9532 ( .A(n7909), .ZN(n7910) );
  INV_X1 U9533 ( .A(n7972), .ZN(n8252) );
  XNOR2_X1 U9534 ( .A(n8426), .B(n7917), .ZN(n7911) );
  XNOR2_X1 U9535 ( .A(n7911), .B(n8244), .ZN(n7968) );
  AOI22_X1 U9536 ( .A1(n7969), .A2(n7968), .B1(n7912), .B2(n7911), .ZN(n8028)
         );
  XNOR2_X1 U9537 ( .A(n8420), .B(n7917), .ZN(n7913) );
  XNOR2_X1 U9538 ( .A(n7913), .B(n8208), .ZN(n8027) );
  INV_X1 U9539 ( .A(n7913), .ZN(n7914) );
  XNOR2_X1 U9540 ( .A(n8213), .B(n7917), .ZN(n7940) );
  XNOR2_X1 U9541 ( .A(n8005), .B(n7917), .ZN(n7915) );
  XNOR2_X1 U9542 ( .A(n7915), .B(n8071), .ZN(n8001) );
  XNOR2_X1 U9543 ( .A(n7981), .B(n7917), .ZN(n7916) );
  XNOR2_X1 U9544 ( .A(n7916), .B(n8194), .ZN(n7977) );
  XNOR2_X1 U9545 ( .A(n8398), .B(n7917), .ZN(n7918) );
  XNOR2_X1 U9546 ( .A(n7920), .B(n7918), .ZN(n8041) );
  NAND2_X1 U9547 ( .A1(n8041), .A2(n8183), .ZN(n7922) );
  INV_X1 U9548 ( .A(n7918), .ZN(n7919) );
  NAND2_X1 U9549 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  NAND2_X1 U9550 ( .A1(n7922), .A2(n7921), .ZN(n7925) );
  XNOR2_X1 U9551 ( .A(n8163), .B(n7960), .ZN(n7923) );
  NAND2_X1 U9552 ( .A1(n7923), .A2(n8069), .ZN(n7957) );
  OAI21_X1 U9553 ( .B1(n7923), .B2(n8069), .A(n7957), .ZN(n7924) );
  AOI21_X1 U9554 ( .B1(n7925), .B2(n7924), .A(n8050), .ZN(n7926) );
  NAND2_X1 U9555 ( .A1(n7926), .A2(n7958), .ZN(n7930) );
  AOI22_X1 U9556 ( .A1(n8161), .A2(n8062), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7927) );
  OAI21_X1 U9557 ( .B1(n8183), .B2(n8045), .A(n7927), .ZN(n7928) );
  AOI21_X1 U9558 ( .B1(n8068), .B2(n8042), .A(n7928), .ZN(n7929) );
  OAI211_X1 U9559 ( .C1(n8163), .C2(n8065), .A(n7930), .B(n7929), .ZN(P2_U3154) );
  INV_X1 U9560 ( .A(n8462), .ZN(n8317) );
  AND3_X1 U9561 ( .A1(n8016), .A2(n7932), .A3(n7931), .ZN(n7933) );
  OAI21_X1 U9562 ( .B1(n7934), .B2(n7933), .A(n8052), .ZN(n7939) );
  NAND2_X1 U9563 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9794) );
  OAI21_X1 U9564 ( .B1(n7935), .B2(n8059), .A(n9794), .ZN(n7937) );
  NOR2_X1 U9565 ( .A1(n7989), .A2(n8316), .ZN(n7936) );
  AOI211_X1 U9566 ( .C1(n8057), .C2(n8313), .A(n7937), .B(n7936), .ZN(n7938)
         );
  OAI211_X1 U9567 ( .C1(n8317), .C2(n8065), .A(n7939), .B(n7938), .ZN(P2_U3155) );
  XNOR2_X1 U9568 ( .A(n7940), .B(n8193), .ZN(n7941) );
  XNOR2_X1 U9569 ( .A(n7942), .B(n7941), .ZN(n7948) );
  INV_X1 U9570 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7943) );
  OAI22_X1 U9571 ( .A1(n8208), .A2(n8045), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7943), .ZN(n7945) );
  NOR2_X1 U9572 ( .A1(n8209), .A2(n8059), .ZN(n7944) );
  AOI211_X1 U9573 ( .C1(n8212), .C2(n8062), .A(n7945), .B(n7944), .ZN(n7947)
         );
  NAND2_X1 U9574 ( .A1(n8213), .A2(n8047), .ZN(n7946) );
  OAI211_X1 U9575 ( .C1(n7948), .C2(n8050), .A(n7947), .B(n7946), .ZN(P2_U3156) );
  NAND2_X1 U9576 ( .A1(n4529), .A2(n7949), .ZN(n7950) );
  XNOR2_X1 U9577 ( .A(n7951), .B(n7950), .ZN(n7956) );
  NAND2_X1 U9578 ( .A1(n8057), .A2(n8277), .ZN(n7952) );
  NAND2_X1 U9579 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8123) );
  OAI211_X1 U9580 ( .C1(n7972), .C2(n8059), .A(n7952), .B(n8123), .ZN(n7953)
         );
  AOI21_X1 U9581 ( .B1(n8256), .B2(n8062), .A(n7953), .ZN(n7955) );
  NAND2_X1 U9582 ( .A1(n8363), .A2(n8047), .ZN(n7954) );
  OAI211_X1 U9583 ( .C1(n7956), .C2(n8050), .A(n7955), .B(n7954), .ZN(P2_U3159) );
  NOR2_X1 U9584 ( .A1(n7961), .A2(n8059), .ZN(n7965) );
  AOI22_X1 U9585 ( .A1(n7962), .A2(n8062), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7963) );
  OAI21_X1 U9586 ( .B1(n8171), .B2(n8045), .A(n7963), .ZN(n7964) );
  AOI211_X1 U9587 ( .C1(n7966), .C2(n8047), .A(n7965), .B(n7964), .ZN(n7967)
         );
  XOR2_X1 U9588 ( .A(n7969), .B(n7968), .Z(n7975) );
  AOI22_X1 U9589 ( .A1(n8233), .A2(n8042), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7971) );
  NAND2_X1 U9590 ( .A1(n8236), .A2(n8062), .ZN(n7970) );
  OAI211_X1 U9591 ( .C1(n7972), .C2(n8045), .A(n7971), .B(n7970), .ZN(n7973)
         );
  AOI21_X1 U9592 ( .B1(n8426), .B2(n8047), .A(n7973), .ZN(n7974) );
  OAI21_X1 U9593 ( .B1(n7975), .B2(n8050), .A(n7974), .ZN(P2_U3163) );
  XOR2_X1 U9594 ( .A(n7977), .B(n7976), .Z(n7983) );
  AOI22_X1 U9595 ( .A1(n8071), .A2(n8057), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7979) );
  NAND2_X1 U9596 ( .A1(n8185), .A2(n8062), .ZN(n7978) );
  OAI211_X1 U9597 ( .C1(n8183), .C2(n8059), .A(n7979), .B(n7978), .ZN(n7980)
         );
  AOI21_X1 U9598 ( .B1(n7981), .B2(n8047), .A(n7980), .ZN(n7982) );
  OAI21_X1 U9599 ( .B1(n7983), .B2(n8050), .A(n7982), .ZN(P2_U3165) );
  XNOR2_X1 U9600 ( .A(n7984), .B(n8060), .ZN(n7985) );
  XNOR2_X1 U9601 ( .A(n7986), .B(n7985), .ZN(n7992) );
  NAND2_X1 U9602 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9827) );
  OAI21_X1 U9603 ( .B1(n8059), .B2(n8284), .A(n9827), .ZN(n7987) );
  AOI21_X1 U9604 ( .B1(n8057), .B2(n8314), .A(n7987), .ZN(n7988) );
  OAI21_X1 U9605 ( .B1(n8292), .B2(n7989), .A(n7988), .ZN(n7990) );
  AOI21_X1 U9606 ( .B1(n8451), .B2(n8047), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9607 ( .B1(n7992), .B2(n8050), .A(n7991), .ZN(P2_U3166) );
  XOR2_X1 U9608 ( .A(n7994), .B(n7993), .Z(n7999) );
  AOI22_X1 U9609 ( .A1(n8042), .A2(n8277), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n7996) );
  NAND2_X1 U9610 ( .A1(n8062), .A2(n8280), .ZN(n7995) );
  OAI211_X1 U9611 ( .C1(n8060), .C2(n8045), .A(n7996), .B(n7995), .ZN(n7997)
         );
  AOI21_X1 U9612 ( .B1(n8445), .B2(n8047), .A(n7997), .ZN(n7998) );
  OAI21_X1 U9613 ( .B1(n7999), .B2(n8050), .A(n7998), .ZN(P2_U3168) );
  XOR2_X1 U9614 ( .A(n8001), .B(n8000), .Z(n8007) );
  AOI22_X1 U9615 ( .A1(n8221), .A2(n8057), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8003) );
  NAND2_X1 U9616 ( .A1(n8196), .A2(n8062), .ZN(n8002) );
  OAI211_X1 U9617 ( .C1(n8194), .C2(n8059), .A(n8003), .B(n8002), .ZN(n8004)
         );
  AOI21_X1 U9618 ( .B1(n8005), .B2(n8047), .A(n8004), .ZN(n8006) );
  OAI21_X1 U9619 ( .B1(n8007), .B2(n8050), .A(n8006), .ZN(P2_U3169) );
  XOR2_X1 U9620 ( .A(n8009), .B(n8008), .Z(n8015) );
  AOI22_X1 U9621 ( .A1(n8244), .A2(n8042), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8011) );
  NAND2_X1 U9622 ( .A1(n8062), .A2(n8240), .ZN(n8010) );
  OAI211_X1 U9623 ( .C1(n8012), .C2(n8045), .A(n8011), .B(n8010), .ZN(n8013)
         );
  AOI21_X1 U9624 ( .B1(n8432), .B2(n8047), .A(n8013), .ZN(n8014) );
  OAI21_X1 U9625 ( .B1(n8015), .B2(n8050), .A(n8014), .ZN(P2_U3173) );
  OAI21_X1 U9626 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8019) );
  NAND2_X1 U9627 ( .A1(n8019), .A2(n8052), .ZN(n8026) );
  INV_X1 U9628 ( .A(n8332), .ZN(n8024) );
  NAND2_X1 U9629 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9777) );
  INV_X1 U9630 ( .A(n9777), .ZN(n8020) );
  AOI21_X1 U9631 ( .B1(n8042), .B2(n8327), .A(n8020), .ZN(n8021) );
  OAI21_X1 U9632 ( .B1(n8022), .B2(n8045), .A(n8021), .ZN(n8023) );
  AOI21_X1 U9633 ( .B1(n8024), .B2(n8062), .A(n8023), .ZN(n8025) );
  OAI211_X1 U9634 ( .C1(n8334), .C2(n8065), .A(n8026), .B(n8025), .ZN(P2_U3174) );
  XOR2_X1 U9635 ( .A(n8028), .B(n8027), .Z(n8033) );
  AOI22_X1 U9636 ( .A1(n8244), .A2(n8057), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8030) );
  NAND2_X1 U9637 ( .A1(n8224), .A2(n8062), .ZN(n8029) );
  OAI211_X1 U9638 ( .C1(n8193), .C2(n8059), .A(n8030), .B(n8029), .ZN(n8031)
         );
  AOI21_X1 U9639 ( .B1(n8420), .B2(n8047), .A(n8031), .ZN(n8032) );
  OAI21_X1 U9640 ( .B1(n8033), .B2(n8050), .A(n8032), .ZN(P2_U3175) );
  XOR2_X1 U9641 ( .A(n8035), .B(n8034), .Z(n8040) );
  AOI22_X1 U9642 ( .A1(n8265), .A2(n8042), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8037) );
  NAND2_X1 U9643 ( .A1(n8062), .A2(n8269), .ZN(n8036) );
  OAI211_X1 U9644 ( .C1(n8284), .C2(n8045), .A(n8037), .B(n8036), .ZN(n8038)
         );
  AOI21_X1 U9645 ( .B1(n8439), .B2(n8047), .A(n8038), .ZN(n8039) );
  OAI21_X1 U9646 ( .B1(n8040), .B2(n8050), .A(n8039), .ZN(P2_U3178) );
  XNOR2_X1 U9647 ( .A(n8041), .B(n8070), .ZN(n8051) );
  NAND2_X1 U9648 ( .A1(n8069), .A2(n8042), .ZN(n8044) );
  AOI22_X1 U9649 ( .A1(n8172), .A2(n8062), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8043) );
  OAI211_X1 U9650 ( .C1(n8194), .C2(n8045), .A(n8044), .B(n8043), .ZN(n8046)
         );
  AOI21_X1 U9651 ( .B1(n8048), .B2(n8047), .A(n8046), .ZN(n8049) );
  OAI21_X1 U9652 ( .B1(n8051), .B2(n8050), .A(n8049), .ZN(P2_U3180) );
  INV_X1 U9653 ( .A(n8457), .ZN(n8066) );
  OAI211_X1 U9654 ( .C1(n8055), .C2(n8054), .A(n8053), .B(n8052), .ZN(n8064)
         );
  INV_X1 U9655 ( .A(n8056), .ZN(n8302) );
  NAND2_X1 U9656 ( .A1(n8057), .A2(n8327), .ZN(n8058) );
  NAND2_X1 U9657 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9810) );
  OAI211_X1 U9658 ( .C1(n8060), .C2(n8059), .A(n8058), .B(n9810), .ZN(n8061)
         );
  AOI21_X1 U9659 ( .B1(n8302), .B2(n8062), .A(n8061), .ZN(n8063) );
  OAI211_X1 U9660 ( .C1(n8066), .C2(n8065), .A(n8064), .B(n8063), .ZN(P2_U3181) );
  MUX2_X1 U9661 ( .A(n8067), .B(P2_DATAO_REG_30__SCAN_IN), .S(n9475), .Z(
        P2_U3521) );
  MUX2_X1 U9662 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8068), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9663 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8069), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9664 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8070), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9665 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n4799), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9666 ( .A(n8071), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9475), .Z(
        P2_U3515) );
  MUX2_X1 U9667 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8221), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9668 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8233), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9669 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8244), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9670 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8252), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9671 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8265), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9672 ( .A(n8277), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9475), .Z(
        P2_U3509) );
  INV_X1 U9673 ( .A(n8284), .ZN(n8266) );
  MUX2_X1 U9674 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8266), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9675 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8300), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9676 ( .A(n8314), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9475), .Z(
        P2_U3506) );
  MUX2_X1 U9677 ( .A(n8327), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9475), .Z(
        P2_U3505) );
  MUX2_X1 U9678 ( .A(n8313), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9475), .Z(
        P2_U3504) );
  MUX2_X1 U9679 ( .A(n8329), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9475), .Z(
        P2_U3503) );
  MUX2_X1 U9680 ( .A(n8072), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9475), .Z(
        P2_U3502) );
  MUX2_X1 U9681 ( .A(n8073), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9475), .Z(
        P2_U3501) );
  MUX2_X1 U9682 ( .A(n4657), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9475), .Z(
        P2_U3499) );
  MUX2_X1 U9683 ( .A(n8074), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9475), .Z(
        P2_U3498) );
  MUX2_X1 U9684 ( .A(n8075), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9475), .Z(
        P2_U3496) );
  MUX2_X1 U9685 ( .A(n8076), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9475), .Z(
        P2_U3495) );
  MUX2_X1 U9686 ( .A(n8077), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9475), .Z(
        P2_U3494) );
  MUX2_X1 U9687 ( .A(n8078), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9475), .Z(
        P2_U3493) );
  MUX2_X1 U9688 ( .A(n8079), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9475), .Z(
        P2_U3492) );
  MUX2_X1 U9689 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8080), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI22_X1 U9690 ( .A1(n8082), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8105), .B2(
        n8081), .ZN(n9724) );
  MUX2_X1 U9691 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8083), .S(n9713), .Z(n9723)
         );
  NOR2_X1 U9692 ( .A1(n9724), .A2(n9723), .ZN(n9722) );
  XNOR2_X1 U9693 ( .A(n9730), .B(n8084), .ZN(n9738) );
  NAND2_X1 U9694 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8129), .ZN(n8085) );
  OAI21_X1 U9695 ( .B1(n8129), .B2(P2_REG2_REG_12__SCAN_IN), .A(n8085), .ZN(
        n9757) );
  NOR2_X1 U9696 ( .A1(n9764), .A2(n8086), .ZN(n8087) );
  INV_X1 U9697 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9773) );
  XNOR2_X1 U9698 ( .A(n9764), .B(n8086), .ZN(n9774) );
  NOR2_X1 U9699 ( .A1(n9773), .A2(n9774), .ZN(n9772) );
  NAND2_X1 U9700 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8127), .ZN(n8088) );
  OAI21_X1 U9701 ( .B1(n8127), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8088), .ZN(
        n9790) );
  NOR2_X1 U9702 ( .A1(n9797), .A2(n8089), .ZN(n8090) );
  NAND2_X1 U9703 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8126), .ZN(n8091) );
  OAI21_X1 U9704 ( .B1(n8126), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8091), .ZN(
        n9823) );
  NOR2_X1 U9705 ( .A1(n9824), .A2(n9823), .ZN(n9822) );
  NOR2_X1 U9706 ( .A1(n9831), .A2(n8092), .ZN(n8093) );
  XNOR2_X1 U9707 ( .A(n9831), .B(n8092), .ZN(n9843) );
  NOR2_X1 U9708 ( .A1(n9479), .A2(n8268), .ZN(n8094) );
  AOI21_X1 U9709 ( .B1(n8268), .B2(n9479), .A(n8094), .ZN(n9482) );
  AOI21_X1 U9710 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9479), .A(n9481), .ZN(
        n8095) );
  INV_X1 U9711 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10219) );
  MUX2_X1 U9712 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n10219), .S(n8125), .Z(n8097) );
  XNOR2_X1 U9713 ( .A(n8096), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U9714 ( .A(n8097), .B(n8149), .S(n8118), .Z(n8122) );
  MUX2_X1 U9715 ( .A(n9842), .B(n8369), .S(n8118), .Z(n8117) );
  XNOR2_X1 U9716 ( .A(n8117), .B(n8146), .ZN(n9837) );
  MUX2_X1 U9717 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8118), .Z(n8098) );
  OR2_X1 U9718 ( .A1(n8098), .A2(n8126), .ZN(n8115) );
  XNOR2_X1 U9719 ( .A(n8098), .B(n9813), .ZN(n9819) );
  MUX2_X1 U9720 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8118), .Z(n8099) );
  OR2_X1 U9721 ( .A1(n8099), .A2(n4701), .ZN(n8114) );
  XNOR2_X1 U9722 ( .A(n9797), .B(n8099), .ZN(n9802) );
  MUX2_X1 U9723 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8118), .Z(n8100) );
  OR2_X1 U9724 ( .A1(n8100), .A2(n8127), .ZN(n8113) );
  XNOR2_X1 U9725 ( .A(n9780), .B(n8100), .ZN(n9786) );
  MUX2_X1 U9726 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8118), .Z(n8101) );
  OR2_X1 U9727 ( .A1(n8101), .A2(n8140), .ZN(n8112) );
  XNOR2_X1 U9728 ( .A(n8101), .B(n9764), .ZN(n9769) );
  MUX2_X1 U9729 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8118), .Z(n8102) );
  OR2_X1 U9730 ( .A1(n8102), .A2(n8129), .ZN(n8111) );
  XNOR2_X1 U9731 ( .A(n8102), .B(n9747), .ZN(n9753) );
  MUX2_X1 U9732 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8118), .Z(n8103) );
  OR2_X1 U9733 ( .A1(n8103), .A2(n8136), .ZN(n8110) );
  XNOR2_X1 U9734 ( .A(n8103), .B(n9730), .ZN(n9735) );
  MUX2_X1 U9735 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8118), .Z(n8104) );
  OR2_X1 U9736 ( .A1(n8104), .A2(n8130), .ZN(n8109) );
  XNOR2_X1 U9737 ( .A(n8104), .B(n9713), .ZN(n9715) );
  OAI22_X1 U9738 ( .A1(n8108), .A2(n8107), .B1(n8106), .B2(n8105), .ZN(n9716)
         );
  NAND2_X1 U9739 ( .A1(n9715), .A2(n9716), .ZN(n9714) );
  NAND2_X1 U9740 ( .A1(n8109), .A2(n9714), .ZN(n9734) );
  NAND2_X1 U9741 ( .A1(n9735), .A2(n9734), .ZN(n9733) );
  NAND2_X1 U9742 ( .A1(n8110), .A2(n9733), .ZN(n9752) );
  NAND2_X1 U9743 ( .A1(n9753), .A2(n9752), .ZN(n9751) );
  NAND2_X1 U9744 ( .A1(n8111), .A2(n9751), .ZN(n9768) );
  NAND2_X1 U9745 ( .A1(n9769), .A2(n9768), .ZN(n9767) );
  NAND2_X1 U9746 ( .A1(n8112), .A2(n9767), .ZN(n9785) );
  NAND2_X1 U9747 ( .A1(n9786), .A2(n9785), .ZN(n9784) );
  NAND2_X1 U9748 ( .A1(n8113), .A2(n9784), .ZN(n9801) );
  NAND2_X1 U9749 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  NAND2_X1 U9750 ( .A1(n8114), .A2(n9800), .ZN(n9818) );
  NAND2_X1 U9751 ( .A1(n9819), .A2(n9818), .ZN(n9817) );
  NAND2_X1 U9752 ( .A1(n8115), .A2(n9817), .ZN(n9836) );
  NAND2_X1 U9753 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  INV_X1 U9754 ( .A(n9835), .ZN(n8116) );
  AOI21_X1 U9755 ( .B1(n8117), .B2(n9831), .A(n8116), .ZN(n8120) );
  MUX2_X1 U9756 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8118), .Z(n8119) );
  NAND2_X1 U9757 ( .A1(n8120), .A2(n8119), .ZN(n9473) );
  NOR2_X1 U9758 ( .A1(n8120), .A2(n8119), .ZN(n9472) );
  AOI21_X1 U9759 ( .B1(n9477), .B2(n9473), .A(n9472), .ZN(n8121) );
  XOR2_X1 U9760 ( .A(n8122), .B(n8121), .Z(n8152) );
  NAND2_X1 U9761 ( .A1(n9830), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8124) );
  OAI211_X1 U9762 ( .C1(n9696), .C2(n8125), .A(n8124), .B(n8123), .ZN(n8151)
         );
  AOI22_X1 U9763 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8126), .B1(n9813), .B2(
        n10161), .ZN(n9816) );
  NAND2_X1 U9764 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8127), .ZN(n8143) );
  AOI22_X1 U9765 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8127), .B1(n9780), .B2(
        n10123), .ZN(n9783) );
  NAND2_X1 U9766 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8129), .ZN(n8139) );
  AOI22_X1 U9767 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8129), .B1(n9747), .B2(
        n8128), .ZN(n9750) );
  INV_X1 U9768 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U9769 ( .A1(n9713), .A2(n10256), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n8130), .ZN(n9718) );
  INV_X1 U9770 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8134) );
  INV_X1 U9771 ( .A(n8131), .ZN(n8132) );
  NAND2_X1 U9772 ( .A1(n8136), .A2(n8137), .ZN(n8138) );
  NAND2_X1 U9773 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n9732), .ZN(n9731) );
  NAND2_X1 U9774 ( .A1(n8140), .A2(n8141), .ZN(n8142) );
  NAND2_X1 U9775 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9766), .ZN(n9765) );
  NAND2_X1 U9776 ( .A1(n8142), .A2(n9765), .ZN(n9782) );
  NAND2_X1 U9777 ( .A1(n9783), .A2(n9782), .ZN(n9781) );
  NAND2_X1 U9778 ( .A1(n8143), .A2(n9781), .ZN(n8144) );
  NAND2_X1 U9779 ( .A1(n4701), .A2(n8144), .ZN(n8145) );
  XNOR2_X1 U9780 ( .A(n9797), .B(n8144), .ZN(n9799) );
  NAND2_X1 U9781 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9799), .ZN(n9798) );
  NAND2_X1 U9782 ( .A1(n8145), .A2(n9798), .ZN(n9815) );
  NAND2_X1 U9783 ( .A1(n9816), .A2(n9815), .ZN(n9814) );
  OAI21_X1 U9784 ( .B1(n9813), .B2(n10161), .A(n9814), .ZN(n8147) );
  NAND2_X1 U9785 ( .A1(n8146), .A2(n8147), .ZN(n8148) );
  XNOR2_X1 U9786 ( .A(n9831), .B(n8147), .ZN(n9834) );
  NAND2_X1 U9787 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n9834), .ZN(n9833) );
  NAND2_X1 U9788 ( .A1(n8148), .A2(n9833), .ZN(n9471) );
  XNOR2_X1 U9789 ( .A(n9477), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9470) );
  AOI22_X1 U9790 ( .A1(n9471), .A2(n9470), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9479), .ZN(n8150) );
  NAND2_X1 U9791 ( .A1(n8154), .A2(n8153), .ZN(n8389) );
  AOI21_X1 U9792 ( .B1(n8155), .B2(n8389), .A(n9871), .ZN(n8157) );
  AOI21_X1 U9793 ( .B1(n9871), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8157), .ZN(
        n8156) );
  OAI21_X1 U9794 ( .B1(n8391), .B2(n8176), .A(n8156), .ZN(P2_U3202) );
  INV_X1 U9795 ( .A(n8392), .ZN(n8159) );
  AOI21_X1 U9796 ( .B1(n9871), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8157), .ZN(
        n8158) );
  OAI21_X1 U9797 ( .B1(n8159), .B2(n8176), .A(n8158), .ZN(P2_U3203) );
  INV_X1 U9798 ( .A(n8160), .ZN(n8167) );
  AOI22_X1 U9799 ( .A1(n8161), .A2(n8303), .B1(n9871), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8162) );
  OAI21_X1 U9800 ( .B1(n8163), .B2(n8176), .A(n8162), .ZN(n8164) );
  AOI21_X1 U9801 ( .B1(n8165), .B2(n8260), .A(n8164), .ZN(n8166) );
  OAI21_X1 U9802 ( .B1(n8167), .B2(n9871), .A(n8166), .ZN(P2_U3206) );
  XNOR2_X1 U9803 ( .A(n8169), .B(n8168), .ZN(n8170) );
  OAI222_X1 U9804 ( .A1(n9861), .A2(n8171), .B1(n9860), .B2(n8194), .C1(n9867), 
        .C2(n8170), .ZN(n8397) );
  AOI21_X1 U9805 ( .B1(n8303), .B2(n8172), .A(n8397), .ZN(n8179) );
  XNOR2_X1 U9806 ( .A(n8174), .B(n8173), .ZN(n8345) );
  OAI22_X1 U9807 ( .A1(n8398), .A2(n8176), .B1(n8175), .B2(n8318), .ZN(n8177)
         );
  AOI21_X1 U9808 ( .B1(n8345), .B2(n8260), .A(n8177), .ZN(n8178) );
  OAI21_X1 U9809 ( .B1(n8179), .B2(n9871), .A(n8178), .ZN(P2_U3207) );
  NOR2_X1 U9810 ( .A1(n8403), .A2(n8333), .ZN(n8184) );
  AOI21_X1 U9811 ( .B1(n8186), .B2(n8181), .A(n8180), .ZN(n8182) );
  OAI222_X1 U9812 ( .A1(n9860), .A2(n8209), .B1(n9861), .B2(n8183), .C1(n9867), 
        .C2(n8182), .ZN(n8402) );
  AOI211_X1 U9813 ( .C1(n8303), .C2(n8185), .A(n8184), .B(n8402), .ZN(n8190)
         );
  XNOR2_X1 U9814 ( .A(n8187), .B(n8186), .ZN(n8404) );
  INV_X1 U9815 ( .A(n8404), .ZN(n8188) );
  AOI22_X1 U9816 ( .A1(n8188), .A2(n8260), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9871), .ZN(n8189) );
  OAI21_X1 U9817 ( .B1(n8190), .B2(n9871), .A(n8189), .ZN(P2_U3208) );
  NOR2_X1 U9818 ( .A1(n8408), .A2(n8333), .ZN(n8195) );
  XOR2_X1 U9819 ( .A(n8191), .B(n8200), .Z(n8192) );
  OAI222_X1 U9820 ( .A1(n9861), .A2(n8194), .B1(n9860), .B2(n8193), .C1(n9867), 
        .C2(n8192), .ZN(n8407) );
  AOI211_X1 U9821 ( .C1(n8303), .C2(n8196), .A(n8195), .B(n8407), .ZN(n8203)
         );
  NAND2_X1 U9822 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  XOR2_X1 U9823 ( .A(n8200), .B(n8199), .Z(n8409) );
  INV_X1 U9824 ( .A(n8409), .ZN(n8201) );
  AOI22_X1 U9825 ( .A1(n8201), .A2(n8260), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9871), .ZN(n8202) );
  OAI21_X1 U9826 ( .B1(n8203), .B2(n9871), .A(n8202), .ZN(P2_U3209) );
  XNOR2_X1 U9827 ( .A(n8204), .B(n8205), .ZN(n8415) );
  XNOR2_X1 U9828 ( .A(n8206), .B(n8205), .ZN(n8207) );
  OAI222_X1 U9829 ( .A1(n9861), .A2(n8209), .B1(n9860), .B2(n8208), .C1(n9867), 
        .C2(n8207), .ZN(n8412) );
  INV_X1 U9830 ( .A(n8412), .ZN(n8210) );
  MUX2_X1 U9831 ( .A(n8211), .B(n8210), .S(n8318), .Z(n8215) );
  AOI22_X1 U9832 ( .A1(n8213), .A2(n8304), .B1(n8303), .B2(n8212), .ZN(n8214)
         );
  OAI211_X1 U9833 ( .C1(n8415), .C2(n8339), .A(n8215), .B(n8214), .ZN(P2_U3210) );
  XNOR2_X1 U9834 ( .A(n8216), .B(n8217), .ZN(n8423) );
  INV_X1 U9835 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8223) );
  OR3_X1 U9836 ( .A1(n8228), .A2(n8218), .A3(n8217), .ZN(n8219) );
  NAND2_X1 U9837 ( .A1(n8220), .A2(n8219), .ZN(n8222) );
  AOI222_X1 U9838 ( .A1(n8331), .A2(n8222), .B1(n8244), .B2(n8328), .C1(n8221), 
        .C2(n8326), .ZN(n8418) );
  MUX2_X1 U9839 ( .A(n8223), .B(n8418), .S(n8318), .Z(n8226) );
  AOI22_X1 U9840 ( .A1(n8420), .A2(n8304), .B1(n8303), .B2(n8224), .ZN(n8225)
         );
  OAI211_X1 U9841 ( .C1(n8423), .C2(n8339), .A(n8226), .B(n8225), .ZN(P2_U3211) );
  XNOR2_X1 U9842 ( .A(n8227), .B(n4791), .ZN(n8429) );
  INV_X1 U9843 ( .A(n8228), .ZN(n8232) );
  NAND3_X1 U9844 ( .A1(n8241), .A2(n8230), .A3(n8229), .ZN(n8231) );
  NAND2_X1 U9845 ( .A1(n8232), .A2(n8231), .ZN(n8234) );
  AOI222_X1 U9846 ( .A1(n8331), .A2(n8234), .B1(n8252), .B2(n8328), .C1(n8233), 
        .C2(n8326), .ZN(n8424) );
  MUX2_X1 U9847 ( .A(n8235), .B(n8424), .S(n8318), .Z(n8238) );
  AOI22_X1 U9848 ( .A1(n8426), .A2(n8304), .B1(n8303), .B2(n8236), .ZN(n8237)
         );
  OAI211_X1 U9849 ( .C1(n8429), .C2(n8339), .A(n8238), .B(n8237), .ZN(P2_U3212) );
  XOR2_X1 U9850 ( .A(n8239), .B(n8242), .Z(n8435) );
  INV_X1 U9851 ( .A(n8240), .ZN(n8246) );
  OAI21_X1 U9852 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8245) );
  AOI222_X1 U9853 ( .A1(n8331), .A2(n8245), .B1(n8244), .B2(n8326), .C1(n8265), 
        .C2(n8328), .ZN(n8430) );
  OAI21_X1 U9854 ( .B1(n8246), .B2(n9857), .A(n8430), .ZN(n8247) );
  NAND2_X1 U9855 ( .A1(n8247), .A2(n8318), .ZN(n8249) );
  AOI22_X1 U9856 ( .A1(n8432), .A2(n8304), .B1(n9871), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n8248) );
  OAI211_X1 U9857 ( .C1(n8435), .C2(n8339), .A(n8249), .B(n8248), .ZN(P2_U3213) );
  XNOR2_X1 U9858 ( .A(n8250), .B(n8251), .ZN(n8253) );
  AOI222_X1 U9859 ( .A1(n8331), .A2(n8253), .B1(n8252), .B2(n8326), .C1(n8277), 
        .C2(n8328), .ZN(n8366) );
  XNOR2_X1 U9860 ( .A(n8255), .B(n8254), .ZN(n8364) );
  NAND2_X1 U9861 ( .A1(n8363), .A2(n8304), .ZN(n8258) );
  AOI22_X1 U9862 ( .A1(n9871), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8303), .B2(
        n8256), .ZN(n8257) );
  NAND2_X1 U9863 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  AOI21_X1 U9864 ( .B1(n8364), .B2(n8260), .A(n8259), .ZN(n8261) );
  OAI21_X1 U9865 ( .B1(n8366), .B2(n9871), .A(n8261), .ZN(P2_U3214) );
  OAI21_X1 U9866 ( .B1(n8263), .B2(n4482), .A(n8262), .ZN(n8442) );
  XNOR2_X1 U9867 ( .A(n8264), .B(n4482), .ZN(n8267) );
  AOI222_X1 U9868 ( .A1(n8331), .A2(n8267), .B1(n8266), .B2(n8328), .C1(n8265), 
        .C2(n8326), .ZN(n8437) );
  MUX2_X1 U9869 ( .A(n8268), .B(n8437), .S(n8318), .Z(n8271) );
  AOI22_X1 U9870 ( .A1(n8439), .A2(n8304), .B1(n8303), .B2(n8269), .ZN(n8270)
         );
  OAI211_X1 U9871 ( .C1(n8442), .C2(n8339), .A(n8271), .B(n8270), .ZN(P2_U3215) );
  XNOR2_X1 U9872 ( .A(n8273), .B(n8272), .ZN(n8448) );
  OAI211_X1 U9873 ( .C1(n8276), .C2(n8275), .A(n8274), .B(n8331), .ZN(n8279)
         );
  AOI22_X1 U9874 ( .A1(n8300), .A2(n8328), .B1(n8277), .B2(n8326), .ZN(n8278)
         );
  AND2_X1 U9875 ( .A1(n8279), .A2(n8278), .ZN(n8444) );
  MUX2_X1 U9876 ( .A(n8444), .B(n9842), .S(n9871), .Z(n8282) );
  AOI22_X1 U9877 ( .A1(n8445), .A2(n8304), .B1(n8303), .B2(n8280), .ZN(n8281)
         );
  OAI211_X1 U9878 ( .C1(n8448), .C2(n8339), .A(n8282), .B(n8281), .ZN(P2_U3216) );
  XNOR2_X1 U9879 ( .A(n8283), .B(n8288), .ZN(n8454) );
  NOR2_X1 U9880 ( .A1(n8284), .A2(n9861), .ZN(n8290) );
  INV_X1 U9881 ( .A(n8285), .ZN(n8286) );
  AOI211_X1 U9882 ( .C1(n8288), .C2(n8287), .A(n9867), .B(n8286), .ZN(n8289)
         );
  AOI211_X1 U9883 ( .C1(n8328), .C2(n8314), .A(n8290), .B(n8289), .ZN(n8449)
         );
  MUX2_X1 U9884 ( .A(n8291), .B(n8449), .S(n8318), .Z(n8295) );
  INV_X1 U9885 ( .A(n8292), .ZN(n8293) );
  AOI22_X1 U9886 ( .A1(n8451), .A2(n8304), .B1(n8303), .B2(n8293), .ZN(n8294)
         );
  OAI211_X1 U9887 ( .C1(n8454), .C2(n8339), .A(n8295), .B(n8294), .ZN(P2_U3217) );
  XNOR2_X1 U9888 ( .A(n8297), .B(n8296), .ZN(n8460) );
  XNOR2_X1 U9889 ( .A(n8299), .B(n8298), .ZN(n8301) );
  AOI222_X1 U9890 ( .A1(n8331), .A2(n8301), .B1(n8300), .B2(n8326), .C1(n8327), 
        .C2(n8328), .ZN(n8455) );
  MUX2_X1 U9891 ( .A(n9806), .B(n8455), .S(n8318), .Z(n8306) );
  AOI22_X1 U9892 ( .A1(n8457), .A2(n8304), .B1(n8303), .B2(n8302), .ZN(n8305)
         );
  OAI211_X1 U9893 ( .C1(n8460), .C2(n8339), .A(n8306), .B(n8305), .ZN(P2_U3218) );
  XOR2_X1 U9894 ( .A(n8311), .B(n8307), .Z(n8465) );
  OR2_X1 U9895 ( .A1(n8325), .A2(n8308), .ZN(n8310) );
  NAND2_X1 U9896 ( .A1(n8310), .A2(n8309), .ZN(n8312) );
  XNOR2_X1 U9897 ( .A(n8312), .B(n8311), .ZN(n8315) );
  AOI222_X1 U9898 ( .A1(n8331), .A2(n8315), .B1(n8314), .B2(n8326), .C1(n8313), 
        .C2(n8328), .ZN(n8461) );
  INV_X1 U9899 ( .A(n8461), .ZN(n8320) );
  OAI22_X1 U9900 ( .A1(n8317), .A2(n8333), .B1(n8316), .B2(n9857), .ZN(n8319)
         );
  OAI21_X1 U9901 ( .B1(n8320), .B2(n8319), .A(n8318), .ZN(n8322) );
  NAND2_X1 U9902 ( .A1(n9871), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8321) );
  OAI211_X1 U9903 ( .C1(n8465), .C2(n8339), .A(n8322), .B(n8321), .ZN(P2_U3219) );
  XNOR2_X1 U9904 ( .A(n8323), .B(n8324), .ZN(n8471) );
  XNOR2_X1 U9905 ( .A(n8325), .B(n8324), .ZN(n8330) );
  AOI222_X1 U9906 ( .A1(n8331), .A2(n8330), .B1(n8329), .B2(n8328), .C1(n8327), 
        .C2(n8326), .ZN(n8466) );
  INV_X1 U9907 ( .A(n8466), .ZN(n8336) );
  OAI22_X1 U9908 ( .A1(n8334), .A2(n8333), .B1(n8332), .B2(n9857), .ZN(n8335)
         );
  OAI21_X1 U9909 ( .B1(n8336), .B2(n8335), .A(n8318), .ZN(n8338) );
  NAND2_X1 U9910 ( .A1(n9871), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8337) );
  OAI211_X1 U9911 ( .C1(n8471), .C2(n8339), .A(n8338), .B(n8337), .ZN(P2_U3220) );
  NOR2_X1 U9912 ( .A1(n8389), .A2(n9927), .ZN(n8341) );
  AOI21_X1 U9913 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9927), .A(n8341), .ZN(
        n8340) );
  OAI21_X1 U9914 ( .B1(n8391), .B2(n8352), .A(n8340), .ZN(P2_U3490) );
  INV_X1 U9915 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U9916 ( .A1(n8392), .A2(n6603), .ZN(n8343) );
  INV_X1 U9917 ( .A(n8341), .ZN(n8342) );
  OAI211_X1 U9918 ( .C1(n8378), .C2(n8344), .A(n8343), .B(n8342), .ZN(P2_U3489) );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8397), .S(n8378), .Z(n8347)
         );
  INV_X1 U9920 ( .A(n8345), .ZN(n8399) );
  OAI22_X1 U9921 ( .A1(n8399), .A2(n8381), .B1(n8398), .B2(n8352), .ZN(n8346)
         );
  MUX2_X1 U9922 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8402), .S(n8378), .Z(n8349)
         );
  OAI22_X1 U9923 ( .A1(n8404), .A2(n8381), .B1(n8403), .B2(n8352), .ZN(n8348)
         );
  OR2_X1 U9924 ( .A1(n8349), .A2(n8348), .ZN(P2_U3484) );
  MUX2_X1 U9925 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8407), .S(n9929), .Z(n8351)
         );
  OAI22_X1 U9926 ( .A1(n8409), .A2(n8381), .B1(n8408), .B2(n8352), .ZN(n8350)
         );
  OR2_X1 U9927 ( .A1(n8351), .A2(n8350), .ZN(P2_U3483) );
  MUX2_X1 U9928 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8412), .S(n8378), .Z(n8354)
         );
  OAI22_X1 U9929 ( .A1(n8415), .A2(n8381), .B1(n8414), .B2(n8352), .ZN(n8353)
         );
  OR2_X1 U9930 ( .A1(n8354), .A2(n8353), .ZN(P2_U3482) );
  MUX2_X1 U9931 ( .A(n10124), .B(n8418), .S(n9929), .Z(n8356) );
  NAND2_X1 U9932 ( .A1(n8420), .A2(n6603), .ZN(n8355) );
  OAI211_X1 U9933 ( .C1(n8381), .C2(n8423), .A(n8356), .B(n8355), .ZN(P2_U3481) );
  INV_X1 U9934 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8357) );
  MUX2_X1 U9935 ( .A(n8357), .B(n8424), .S(n9929), .Z(n8359) );
  NAND2_X1 U9936 ( .A1(n8426), .A2(n6603), .ZN(n8358) );
  OAI211_X1 U9937 ( .C1(n8381), .C2(n8429), .A(n8359), .B(n8358), .ZN(P2_U3480) );
  INV_X1 U9938 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8360) );
  MUX2_X1 U9939 ( .A(n8360), .B(n8430), .S(n8378), .Z(n8362) );
  NAND2_X1 U9940 ( .A1(n8432), .A2(n6603), .ZN(n8361) );
  OAI211_X1 U9941 ( .C1(n8435), .C2(n8381), .A(n8362), .B(n8361), .ZN(P2_U3479) );
  AOI22_X1 U9942 ( .A1(n8364), .A2(n9914), .B1(n9907), .B2(n8363), .ZN(n8365)
         );
  NAND2_X1 U9943 ( .A1(n8366), .A2(n8365), .ZN(n8436) );
  MUX2_X1 U9944 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8436), .S(n8378), .Z(
        P2_U3478) );
  MUX2_X1 U9945 ( .A(n10228), .B(n8437), .S(n8378), .Z(n8368) );
  NAND2_X1 U9946 ( .A1(n8439), .A2(n6603), .ZN(n8367) );
  OAI211_X1 U9947 ( .C1(n8381), .C2(n8442), .A(n8368), .B(n8367), .ZN(P2_U3477) );
  MUX2_X1 U9948 ( .A(n8369), .B(n8444), .S(n8378), .Z(n8371) );
  NAND2_X1 U9949 ( .A1(n8445), .A2(n6603), .ZN(n8370) );
  OAI211_X1 U9950 ( .C1(n8448), .C2(n8381), .A(n8371), .B(n8370), .ZN(P2_U3476) );
  MUX2_X1 U9951 ( .A(n10161), .B(n8449), .S(n9929), .Z(n8373) );
  NAND2_X1 U9952 ( .A1(n8451), .A2(n6603), .ZN(n8372) );
  OAI211_X1 U9953 ( .C1(n8454), .C2(n8381), .A(n8373), .B(n8372), .ZN(P2_U3475) );
  MUX2_X1 U9954 ( .A(n10060), .B(n8455), .S(n8378), .Z(n8375) );
  NAND2_X1 U9955 ( .A1(n8457), .A2(n6603), .ZN(n8374) );
  OAI211_X1 U9956 ( .C1(n8381), .C2(n8460), .A(n8375), .B(n8374), .ZN(P2_U3474) );
  MUX2_X1 U9957 ( .A(n10123), .B(n8461), .S(n9929), .Z(n8377) );
  NAND2_X1 U9958 ( .A1(n8462), .A2(n6603), .ZN(n8376) );
  OAI211_X1 U9959 ( .C1(n8465), .C2(n8381), .A(n8377), .B(n8376), .ZN(P2_U3473) );
  MUX2_X1 U9960 ( .A(n10242), .B(n8466), .S(n8378), .Z(n8380) );
  NAND2_X1 U9961 ( .A1(n8467), .A2(n6603), .ZN(n8379) );
  OAI211_X1 U9962 ( .C1(n8381), .C2(n8471), .A(n8380), .B(n8379), .ZN(P2_U3472) );
  INV_X1 U9963 ( .A(n8382), .ZN(n8387) );
  NAND3_X1 U9964 ( .A1(n8384), .A2(n8383), .A3(n9914), .ZN(n8385) );
  OAI211_X1 U9965 ( .C1(n8387), .C2(n9909), .A(n8386), .B(n8385), .ZN(n8472)
         );
  MUX2_X1 U9966 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8472), .S(n9929), .Z(
        P2_U3471) );
  MUX2_X1 U9967 ( .A(n8388), .B(P2_REG1_REG_0__SCAN_IN), .S(n9927), .Z(
        P2_U3459) );
  NOR2_X1 U9968 ( .A1(n8389), .A2(n9917), .ZN(n8393) );
  AOI21_X1 U9969 ( .B1(n9917), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8393), .ZN(
        n8390) );
  OAI21_X1 U9970 ( .B1(n8391), .B2(n8413), .A(n8390), .ZN(P2_U3458) );
  INV_X1 U9971 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U9972 ( .A1(n8392), .A2(n6608), .ZN(n8395) );
  INV_X1 U9973 ( .A(n8393), .ZN(n8394) );
  OAI211_X1 U9974 ( .C1(n8396), .C2(n9915), .A(n8395), .B(n8394), .ZN(P2_U3457) );
  MUX2_X1 U9975 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8397), .S(n9915), .Z(n8401)
         );
  OAI22_X1 U9976 ( .A1(n8399), .A2(n8470), .B1(n8398), .B2(n8413), .ZN(n8400)
         );
  MUX2_X1 U9977 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8402), .S(n9915), .Z(n8406)
         );
  OAI22_X1 U9978 ( .A1(n8404), .A2(n8470), .B1(n8403), .B2(n8413), .ZN(n8405)
         );
  OR2_X1 U9979 ( .A1(n8406), .A2(n8405), .ZN(P2_U3452) );
  MUX2_X1 U9980 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8407), .S(n9915), .Z(n8411)
         );
  OAI22_X1 U9981 ( .A1(n8409), .A2(n8470), .B1(n8408), .B2(n8413), .ZN(n8410)
         );
  OR2_X1 U9982 ( .A1(n8411), .A2(n8410), .ZN(P2_U3451) );
  MUX2_X1 U9983 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8412), .S(n9915), .Z(n8417)
         );
  OAI22_X1 U9984 ( .A1(n8415), .A2(n8470), .B1(n8414), .B2(n8413), .ZN(n8416)
         );
  OR2_X1 U9985 ( .A1(n8417), .A2(n8416), .ZN(P2_U3450) );
  INV_X1 U9986 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8419) );
  MUX2_X1 U9987 ( .A(n8419), .B(n8418), .S(n9915), .Z(n8422) );
  NAND2_X1 U9988 ( .A1(n8420), .A2(n6608), .ZN(n8421) );
  OAI211_X1 U9989 ( .C1(n8423), .C2(n8470), .A(n8422), .B(n8421), .ZN(P2_U3449) );
  INV_X1 U9990 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8425) );
  MUX2_X1 U9991 ( .A(n8425), .B(n8424), .S(n9915), .Z(n8428) );
  NAND2_X1 U9992 ( .A1(n8426), .A2(n6608), .ZN(n8427) );
  OAI211_X1 U9993 ( .C1(n8429), .C2(n8470), .A(n8428), .B(n8427), .ZN(P2_U3448) );
  INV_X1 U9994 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8431) );
  MUX2_X1 U9995 ( .A(n8431), .B(n8430), .S(n9915), .Z(n8434) );
  NAND2_X1 U9996 ( .A1(n8432), .A2(n6608), .ZN(n8433) );
  OAI211_X1 U9997 ( .C1(n8435), .C2(n8470), .A(n8434), .B(n8433), .ZN(P2_U3447) );
  MUX2_X1 U9998 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8436), .S(n9915), .Z(
        P2_U3446) );
  INV_X1 U9999 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8438) );
  MUX2_X1 U10000 ( .A(n8438), .B(n8437), .S(n9915), .Z(n8441) );
  NAND2_X1 U10001 ( .A1(n8439), .A2(n6608), .ZN(n8440) );
  OAI211_X1 U10002 ( .C1(n8442), .C2(n8470), .A(n8441), .B(n8440), .ZN(
        P2_U3444) );
  MUX2_X1 U10003 ( .A(n8444), .B(n8443), .S(n9917), .Z(n8447) );
  NAND2_X1 U10004 ( .A1(n8445), .A2(n6608), .ZN(n8446) );
  OAI211_X1 U10005 ( .C1(n8448), .C2(n8470), .A(n8447), .B(n8446), .ZN(
        P2_U3441) );
  INV_X1 U10006 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8450) );
  MUX2_X1 U10007 ( .A(n8450), .B(n8449), .S(n9915), .Z(n8453) );
  NAND2_X1 U10008 ( .A1(n8451), .A2(n6608), .ZN(n8452) );
  OAI211_X1 U10009 ( .C1(n8454), .C2(n8470), .A(n8453), .B(n8452), .ZN(
        P2_U3438) );
  INV_X1 U10010 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8456) );
  MUX2_X1 U10011 ( .A(n8456), .B(n8455), .S(n9915), .Z(n8459) );
  NAND2_X1 U10012 ( .A1(n8457), .A2(n6608), .ZN(n8458) );
  OAI211_X1 U10013 ( .C1(n8460), .C2(n8470), .A(n8459), .B(n8458), .ZN(
        P2_U3435) );
  MUX2_X1 U10014 ( .A(n10169), .B(n8461), .S(n9915), .Z(n8464) );
  NAND2_X1 U10015 ( .A1(n8462), .A2(n6608), .ZN(n8463) );
  OAI211_X1 U10016 ( .C1(n8465), .C2(n8470), .A(n8464), .B(n8463), .ZN(
        P2_U3432) );
  MUX2_X1 U10017 ( .A(n10217), .B(n8466), .S(n9915), .Z(n8469) );
  NAND2_X1 U10018 ( .A1(n8467), .A2(n6608), .ZN(n8468) );
  OAI211_X1 U10019 ( .C1(n8471), .C2(n8470), .A(n8469), .B(n8468), .ZN(
        P2_U3429) );
  MUX2_X1 U10020 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8472), .S(n9915), .Z(
        P2_U3426) );
  INV_X1 U10021 ( .A(n8760), .ZN(n9456) );
  NOR4_X1 U10022 ( .A1(n8474), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8473), .ZN(n8475) );
  AOI21_X1 U10023 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n8489), .A(n8475), .ZN(
        n8476) );
  OAI21_X1 U10024 ( .B1(n9456), .B2(n6677), .A(n8476), .ZN(P2_U3264) );
  INV_X1 U10025 ( .A(n8755), .ZN(n9458) );
  AOI22_X1 U10026 ( .A1(n8477), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8489), .ZN(n8478) );
  OAI21_X1 U10027 ( .B1(n9458), .B2(n6677), .A(n8478), .ZN(P2_U3265) );
  OAI222_X1 U10028 ( .A1(n8483), .A2(n8482), .B1(P2_U3151), .B2(n8479), .C1(
        n10095), .C2(n8480), .ZN(P2_U3266) );
  INV_X1 U10029 ( .A(n8484), .ZN(n9461) );
  AOI21_X1 U10030 ( .B1(n8489), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8485), .ZN(
        n8486) );
  OAI21_X1 U10031 ( .B1(n9461), .B2(n6677), .A(n8486), .ZN(P2_U3267) );
  INV_X1 U10032 ( .A(n8487), .ZN(n9465) );
  AOI21_X1 U10033 ( .B1(n8489), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8488), .ZN(
        n8490) );
  OAI21_X1 U10034 ( .B1(n9465), .B2(n6677), .A(n8490), .ZN(P2_U3268) );
  MUX2_X1 U10035 ( .A(n8491), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10036 ( .A1(n8493), .A2(n8492), .ZN(n8494) );
  XOR2_X1 U10037 ( .A(n8495), .B(n8494), .Z(n8503) );
  OAI22_X1 U10038 ( .A1(n8497), .A2(n9489), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8496), .ZN(n8500) );
  NOR2_X1 U10039 ( .A1(n8498), .A2(n8651), .ZN(n8499) );
  AOI211_X1 U10040 ( .C1(n8501), .C2(n8656), .A(n8500), .B(n8499), .ZN(n8502)
         );
  OAI21_X1 U10041 ( .B1(n8503), .B2(n9493), .A(n8502), .ZN(P1_U3215) );
  AOI21_X1 U10042 ( .B1(n8505), .B2(n8507), .A(n8504), .ZN(n8506) );
  AOI21_X1 U10043 ( .B1(n4491), .B2(n8507), .A(n8506), .ZN(n8513) );
  NOR2_X1 U10044 ( .A1(n9044), .A2(n8508), .ZN(n8509) );
  AOI21_X1 U10045 ( .B1(n9048), .B2(n9012), .A(n8509), .ZN(n9177) );
  AOI22_X1 U10046 ( .A1(n9171), .A2(n8656), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        n4437), .ZN(n8510) );
  OAI21_X1 U10047 ( .B1(n9177), .B2(n9489), .A(n8510), .ZN(n8511) );
  AOI21_X1 U10048 ( .B1(n9332), .B2(n9497), .A(n8511), .ZN(n8512) );
  OAI21_X1 U10049 ( .B1(n8513), .B2(n9493), .A(n8512), .ZN(P1_U3216) );
  OAI21_X1 U10050 ( .B1(n8516), .B2(n8515), .A(n8514), .ZN(n8517) );
  NAND2_X1 U10051 ( .A1(n8517), .A2(n8634), .ZN(n8522) );
  AOI22_X1 U10052 ( .A1(n8519), .A2(n8636), .B1(n8518), .B2(n9497), .ZN(n8521)
         );
  MUX2_X1 U10053 ( .A(n9501), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n8520) );
  NAND3_X1 U10054 ( .A1(n8522), .A2(n8521), .A3(n8520), .ZN(P1_U3218) );
  XNOR2_X1 U10055 ( .A(n8523), .B(n8535), .ZN(n8621) );
  OAI22_X1 U10056 ( .A1(n8621), .A2(n8536), .B1(n8523), .B2(n8535), .ZN(n8527)
         );
  OR2_X1 U10057 ( .A1(n8525), .A2(n8524), .ZN(n8534) );
  NAND2_X1 U10058 ( .A1(n8540), .A2(n8534), .ZN(n8526) );
  XNOR2_X1 U10059 ( .A(n8527), .B(n8526), .ZN(n8533) );
  NOR2_X1 U10060 ( .A1(n9501), .A2(n9237), .ZN(n8531) );
  AND2_X1 U10061 ( .A1(n9029), .A2(n8595), .ZN(n8528) );
  AOI21_X1 U10062 ( .B1(n9038), .B2(n9012), .A(n8528), .ZN(n9230) );
  OAI22_X1 U10063 ( .A1(n9230), .A2(n9489), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8529), .ZN(n8530) );
  AOI211_X1 U10064 ( .C1(n9429), .C2(n9497), .A(n8531), .B(n8530), .ZN(n8532)
         );
  OAI21_X1 U10065 ( .B1(n8533), .B2(n9493), .A(n8532), .ZN(P1_U3219) );
  INV_X1 U10066 ( .A(n8523), .ZN(n8539) );
  INV_X1 U10067 ( .A(n8534), .ZN(n8538) );
  AOI21_X1 U10068 ( .B1(n8523), .B2(n8536), .A(n8535), .ZN(n8537) );
  AOI211_X1 U10069 ( .C1(n8620), .C2(n8539), .A(n8538), .B(n8537), .ZN(n8591)
         );
  INV_X1 U10070 ( .A(n8540), .ZN(n8590) );
  NAND2_X1 U10071 ( .A1(n8541), .A2(n8542), .ZN(n8594) );
  NOR3_X1 U10072 ( .A1(n8591), .A2(n8590), .A3(n8594), .ZN(n8592) );
  INV_X1 U10073 ( .A(n8542), .ZN(n8544) );
  NOR3_X1 U10074 ( .A1(n8592), .A2(n8544), .A3(n8543), .ZN(n8547) );
  INV_X1 U10075 ( .A(n8545), .ZN(n8546) );
  OAI21_X1 U10076 ( .B1(n8547), .B2(n8546), .A(n8634), .ZN(n8554) );
  OR2_X1 U10077 ( .A1(n9044), .A2(n8548), .ZN(n8550) );
  NAND2_X1 U10078 ( .A1(n9038), .A2(n8595), .ZN(n8549) );
  NAND2_X1 U10079 ( .A1(n8550), .A2(n8549), .ZN(n9202) );
  INV_X1 U10080 ( .A(n9206), .ZN(n8551) );
  INV_X1 U10081 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10078) );
  OAI22_X1 U10082 ( .A1(n8551), .A2(n9501), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10078), .ZN(n8552) );
  AOI21_X1 U10083 ( .B1(n9202), .B2(n8636), .A(n8552), .ZN(n8553) );
  OAI211_X1 U10084 ( .C1(n5019), .C2(n8651), .A(n8554), .B(n8553), .ZN(
        P1_U3223) );
  XNOR2_X1 U10085 ( .A(n8555), .B(n8556), .ZN(n8557) );
  NAND2_X1 U10086 ( .A1(n8557), .A2(n8634), .ZN(n8562) );
  NAND2_X1 U10087 ( .A1(n8922), .A2(n9012), .ZN(n8559) );
  NAND2_X1 U10088 ( .A1(n9048), .A2(n8595), .ZN(n8558) );
  NAND2_X1 U10089 ( .A1(n8559), .A2(n8558), .ZN(n9141) );
  INV_X1 U10090 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10129) );
  OAI22_X1 U10091 ( .A1(n9146), .A2(n9501), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10129), .ZN(n8560) );
  AOI21_X1 U10092 ( .B1(n9141), .B2(n8636), .A(n8560), .ZN(n8561) );
  OAI211_X1 U10093 ( .C1(n9144), .C2(n8651), .A(n8562), .B(n8561), .ZN(
        P1_U3225) );
  INV_X1 U10094 ( .A(n9370), .ZN(n9291) );
  OAI21_X1 U10095 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8566) );
  NAND2_X1 U10096 ( .A1(n8566), .A2(n8634), .ZN(n8571) );
  AND2_X1 U10097 ( .A1(n4437), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U10098 ( .A1(n9028), .A2(n9012), .ZN(n8568) );
  NAND2_X1 U10099 ( .A1(n9023), .A2(n8595), .ZN(n8567) );
  AND2_X1 U10100 ( .A1(n8568), .A2(n8567), .ZN(n9282) );
  NOR2_X1 U10101 ( .A1(n9282), .A2(n9489), .ZN(n8569) );
  AOI211_X1 U10102 ( .C1(n9288), .C2(n8656), .A(n9546), .B(n8569), .ZN(n8570)
         );
  OAI211_X1 U10103 ( .C1(n9291), .C2(n8651), .A(n8571), .B(n8570), .ZN(
        P1_U3226) );
  INV_X1 U10104 ( .A(n9267), .ZN(n9445) );
  AND2_X1 U10105 ( .A1(n8563), .A2(n8572), .ZN(n8575) );
  OAI211_X1 U10106 ( .C1(n8575), .C2(n8574), .A(n8634), .B(n8573), .ZN(n8579)
         );
  INV_X1 U10107 ( .A(n8576), .ZN(n9268) );
  AOI22_X1 U10108 ( .A1(n9029), .A2(n9012), .B1(n8595), .B2(n9027), .ZN(n9263)
         );
  NAND2_X1 U10109 ( .A1(n4437), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9567) );
  OAI21_X1 U10110 ( .B1(n9263), .B2(n9489), .A(n9567), .ZN(n8577) );
  AOI21_X1 U10111 ( .B1(n9268), .B2(n8656), .A(n8577), .ZN(n8578) );
  OAI211_X1 U10112 ( .C1(n9445), .C2(n8651), .A(n8579), .B(n8578), .ZN(
        P1_U3228) );
  OAI21_X1 U10113 ( .B1(n8582), .B2(n8581), .A(n8580), .ZN(n8583) );
  NAND2_X1 U10114 ( .A1(n8583), .A2(n8634), .ZN(n8589) );
  NAND2_X1 U10115 ( .A1(n9052), .A2(n9012), .ZN(n8585) );
  NAND2_X1 U10116 ( .A1(n9045), .A2(n8595), .ZN(n8584) );
  NAND2_X1 U10117 ( .A1(n8585), .A2(n8584), .ZN(n9157) );
  INV_X1 U10118 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8586) );
  OAI22_X1 U10119 ( .A1(n9161), .A2(n9501), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8586), .ZN(n8587) );
  AOI21_X1 U10120 ( .B1(n9157), .B2(n8636), .A(n8587), .ZN(n8588) );
  OAI211_X1 U10121 ( .C1(n9165), .C2(n8651), .A(n8589), .B(n8588), .ZN(
        P1_U3229) );
  OR2_X1 U10122 ( .A1(n8591), .A2(n8590), .ZN(n8593) );
  AOI21_X1 U10123 ( .B1(n8594), .B2(n8593), .A(n8592), .ZN(n8601) );
  NAND2_X1 U10124 ( .A1(n9042), .A2(n9012), .ZN(n8597) );
  NAND2_X1 U10125 ( .A1(n9032), .A2(n8595), .ZN(n8596) );
  NAND2_X1 U10126 ( .A1(n8597), .A2(n8596), .ZN(n9218) );
  AOI22_X1 U10127 ( .A1(n9218), .A2(n8636), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        n4437), .ZN(n8598) );
  OAI21_X1 U10128 ( .B1(n9501), .B2(n9221), .A(n8598), .ZN(n8599) );
  AOI21_X1 U10129 ( .B1(n9348), .B2(n9497), .A(n8599), .ZN(n8600) );
  OAI21_X1 U10130 ( .B1(n8601), .B2(n9493), .A(n8600), .ZN(P1_U3233) );
  INV_X1 U10131 ( .A(n8602), .ZN(n8606) );
  NOR3_X1 U10132 ( .A1(n4526), .A2(n8604), .A3(n8603), .ZN(n8605) );
  OAI21_X1 U10133 ( .B1(n8606), .B2(n8605), .A(n8634), .ZN(n8611) );
  NAND2_X1 U10134 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9511) );
  OAI21_X1 U10135 ( .B1(n8607), .B2(n9489), .A(n9511), .ZN(n8608) );
  AOI21_X1 U10136 ( .B1(n8609), .B2(n8656), .A(n8608), .ZN(n8610) );
  OAI211_X1 U10137 ( .C1(n8612), .C2(n8651), .A(n8611), .B(n8610), .ZN(
        P1_U3234) );
  AOI21_X1 U10138 ( .B1(n8614), .B2(n8613), .A(n4490), .ZN(n8619) );
  AND2_X1 U10139 ( .A1(n9042), .A2(n8595), .ZN(n8615) );
  AOI21_X1 U10140 ( .B1(n9045), .B2(n9012), .A(n8615), .ZN(n9188) );
  AOI22_X1 U10141 ( .A1(n9193), .A2(n8656), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8616) );
  OAI21_X1 U10142 ( .B1(n9188), .B2(n9489), .A(n8616), .ZN(n8617) );
  AOI21_X1 U10143 ( .B1(n4671), .B2(n9497), .A(n8617), .ZN(n8618) );
  OAI21_X1 U10144 ( .B1(n8619), .B2(n9493), .A(n8618), .ZN(P1_U3235) );
  XNOR2_X1 U10145 ( .A(n8621), .B(n8620), .ZN(n8626) );
  NOR2_X1 U10146 ( .A1(n9501), .A2(n9252), .ZN(n8624) );
  AOI22_X1 U10147 ( .A1(n9032), .A2(n9012), .B1(n8595), .B2(n9028), .ZN(n9250)
         );
  OAI22_X1 U10148 ( .A1(n9250), .A2(n9489), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8622), .ZN(n8623) );
  AOI211_X1 U10149 ( .C1(n9358), .C2(n9497), .A(n8624), .B(n8623), .ZN(n8625)
         );
  OAI21_X1 U10150 ( .B1(n8626), .B2(n9493), .A(n8625), .ZN(P1_U3238) );
  INV_X1 U10151 ( .A(n8627), .ZN(n8628) );
  NOR2_X1 U10152 ( .A1(n8629), .A2(n8628), .ZN(n8633) );
  NAND2_X1 U10153 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  XNOR2_X1 U10154 ( .A(n8633), .B(n8632), .ZN(n8635) );
  NAND2_X1 U10155 ( .A1(n8635), .A2(n8634), .ZN(n8642) );
  AOI22_X1 U10156 ( .A1(n8637), .A2(n8636), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n8641) );
  NAND2_X1 U10157 ( .A1(n8674), .A2(n9497), .ZN(n8640) );
  NAND2_X1 U10158 ( .A1(n8656), .A2(n8638), .ZN(n8639) );
  NAND4_X1 U10159 ( .A1(n8642), .A2(n8641), .A3(n8640), .A4(n8639), .ZN(
        P1_U3239) );
  AOI21_X1 U10160 ( .B1(n8643), .B2(n8644), .A(n9493), .ZN(n8646) );
  NAND2_X1 U10161 ( .A1(n8646), .A2(n8645), .ZN(n8650) );
  NOR2_X1 U10162 ( .A1(n9123), .A2(n9501), .ZN(n8648) );
  AOI22_X1 U10163 ( .A1(n8921), .A2(n9012), .B1(n8595), .B2(n9052), .ZN(n9129)
         );
  NOR2_X1 U10164 ( .A1(n9129), .A2(n9489), .ZN(n8647) );
  AOI211_X1 U10165 ( .C1(P1_REG3_REG_26__SCAN_IN), .C2(P1_U3086), .A(n8648), 
        .B(n8647), .ZN(n8649) );
  OAI211_X1 U10166 ( .C1(n9126), .C2(n8651), .A(n8650), .B(n8649), .ZN(
        P1_U3240) );
  NOR2_X1 U10167 ( .A1(n8654), .A2(n8653), .ZN(n8652) );
  AOI21_X1 U10168 ( .B1(n8654), .B2(n8653), .A(n8652), .ZN(n8661) );
  NAND2_X1 U10169 ( .A1(n8656), .A2(n8655), .ZN(n8657) );
  NAND2_X1 U10170 ( .A1(n4437), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9538) );
  OAI211_X1 U10171 ( .C1(n8658), .C2(n9489), .A(n8657), .B(n9538), .ZN(n8659)
         );
  AOI21_X1 U10172 ( .B1(n9024), .B2(n9497), .A(n8659), .ZN(n8660) );
  OAI21_X1 U10173 ( .B1(n8661), .B2(n9493), .A(n8660), .ZN(P1_U3241) );
  INV_X1 U10174 ( .A(n9027), .ZN(n8694) );
  INV_X1 U10175 ( .A(n8770), .ZN(n8758) );
  NOR4_X1 U10176 ( .A1(n8669), .A2(n8668), .A3(n8770), .A4(n8933), .ZN(n8680)
         );
  NOR4_X1 U10177 ( .A1(n8789), .A2(n8671), .A3(n8758), .A4(n8670), .ZN(n8679)
         );
  AOI21_X1 U10178 ( .B1(n8673), .B2(n8758), .A(n8672), .ZN(n8676) );
  AOI21_X1 U10179 ( .B1(n8770), .B2(n8932), .A(n8674), .ZN(n8675) );
  NOR2_X1 U10180 ( .A1(n8676), .A2(n8675), .ZN(n8678) );
  NOR4_X1 U10181 ( .A1(n8680), .A2(n8679), .A3(n8678), .A4(n8677), .ZN(n8681)
         );
  NAND2_X1 U10182 ( .A1(n8699), .A2(n8687), .ZN(n8690) );
  AND2_X1 U10183 ( .A1(n8701), .A2(n8688), .ZN(n8865) );
  INV_X1 U10184 ( .A(n8865), .ZN(n8689) );
  AOI21_X1 U10185 ( .B1(n8690), .B2(n8861), .A(n8689), .ZN(n8691) );
  NAND2_X1 U10186 ( .A1(n8704), .A2(n8700), .ZN(n8864) );
  OAI21_X1 U10187 ( .B1(n8691), .B2(n8864), .A(n8867), .ZN(n8692) );
  AOI211_X1 U10188 ( .C1(n8692), .C2(n8870), .A(n8797), .B(n4722), .ZN(n8696)
         );
  OR2_X1 U10189 ( .A1(n9375), .A2(n8693), .ZN(n8869) );
  NAND3_X1 U10190 ( .A1(n8876), .A2(n8770), .A3(n8869), .ZN(n8695) );
  NAND2_X1 U10191 ( .A1(n9370), .A2(n8694), .ZN(n8878) );
  AOI21_X1 U10192 ( .B1(n8878), .B2(n9023), .A(n8770), .ZN(n8710) );
  OAI22_X1 U10193 ( .A1(n8696), .A2(n8695), .B1(n8710), .B2(n8708), .ZN(n8713)
         );
  AOI21_X1 U10194 ( .B1(n8699), .B2(n8698), .A(n8697), .ZN(n8703) );
  NAND2_X1 U10195 ( .A1(n8700), .A2(n8861), .ZN(n8702) );
  OAI211_X1 U10196 ( .C1(n8703), .C2(n8702), .A(n8867), .B(n8701), .ZN(n8705)
         );
  NAND2_X1 U10197 ( .A1(n8706), .A2(n8870), .ZN(n8709) );
  AND2_X1 U10198 ( .A1(n8708), .A2(n8707), .ZN(n8874) );
  INV_X1 U10199 ( .A(n8878), .ZN(n8711) );
  AOI21_X1 U10200 ( .B1(n8877), .B2(n8713), .A(n8712), .ZN(n8716) );
  INV_X1 U10201 ( .A(n9028), .ZN(n8714) );
  NAND2_X1 U10202 ( .A1(n9267), .A2(n8714), .ZN(n8718) );
  INV_X1 U10203 ( .A(n9261), .ZN(n8715) );
  INV_X1 U10204 ( .A(n9029), .ZN(n9030) );
  AND2_X1 U10205 ( .A1(n9228), .A2(n8837), .ZN(n8882) );
  INV_X1 U10206 ( .A(n8882), .ZN(n8717) );
  NAND2_X1 U10207 ( .A1(n9358), .A2(n9030), .ZN(n8776) );
  INV_X1 U10208 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U10209 ( .A1(n9429), .A2(n9033), .ZN(n8883) );
  OAI211_X1 U10210 ( .C1(n8720), .C2(n8717), .A(n8776), .B(n8883), .ZN(n8721)
         );
  NAND2_X1 U10211 ( .A1(n8776), .A2(n8718), .ZN(n8880) );
  OR2_X1 U10212 ( .A1(n9429), .A2(n9033), .ZN(n8775) );
  NAND2_X1 U10213 ( .A1(n8775), .A2(n9228), .ZN(n8884) );
  INV_X1 U10214 ( .A(n8884), .ZN(n8719) );
  INV_X1 U10215 ( .A(n9038), .ZN(n9036) );
  NAND2_X1 U10216 ( .A1(n9348), .A2(n9036), .ZN(n8774) );
  INV_X1 U10217 ( .A(n9061), .ZN(n8723) );
  INV_X1 U10218 ( .A(n8775), .ZN(n8722) );
  OAI21_X1 U10219 ( .B1(n8723), .B2(n8722), .A(n8758), .ZN(n8726) );
  INV_X1 U10220 ( .A(n9042), .ZN(n9041) );
  NAND2_X1 U10221 ( .A1(n9421), .A2(n9041), .ZN(n9062) );
  NAND2_X1 U10222 ( .A1(n9062), .A2(n8774), .ZN(n8816) );
  OR2_X1 U10223 ( .A1(n9421), .A2(n9041), .ZN(n8815) );
  AND2_X1 U10224 ( .A1(n8815), .A2(n9061), .ZN(n8826) );
  INV_X1 U10225 ( .A(n8826), .ZN(n8724) );
  MUX2_X1 U10226 ( .A(n8816), .B(n8724), .S(n8770), .Z(n8725) );
  AOI21_X1 U10227 ( .B1(n8727), .B2(n8726), .A(n8725), .ZN(n8730) );
  INV_X1 U10228 ( .A(n8815), .ZN(n8728) );
  MUX2_X1 U10229 ( .A(n8728), .B(n4747), .S(n8770), .Z(n8729) );
  INV_X1 U10230 ( .A(n9044), .ZN(n8923) );
  NAND2_X1 U10231 ( .A1(n9196), .A2(n8923), .ZN(n8731) );
  OAI21_X1 U10232 ( .B1(n8730), .B2(n8729), .A(n9185), .ZN(n8738) );
  INV_X1 U10233 ( .A(n9045), .ZN(n8732) );
  OR2_X1 U10234 ( .A1(n9332), .A2(n8732), .ZN(n8773) );
  NAND2_X1 U10235 ( .A1(n8773), .A2(n8731), .ZN(n8810) );
  INV_X1 U10236 ( .A(n8810), .ZN(n8734) );
  INV_X1 U10237 ( .A(n9063), .ZN(n8733) );
  NOR2_X1 U10238 ( .A1(n9060), .A2(n8733), .ZN(n8819) );
  MUX2_X1 U10239 ( .A(n8734), .B(n8819), .S(n8770), .Z(n8737) );
  INV_X1 U10240 ( .A(n8773), .ZN(n8735) );
  MUX2_X1 U10241 ( .A(n9060), .B(n8735), .S(n8770), .Z(n8736) );
  OR2_X1 U10242 ( .A1(n9329), .A2(n9050), .ZN(n9136) );
  NAND2_X1 U10243 ( .A1(n9329), .A2(n9050), .ZN(n8818) );
  NAND2_X1 U10244 ( .A1(n9136), .A2(n8818), .ZN(n9153) );
  INV_X1 U10245 ( .A(n9136), .ZN(n8740) );
  INV_X1 U10246 ( .A(n8818), .ZN(n8739) );
  MUX2_X1 U10247 ( .A(n8740), .B(n8739), .S(n8770), .Z(n8741) );
  INV_X1 U10248 ( .A(n9052), .ZN(n9051) );
  OR2_X1 U10249 ( .A1(n9408), .A2(n9051), .ZN(n8813) );
  NAND2_X1 U10250 ( .A1(n9408), .A2(n9051), .ZN(n9066) );
  INV_X1 U10251 ( .A(n9066), .ZN(n8820) );
  NAND2_X1 U10252 ( .A1(n9318), .A2(n9054), .ZN(n9067) );
  INV_X1 U10253 ( .A(n9067), .ZN(n9106) );
  OR2_X1 U10254 ( .A1(n9318), .A2(n9054), .ZN(n8828) );
  NAND2_X1 U10255 ( .A1(n8830), .A2(n8828), .ZN(n8823) );
  INV_X1 U10256 ( .A(n9077), .ZN(n9058) );
  NAND2_X1 U10257 ( .A1(n9113), .A2(n9055), .ZN(n9069) );
  NAND2_X1 U10258 ( .A1(n9070), .A2(n9069), .ZN(n8825) );
  OAI21_X1 U10259 ( .B1(n8742), .B2(n8825), .A(n8829), .ZN(n8749) );
  INV_X1 U10260 ( .A(n8743), .ZN(n8744) );
  OAI211_X1 U10261 ( .C1(n8744), .C2(n8820), .A(n8828), .B(n8813), .ZN(n8745)
         );
  NAND3_X1 U10262 ( .A1(n8745), .A2(n9069), .A3(n9067), .ZN(n8746) );
  NAND3_X1 U10263 ( .A1(n8746), .A2(n8830), .A3(n8829), .ZN(n8747) );
  NAND2_X1 U10264 ( .A1(n8747), .A2(n9070), .ZN(n8748) );
  NAND2_X1 U10265 ( .A1(n7888), .A2(n8759), .ZN(n8751) );
  NAND2_X1 U10266 ( .A1(n8761), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8750) );
  NAND2_X2 U10267 ( .A1(n8751), .A2(n8750), .ZN(n9301) );
  INV_X1 U10268 ( .A(n8920), .ZN(n8752) );
  NAND2_X1 U10269 ( .A1(n9301), .A2(n8752), .ZN(n8841) );
  INV_X1 U10270 ( .A(n9059), .ZN(n9073) );
  MUX2_X1 U10271 ( .A(n8841), .B(n8833), .S(n8770), .Z(n8753) );
  NAND2_X1 U10272 ( .A1(n8755), .A2(n8759), .ZN(n8757) );
  NAND2_X1 U10273 ( .A1(n8761), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U10274 ( .A1(n8760), .A2(n8759), .ZN(n8763) );
  NAND2_X1 U10275 ( .A1(n8761), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8762) );
  AND2_X1 U10276 ( .A1(n9389), .A2(n9013), .ZN(n8806) );
  NAND2_X1 U10277 ( .A1(n8764), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U10278 ( .A1(n8765), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U10279 ( .A1(n8766), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8767) );
  NAND3_X1 U10280 ( .A1(n8769), .A2(n8768), .A3(n8767), .ZN(n9076) );
  NAND2_X1 U10281 ( .A1(n9076), .A2(n9013), .ZN(n8843) );
  INV_X1 U10282 ( .A(n9389), .ZN(n8772) );
  INV_X1 U10283 ( .A(n9013), .ZN(n8771) );
  INV_X1 U10284 ( .A(n8893), .ZN(n8909) );
  AOI21_X1 U10285 ( .B1(n8908), .B2(n8911), .A(n6522), .ZN(n8919) );
  XOR2_X1 U10286 ( .A(n9076), .B(n9009), .Z(n8807) );
  NAND2_X1 U10287 ( .A1(n8830), .A2(n9069), .ZN(n9102) );
  INV_X1 U10288 ( .A(n9102), .ZN(n9105) );
  INV_X1 U10289 ( .A(n9127), .ZN(n8803) );
  AND2_X1 U10290 ( .A1(n8813), .A2(n9066), .ZN(n9065) );
  NAND2_X1 U10291 ( .A1(n9061), .A2(n8774), .ZN(n9217) );
  NAND2_X1 U10292 ( .A1(n8775), .A2(n8883), .ZN(n9233) );
  INV_X1 U10293 ( .A(n8777), .ZN(n8793) );
  INV_X1 U10294 ( .A(n8778), .ZN(n8782) );
  INV_X1 U10295 ( .A(n8779), .ZN(n8781) );
  NAND4_X1 U10296 ( .A1(n8782), .A2(n8781), .A3(n6522), .A4(n8780), .ZN(n8786)
         );
  OR4_X1 U10297 ( .A1(n8786), .A2(n8785), .A3(n8784), .A4(n8783), .ZN(n8790)
         );
  NOR4_X1 U10298 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n8791)
         );
  NAND4_X1 U10299 ( .A1(n8794), .A2(n8793), .A3(n8792), .A4(n8791), .ZN(n8795)
         );
  NOR4_X1 U10300 ( .A1(n8798), .A2(n8797), .A3(n8796), .A4(n8795), .ZN(n8799)
         );
  NAND4_X1 U10301 ( .A1(n9249), .A2(n9261), .A3(n9280), .A4(n8799), .ZN(n8800)
         );
  NOR3_X1 U10302 ( .A1(n9217), .A2(n9233), .A3(n8800), .ZN(n8801) );
  XNOR2_X1 U10303 ( .A(n9421), .B(n9041), .ZN(n9200) );
  INV_X1 U10304 ( .A(n9200), .ZN(n9199) );
  NAND4_X1 U10305 ( .A1(n9176), .A2(n9185), .A3(n8801), .A4(n9199), .ZN(n8802)
         );
  NOR4_X1 U10306 ( .A1(n8803), .A2(n9137), .A3(n9153), .A4(n8802), .ZN(n8804)
         );
  NAND4_X1 U10307 ( .A1(n9059), .A2(n9088), .A3(n9105), .A4(n8804), .ZN(n8805)
         );
  INV_X1 U10308 ( .A(n8849), .ZN(n8809) );
  NOR2_X1 U10309 ( .A1(n8912), .A2(n8808), .ZN(n8847) );
  NAND3_X1 U10310 ( .A1(n8809), .A2(n9002), .A3(n8847), .ZN(n8918) );
  NAND2_X1 U10311 ( .A1(n9155), .A2(n8810), .ZN(n8811) );
  NAND2_X1 U10312 ( .A1(n8811), .A2(n9136), .ZN(n8812) );
  NAND2_X1 U10313 ( .A1(n8812), .A2(n8818), .ZN(n8814) );
  AND2_X1 U10314 ( .A1(n8814), .A2(n8813), .ZN(n8827) );
  NAND2_X1 U10315 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  NAND3_X1 U10316 ( .A1(n8819), .A2(n8818), .A3(n8817), .ZN(n8821) );
  AOI21_X1 U10317 ( .B1(n8827), .B2(n8821), .A(n8820), .ZN(n8822) );
  NOR2_X1 U10318 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  OR2_X1 U10319 ( .A1(n8825), .A2(n8824), .ZN(n8831) );
  OR2_X1 U10320 ( .A1(n8831), .A2(n9106), .ZN(n8887) );
  AND3_X1 U10321 ( .A1(n8828), .A2(n8827), .A3(n8826), .ZN(n8835) );
  OAI21_X1 U10322 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8832) );
  INV_X1 U10323 ( .A(n8832), .ZN(n8834) );
  OAI211_X1 U10324 ( .C1(n8887), .C2(n8835), .A(n8834), .B(n8833), .ZN(n8889)
         );
  NAND2_X1 U10325 ( .A1(n9279), .A2(n8877), .ZN(n9262) );
  INV_X1 U10326 ( .A(n9228), .ZN(n8838) );
  NOR2_X1 U10327 ( .A1(n9233), .A2(n8838), .ZN(n8839) );
  NOR2_X1 U10328 ( .A1(n8887), .A2(n9216), .ZN(n8840) );
  OAI22_X1 U10329 ( .A1(n8889), .A2(n8840), .B1(n4567), .B2(n9013), .ZN(n8844)
         );
  INV_X1 U10330 ( .A(n9076), .ZN(n8890) );
  NAND2_X1 U10331 ( .A1(n9009), .A2(n8890), .ZN(n8842) );
  NAND2_X1 U10332 ( .A1(n8842), .A2(n8841), .ZN(n8891) );
  OAI22_X1 U10333 ( .A1(n8844), .A2(n8891), .B1(n9009), .B2(n8843), .ZN(n8846)
         );
  AOI211_X1 U10334 ( .C1(n8846), .C2(n8915), .A(n8845), .B(n8893), .ZN(n8848)
         );
  OAI211_X1 U10335 ( .C1(n8849), .C2(n8848), .A(n8847), .B(n6345), .ZN(n8907)
         );
  NAND2_X1 U10336 ( .A1(n7022), .A2(n8850), .ZN(n8854) );
  NAND2_X1 U10337 ( .A1(n8936), .A2(n8851), .ZN(n8853) );
  AND4_X1 U10338 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .ZN(n8858)
         );
  AND4_X1 U10339 ( .A1(n8859), .A2(n8858), .A3(n8857), .A4(n8856), .ZN(n8862)
         );
  OAI211_X1 U10340 ( .C1(n8863), .C2(n8862), .A(n8861), .B(n8860), .ZN(n8866)
         );
  AOI21_X1 U10341 ( .B1(n8866), .B2(n8865), .A(n8864), .ZN(n8872) );
  NAND2_X1 U10342 ( .A1(n8868), .A2(n8867), .ZN(n8871) );
  OAI211_X1 U10343 ( .C1(n8872), .C2(n8871), .A(n8870), .B(n8869), .ZN(n8873)
         );
  NAND2_X1 U10344 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  NAND3_X1 U10345 ( .A1(n8877), .A2(n8876), .A3(n8875), .ZN(n8879) );
  NAND2_X1 U10346 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  AOI21_X1 U10347 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n8885) );
  OAI21_X1 U10348 ( .B1(n8885), .B2(n8884), .A(n8883), .ZN(n8886) );
  NOR2_X1 U10349 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  NOR2_X1 U10350 ( .A1(n8889), .A2(n8888), .ZN(n8892) );
  OAI22_X1 U10351 ( .A1(n8892), .A2(n8891), .B1(n8890), .B2(n9009), .ZN(n8894)
         );
  AOI21_X1 U10352 ( .B1(n8894), .B2(n8915), .A(n8893), .ZN(n8903) );
  OR4_X1 U10353 ( .A1(n8903), .A2(n8895), .A3(n6345), .A4(n8912), .ZN(n8906)
         );
  NAND2_X1 U10354 ( .A1(n8902), .A2(n8896), .ZN(n8897) );
  OAI211_X1 U10355 ( .C1(n8899), .C2(n8898), .A(P1_B_REG_SCAN_IN), .B(n8897), 
        .ZN(n8905) );
  INV_X1 U10356 ( .A(n8900), .ZN(n8901) );
  NAND3_X1 U10357 ( .A1(n8903), .A2(n8902), .A3(n8901), .ZN(n8904) );
  AND4_X1 U10358 ( .A1(n8907), .A2(n8906), .A3(n8905), .A4(n8904), .ZN(n8917)
         );
  OAI21_X1 U10359 ( .B1(n8909), .B2(n6345), .A(n8908), .ZN(n8914) );
  NOR3_X1 U10360 ( .A1(n8912), .A2(n8911), .A3(n8910), .ZN(n8913) );
  OAI211_X1 U10361 ( .C1(n8915), .C2(n6345), .A(n8914), .B(n8913), .ZN(n8916)
         );
  OAI211_X1 U10362 ( .C1(n8919), .C2(n8918), .A(n8917), .B(n8916), .ZN(
        P1_U3242) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9076), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8920), .S(n8935), .Z(
        P1_U3583) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9077), .S(n8935), .Z(
        P1_U3582) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8921), .S(n8935), .Z(
        P1_U3581) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8922), .S(n8935), .Z(
        P1_U3580) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9052), .S(n8935), .Z(
        P1_U3579) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9048), .S(n8935), .Z(
        P1_U3578) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9045), .S(n8935), .Z(
        P1_U3577) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8923), .S(n8935), .Z(
        P1_U3576) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9042), .S(n8935), .Z(
        P1_U3575) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9038), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9032), .S(n8935), .Z(
        P1_U3573) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9029), .S(n8935), .Z(
        P1_U3572) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9028), .S(n8935), .Z(
        P1_U3571) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9027), .S(n8935), .Z(
        P1_U3570) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9023), .S(n8935), .Z(
        P1_U3569) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8924), .S(n8935), .Z(
        P1_U3568) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8925), .S(n8935), .Z(
        P1_U3567) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8926), .S(n8935), .Z(
        P1_U3566) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8927), .S(n8935), .Z(
        P1_U3565) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8928), .S(n8935), .Z(
        P1_U3564) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8929), .S(n8935), .Z(
        P1_U3563) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8930), .S(n8935), .Z(
        P1_U3562) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8931), .S(n8935), .Z(
        P1_U3561) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8932), .S(n8935), .Z(
        P1_U3560) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8933), .S(n8935), .Z(
        P1_U3559) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8934), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6046), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7022), .S(n8935), .Z(
        P1_U3555) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8936), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10393 ( .C1(n8939), .C2(n8938), .A(n9570), .B(n8937), .ZN(n8947)
         );
  OAI211_X1 U10394 ( .C1(n8942), .C2(n8941), .A(n9560), .B(n8940), .ZN(n8946)
         );
  AOI22_X1 U10395 ( .A1(n9547), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n4437), .ZN(n8945) );
  NAND2_X1 U10396 ( .A1(n9577), .A2(n8943), .ZN(n8944) );
  NAND4_X1 U10397 ( .A1(n8947), .A2(n8946), .A3(n8945), .A4(n8944), .ZN(
        P1_U3244) );
  INV_X1 U10398 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U10399 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n4437), .ZN(n8948) );
  OAI21_X1 U10400 ( .B1(n9585), .B2(n10259), .A(n8948), .ZN(n8949) );
  AOI21_X1 U10401 ( .B1(n8950), .B2(n9577), .A(n8949), .ZN(n8959) );
  OAI211_X1 U10402 ( .C1(n8953), .C2(n8952), .A(n9570), .B(n8951), .ZN(n8958)
         );
  OAI211_X1 U10403 ( .C1(n8956), .C2(n8955), .A(n9560), .B(n8954), .ZN(n8957)
         );
  NAND3_X1 U10404 ( .A1(n8959), .A2(n8958), .A3(n8957), .ZN(P1_U3246) );
  INV_X1 U10405 ( .A(n8960), .ZN(n8975) );
  NAND2_X1 U10406 ( .A1(n9547), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n8961) );
  OAI211_X1 U10407 ( .C1(n9565), .C2(n8963), .A(n8962), .B(n8961), .ZN(n8964)
         );
  INV_X1 U10408 ( .A(n8964), .ZN(n8974) );
  OAI211_X1 U10409 ( .C1(n8967), .C2(n8966), .A(n9570), .B(n8965), .ZN(n8973)
         );
  INV_X1 U10410 ( .A(n8968), .ZN(n8969) );
  OAI211_X1 U10411 ( .C1(n8971), .C2(n8970), .A(n9560), .B(n8969), .ZN(n8972)
         );
  NAND4_X1 U10412 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(
        P1_U3247) );
  XNOR2_X1 U10413 ( .A(n9510), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9506) );
  OAI21_X1 U10414 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n8985), .A(n8976), .ZN(
        n9507) );
  NOR2_X1 U10415 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  XNOR2_X1 U10416 ( .A(n8987), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9519) );
  NOR2_X1 U10417 ( .A1(n9520), .A2(n9519), .ZN(n9518) );
  NOR2_X1 U10418 ( .A1(n8977), .A2(n8989), .ZN(n8978) );
  INV_X1 U10419 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9530) );
  XNOR2_X1 U10420 ( .A(n8989), .B(n8977), .ZN(n9531) );
  NOR2_X1 U10421 ( .A1(n9530), .A2(n9531), .ZN(n9529) );
  INV_X1 U10422 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10192) );
  XNOR2_X1 U10423 ( .A(n9550), .B(n10192), .ZN(n9548) );
  NOR2_X1 U10424 ( .A1(n9550), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U10425 ( .A(n8993), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9558) );
  OAI22_X1 U10426 ( .A1(n9559), .A2(n9558), .B1(n8993), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U10427 ( .A1(n9578), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8980) );
  OAI21_X1 U10428 ( .B1(n9578), .B2(P1_REG1_REG_18__SCAN_IN), .A(n8980), .ZN(
        n9575) );
  OR2_X1 U10429 ( .A1(n9576), .A2(n9575), .ZN(n9579) );
  NAND2_X1 U10430 ( .A1(n9579), .A2(n8980), .ZN(n8981) );
  XOR2_X1 U10431 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n8981), .Z(n8999) );
  INV_X1 U10432 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8983) );
  AOI22_X1 U10433 ( .A1(n9510), .A2(n8983), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n8982), .ZN(n9503) );
  OAI21_X1 U10434 ( .B1(n8985), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8984), .ZN(
        n9504) );
  NOR2_X1 U10435 ( .A1(n9503), .A2(n9504), .ZN(n9502) );
  INV_X1 U10436 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8986) );
  AOI22_X1 U10437 ( .A1(n8987), .A2(n8986), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n9524), .ZN(n9516) );
  NOR2_X1 U10438 ( .A1(n9515), .A2(n9516), .ZN(n9514) );
  NOR2_X1 U10439 ( .A1(n8988), .A2(n8989), .ZN(n8990) );
  INV_X1 U10440 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9533) );
  XNOR2_X1 U10441 ( .A(n8989), .B(n8988), .ZN(n9534) );
  NOR2_X1 U10442 ( .A1(n9533), .A2(n9534), .ZN(n9532) );
  XNOR2_X1 U10443 ( .A(n9550), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U10444 ( .A1(n9550), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8991) );
  XNOR2_X1 U10445 ( .A(n8993), .B(n8992), .ZN(n9556) );
  NAND2_X1 U10446 ( .A1(n9555), .A2(n9556), .ZN(n9554) );
  OR2_X1 U10447 ( .A1(n8993), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U10448 ( .A1(n9578), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8996) );
  OAI21_X1 U10449 ( .B1(n9578), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8996), .ZN(
        n8995) );
  INV_X1 U10450 ( .A(n8995), .ZN(n9572) );
  NAND2_X1 U10451 ( .A1(n9573), .A2(n9572), .ZN(n9571) );
  NAND2_X1 U10452 ( .A1(n9571), .A2(n8996), .ZN(n8997) );
  XNOR2_X1 U10453 ( .A(n8997), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9001) );
  INV_X1 U10454 ( .A(n9001), .ZN(n8998) );
  AOI22_X1 U10455 ( .A1(n9560), .A2(n8999), .B1(n8998), .B2(n9570), .ZN(n9004)
         );
  OAI21_X1 U10456 ( .B1(n8999), .B2(n9574), .A(n9565), .ZN(n9000) );
  AOI21_X1 U10457 ( .B1(n9570), .B2(n9001), .A(n9000), .ZN(n9003) );
  MUX2_X1 U10458 ( .A(n9004), .B(n9003), .S(n9002), .Z(n9006) );
  NAND2_X1 U10459 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9005) );
  OAI211_X1 U10460 ( .C1(n9007), .C2(n9585), .A(n9006), .B(n9005), .ZN(
        P1_U3262) );
  INV_X1 U10461 ( .A(n9429), .ZN(n9240) );
  OR2_X1 U10462 ( .A1(n9348), .A2(n9239), .ZN(n9204) );
  NOR2_X2 U10463 ( .A1(n9421), .A2(n9204), .ZN(n9190) );
  NOR2_X2 U10464 ( .A1(n9121), .A2(n9113), .ZN(n9093) );
  NAND2_X1 U10465 ( .A1(n9295), .A2(n9596), .ZN(n9015) );
  NAND2_X1 U10466 ( .A1(n9463), .A2(P1_B_REG_SCAN_IN), .ZN(n9011) );
  AND2_X1 U10467 ( .A1(n9012), .A2(n9011), .ZN(n9075) );
  AND2_X1 U10468 ( .A1(n9272), .A2(n9298), .ZN(n9017) );
  AOI21_X1 U10469 ( .B1(n9609), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9017), .ZN(
        n9014) );
  OAI211_X1 U10470 ( .C1(n9389), .C2(n9602), .A(n9015), .B(n9014), .ZN(
        P1_U3263) );
  XNOR2_X1 U10471 ( .A(n9080), .B(n4567), .ZN(n9299) );
  NAND2_X1 U10472 ( .A1(n9299), .A2(n9182), .ZN(n9019) );
  AND2_X1 U10473 ( .A1(n9609), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9016) );
  NOR2_X1 U10474 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  OAI211_X1 U10475 ( .C1(n4567), .C2(n9602), .A(n9019), .B(n9018), .ZN(
        P1_U3264) );
  NAND2_X1 U10476 ( .A1(n9022), .A2(n5049), .ZN(n9026) );
  NAND2_X1 U10477 ( .A1(n9026), .A2(n9025), .ZN(n9276) );
  NOR2_X1 U10478 ( .A1(n9358), .A2(n9029), .ZN(n9031) );
  AOI21_X1 U10479 ( .B1(n9429), .B2(n9032), .A(n9234), .ZN(n9035) );
  NOR2_X1 U10480 ( .A1(n9035), .A2(n9034), .ZN(n9212) );
  INV_X1 U10481 ( .A(n9348), .ZN(n9225) );
  NAND2_X1 U10482 ( .A1(n9225), .A2(n9036), .ZN(n9037) );
  NAND2_X1 U10483 ( .A1(n9212), .A2(n9037), .ZN(n9040) );
  NAND2_X1 U10484 ( .A1(n9332), .A2(n9045), .ZN(n9047) );
  NOR2_X1 U10485 ( .A1(n9332), .A2(n9045), .ZN(n9046) );
  AOI21_X1 U10486 ( .B1(n9168), .B2(n9047), .A(n9046), .ZN(n9152) );
  OAI21_X1 U10487 ( .B1(n9048), .B2(n9329), .A(n9152), .ZN(n9049) );
  NOR2_X1 U10488 ( .A1(n9144), .A2(n9051), .ZN(n9053) );
  NAND2_X1 U10489 ( .A1(n9103), .A2(n9102), .ZN(n9057) );
  NAND2_X1 U10490 ( .A1(n9404), .A2(n9055), .ZN(n9056) );
  NAND2_X1 U10491 ( .A1(n9057), .A2(n9056), .ZN(n9087) );
  INV_X1 U10492 ( .A(n9311), .ZN(n9099) );
  NOR2_X1 U10493 ( .A1(n9153), .A2(n9060), .ZN(n9064) );
  NAND2_X1 U10494 ( .A1(n9213), .A2(n9061), .ZN(n9201) );
  NAND2_X1 U10495 ( .A1(n9175), .A2(n9176), .ZN(n9174) );
  NAND2_X1 U10496 ( .A1(n9064), .A2(n9174), .ZN(n9156) );
  NAND3_X1 U10497 ( .A1(n9156), .A2(n9065), .A3(n9136), .ZN(n9139) );
  NAND2_X1 U10498 ( .A1(n9139), .A2(n9066), .ZN(n9128) );
  NAND2_X1 U10499 ( .A1(n9128), .A2(n9127), .ZN(n9108) );
  NAND2_X1 U10500 ( .A1(n9108), .A2(n9067), .ZN(n9068) );
  NAND2_X1 U10501 ( .A1(n9068), .A2(n9105), .ZN(n9104) );
  INV_X1 U10502 ( .A(n9070), .ZN(n9071) );
  AOI21_X1 U10503 ( .B1(n9089), .B2(n9088), .A(n9071), .ZN(n9072) );
  XNOR2_X1 U10504 ( .A(n9073), .B(n9072), .ZN(n9074) );
  NAND2_X1 U10505 ( .A1(n9074), .A2(n9278), .ZN(n9079) );
  AOI22_X1 U10506 ( .A1(n8595), .A2(n9077), .B1(n9076), .B2(n9075), .ZN(n9078)
         );
  AOI21_X1 U10507 ( .B1(n9301), .B2(n9094), .A(n9286), .ZN(n9081) );
  NAND2_X1 U10508 ( .A1(n9081), .A2(n9080), .ZN(n9302) );
  AOI22_X1 U10509 ( .A1(n9609), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9598), .B2(
        n9082), .ZN(n9084) );
  NAND2_X1 U10510 ( .A1(n9301), .A2(n9587), .ZN(n9083) );
  OAI211_X1 U10511 ( .C1(n9302), .C2(n9241), .A(n9084), .B(n9083), .ZN(n9085)
         );
  AOI21_X1 U10512 ( .B1(n9305), .B2(n9272), .A(n9085), .ZN(n9086) );
  XNOR2_X1 U10513 ( .A(n9087), .B(n9088), .ZN(n9398) );
  XNOR2_X1 U10514 ( .A(n9089), .B(n9088), .ZN(n9090) );
  NAND2_X1 U10515 ( .A1(n9090), .A2(n9278), .ZN(n9092) );
  INV_X1 U10516 ( .A(n9094), .ZN(n9095) );
  AOI211_X1 U10517 ( .C1(n9311), .C2(n9112), .A(n9286), .B(n9095), .ZN(n9310)
         );
  NAND2_X1 U10518 ( .A1(n9310), .A2(n9596), .ZN(n9098) );
  AOI22_X1 U10519 ( .A1(n9609), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9096), .B2(
        n9598), .ZN(n9097) );
  OAI211_X1 U10520 ( .C1(n9099), .C2(n9602), .A(n9098), .B(n9097), .ZN(n9100)
         );
  AOI21_X1 U10521 ( .B1(n9272), .B2(n9309), .A(n9100), .ZN(n9101) );
  OAI21_X1 U10522 ( .B1(n9398), .B2(n9294), .A(n9101), .ZN(P1_U3265) );
  XNOR2_X1 U10523 ( .A(n9103), .B(n9102), .ZN(n9399) );
  INV_X1 U10524 ( .A(n9399), .ZN(n9119) );
  INV_X1 U10525 ( .A(n9104), .ZN(n9109) );
  OAI21_X1 U10526 ( .B1(n9106), .B2(n9105), .A(n9104), .ZN(n9107) );
  OAI211_X1 U10527 ( .C1(n9109), .C2(n9108), .A(n9278), .B(n9107), .ZN(n9111)
         );
  NAND2_X1 U10528 ( .A1(n9111), .A2(n9110), .ZN(n9314) );
  AOI211_X1 U10529 ( .C1(n9113), .C2(n9121), .A(n9286), .B(n9093), .ZN(n9313)
         );
  NAND2_X1 U10530 ( .A1(n9313), .A2(n9596), .ZN(n9116) );
  AOI22_X1 U10531 ( .A1(n9114), .A2(n9598), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9609), .ZN(n9115) );
  OAI211_X1 U10532 ( .C1(n9404), .C2(n9602), .A(n9116), .B(n9115), .ZN(n9117)
         );
  AOI21_X1 U10533 ( .B1(n9272), .B2(n9314), .A(n9117), .ZN(n9118) );
  OAI21_X1 U10534 ( .B1(n9119), .B2(n9294), .A(n9118), .ZN(P1_U3266) );
  XNOR2_X1 U10535 ( .A(n9120), .B(n9127), .ZN(n9322) );
  INV_X1 U10536 ( .A(n9121), .ZN(n9122) );
  AOI21_X1 U10537 ( .B1(n9318), .B2(n9143), .A(n9122), .ZN(n9319) );
  INV_X1 U10538 ( .A(n9123), .ZN(n9124) );
  AOI22_X1 U10539 ( .A1(n9124), .A2(n9598), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9609), .ZN(n9125) );
  OAI21_X1 U10540 ( .B1(n9126), .B2(n9602), .A(n9125), .ZN(n9133) );
  XNOR2_X1 U10541 ( .A(n9128), .B(n9127), .ZN(n9131) );
  INV_X1 U10542 ( .A(n9129), .ZN(n9130) );
  AOI21_X1 U10543 ( .B1(n9131), .B2(n9278), .A(n9130), .ZN(n9321) );
  NOR2_X1 U10544 ( .A1(n9321), .A2(n9609), .ZN(n9132) );
  AOI211_X1 U10545 ( .C1(n9182), .C2(n9319), .A(n9133), .B(n9132), .ZN(n9134)
         );
  OAI21_X1 U10546 ( .B1(n9322), .B2(n9294), .A(n9134), .ZN(P1_U3267) );
  XNOR2_X1 U10547 ( .A(n9135), .B(n9137), .ZN(n9410) );
  NAND2_X1 U10548 ( .A1(n9156), .A2(n9136), .ZN(n9138) );
  NAND2_X1 U10549 ( .A1(n9138), .A2(n9137), .ZN(n9140) );
  NAND2_X1 U10550 ( .A1(n9140), .A2(n9139), .ZN(n9142) );
  AOI21_X1 U10551 ( .B1(n9142), .B2(n9278), .A(n9141), .ZN(n9324) );
  INV_X1 U10552 ( .A(n9324), .ZN(n9150) );
  OAI211_X1 U10553 ( .C1(n9144), .C2(n4464), .A(n9333), .B(n9143), .ZN(n9323)
         );
  INV_X1 U10554 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9145) );
  OAI22_X1 U10555 ( .A1(n9146), .A2(n9236), .B1(n9145), .B2(n9272), .ZN(n9147)
         );
  AOI21_X1 U10556 ( .B1(n9408), .B2(n9587), .A(n9147), .ZN(n9148) );
  OAI21_X1 U10557 ( .B1(n9323), .B2(n9241), .A(n9148), .ZN(n9149) );
  AOI21_X1 U10558 ( .B1(n9150), .B2(n9272), .A(n9149), .ZN(n9151) );
  OAI21_X1 U10559 ( .B1(n9410), .B2(n9294), .A(n9151), .ZN(P1_U3268) );
  XNOR2_X1 U10560 ( .A(n9152), .B(n9153), .ZN(n9414) );
  INV_X1 U10561 ( .A(n9153), .ZN(n9154) );
  AOI21_X1 U10562 ( .B1(n9174), .B2(n9155), .A(n9154), .ZN(n9160) );
  NAND2_X1 U10563 ( .A1(n9156), .A2(n9278), .ZN(n9159) );
  INV_X1 U10564 ( .A(n9157), .ZN(n9158) );
  OAI21_X1 U10565 ( .B1(n9160), .B2(n9159), .A(n9158), .ZN(n9327) );
  AOI211_X1 U10566 ( .C1(n9329), .C2(n9169), .A(n9286), .B(n4464), .ZN(n9328)
         );
  NAND2_X1 U10567 ( .A1(n9328), .A2(n9596), .ZN(n9164) );
  INV_X1 U10568 ( .A(n9161), .ZN(n9162) );
  AOI22_X1 U10569 ( .A1(n9162), .A2(n9598), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9609), .ZN(n9163) );
  OAI211_X1 U10570 ( .C1(n9165), .C2(n9602), .A(n9164), .B(n9163), .ZN(n9166)
         );
  AOI21_X1 U10571 ( .B1(n9272), .B2(n9327), .A(n9166), .ZN(n9167) );
  OAI21_X1 U10572 ( .B1(n9414), .B2(n9294), .A(n9167), .ZN(P1_U3269) );
  XNOR2_X1 U10573 ( .A(n9168), .B(n9176), .ZN(n9337) );
  INV_X1 U10574 ( .A(n9169), .ZN(n9170) );
  AOI21_X1 U10575 ( .B1(n9332), .B2(n9191), .A(n9170), .ZN(n9334) );
  INV_X1 U10576 ( .A(n9332), .ZN(n9173) );
  AOI22_X1 U10577 ( .A1(n9171), .A2(n9598), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9609), .ZN(n9172) );
  OAI21_X1 U10578 ( .B1(n9173), .B2(n9602), .A(n9172), .ZN(n9181) );
  OAI21_X1 U10579 ( .B1(n9176), .B2(n9175), .A(n9174), .ZN(n9179) );
  INV_X1 U10580 ( .A(n9177), .ZN(n9178) );
  AOI21_X1 U10581 ( .B1(n9179), .B2(n9278), .A(n9178), .ZN(n9336) );
  NOR2_X1 U10582 ( .A1(n9336), .A2(n9609), .ZN(n9180) );
  AOI211_X1 U10583 ( .C1(n9334), .C2(n9182), .A(n9181), .B(n9180), .ZN(n9183)
         );
  OAI21_X1 U10584 ( .B1(n9337), .B2(n9294), .A(n9183), .ZN(P1_U3270) );
  XNOR2_X1 U10585 ( .A(n9184), .B(n9185), .ZN(n9418) );
  XNOR2_X1 U10586 ( .A(n9186), .B(n9185), .ZN(n9187) );
  NAND2_X1 U10587 ( .A1(n9187), .A2(n9278), .ZN(n9189) );
  NAND2_X1 U10588 ( .A1(n9189), .A2(n9188), .ZN(n9338) );
  INV_X1 U10589 ( .A(n9190), .ZN(n9205) );
  INV_X1 U10590 ( .A(n9191), .ZN(n9192) );
  AOI211_X1 U10591 ( .C1(n4671), .C2(n9205), .A(n9286), .B(n9192), .ZN(n9339)
         );
  NAND2_X1 U10592 ( .A1(n9339), .A2(n9596), .ZN(n9195) );
  AOI22_X1 U10593 ( .A1(n9193), .A2(n9598), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9609), .ZN(n9194) );
  OAI211_X1 U10594 ( .C1(n9196), .C2(n9602), .A(n9195), .B(n9194), .ZN(n9197)
         );
  AOI21_X1 U10595 ( .B1(n9272), .B2(n9338), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10596 ( .B1(n9418), .B2(n9294), .A(n9198), .ZN(P1_U3271) );
  XNOR2_X1 U10597 ( .A(n4474), .B(n9199), .ZN(n9423) );
  XNOR2_X1 U10598 ( .A(n9201), .B(n9200), .ZN(n9203) );
  AOI21_X1 U10599 ( .B1(n9203), .B2(n9278), .A(n9202), .ZN(n9343) );
  INV_X1 U10600 ( .A(n9343), .ZN(n9210) );
  INV_X1 U10601 ( .A(n9204), .ZN(n9220) );
  OAI211_X1 U10602 ( .C1(n5019), .C2(n9220), .A(n9205), .B(n9333), .ZN(n9342)
         );
  AOI22_X1 U10603 ( .A1(n9206), .A2(n9598), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9609), .ZN(n9208) );
  NAND2_X1 U10604 ( .A1(n9421), .A2(n9587), .ZN(n9207) );
  OAI211_X1 U10605 ( .C1(n9342), .C2(n9241), .A(n9208), .B(n9207), .ZN(n9209)
         );
  AOI21_X1 U10606 ( .B1(n9210), .B2(n9272), .A(n9209), .ZN(n9211) );
  OAI21_X1 U10607 ( .B1(n9423), .B2(n9294), .A(n9211), .ZN(P1_U3272) );
  XNOR2_X1 U10608 ( .A(n9212), .B(n9217), .ZN(n9426) );
  INV_X1 U10609 ( .A(n9213), .ZN(n9214) );
  AOI211_X1 U10610 ( .C1(n9217), .C2(n9216), .A(n9215), .B(n9214), .ZN(n9219)
         );
  OR2_X1 U10611 ( .A1(n9219), .A2(n9218), .ZN(n9346) );
  AOI211_X1 U10612 ( .C1(n9348), .C2(n9239), .A(n9286), .B(n9220), .ZN(n9347)
         );
  NAND2_X1 U10613 ( .A1(n9347), .A2(n9596), .ZN(n9224) );
  INV_X1 U10614 ( .A(n9221), .ZN(n9222) );
  AOI22_X1 U10615 ( .A1(n9222), .A2(n9598), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9609), .ZN(n9223) );
  OAI211_X1 U10616 ( .C1(n9225), .C2(n9602), .A(n9224), .B(n9223), .ZN(n9226)
         );
  AOI21_X1 U10617 ( .B1(n9346), .B2(n9272), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10618 ( .B1(n9426), .B2(n9294), .A(n9227), .ZN(P1_U3273) );
  NAND2_X1 U10619 ( .A1(n9247), .A2(n9228), .ZN(n9229) );
  XNOR2_X1 U10620 ( .A(n9229), .B(n9233), .ZN(n9232) );
  INV_X1 U10621 ( .A(n9230), .ZN(n9231) );
  AOI21_X1 U10622 ( .B1(n9232), .B2(n9278), .A(n9231), .ZN(n9352) );
  XNOR2_X1 U10623 ( .A(n9234), .B(n9233), .ZN(n9432) );
  INV_X1 U10624 ( .A(n9432), .ZN(n9235) );
  NAND2_X1 U10625 ( .A1(n9235), .A2(n9606), .ZN(n9245) );
  INV_X1 U10626 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9238) );
  OAI22_X1 U10627 ( .A1(n9272), .A2(n9238), .B1(n9237), .B2(n9236), .ZN(n9243)
         );
  OAI211_X1 U10628 ( .C1(n9240), .C2(n4525), .A(n9239), .B(n9333), .ZN(n9351)
         );
  NOR2_X1 U10629 ( .A1(n9351), .A2(n9241), .ZN(n9242) );
  AOI211_X1 U10630 ( .C1(n9587), .C2(n9429), .A(n9243), .B(n9242), .ZN(n9244)
         );
  OAI211_X1 U10631 ( .C1(n9609), .C2(n9352), .A(n9245), .B(n9244), .ZN(
        P1_U3274) );
  XNOR2_X1 U10632 ( .A(n9246), .B(n9249), .ZN(n9436) );
  OAI211_X1 U10633 ( .C1(n9249), .C2(n9248), .A(n9247), .B(n9278), .ZN(n9251)
         );
  NAND2_X1 U10634 ( .A1(n9251), .A2(n9250), .ZN(n9356) );
  AOI211_X1 U10635 ( .C1(n9358), .C2(n9265), .A(n9286), .B(n4525), .ZN(n9357)
         );
  NAND2_X1 U10636 ( .A1(n9357), .A2(n9596), .ZN(n9255) );
  INV_X1 U10637 ( .A(n9252), .ZN(n9253) );
  AOI22_X1 U10638 ( .A1(n9609), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9253), .B2(
        n9598), .ZN(n9254) );
  OAI211_X1 U10639 ( .C1(n4672), .C2(n9602), .A(n9255), .B(n9254), .ZN(n9256)
         );
  AOI21_X1 U10640 ( .B1(n9272), .B2(n9356), .A(n9256), .ZN(n9257) );
  OAI21_X1 U10641 ( .B1(n9436), .B2(n9294), .A(n9257), .ZN(P1_U3275) );
  AOI21_X1 U10642 ( .B1(n9259), .B2(n9261), .A(n9258), .ZN(n9438) );
  INV_X1 U10643 ( .A(n9438), .ZN(n9274) );
  OAI211_X1 U10644 ( .C1(n9262), .C2(n9261), .A(n9260), .B(n9278), .ZN(n9264)
         );
  NAND2_X1 U10645 ( .A1(n9264), .A2(n9263), .ZN(n9363) );
  INV_X1 U10646 ( .A(n9265), .ZN(n9266) );
  AOI211_X1 U10647 ( .C1(n9267), .C2(n9284), .A(n9286), .B(n9266), .ZN(n9362)
         );
  NAND2_X1 U10648 ( .A1(n9362), .A2(n9596), .ZN(n9270) );
  AOI22_X1 U10649 ( .A1(n9609), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9268), .B2(
        n9598), .ZN(n9269) );
  OAI211_X1 U10650 ( .C1(n9445), .C2(n9602), .A(n9270), .B(n9269), .ZN(n9271)
         );
  AOI21_X1 U10651 ( .B1(n9272), .B2(n9363), .A(n9271), .ZN(n9273) );
  OAI21_X1 U10652 ( .B1(n9274), .B2(n9294), .A(n9273), .ZN(P1_U3276) );
  AOI21_X1 U10653 ( .B1(n9280), .B2(n9276), .A(n9275), .ZN(n9277) );
  INV_X1 U10654 ( .A(n9277), .ZN(n9450) );
  OAI211_X1 U10655 ( .C1(n9281), .C2(n9280), .A(n9279), .B(n9278), .ZN(n9283)
         );
  NAND2_X1 U10656 ( .A1(n9283), .A2(n9282), .ZN(n9368) );
  INV_X1 U10657 ( .A(n9284), .ZN(n9285) );
  AOI211_X1 U10658 ( .C1(n9370), .C2(n9287), .A(n9286), .B(n9285), .ZN(n9369)
         );
  NAND2_X1 U10659 ( .A1(n9369), .A2(n9596), .ZN(n9290) );
  AOI22_X1 U10660 ( .A1(n9609), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9288), .B2(
        n9598), .ZN(n9289) );
  OAI211_X1 U10661 ( .C1(n9291), .C2(n9602), .A(n9290), .B(n9289), .ZN(n9292)
         );
  AOI21_X1 U10662 ( .B1(n9272), .B2(n9368), .A(n9292), .ZN(n9293) );
  OAI21_X1 U10663 ( .B1(n9450), .B2(n9294), .A(n9293), .ZN(P1_U3277) );
  INV_X1 U10664 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9296) );
  NOR2_X1 U10665 ( .A1(n9295), .A2(n9298), .ZN(n9387) );
  MUX2_X1 U10666 ( .A(n9296), .B(n9387), .S(n9667), .Z(n9297) );
  OAI21_X1 U10667 ( .B1(n9389), .B2(n9367), .A(n9297), .ZN(P1_U3553) );
  INV_X1 U10668 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10159) );
  AOI21_X1 U10669 ( .B1(n9299), .B2(n9333), .A(n9298), .ZN(n9390) );
  MUX2_X1 U10670 ( .A(n10159), .B(n9390), .S(n9667), .Z(n9300) );
  OAI21_X1 U10671 ( .B1(n4567), .B2(n9367), .A(n9300), .ZN(P1_U3552) );
  NAND2_X1 U10672 ( .A1(n9392), .A2(n9361), .ZN(n9308) );
  INV_X1 U10673 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9306) );
  INV_X1 U10674 ( .A(n9301), .ZN(n9303) );
  OAI21_X1 U10675 ( .B1(n9303), .B2(n9654), .A(n9302), .ZN(n9304) );
  MUX2_X1 U10676 ( .A(n9306), .B(n9393), .S(n9667), .Z(n9307) );
  NAND2_X1 U10677 ( .A1(n9308), .A2(n9307), .ZN(P1_U3551) );
  INV_X1 U10678 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10247) );
  MUX2_X1 U10679 ( .A(n10247), .B(n9395), .S(n9667), .Z(n9312) );
  NAND2_X1 U10680 ( .A1(n9399), .A2(n9361), .ZN(n9317) );
  NOR2_X1 U10681 ( .A1(n9314), .A2(n9313), .ZN(n9400) );
  MUX2_X1 U10682 ( .A(n9315), .B(n9400), .S(n9667), .Z(n9316) );
  OAI211_X1 U10683 ( .C1(n9404), .C2(n9367), .A(n9317), .B(n9316), .ZN(
        P1_U3549) );
  AOI22_X1 U10684 ( .A1(n9319), .A2(n9333), .B1(n9382), .B2(n9318), .ZN(n9320)
         );
  OAI211_X1 U10685 ( .C1(n9322), .C2(n9384), .A(n9321), .B(n9320), .ZN(n9405)
         );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9405), .S(n9667), .Z(
        P1_U3548) );
  NAND2_X1 U10687 ( .A1(n9324), .A2(n9323), .ZN(n9406) );
  MUX2_X1 U10688 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9406), .S(n9667), .Z(n9325) );
  AOI21_X1 U10689 ( .B1(n9354), .B2(n9408), .A(n9325), .ZN(n9326) );
  OAI21_X1 U10690 ( .B1(n9410), .B2(n9372), .A(n9326), .ZN(P1_U3547) );
  AOI211_X1 U10691 ( .C1(n9382), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9411)
         );
  MUX2_X1 U10692 ( .A(n9330), .B(n9411), .S(n9667), .Z(n9331) );
  OAI21_X1 U10693 ( .B1(n9414), .B2(n9372), .A(n9331), .ZN(P1_U3546) );
  AOI22_X1 U10694 ( .A1(n9334), .A2(n9333), .B1(n9382), .B2(n9332), .ZN(n9335)
         );
  OAI211_X1 U10695 ( .C1(n9337), .C2(n9384), .A(n9336), .B(n9335), .ZN(n9415)
         );
  MUX2_X1 U10696 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9415), .S(n9667), .Z(
        P1_U3545) );
  INV_X1 U10697 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9340) );
  AOI211_X1 U10698 ( .C1(n9382), .C2(n4671), .A(n9339), .B(n9338), .ZN(n9416)
         );
  MUX2_X1 U10699 ( .A(n9340), .B(n9416), .S(n9667), .Z(n9341) );
  OAI21_X1 U10700 ( .B1(n9418), .B2(n9372), .A(n9341), .ZN(P1_U3544) );
  NAND2_X1 U10701 ( .A1(n9343), .A2(n9342), .ZN(n9419) );
  MUX2_X1 U10702 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9419), .S(n9667), .Z(n9344) );
  AOI21_X1 U10703 ( .B1(n9354), .B2(n9421), .A(n9344), .ZN(n9345) );
  OAI21_X1 U10704 ( .B1(n9423), .B2(n9372), .A(n9345), .ZN(P1_U3543) );
  INV_X1 U10705 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9349) );
  AOI211_X1 U10706 ( .C1(n9382), .C2(n9348), .A(n9347), .B(n9346), .ZN(n9424)
         );
  MUX2_X1 U10707 ( .A(n9349), .B(n9424), .S(n9667), .Z(n9350) );
  OAI21_X1 U10708 ( .B1(n9426), .B2(n9372), .A(n9350), .ZN(P1_U3542) );
  NAND2_X1 U10709 ( .A1(n9352), .A2(n9351), .ZN(n9427) );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9427), .S(n9667), .Z(n9353) );
  AOI21_X1 U10711 ( .B1(n9354), .B2(n9429), .A(n9353), .ZN(n9355) );
  OAI21_X1 U10712 ( .B1(n9432), .B2(n9372), .A(n9355), .ZN(P1_U3541) );
  INV_X1 U10713 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9359) );
  AOI211_X1 U10714 ( .C1(n9382), .C2(n9358), .A(n9357), .B(n9356), .ZN(n9433)
         );
  MUX2_X1 U10715 ( .A(n9359), .B(n9433), .S(n9667), .Z(n9360) );
  OAI21_X1 U10716 ( .B1(n9436), .B2(n9372), .A(n9360), .ZN(P1_U3540) );
  NAND2_X1 U10717 ( .A1(n9438), .A2(n9361), .ZN(n9366) );
  NOR2_X1 U10718 ( .A1(n9363), .A2(n9362), .ZN(n9440) );
  MUX2_X1 U10719 ( .A(n9364), .B(n9440), .S(n9667), .Z(n9365) );
  OAI211_X1 U10720 ( .C1(n9445), .C2(n9367), .A(n9366), .B(n9365), .ZN(
        P1_U3539) );
  AOI211_X1 U10721 ( .C1(n9382), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9446)
         );
  MUX2_X1 U10722 ( .A(n10192), .B(n9446), .S(n9667), .Z(n9371) );
  OAI21_X1 U10723 ( .B1(n9450), .B2(n9372), .A(n9371), .ZN(P1_U3538) );
  INV_X1 U10724 ( .A(n9373), .ZN(n9378) );
  AOI21_X1 U10725 ( .B1(n9382), .B2(n9375), .A(n9374), .ZN(n9376) );
  OAI211_X1 U10726 ( .C1(n9652), .C2(n9378), .A(n9377), .B(n9376), .ZN(n9451)
         );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9451), .S(n9667), .Z(
        P1_U3536) );
  AOI211_X1 U10728 ( .C1(n9382), .C2(n9381), .A(n9380), .B(n9379), .ZN(n9383)
         );
  OAI21_X1 U10729 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9452) );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9452), .S(n9667), .Z(
        P1_U3535) );
  MUX2_X1 U10731 ( .A(n9386), .B(P1_REG1_REG_0__SCAN_IN), .S(n9665), .Z(
        P1_U3522) );
  INV_X1 U10732 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10244) );
  MUX2_X1 U10733 ( .A(n10244), .B(n9387), .S(n9439), .Z(n9388) );
  OAI21_X1 U10734 ( .B1(n9389), .B2(n9444), .A(n9388), .ZN(P1_U3521) );
  INV_X1 U10735 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10231) );
  MUX2_X1 U10736 ( .A(n10231), .B(n9390), .S(n9439), .Z(n9391) );
  OAI21_X1 U10737 ( .B1(n4567), .B2(n9444), .A(n9391), .ZN(P1_U3520) );
  NAND2_X1 U10738 ( .A1(n9392), .A2(n9437), .ZN(n9394) );
  INV_X1 U10739 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10044) );
  INV_X1 U10740 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9396) );
  MUX2_X1 U10741 ( .A(n9396), .B(n9395), .S(n9439), .Z(n9397) );
  NAND2_X1 U10742 ( .A1(n9399), .A2(n9437), .ZN(n9403) );
  INV_X1 U10743 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9401) );
  MUX2_X1 U10744 ( .A(n9401), .B(n9400), .S(n9439), .Z(n9402) );
  OAI211_X1 U10745 ( .C1(n9404), .C2(n9444), .A(n9403), .B(n9402), .ZN(
        P1_U3517) );
  MUX2_X1 U10746 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9405), .S(n9439), .Z(
        P1_U3516) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9406), .S(n9439), .Z(n9407) );
  AOI21_X1 U10748 ( .B1(n9430), .B2(n9408), .A(n9407), .ZN(n9409) );
  OAI21_X1 U10749 ( .B1(n9410), .B2(n9449), .A(n9409), .ZN(P1_U3515) );
  INV_X1 U10750 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9412) );
  MUX2_X1 U10751 ( .A(n9412), .B(n9411), .S(n9439), .Z(n9413) );
  OAI21_X1 U10752 ( .B1(n9414), .B2(n9449), .A(n9413), .ZN(P1_U3514) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9415), .S(n9439), .Z(
        P1_U3513) );
  MUX2_X1 U10754 ( .A(n10096), .B(n9416), .S(n9439), .Z(n9417) );
  OAI21_X1 U10755 ( .B1(n9418), .B2(n9449), .A(n9417), .ZN(P1_U3512) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9419), .S(n9439), .Z(n9420) );
  AOI21_X1 U10757 ( .B1(n9430), .B2(n9421), .A(n9420), .ZN(n9422) );
  OAI21_X1 U10758 ( .B1(n9423), .B2(n9449), .A(n9422), .ZN(P1_U3511) );
  MUX2_X1 U10759 ( .A(n10168), .B(n9424), .S(n9439), .Z(n9425) );
  OAI21_X1 U10760 ( .B1(n9426), .B2(n9449), .A(n9425), .ZN(P1_U3510) );
  MUX2_X1 U10761 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9427), .S(n9439), .Z(n9428) );
  AOI21_X1 U10762 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9431) );
  OAI21_X1 U10763 ( .B1(n9432), .B2(n9449), .A(n9431), .ZN(P1_U3509) );
  INV_X1 U10764 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9434) );
  MUX2_X1 U10765 ( .A(n9434), .B(n9433), .S(n9439), .Z(n9435) );
  OAI21_X1 U10766 ( .B1(n9436), .B2(n9449), .A(n9435), .ZN(P1_U3507) );
  NAND2_X1 U10767 ( .A1(n9438), .A2(n9437), .ZN(n9443) );
  MUX2_X1 U10768 ( .A(n9441), .B(n9440), .S(n9439), .Z(n9442) );
  OAI211_X1 U10769 ( .C1(n9445), .C2(n9444), .A(n9443), .B(n9442), .ZN(
        P1_U3504) );
  INV_X1 U10770 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9447) );
  MUX2_X1 U10771 ( .A(n9447), .B(n9446), .S(n9439), .Z(n9448) );
  OAI21_X1 U10772 ( .B1(n9450), .B2(n9449), .A(n9448), .ZN(P1_U3501) );
  MUX2_X1 U10773 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9451), .S(n9439), .Z(
        P1_U3495) );
  MUX2_X1 U10774 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9452), .S(n9439), .Z(
        P1_U3492) );
  NOR4_X1 U10775 ( .A1(n9453), .A2(P1_IR_REG_30__SCAN_IN), .A3(n6198), .A4(
        P1_U3086), .ZN(n9454) );
  AOI21_X1 U10776 ( .B1(n9462), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9454), .ZN(
        n9455) );
  OAI21_X1 U10777 ( .B1(n9456), .B2(n7778), .A(n9455), .ZN(P1_U3324) );
  AOI22_X1 U10778 ( .A1(n5981), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9462), .ZN(n9457) );
  OAI21_X1 U10779 ( .B1(n9458), .B2(n7778), .A(n9457), .ZN(P1_U3325) );
  AOI22_X1 U10780 ( .A1(n9459), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9462), .ZN(n9460) );
  OAI21_X1 U10781 ( .B1(n9461), .B2(n7778), .A(n9460), .ZN(P1_U3327) );
  AOI22_X1 U10782 ( .A1(n9463), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9462), .ZN(n9464) );
  OAI21_X1 U10783 ( .B1(n9465), .B2(n7778), .A(n9464), .ZN(P1_U3328) );
  OAI222_X1 U10784 ( .A1(n9468), .A2(n4437), .B1(n7778), .B2(n9467), .C1(
        n10183), .C2(n9466), .ZN(P1_U3329) );
  MUX2_X1 U10785 ( .A(n9469), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI22_X1 U10786 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9830), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(P2_U3151), .ZN(n9487) );
  XNOR2_X1 U10787 ( .A(n9471), .B(n9470), .ZN(n9478) );
  INV_X1 U10788 ( .A(n9472), .ZN(n9474) );
  NAND2_X1 U10789 ( .A1(n9474), .A2(n9473), .ZN(n9480) );
  OAI21_X1 U10790 ( .B1(n9480), .B2(n9475), .A(n9696), .ZN(n9476) );
  AOI22_X1 U10791 ( .A1(n9478), .A2(n9839), .B1(n9477), .B2(n9476), .ZN(n9486)
         );
  NAND3_X1 U10792 ( .A1(n9480), .A2(n6714), .A3(n9479), .ZN(n9485) );
  OR2_X1 U10793 ( .A1(n9483), .A2(n9845), .ZN(n9484) );
  NAND4_X1 U10794 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(
        P2_U3200) );
  OAI21_X1 U10795 ( .B1(n9490), .B2(n9489), .A(n9488), .ZN(n9496) );
  AOI21_X1 U10796 ( .B1(n9492), .B2(n9491), .A(n7828), .ZN(n9494) );
  NOR2_X1 U10797 ( .A1(n9494), .A2(n9493), .ZN(n9495) );
  AOI211_X1 U10798 ( .C1(n9498), .C2(n9497), .A(n9496), .B(n9495), .ZN(n9499)
         );
  OAI21_X1 U10799 ( .B1(n9501), .B2(n9500), .A(n9499), .ZN(P1_U3217) );
  XNOR2_X1 U10800 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10801 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10802 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9513) );
  AOI211_X1 U10803 ( .C1(n9504), .C2(n9503), .A(n9502), .B(n9541), .ZN(n9509)
         );
  AOI211_X1 U10804 ( .C1(n9507), .C2(n9506), .A(n9505), .B(n9574), .ZN(n9508)
         );
  AOI211_X1 U10805 ( .C1(n9577), .C2(n9510), .A(n9509), .B(n9508), .ZN(n9512)
         );
  OAI211_X1 U10806 ( .C1(n9585), .C2(n9513), .A(n9512), .B(n9511), .ZN(
        P1_U3256) );
  INV_X1 U10807 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9528) );
  AOI21_X1 U10808 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(n9517) );
  NAND2_X1 U10809 ( .A1(n9570), .A2(n9517), .ZN(n9523) );
  AOI21_X1 U10810 ( .B1(n9520), .B2(n9519), .A(n9518), .ZN(n9521) );
  NAND2_X1 U10811 ( .A1(n9560), .A2(n9521), .ZN(n9522) );
  OAI211_X1 U10812 ( .C1(n9565), .C2(n9524), .A(n9523), .B(n9522), .ZN(n9525)
         );
  INV_X1 U10813 ( .A(n9525), .ZN(n9527) );
  NAND2_X1 U10814 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9526) );
  OAI211_X1 U10815 ( .C1(n9585), .C2(n9528), .A(n9527), .B(n9526), .ZN(
        P1_U3257) );
  INV_X1 U10816 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10079) );
  AOI211_X1 U10817 ( .C1(n9531), .C2(n9530), .A(n9529), .B(n9574), .ZN(n9536)
         );
  AOI211_X1 U10818 ( .C1(n9534), .C2(n9533), .A(n9532), .B(n9541), .ZN(n9535)
         );
  AOI211_X1 U10819 ( .C1(n9577), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9539)
         );
  OAI211_X1 U10820 ( .C1(n9585), .C2(n10079), .A(n9539), .B(n9538), .ZN(
        P1_U3258) );
  INV_X1 U10821 ( .A(n9540), .ZN(n9542) );
  AOI211_X1 U10822 ( .C1(n9544), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9545)
         );
  AOI211_X1 U10823 ( .C1(n9547), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9546), .B(
        n9545), .ZN(n9553) );
  XNOR2_X1 U10824 ( .A(n9549), .B(n9548), .ZN(n9551) );
  AOI22_X1 U10825 ( .A1(n9551), .A2(n9560), .B1(n9550), .B2(n9577), .ZN(n9552)
         );
  NAND2_X1 U10826 ( .A1(n9553), .A2(n9552), .ZN(P1_U3259) );
  INV_X1 U10827 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9569) );
  OAI21_X1 U10828 ( .B1(n9556), .B2(n9555), .A(n9554), .ZN(n9557) );
  NAND2_X1 U10829 ( .A1(n9557), .A2(n9570), .ZN(n9563) );
  XNOR2_X1 U10830 ( .A(n9559), .B(n9558), .ZN(n9561) );
  NAND2_X1 U10831 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  OAI211_X1 U10832 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9566)
         );
  INV_X1 U10833 ( .A(n9566), .ZN(n9568) );
  OAI211_X1 U10834 ( .C1(n9585), .C2(n9569), .A(n9568), .B(n9567), .ZN(
        P1_U3260) );
  OAI211_X1 U10835 ( .C1(n9573), .C2(n9572), .A(n9571), .B(n9570), .ZN(n9582)
         );
  AOI21_X1 U10836 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9580) );
  AOI22_X1 U10837 ( .A1(n9580), .A2(n9579), .B1(n9578), .B2(n9577), .ZN(n9581)
         );
  AND2_X1 U10838 ( .A1(n9582), .A2(n9581), .ZN(n9584) );
  NAND2_X1 U10839 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(n4437), .ZN(n9583) );
  OAI211_X1 U10840 ( .C1(n9585), .C2(n9936), .A(n9584), .B(n9583), .ZN(
        P1_U3261) );
  AOI222_X1 U10841 ( .A1(n9588), .A2(n9587), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9609), .C1(n9586), .C2(n9598), .ZN(n9594) );
  INV_X1 U10842 ( .A(n9589), .ZN(n9590) );
  AOI22_X1 U10843 ( .A1(n9592), .A2(n9591), .B1(n9596), .B2(n9590), .ZN(n9593)
         );
  OAI211_X1 U10844 ( .C1(n9609), .C2(n9595), .A(n9594), .B(n9593), .ZN(
        P1_U3286) );
  NAND2_X1 U10845 ( .A1(n9597), .A2(n9596), .ZN(n9601) );
  AOI22_X1 U10846 ( .A1(n9609), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9599), .B2(
        n9598), .ZN(n9600) );
  OAI211_X1 U10847 ( .C1(n9603), .C2(n9602), .A(n9601), .B(n9600), .ZN(n9604)
         );
  AOI21_X1 U10848 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  OAI21_X1 U10849 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(P1_U3289) );
  INV_X1 U10850 ( .A(n9610), .ZN(n9611) );
  NOR2_X4 U10851 ( .A1(n9612), .A2(n9611), .ZN(n9635) );
  INV_X1 U10852 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9613) );
  NOR2_X1 U10853 ( .A1(n9635), .A2(n9613), .ZN(P1_U3294) );
  INV_X1 U10854 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9614) );
  NOR2_X1 U10855 ( .A1(n9635), .A2(n9614), .ZN(P1_U3295) );
  INV_X1 U10856 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9615) );
  NOR2_X1 U10857 ( .A1(n9635), .A2(n9615), .ZN(P1_U3296) );
  INV_X1 U10858 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9616) );
  NOR2_X1 U10859 ( .A1(n9635), .A2(n9616), .ZN(P1_U3297) );
  INV_X1 U10860 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U10861 ( .A1(n9635), .A2(n10112), .ZN(P1_U3298) );
  INV_X1 U10862 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9617) );
  NOR2_X1 U10863 ( .A1(n9635), .A2(n9617), .ZN(P1_U3299) );
  INV_X1 U10864 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9618) );
  NOR2_X1 U10865 ( .A1(n9635), .A2(n9618), .ZN(P1_U3300) );
  INV_X1 U10866 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9619) );
  NOR2_X1 U10867 ( .A1(n9635), .A2(n9619), .ZN(P1_U3301) );
  INV_X1 U10868 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9620) );
  NOR2_X1 U10869 ( .A1(n9635), .A2(n9620), .ZN(P1_U3302) );
  INV_X1 U10870 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9621) );
  NOR2_X1 U10871 ( .A1(n9635), .A2(n9621), .ZN(P1_U3303) );
  INV_X1 U10872 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9622) );
  NOR2_X1 U10873 ( .A1(n9635), .A2(n9622), .ZN(P1_U3304) );
  INV_X1 U10874 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9623) );
  NOR2_X1 U10875 ( .A1(n9635), .A2(n9623), .ZN(P1_U3305) );
  INV_X1 U10876 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9624) );
  NOR2_X1 U10877 ( .A1(n9635), .A2(n9624), .ZN(P1_U3306) );
  INV_X1 U10878 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9625) );
  NOR2_X1 U10879 ( .A1(n9635), .A2(n9625), .ZN(P1_U3307) );
  INV_X1 U10880 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9626) );
  NOR2_X1 U10881 ( .A1(n9635), .A2(n9626), .ZN(P1_U3308) );
  INV_X1 U10882 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9627) );
  NOR2_X1 U10883 ( .A1(n9635), .A2(n9627), .ZN(P1_U3309) );
  INV_X1 U10884 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U10885 ( .A1(n9635), .A2(n10115), .ZN(P1_U3310) );
  INV_X1 U10886 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9628) );
  NOR2_X1 U10887 ( .A1(n9635), .A2(n9628), .ZN(P1_U3311) );
  INV_X1 U10888 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9629) );
  NOR2_X1 U10889 ( .A1(n9635), .A2(n9629), .ZN(P1_U3312) );
  INV_X1 U10890 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U10891 ( .A1(n9635), .A2(n9630), .ZN(P1_U3313) );
  INV_X1 U10892 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U10893 ( .A1(n9635), .A2(n10028), .ZN(P1_U3314) );
  INV_X1 U10894 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U10895 ( .A1(n9635), .A2(n9631), .ZN(P1_U3315) );
  INV_X1 U10896 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9632) );
  NOR2_X1 U10897 ( .A1(n9635), .A2(n9632), .ZN(P1_U3316) );
  INV_X1 U10898 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9633) );
  NOR2_X1 U10899 ( .A1(n9635), .A2(n9633), .ZN(P1_U3317) );
  INV_X1 U10900 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U10901 ( .A1(n9635), .A2(n10184), .ZN(P1_U3318) );
  INV_X1 U10902 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9634) );
  NOR2_X1 U10903 ( .A1(n9635), .A2(n9634), .ZN(P1_U3319) );
  INV_X1 U10904 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10089) );
  NOR2_X1 U10905 ( .A1(n9635), .A2(n10089), .ZN(P1_U3320) );
  INV_X1 U10906 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10260) );
  NOR2_X1 U10907 ( .A1(n9635), .A2(n10260), .ZN(P1_U3321) );
  INV_X1 U10908 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U10909 ( .A1(n9635), .A2(n10034), .ZN(P1_U3322) );
  INV_X1 U10910 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U10911 ( .A1(n9635), .A2(n10058), .ZN(P1_U3323) );
  INV_X1 U10912 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9637) );
  OAI21_X1 U10913 ( .B1(n9638), .B2(n9637), .A(n9636), .ZN(P1_U3439) );
  OAI21_X1 U10914 ( .B1(n9640), .B2(n9654), .A(n9639), .ZN(n9642) );
  AOI211_X1 U10915 ( .C1(n9650), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9662)
         );
  INV_X1 U10916 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9644) );
  AOI22_X1 U10917 ( .A1(n9439), .A2(n9662), .B1(n9644), .B2(n9661), .ZN(
        P1_U3462) );
  OAI21_X1 U10918 ( .B1(n9646), .B2(n9654), .A(n9645), .ZN(n9648) );
  AOI211_X1 U10919 ( .C1(n9650), .C2(n9649), .A(n9648), .B(n9647), .ZN(n9664)
         );
  INV_X1 U10920 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9651) );
  AOI22_X1 U10921 ( .A1(n9439), .A2(n9664), .B1(n9651), .B2(n9661), .ZN(
        P1_U3477) );
  INV_X1 U10922 ( .A(n9652), .ZN(n9657) );
  OAI21_X1 U10923 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9656) );
  AOI21_X1 U10924 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9659) );
  AND2_X1 U10925 ( .A1(n9660), .A2(n9659), .ZN(n9666) );
  INV_X1 U10926 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U10927 ( .A1(n9439), .A2(n9666), .B1(n10257), .B2(n9661), .ZN(
        P1_U3486) );
  AOI22_X1 U10928 ( .A1(n9667), .A2(n9662), .B1(n6799), .B2(n9665), .ZN(
        P1_U3525) );
  INV_X1 U10929 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U10930 ( .A1(n9667), .A2(n9664), .B1(n9663), .B2(n9665), .ZN(
        P1_U3530) );
  AOI22_X1 U10931 ( .A1(n9667), .A2(n9666), .B1(n7013), .B2(n9665), .ZN(
        P1_U3533) );
  AOI22_X1 U10932 ( .A1(n9832), .A2(P2_IR_REG_0__SCAN_IN), .B1(n9830), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n9673) );
  INV_X1 U10933 ( .A(n9668), .ZN(n9671) );
  XNOR2_X1 U10934 ( .A(n9669), .B(P2_IR_REG_0__SCAN_IN), .ZN(n9670) );
  OAI21_X1 U10935 ( .B1(n6714), .B2(n9671), .A(n9670), .ZN(n9672) );
  OAI211_X1 U10936 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10057), .A(n9673), .B(
        n9672), .ZN(P2_U3182) );
  INV_X1 U10937 ( .A(n9674), .ZN(n9675) );
  AOI21_X1 U10938 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9682) );
  XNOR2_X1 U10939 ( .A(n9678), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U10940 ( .A1(n9839), .A2(n9679), .ZN(n9681) );
  OAI211_X1 U10941 ( .C1(n9682), .C2(n9845), .A(n9681), .B(n9680), .ZN(n9683)
         );
  AOI21_X1 U10942 ( .B1(n9684), .B2(n9832), .A(n9683), .ZN(n9691) );
  AOI21_X1 U10943 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9688) );
  NOR2_X1 U10944 ( .A1(n9688), .A2(n9708), .ZN(n9689) );
  AOI21_X1 U10945 ( .B1(n9830), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n9689), .ZN(
        n9690) );
  NAND2_X1 U10946 ( .A1(n9691), .A2(n9690), .ZN(P2_U3185) );
  OAI21_X1 U10947 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9704) );
  OAI21_X1 U10948 ( .B1(n9696), .B2(n4622), .A(n9695), .ZN(n9703) );
  NAND2_X1 U10949 ( .A1(n9698), .A2(n9697), .ZN(n9700) );
  AOI21_X1 U10950 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9702) );
  AOI211_X1 U10951 ( .C1(n9740), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9712)
         );
  AOI21_X1 U10952 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9709) );
  NOR2_X1 U10953 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  AOI21_X1 U10954 ( .B1(n9830), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9710), .ZN(
        n9711) );
  NAND2_X1 U10955 ( .A1(n9712), .A2(n9711), .ZN(P2_U3188) );
  AOI22_X1 U10956 ( .A1(n9832), .A2(n9713), .B1(n9830), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n9729) );
  OAI21_X1 U10957 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9721) );
  OAI21_X1 U10958 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9720) );
  AOI22_X1 U10959 ( .A1(n9721), .A2(n6714), .B1(n9839), .B2(n9720), .ZN(n9728)
         );
  AOI21_X1 U10960 ( .B1(n9724), .B2(n9723), .A(n9722), .ZN(n9725) );
  OR2_X1 U10961 ( .A1(n9725), .A2(n9845), .ZN(n9726) );
  NAND4_X1 U10962 ( .A1(n9729), .A2(n9728), .A3(n9727), .A4(n9726), .ZN(
        P2_U3192) );
  AOI22_X1 U10963 ( .A1(n9832), .A2(n9730), .B1(n9830), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n9746) );
  OAI21_X1 U10964 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n9732), .A(n9731), .ZN(
        n9737) );
  OAI21_X1 U10965 ( .B1(n9735), .B2(n9734), .A(n9733), .ZN(n9736) );
  AOI22_X1 U10966 ( .A1(n9737), .A2(n9839), .B1(n6714), .B2(n9736), .ZN(n9745)
         );
  INV_X1 U10967 ( .A(n9738), .ZN(n9739) );
  NOR2_X1 U10968 ( .A1(n9739), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9741) );
  OAI21_X1 U10969 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9743) );
  NAND4_X1 U10970 ( .A1(n9746), .A2(n9745), .A3(n9744), .A4(n9743), .ZN(
        P2_U3193) );
  AOI22_X1 U10971 ( .A1(n9832), .A2(n9747), .B1(n9830), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9763) );
  OAI21_X1 U10972 ( .B1(n9750), .B2(n9749), .A(n9748), .ZN(n9755) );
  OAI21_X1 U10973 ( .B1(n9753), .B2(n9752), .A(n9751), .ZN(n9754) );
  AOI22_X1 U10974 ( .A1(n9755), .A2(n9839), .B1(n6714), .B2(n9754), .ZN(n9762)
         );
  AOI21_X1 U10975 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9759) );
  OR2_X1 U10976 ( .A1(n9759), .A2(n9845), .ZN(n9760) );
  NAND4_X1 U10977 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(
        P2_U3194) );
  AOI22_X1 U10978 ( .A1(n9832), .A2(n9764), .B1(n9830), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9779) );
  OAI21_X1 U10979 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9766), .A(n9765), .ZN(
        n9771) );
  OAI21_X1 U10980 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  AOI22_X1 U10981 ( .A1(n9771), .A2(n9839), .B1(n6714), .B2(n9770), .ZN(n9778)
         );
  AOI21_X1 U10982 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9775) );
  OR2_X1 U10983 ( .A1(n9775), .A2(n9845), .ZN(n9776) );
  NAND4_X1 U10984 ( .A1(n9779), .A2(n9778), .A3(n9777), .A4(n9776), .ZN(
        P2_U3195) );
  AOI22_X1 U10985 ( .A1(n9832), .A2(n9780), .B1(n9830), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9796) );
  OAI21_X1 U10986 ( .B1(n9783), .B2(n9782), .A(n9781), .ZN(n9788) );
  OAI21_X1 U10987 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(n9787) );
  AOI22_X1 U10988 ( .A1(n9788), .A2(n9839), .B1(n6714), .B2(n9787), .ZN(n9795)
         );
  AOI21_X1 U10989 ( .B1(n9791), .B2(n9790), .A(n9789), .ZN(n9792) );
  OR2_X1 U10990 ( .A1(n9792), .A2(n9845), .ZN(n9793) );
  NAND4_X1 U10991 ( .A1(n9796), .A2(n9795), .A3(n9794), .A4(n9793), .ZN(
        P2_U3196) );
  AOI22_X1 U10992 ( .A1(n9832), .A2(n9797), .B1(n9830), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9812) );
  OAI21_X1 U10993 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9799), .A(n9798), .ZN(
        n9804) );
  OAI21_X1 U10994 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(n9803) );
  AOI22_X1 U10995 ( .A1(n9804), .A2(n9839), .B1(n6714), .B2(n9803), .ZN(n9811)
         );
  AOI21_X1 U10996 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9808) );
  OR2_X1 U10997 ( .A1(n9808), .A2(n9845), .ZN(n9809) );
  NAND4_X1 U10998 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(
        P2_U3197) );
  AOI22_X1 U10999 ( .A1(n9832), .A2(n9813), .B1(n9830), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n9829) );
  OAI21_X1 U11000 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9821) );
  OAI21_X1 U11001 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(n9820) );
  AOI22_X1 U11002 ( .A1(n9821), .A2(n9839), .B1(n6714), .B2(n9820), .ZN(n9828)
         );
  AOI21_X1 U11003 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9825) );
  OR2_X1 U11004 ( .A1(n9825), .A2(n9845), .ZN(n9826) );
  NAND4_X1 U11005 ( .A1(n9829), .A2(n9828), .A3(n9827), .A4(n9826), .ZN(
        P2_U3198) );
  AOI22_X1 U11006 ( .A1(n9832), .A2(n9831), .B1(n9830), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9849) );
  OAI21_X1 U11007 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9834), .A(n9833), .ZN(
        n9840) );
  OAI21_X1 U11008 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9838) );
  AOI22_X1 U11009 ( .A1(n9840), .A2(n9839), .B1(n6714), .B2(n9838), .ZN(n9848)
         );
  NAND2_X1 U11010 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n9847) );
  AOI21_X1 U11011 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9844) );
  OR2_X1 U11012 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  NAND4_X1 U11013 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(
        P2_U3199) );
  OAI21_X1 U11014 ( .B1(n9851), .B2(n9859), .A(n9850), .ZN(n9874) );
  AND2_X1 U11015 ( .A1(n9852), .A2(n9907), .ZN(n9873) );
  INV_X1 U11016 ( .A(n9853), .ZN(n9854) );
  NAND2_X1 U11017 ( .A1(n9873), .A2(n9854), .ZN(n9855) );
  OAI21_X1 U11018 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9868) );
  XNOR2_X1 U11019 ( .A(n9858), .B(n9859), .ZN(n9866) );
  OAI22_X1 U11020 ( .A1(n9862), .A2(n9861), .B1(n5881), .B2(n9860), .ZN(n9863)
         );
  AOI21_X1 U11021 ( .B1(n9874), .B2(n9864), .A(n9863), .ZN(n9865) );
  OAI21_X1 U11022 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(n9872) );
  AOI211_X1 U11023 ( .C1(n9869), .C2(n9874), .A(n9868), .B(n9872), .ZN(n9870)
         );
  AOI22_X1 U11024 ( .A1(n9871), .A2(n6762), .B1(n9870), .B2(n8318), .ZN(
        P2_U3231) );
  INV_X1 U11025 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9876) );
  INV_X1 U11026 ( .A(n9902), .ZN(n9875) );
  AOI211_X1 U11027 ( .C1(n9875), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9918)
         );
  AOI22_X1 U11028 ( .A1(n9917), .A2(n9876), .B1(n9918), .B2(n9915), .ZN(
        P2_U3396) );
  INV_X1 U11029 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9882) );
  INV_X1 U11030 ( .A(n9877), .ZN(n9881) );
  OAI21_X1 U11031 ( .B1(n9879), .B2(n9909), .A(n9878), .ZN(n9880) );
  AOI21_X1 U11032 ( .B1(n9881), .B2(n9914), .A(n9880), .ZN(n9919) );
  AOI22_X1 U11033 ( .A1(n9917), .A2(n9882), .B1(n9919), .B2(n9915), .ZN(
        P2_U3402) );
  OAI22_X1 U11034 ( .A1(n9884), .A2(n9902), .B1(n9883), .B2(n9909), .ZN(n9885)
         );
  NOR2_X1 U11035 ( .A1(n9886), .A2(n9885), .ZN(n9921) );
  AOI22_X1 U11036 ( .A1(n9917), .A2(n5346), .B1(n9921), .B2(n9915), .ZN(
        P2_U3405) );
  NOR2_X1 U11037 ( .A1(n9888), .A2(n9887), .ZN(n9891) );
  INV_X1 U11038 ( .A(n9889), .ZN(n9890) );
  AOI211_X1 U11039 ( .C1(n9907), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9923)
         );
  AOI22_X1 U11040 ( .A1(n9917), .A2(n5368), .B1(n9923), .B2(n9915), .ZN(
        P2_U3408) );
  NOR2_X1 U11041 ( .A1(n9893), .A2(n9902), .ZN(n9895) );
  AOI211_X1 U11042 ( .C1(n9907), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9924)
         );
  AOI22_X1 U11043 ( .A1(n9917), .A2(n5393), .B1(n9924), .B2(n9915), .ZN(
        P2_U3411) );
  INV_X1 U11044 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9901) );
  NOR2_X1 U11045 ( .A1(n9897), .A2(n9909), .ZN(n9899) );
  AOI211_X1 U11046 ( .C1(n9914), .C2(n9900), .A(n9899), .B(n9898), .ZN(n9925)
         );
  AOI22_X1 U11047 ( .A1(n9917), .A2(n9901), .B1(n9925), .B2(n9915), .ZN(
        P2_U3414) );
  INV_X1 U11048 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U11049 ( .A1(n9903), .A2(n9902), .ZN(n9905) );
  AOI211_X1 U11050 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9926)
         );
  AOI22_X1 U11051 ( .A1(n9917), .A2(n9908), .B1(n9926), .B2(n9915), .ZN(
        P2_U3417) );
  INV_X1 U11052 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U11053 ( .A1(n9910), .A2(n9909), .ZN(n9912) );
  AOI211_X1 U11054 ( .C1(n9914), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9928)
         );
  AOI22_X1 U11055 ( .A1(n9917), .A2(n9916), .B1(n9928), .B2(n9915), .ZN(
        P2_U3420) );
  AOI22_X1 U11056 ( .A1(n9929), .A2(n9918), .B1(n6732), .B2(n9927), .ZN(
        P2_U3461) );
  AOI22_X1 U11057 ( .A1(n9929), .A2(n9919), .B1(n6758), .B2(n9927), .ZN(
        P2_U3463) );
  INV_X1 U11058 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U11059 ( .A1(n9929), .A2(n9921), .B1(n9920), .B2(n9927), .ZN(
        P2_U3464) );
  AOI22_X1 U11060 ( .A1(n9929), .A2(n9923), .B1(n9922), .B2(n9927), .ZN(
        P2_U3465) );
  AOI22_X1 U11061 ( .A1(n9929), .A2(n9924), .B1(n7234), .B2(n9927), .ZN(
        P2_U3466) );
  AOI22_X1 U11062 ( .A1(n9929), .A2(n9925), .B1(n7230), .B2(n9927), .ZN(
        P2_U3467) );
  AOI22_X1 U11063 ( .A1(n9929), .A2(n9926), .B1(n8134), .B2(n9927), .ZN(
        P2_U3468) );
  AOI22_X1 U11064 ( .A1(n9929), .A2(n9928), .B1(n10256), .B2(n9927), .ZN(
        P2_U3469) );
  OAI222_X1 U11065 ( .A1(n9934), .A2(n9933), .B1(n9934), .B2(n9932), .C1(n9931), .C2(n9930), .ZN(ADD_1068_U5) );
  XOR2_X1 U11066 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11067 ( .B1(n9937), .B2(n9936), .A(n9935), .ZN(n9938) );
  XNOR2_X1 U11068 ( .A(n9938), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11069 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(ADD_1068_U56) );
  OAI21_X1 U11070 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(ADD_1068_U57) );
  OAI21_X1 U11071 ( .B1(n9947), .B2(n9946), .A(n9945), .ZN(ADD_1068_U58) );
  OAI21_X1 U11072 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(ADD_1068_U59) );
  OAI21_X1 U11073 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(ADD_1068_U60) );
  OAI21_X1 U11074 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(ADD_1068_U61) );
  OAI21_X1 U11075 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(ADD_1068_U62) );
  OAI21_X1 U11076 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(ADD_1068_U63) );
  NAND2_X1 U11077 ( .A1(n9963), .A2(P2_D_REG_30__SCAN_IN), .ZN(n10284) );
  INV_X1 U11078 ( .A(keyinput40), .ZN(n9964) );
  NOR4_X1 U11079 ( .A1(keyinput58), .A2(keyinput16), .A3(keyinput125), .A4(
        n9964), .ZN(n9966) );
  INV_X1 U11080 ( .A(keyinput114), .ZN(n9965) );
  NAND4_X1 U11081 ( .A1(keyinput74), .A2(keyinput122), .A3(n9966), .A4(n9965), 
        .ZN(n9978) );
  NOR2_X1 U11082 ( .A1(keyinput49), .A2(keyinput103), .ZN(n9967) );
  NAND3_X1 U11083 ( .A1(keyinput18), .A2(keyinput118), .A3(n9967), .ZN(n9977)
         );
  INV_X1 U11084 ( .A(keyinput96), .ZN(n10264) );
  NAND4_X1 U11085 ( .A1(keyinput59), .A2(keyinput26), .A3(keyinput105), .A4(
        n10264), .ZN(n9976) );
  NAND2_X1 U11086 ( .A1(keyinput87), .A2(keyinput41), .ZN(n9968) );
  NOR3_X1 U11087 ( .A1(keyinput7), .A2(keyinput42), .A3(n9968), .ZN(n9974) );
  NOR4_X1 U11088 ( .A1(keyinput1), .A2(keyinput116), .A3(keyinput126), .A4(
        keyinput106), .ZN(n9973) );
  INV_X1 U11089 ( .A(keyinput69), .ZN(n9969) );
  NOR4_X1 U11090 ( .A1(keyinput43), .A2(keyinput111), .A3(keyinput12), .A4(
        n9969), .ZN(n9972) );
  NAND3_X1 U11091 ( .A1(keyinput6), .A2(keyinput14), .A3(keyinput2), .ZN(n9970) );
  NOR2_X1 U11092 ( .A1(keyinput72), .A2(n9970), .ZN(n9971) );
  NAND4_X1 U11093 ( .A1(n9974), .A2(n9973), .A3(n9972), .A4(n9971), .ZN(n9975)
         );
  NOR4_X1 U11094 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n10026)
         );
  INV_X1 U11095 ( .A(keyinput11), .ZN(n9979) );
  NAND4_X1 U11096 ( .A1(keyinput76), .A2(keyinput119), .A3(keyinput124), .A4(
        n9979), .ZN(n9985) );
  NOR3_X1 U11097 ( .A1(keyinput64), .A2(keyinput54), .A3(keyinput113), .ZN(
        n9980) );
  NAND2_X1 U11098 ( .A1(keyinput99), .A2(n9980), .ZN(n9984) );
  NAND4_X1 U11099 ( .A1(keyinput33), .A2(keyinput70), .A3(keyinput29), .A4(
        keyinput45), .ZN(n9983) );
  NOR3_X1 U11100 ( .A1(keyinput34), .A2(keyinput60), .A3(keyinput107), .ZN(
        n9981) );
  NAND2_X1 U11101 ( .A1(keyinput61), .A2(n9981), .ZN(n9982) );
  NOR4_X1 U11102 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n10025)
         );
  INV_X1 U11103 ( .A(keyinput19), .ZN(n9986) );
  NAND4_X1 U11104 ( .A1(keyinput5), .A2(keyinput15), .A3(keyinput98), .A4(
        n9986), .ZN(n9992) );
  NOR2_X1 U11105 ( .A1(keyinput75), .A2(keyinput22), .ZN(n9987) );
  NAND3_X1 U11106 ( .A1(keyinput27), .A2(keyinput9), .A3(n9987), .ZN(n9991) );
  NAND4_X1 U11107 ( .A1(keyinput73), .A2(keyinput17), .A3(keyinput4), .A4(
        keyinput21), .ZN(n9990) );
  NOR3_X1 U11108 ( .A1(keyinput55), .A2(keyinput53), .A3(keyinput71), .ZN(
        n9988) );
  NAND2_X1 U11109 ( .A1(keyinput121), .A2(n9988), .ZN(n9989) );
  NOR4_X1 U11110 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(n10024)
         );
  INV_X1 U11111 ( .A(keyinput89), .ZN(n9993) );
  NAND4_X1 U11112 ( .A1(keyinput102), .A2(keyinput101), .A3(keyinput56), .A4(
        n9993), .ZN(n10022) );
  NOR2_X1 U11113 ( .A1(keyinput86), .A2(keyinput44), .ZN(n9994) );
  NAND3_X1 U11114 ( .A1(keyinput47), .A2(keyinput62), .A3(n9994), .ZN(n10021)
         );
  NOR2_X1 U11115 ( .A1(keyinput92), .A2(keyinput83), .ZN(n9995) );
  NAND3_X1 U11116 ( .A1(keyinput68), .A2(keyinput30), .A3(n9995), .ZN(n9996)
         );
  NOR3_X1 U11117 ( .A1(keyinput94), .A2(keyinput63), .A3(n9996), .ZN(n10004)
         );
  INV_X1 U11118 ( .A(keyinput97), .ZN(n9997) );
  NAND4_X1 U11119 ( .A1(keyinput36), .A2(keyinput31), .A3(keyinput24), .A4(
        n9997), .ZN(n10002) );
  NAND4_X1 U11120 ( .A1(keyinput37), .A2(keyinput109), .A3(keyinput79), .A4(
        keyinput100), .ZN(n10001) );
  NAND4_X1 U11121 ( .A1(keyinput38), .A2(keyinput85), .A3(keyinput77), .A4(
        keyinput48), .ZN(n10000) );
  INV_X1 U11122 ( .A(keyinput3), .ZN(n9998) );
  NAND4_X1 U11123 ( .A1(keyinput115), .A2(keyinput32), .A3(keyinput120), .A4(
        n9998), .ZN(n9999) );
  NOR4_X1 U11124 ( .A1(n10002), .A2(n10001), .A3(n10000), .A4(n9999), .ZN(
        n10003) );
  NAND4_X1 U11125 ( .A1(keyinput93), .A2(keyinput80), .A3(n10004), .A4(n10003), 
        .ZN(n10020) );
  NAND2_X1 U11126 ( .A1(keyinput57), .A2(keyinput20), .ZN(n10005) );
  NOR3_X1 U11127 ( .A1(keyinput39), .A2(keyinput90), .A3(n10005), .ZN(n10018)
         );
  NOR4_X1 U11128 ( .A1(keyinput110), .A2(keyinput108), .A3(keyinput52), .A4(
        keyinput28), .ZN(n10017) );
  NAND2_X1 U11129 ( .A1(keyinput23), .A2(keyinput78), .ZN(n10006) );
  NOR3_X1 U11130 ( .A1(keyinput46), .A2(keyinput65), .A3(n10006), .ZN(n10007)
         );
  NAND3_X1 U11131 ( .A1(keyinput112), .A2(keyinput88), .A3(n10007), .ZN(n10008) );
  NOR3_X1 U11132 ( .A1(keyinput81), .A2(keyinput13), .A3(n10008), .ZN(n10016)
         );
  NAND4_X1 U11133 ( .A1(keyinput123), .A2(keyinput66), .A3(keyinput84), .A4(
        keyinput10), .ZN(n10014) );
  INV_X1 U11134 ( .A(keyinput91), .ZN(n10009) );
  NAND4_X1 U11135 ( .A1(keyinput127), .A2(keyinput95), .A3(keyinput0), .A4(
        n10009), .ZN(n10013) );
  NOR3_X1 U11136 ( .A1(keyinput50), .A2(keyinput82), .A3(keyinput67), .ZN(
        n10010) );
  NAND2_X1 U11137 ( .A1(keyinput117), .A2(n10010), .ZN(n10012) );
  NAND4_X1 U11138 ( .A1(keyinput35), .A2(keyinput104), .A3(keyinput8), .A4(
        keyinput51), .ZN(n10011) );
  NOR4_X1 U11139 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10015) );
  NAND4_X1 U11140 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n10019) );
  NOR4_X1 U11141 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10023) );
  NAND4_X1 U11142 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10281) );
  AOI22_X1 U11143 ( .A1(n10029), .A2(keyinput83), .B1(keyinput86), .B2(n10028), 
        .ZN(n10027) );
  OAI221_X1 U11144 ( .B1(n10029), .B2(keyinput83), .C1(n10028), .C2(keyinput86), .A(n10027), .ZN(n10042) );
  AOI22_X1 U11145 ( .A1(n10032), .A2(keyinput63), .B1(n10031), .B2(keyinput30), 
        .ZN(n10030) );
  OAI221_X1 U11146 ( .B1(n10032), .B2(keyinput63), .C1(n10031), .C2(keyinput30), .A(n10030), .ZN(n10041) );
  INV_X1 U11147 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U11148 ( .A1(n10035), .A2(keyinput80), .B1(n10034), .B2(keyinput94), 
        .ZN(n10033) );
  OAI221_X1 U11149 ( .B1(n10035), .B2(keyinput80), .C1(n10034), .C2(keyinput94), .A(n10033), .ZN(n10040) );
  INV_X1 U11150 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10036) );
  XOR2_X1 U11151 ( .A(n10036), .B(keyinput92), .Z(n10038) );
  XNOR2_X1 U11152 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput93), .ZN(n10037) );
  NAND2_X1 U11153 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  NOR4_X1 U11154 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10087) );
  AOI22_X1 U11155 ( .A1(n6801), .A2(keyinput44), .B1(n10044), .B2(keyinput89), 
        .ZN(n10043) );
  OAI221_X1 U11156 ( .B1(n6801), .B2(keyinput44), .C1(n10044), .C2(keyinput89), 
        .A(n10043), .ZN(n10052) );
  XOR2_X1 U11157 ( .A(P2_REG2_REG_30__SCAN_IN), .B(keyinput37), .Z(n10051) );
  XOR2_X1 U11158 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput56), .Z(n10050) );
  XNOR2_X1 U11159 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput62), .ZN(n10048) );
  XNOR2_X1 U11160 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput47), .ZN(n10047)
         );
  XNOR2_X1 U11161 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput101), .ZN(n10046) );
  XNOR2_X1 U11162 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput102), .ZN(n10045)
         );
  NAND4_X1 U11163 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10049) );
  NOR4_X1 U11164 ( .A1(n10052), .A2(n10051), .A3(n10050), .A4(n10049), .ZN(
        n10086) );
  AOI22_X1 U11165 ( .A1(n10055), .A2(keyinput24), .B1(keyinput115), .B2(n10054), .ZN(n10053) );
  OAI221_X1 U11166 ( .B1(n10055), .B2(keyinput24), .C1(n10054), .C2(
        keyinput115), .A(n10053), .ZN(n10068) );
  AOI22_X1 U11167 ( .A1(n10058), .A2(keyinput100), .B1(n10057), .B2(keyinput31), .ZN(n10056) );
  OAI221_X1 U11168 ( .B1(n10058), .B2(keyinput100), .C1(n10057), .C2(
        keyinput31), .A(n10056), .ZN(n10067) );
  AOI22_X1 U11169 ( .A1(n10061), .A2(keyinput109), .B1(keyinput79), .B2(n10060), .ZN(n10059) );
  OAI221_X1 U11170 ( .B1(n10061), .B2(keyinput109), .C1(n10060), .C2(
        keyinput79), .A(n10059), .ZN(n10066) );
  XOR2_X1 U11171 ( .A(n10062), .B(keyinput97), .Z(n10064) );
  XNOR2_X1 U11172 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput36), .ZN(n10063)
         );
  NAND2_X1 U11173 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  NOR4_X1 U11174 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(
        n10085) );
  AOI22_X1 U11175 ( .A1(n10071), .A2(keyinput3), .B1(n10070), .B2(keyinput32), 
        .ZN(n10069) );
  OAI221_X1 U11176 ( .B1(n10071), .B2(keyinput3), .C1(n10070), .C2(keyinput32), 
        .A(n10069), .ZN(n10083) );
  AOI22_X1 U11177 ( .A1(n5094), .A2(keyinput120), .B1(keyinput38), .B2(n10073), 
        .ZN(n10072) );
  OAI221_X1 U11178 ( .B1(n5094), .B2(keyinput120), .C1(n10073), .C2(keyinput38), .A(n10072), .ZN(n10082) );
  AOI22_X1 U11179 ( .A1(n10076), .A2(keyinput85), .B1(n10075), .B2(keyinput77), 
        .ZN(n10074) );
  OAI221_X1 U11180 ( .B1(n10076), .B2(keyinput85), .C1(n10075), .C2(keyinput77), .A(n10074), .ZN(n10081) );
  AOI22_X1 U11181 ( .A1(n10079), .A2(keyinput48), .B1(n10078), .B2(keyinput95), 
        .ZN(n10077) );
  OAI221_X1 U11182 ( .B1(n10079), .B2(keyinput48), .C1(n10078), .C2(keyinput95), .A(n10077), .ZN(n10080) );
  NOR4_X1 U11183 ( .A1(n10083), .A2(n10082), .A3(n10081), .A4(n10080), .ZN(
        n10084) );
  NAND4_X1 U11184 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10279) );
  AOI22_X1 U11185 ( .A1(n10090), .A2(keyinput66), .B1(n10089), .B2(keyinput84), 
        .ZN(n10088) );
  OAI221_X1 U11186 ( .B1(n10090), .B2(keyinput66), .C1(n10089), .C2(keyinput84), .A(n10088), .ZN(n10103) );
  INV_X1 U11187 ( .A(SI_29_), .ZN(n10093) );
  AOI22_X1 U11188 ( .A1(n10093), .A2(keyinput127), .B1(n10092), .B2(keyinput91), .ZN(n10091) );
  OAI221_X1 U11189 ( .B1(n10093), .B2(keyinput127), .C1(n10092), .C2(
        keyinput91), .A(n10091), .ZN(n10102) );
  AOI22_X1 U11190 ( .A1(n10096), .A2(keyinput0), .B1(n10095), .B2(keyinput123), 
        .ZN(n10094) );
  OAI221_X1 U11191 ( .B1(n10096), .B2(keyinput0), .C1(n10095), .C2(keyinput123), .A(n10094), .ZN(n10101) );
  INV_X1 U11192 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10097) );
  XOR2_X1 U11193 ( .A(n10097), .B(keyinput110), .Z(n10099) );
  XNOR2_X1 U11194 ( .A(SI_7_), .B(keyinput10), .ZN(n10098) );
  NAND2_X1 U11195 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NOR4_X1 U11196 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10151) );
  AOI22_X1 U11197 ( .A1(n10105), .A2(keyinput108), .B1(n6629), .B2(keyinput52), 
        .ZN(n10104) );
  OAI221_X1 U11198 ( .B1(n10105), .B2(keyinput108), .C1(n6629), .C2(keyinput52), .A(n10104), .ZN(n10109) );
  XNOR2_X1 U11199 ( .A(n10106), .B(keyinput90), .ZN(n10108) );
  XOR2_X1 U11200 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput39), .Z(n10107) );
  OR3_X1 U11201 ( .A1(n10109), .A2(n10108), .A3(n10107), .ZN(n10118) );
  AOI22_X1 U11202 ( .A1(n10112), .A2(keyinput57), .B1(n10111), .B2(keyinput35), 
        .ZN(n10110) );
  OAI221_X1 U11203 ( .B1(n10112), .B2(keyinput57), .C1(n10111), .C2(keyinput35), .A(n10110), .ZN(n10117) );
  AOI22_X1 U11204 ( .A1(n10115), .A2(keyinput28), .B1(n10114), .B2(keyinput20), 
        .ZN(n10113) );
  OAI221_X1 U11205 ( .B1(n10115), .B2(keyinput28), .C1(n10114), .C2(keyinput20), .A(n10113), .ZN(n10116) );
  NOR3_X1 U11206 ( .A1(n10118), .A2(n10117), .A3(n10116), .ZN(n10150) );
  AOI22_X1 U11207 ( .A1(n10121), .A2(keyinput104), .B1(keyinput50), .B2(n10120), .ZN(n10119) );
  OAI221_X1 U11208 ( .B1(n10121), .B2(keyinput104), .C1(n10120), .C2(
        keyinput50), .A(n10119), .ZN(n10133) );
  AOI22_X1 U11209 ( .A1(n10124), .A2(keyinput67), .B1(keyinput8), .B2(n10123), 
        .ZN(n10122) );
  OAI221_X1 U11210 ( .B1(n10124), .B2(keyinput67), .C1(n10123), .C2(keyinput8), 
        .A(n10122), .ZN(n10132) );
  AOI22_X1 U11211 ( .A1(n10126), .A2(keyinput51), .B1(n8083), .B2(keyinput82), 
        .ZN(n10125) );
  OAI221_X1 U11212 ( .B1(n10126), .B2(keyinput51), .C1(n8083), .C2(keyinput82), 
        .A(n10125), .ZN(n10131) );
  AOI22_X1 U11213 ( .A1(n10129), .A2(keyinput117), .B1(n10128), .B2(keyinput46), .ZN(n10127) );
  OAI221_X1 U11214 ( .B1(n10129), .B2(keyinput117), .C1(n10128), .C2(
        keyinput46), .A(n10127), .ZN(n10130) );
  NOR4_X1 U11215 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10149) );
  INV_X1 U11216 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10136) );
  INV_X1 U11217 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U11218 ( .A1(n10136), .A2(keyinput122), .B1(n10135), .B2(keyinput13), .ZN(n10134) );
  OAI221_X1 U11219 ( .B1(n10136), .B2(keyinput122), .C1(n10135), .C2(
        keyinput13), .A(n10134), .ZN(n10147) );
  AOI22_X1 U11220 ( .A1(n10139), .A2(keyinput88), .B1(n10138), .B2(keyinput65), 
        .ZN(n10137) );
  OAI221_X1 U11221 ( .B1(n10139), .B2(keyinput88), .C1(n10138), .C2(keyinput65), .A(n10137), .ZN(n10146) );
  INV_X1 U11222 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10140) );
  XOR2_X1 U11223 ( .A(n10140), .B(keyinput112), .Z(n10144) );
  XNOR2_X1 U11224 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput78), .ZN(n10143) );
  XNOR2_X1 U11225 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput23), .ZN(n10142) );
  XNOR2_X1 U11226 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput81), .ZN(n10141)
         );
  NAND4_X1 U11227 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10145) );
  NOR3_X1 U11228 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10148) );
  NAND4_X1 U11229 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10278) );
  AOI22_X1 U11230 ( .A1(n10154), .A2(keyinput17), .B1(n10153), .B2(keyinput4), 
        .ZN(n10152) );
  OAI221_X1 U11231 ( .B1(n10154), .B2(keyinput17), .C1(n10153), .C2(keyinput4), 
        .A(n10152), .ZN(n10166) );
  AOI22_X1 U11232 ( .A1(n10156), .A2(keyinput121), .B1(n5210), .B2(keyinput73), 
        .ZN(n10155) );
  OAI221_X1 U11233 ( .B1(n10156), .B2(keyinput121), .C1(n5210), .C2(keyinput73), .A(n10155), .ZN(n10165) );
  AOI22_X1 U11234 ( .A1(n10159), .A2(keyinput53), .B1(n10158), .B2(keyinput99), 
        .ZN(n10157) );
  OAI221_X1 U11235 ( .B1(n10159), .B2(keyinput53), .C1(n10158), .C2(keyinput99), .A(n10157), .ZN(n10164) );
  AOI22_X1 U11236 ( .A1(n10162), .A2(keyinput21), .B1(n10161), .B2(keyinput71), 
        .ZN(n10160) );
  OAI221_X1 U11237 ( .B1(n10162), .B2(keyinput21), .C1(n10161), .C2(keyinput71), .A(n10160), .ZN(n10163) );
  NOR4_X1 U11238 ( .A1(n10166), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10215) );
  AOI22_X1 U11239 ( .A1(n10169), .A2(keyinput9), .B1(keyinput15), .B2(n10168), 
        .ZN(n10167) );
  OAI221_X1 U11240 ( .B1(n10169), .B2(keyinput9), .C1(n10168), .C2(keyinput15), 
        .A(n10167), .ZN(n10180) );
  AOI22_X1 U11241 ( .A1(n10171), .A2(keyinput27), .B1(n5393), .B2(keyinput22), 
        .ZN(n10170) );
  OAI221_X1 U11242 ( .B1(n10171), .B2(keyinput27), .C1(n5393), .C2(keyinput22), 
        .A(n10170), .ZN(n10179) );
  INV_X1 U11243 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U11244 ( .A1(n7806), .A2(keyinput98), .B1(keyinput55), .B2(n10173), 
        .ZN(n10172) );
  OAI221_X1 U11245 ( .B1(n7806), .B2(keyinput98), .C1(n10173), .C2(keyinput55), 
        .A(n10172), .ZN(n10178) );
  AOI22_X1 U11246 ( .A1(n10176), .A2(keyinput5), .B1(n10175), .B2(keyinput19), 
        .ZN(n10174) );
  OAI221_X1 U11247 ( .B1(n10176), .B2(keyinput5), .C1(n10175), .C2(keyinput19), 
        .A(n10174), .ZN(n10177) );
  NOR4_X1 U11248 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10214) );
  AOI22_X1 U11249 ( .A1(n10183), .A2(keyinput45), .B1(keyinput107), .B2(n10182), .ZN(n10181) );
  OAI221_X1 U11250 ( .B1(n10183), .B2(keyinput45), .C1(n10182), .C2(
        keyinput107), .A(n10181), .ZN(n10187) );
  XNOR2_X1 U11251 ( .A(n10184), .B(keyinput60), .ZN(n10186) );
  XOR2_X1 U11252 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput68), .Z(n10185) );
  OR3_X1 U11253 ( .A1(n10187), .A2(n10186), .A3(n10185), .ZN(n10196) );
  INV_X1 U11254 ( .A(keyinput33), .ZN(n10189) );
  AOI22_X1 U11255 ( .A1(n10190), .A2(keyinput61), .B1(P2_WR_REG_SCAN_IN), .B2(
        n10189), .ZN(n10188) );
  OAI221_X1 U11256 ( .B1(n10190), .B2(keyinput61), .C1(n10189), .C2(
        P2_WR_REG_SCAN_IN), .A(n10188), .ZN(n10195) );
  AOI22_X1 U11257 ( .A1(n10193), .A2(keyinput70), .B1(keyinput29), .B2(n10192), 
        .ZN(n10191) );
  OAI221_X1 U11258 ( .B1(n10193), .B2(keyinput70), .C1(n10192), .C2(keyinput29), .A(n10191), .ZN(n10194) );
  NOR3_X1 U11259 ( .A1(n10196), .A2(n10195), .A3(n10194), .ZN(n10213) );
  INV_X1 U11260 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U11261 ( .A1(n10199), .A2(keyinput54), .B1(n10198), .B2(keyinput76), 
        .ZN(n10197) );
  OAI221_X1 U11262 ( .B1(n10199), .B2(keyinput54), .C1(n10198), .C2(keyinput76), .A(n10197), .ZN(n10211) );
  INV_X1 U11263 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U11264 ( .A1(n10202), .A2(keyinput11), .B1(n10201), .B2(keyinput119), .ZN(n10200) );
  OAI221_X1 U11265 ( .B1(n10202), .B2(keyinput11), .C1(n10201), .C2(
        keyinput119), .A(n10200), .ZN(n10210) );
  AOI22_X1 U11266 ( .A1(n10205), .A2(keyinput124), .B1(n10204), .B2(keyinput34), .ZN(n10203) );
  OAI221_X1 U11267 ( .B1(n10205), .B2(keyinput124), .C1(n10204), .C2(
        keyinput34), .A(n10203), .ZN(n10209) );
  XNOR2_X1 U11268 ( .A(P1_REG0_REG_15__SCAN_IN), .B(keyinput113), .ZN(n10207)
         );
  XNOR2_X1 U11269 ( .A(SI_1_), .B(keyinput64), .ZN(n10206) );
  NAND2_X1 U11270 ( .A1(n10207), .A2(n10206), .ZN(n10208) );
  NOR4_X1 U11271 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10212) );
  NAND4_X1 U11272 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10277) );
  AOI22_X1 U11273 ( .A1(n10217), .A2(keyinput106), .B1(keyinput87), .B2(n8586), 
        .ZN(n10216) );
  OAI221_X1 U11274 ( .B1(n10217), .B2(keyinput106), .C1(n8586), .C2(keyinput87), .A(n10216), .ZN(n10226) );
  AOI22_X1 U11275 ( .A1(n8496), .A2(keyinput42), .B1(n10219), .B2(keyinput59), 
        .ZN(n10218) );
  OAI221_X1 U11276 ( .B1(n8496), .B2(keyinput42), .C1(n10219), .C2(keyinput59), 
        .A(n10218), .ZN(n10225) );
  XNOR2_X1 U11277 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput126), .ZN(n10223)
         );
  XNOR2_X1 U11278 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput41), .ZN(n10222)
         );
  XNOR2_X1 U11279 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput116), .ZN(n10221) );
  XNOR2_X1 U11280 ( .A(keyinput7), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n10220) );
  NAND4_X1 U11281 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10224) );
  NOR3_X1 U11282 ( .A1(n10226), .A2(n10225), .A3(n10224), .ZN(n10275) );
  AOI22_X1 U11283 ( .A1(n10228), .A2(keyinput74), .B1(keyinput114), .B2(n6839), 
        .ZN(n10227) );
  OAI221_X1 U11284 ( .B1(n10228), .B2(keyinput74), .C1(n6839), .C2(keyinput114), .A(n10227), .ZN(n10239) );
  INV_X1 U11285 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U11286 ( .A1(n10231), .A2(keyinput16), .B1(keyinput58), .B2(n10230), 
        .ZN(n10229) );
  OAI221_X1 U11287 ( .B1(n10231), .B2(keyinput16), .C1(n10230), .C2(keyinput58), .A(n10229), .ZN(n10238) );
  INV_X1 U11288 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11289 ( .A1(keyinput40), .A2(n10233), .B1(keyinput25), .B2(n10282), 
        .ZN(n10232) );
  OAI21_X1 U11290 ( .B1(n10233), .B2(keyinput40), .A(n10232), .ZN(n10237) );
  XNOR2_X1 U11291 ( .A(P1_REG3_REG_26__SCAN_IN), .B(keyinput1), .ZN(n10235) );
  XNOR2_X1 U11292 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput125), .ZN(n10234)
         );
  NAND2_X1 U11293 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  NOR4_X1 U11294 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10274) );
  AOI22_X1 U11295 ( .A1(n10242), .A2(keyinput72), .B1(n10241), .B2(keyinput43), 
        .ZN(n10240) );
  OAI221_X1 U11296 ( .B1(n10242), .B2(keyinput72), .C1(n10241), .C2(keyinput43), .A(n10240), .ZN(n10254) );
  INV_X1 U11297 ( .A(SI_24_), .ZN(n10245) );
  AOI22_X1 U11298 ( .A1(n10245), .A2(keyinput2), .B1(keyinput6), .B2(n10244), 
        .ZN(n10243) );
  OAI221_X1 U11299 ( .B1(n10245), .B2(keyinput2), .C1(n10244), .C2(keyinput6), 
        .A(n10243), .ZN(n10253) );
  AOI22_X1 U11300 ( .A1(n10248), .A2(keyinput12), .B1(keyinput75), .B2(n10247), 
        .ZN(n10246) );
  OAI221_X1 U11301 ( .B1(n10248), .B2(keyinput12), .C1(n10247), .C2(keyinput75), .A(n10246), .ZN(n10252) );
  AOI22_X1 U11302 ( .A1(n5224), .A2(keyinput111), .B1(keyinput69), .B2(n10250), 
        .ZN(n10249) );
  OAI221_X1 U11303 ( .B1(n5224), .B2(keyinput111), .C1(n10250), .C2(keyinput69), .A(n10249), .ZN(n10251) );
  NOR4_X1 U11304 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n10273) );
  AOI22_X1 U11305 ( .A1(n10257), .A2(keyinput103), .B1(n10256), .B2(keyinput14), .ZN(n10255) );
  OAI221_X1 U11306 ( .B1(n10257), .B2(keyinput103), .C1(n10256), .C2(
        keyinput14), .A(n10255), .ZN(n10271) );
  AOI22_X1 U11307 ( .A1(n10260), .A2(keyinput105), .B1(keyinput18), .B2(n10259), .ZN(n10258) );
  OAI221_X1 U11308 ( .B1(n10260), .B2(keyinput105), .C1(n10259), .C2(
        keyinput18), .A(n10258), .ZN(n10270) );
  AOI22_X1 U11309 ( .A1(n10263), .A2(keyinput49), .B1(keyinput118), .B2(n10262), .ZN(n10261) );
  OAI221_X1 U11310 ( .B1(n10263), .B2(keyinput49), .C1(n10262), .C2(
        keyinput118), .A(n10261), .ZN(n10268) );
  XNOR2_X1 U11311 ( .A(n10264), .B(P1_WR_REG_SCAN_IN), .ZN(n10267) );
  XNOR2_X1 U11312 ( .A(n10265), .B(keyinput26), .ZN(n10266) );
  OR3_X1 U11313 ( .A1(n10268), .A2(n10267), .A3(n10266), .ZN(n10269) );
  NOR3_X1 U11314 ( .A1(n10271), .A2(n10270), .A3(n10269), .ZN(n10272) );
  NAND4_X1 U11315 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10276) );
  NOR4_X1 U11316 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  OAI221_X1 U11317 ( .B1(keyinput25), .B2(n10282), .C1(keyinput25), .C2(n10281), .A(n10280), .ZN(n10283) );
  XOR2_X1 U11318 ( .A(n10284), .B(n10283), .Z(P2_U3235) );
  OAI21_X1 U11319 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(ADD_1068_U50) );
  OAI21_X1 U11320 ( .B1(n10290), .B2(n10289), .A(n10288), .ZN(ADD_1068_U51) );
  OAI21_X1 U11321 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(ADD_1068_U47) );
  OAI21_X1 U11322 ( .B1(n10296), .B2(n10295), .A(n10294), .ZN(ADD_1068_U49) );
  OAI21_X1 U11323 ( .B1(n10299), .B2(n10298), .A(n10297), .ZN(ADD_1068_U48) );
  AOI21_X1 U11324 ( .B1(n10302), .B2(n10301), .A(n10300), .ZN(ADD_1068_U54) );
  AOI21_X1 U11325 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(ADD_1068_U53) );
  OAI21_X1 U11326 ( .B1(n10308), .B2(n10307), .A(n10306), .ZN(ADD_1068_U52) );
  INV_X2 U4998 ( .A(n6484), .ZN(n6497) );
  CLKBUF_X1 U5160 ( .A(n7960), .Z(n7917) );
endmodule

